

module b17_C_AntiSAT_k_128_3 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9650, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076;

  NAND2_X1 U11094 ( .A1(n15238), .A2(n15237), .ZN(n15236) );
  NAND2_X1 U11095 ( .A1(n10886), .A2(n10013), .ZN(n15390) );
  AOI21_X1 U11096 ( .B1(n19052), .B2(n19055), .A(n19051), .ZN(n19047) );
  CLKBUF_X1 U11097 ( .A(n11983), .Z(n14356) );
  INV_X1 U11098 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20697) );
  OR3_X1 U11099 ( .A1(n10458), .A2(n11439), .A3(n10450), .ZN(n10684) );
  OR2_X1 U11100 ( .A1(n10454), .A2(n15894), .ZN(n10628) );
  INV_X1 U11102 ( .A(n14037), .ZN(n16041) );
  CLKBUF_X2 U11103 ( .A(n13963), .Z(n17489) );
  INV_X1 U11104 ( .A(n17538), .ZN(n17571) );
  INV_X1 U11105 ( .A(n9720), .ZN(n17441) );
  CLKBUF_X1 U11106 ( .A(n13950), .Z(n17554) );
  INV_X1 U11107 ( .A(n10582), .ZN(n11007) );
  CLKBUF_X1 U11109 ( .A(n13963), .Z(n17580) );
  INV_X1 U11110 ( .A(n17458), .ZN(n16022) );
  INV_X1 U11111 ( .A(n17538), .ZN(n17524) );
  NOR2_X1 U11112 ( .A1(n13884), .A2(n13883), .ZN(n13964) );
  NOR2_X1 U11113 ( .A1(n13881), .A2(n13883), .ZN(n13950) );
  CLKBUF_X2 U11114 ( .A(n12218), .Z(n9670) );
  CLKBUF_X2 U11115 ( .A(n12212), .Z(n11948) );
  AND3_X1 U11116 ( .A1(n11944), .A2(n11943), .A3(n11942), .ZN(n11945) );
  NAND2_X2 U11117 ( .A1(n19232), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13881) );
  INV_X2 U11118 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19227) );
  AND2_X1 U11119 ( .A1(n11674), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10515) );
  AND2_X1 U11120 ( .A1(n11666), .A2(n9802), .ZN(n11201) );
  AND2_X1 U11121 ( .A1(n11587), .A2(n10476), .ZN(n11618) );
  AND2_X1 U11122 ( .A1(n11587), .A2(n10477), .ZN(n11464) );
  INV_X1 U11123 ( .A(n9718), .ZN(n11288) );
  INV_X1 U11124 ( .A(n9715), .ZN(n11617) );
  CLKBUF_X2 U11125 ( .A(n11947), .Z(n14366) );
  INV_X2 U11126 ( .A(n20279), .ZN(n11070) );
  CLKBUF_X3 U11127 ( .A(n11947), .Z(n14338) );
  AND2_X1 U11128 ( .A1(n11878), .A2(n11881), .ZN(n12211) );
  AND2_X1 U11129 ( .A1(n11880), .A2(n11879), .ZN(n12212) );
  NAND2_X2 U11130 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19219), .ZN(
        n13882) );
  CLKBUF_X1 U11132 ( .A(n12656), .Z(n9650) );
  NOR2_X1 U11133 ( .A1(n14482), .A2(n14888), .ZN(n12656) );
  NOR2_X1 U11134 ( .A1(n21075), .A2(n21076), .ZN(n17333) );
  INV_X2 U11139 ( .A(n18476), .ZN(n18481) );
  CLKBUF_X1 U11140 ( .A(n18785), .Z(n9655) );
  NOR2_X1 U11141 ( .A1(n19075), .A2(n18772), .ZN(n18785) );
  CLKBUF_X1 U11142 ( .A(n12909), .Z(n9656) );
  NOR2_X1 U11143 ( .A1(n14888), .A2(n14475), .ZN(n12909) );
  OR2_X1 U11144 ( .A1(n19543), .A2(n19544), .ZN(n19584) );
  INV_X1 U11145 ( .A(n19584), .ZN(n9657) );
  AND2_X1 U11146 ( .A1(n10657), .A2(n10656), .ZN(n10669) );
  NOR2_X2 U11147 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11881) );
  INV_X1 U11148 ( .A(n11585), .ZN(n10485) );
  AND2_X1 U11149 ( .A1(n13592), .A2(n10135), .ZN(n9881) );
  AND2_X2 U11150 ( .A1(n15883), .A2(n10572), .ZN(n10484) );
  AND2_X1 U11151 ( .A1(n12800), .A2(n11882), .ZN(n12200) );
  INV_X1 U11152 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U11153 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19207), .ZN(
        n13883) );
  INV_X1 U11154 ( .A(n17405), .ZN(n16040) );
  INV_X1 U11155 ( .A(n10251), .ZN(n16010) );
  NAND2_X1 U11156 ( .A1(n19227), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13884) );
  INV_X1 U11157 ( .A(n13723), .ZN(n14806) );
  INV_X1 U11158 ( .A(n10372), .ZN(n11423) );
  INV_X2 U11159 ( .A(n10582), .ZN(n11821) );
  AND2_X1 U11160 ( .A1(n10350), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11564) );
  BUF_X1 U11161 ( .A(n10902), .Z(n11021) );
  OR2_X1 U11162 ( .A1(n12837), .A2(n12469), .ZN(n12564) );
  XNOR2_X1 U11163 ( .A(n10715), .B(n15846), .ZN(n13592) );
  OR2_X1 U11164 ( .A1(n14551), .A2(n14535), .ZN(n14537) );
  NOR2_X1 U11165 ( .A1(n20370), .A2(n13059), .ZN(n13358) );
  OR2_X2 U11166 ( .A1(n11958), .A2(n11957), .ZN(n13019) );
  NAND2_X1 U11167 ( .A1(n11045), .A2(n13262), .ZN(n11349) );
  OR2_X1 U11168 ( .A1(n12827), .A2(n12826), .ZN(n13094) );
  NAND2_X1 U11169 ( .A1(n15300), .A2(n15299), .ZN(n15302) );
  INV_X1 U11170 ( .A(n18170), .ZN(n18156) );
  AOI221_X1 U11171 ( .B1(n18052), .B2(n18286), .C1(n17942), .C2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n17941), .ZN(n17927) );
  NAND2_X1 U11172 ( .A1(n19055), .A2(n15970), .ZN(n18585) );
  INV_X1 U11173 ( .A(n20322), .ZN(n20384) );
  XNOR2_X1 U11174 ( .A(n11023), .B(n11022), .ZN(n16525) );
  INV_X1 U11175 ( .A(n10437), .ZN(n12104) );
  OR2_X1 U11176 ( .A1(n13882), .A2(n13884), .ZN(n9658) );
  CLKBUF_X3 U11177 ( .A(n11913), .Z(n9675) );
  NAND2_X2 U11178 ( .A1(n13617), .A2(n13616), .ZN(n13619) );
  AND2_X2 U11179 ( .A1(n20452), .A2(n9813), .ZN(n9812) );
  BUF_X4 U11180 ( .A(n16723), .Z(n9659) );
  INV_X2 U11181 ( .A(n20281), .ZN(n16723) );
  NAND2_X4 U11182 ( .A1(n13654), .A2(n13653), .ZN(n13723) );
  CLKBUF_X3 U11183 ( .A(n19047), .Z(n9660) );
  NOR2_X2 U11184 ( .A1(n10659), .A2(n10029), .ZN(n10028) );
  NAND2_X2 U11185 ( .A1(n10588), .A2(n10587), .ZN(n10659) );
  XNOR2_X2 U11186 ( .A(n13629), .B(n13725), .ZN(n16385) );
  NAND2_X2 U11187 ( .A1(n20451), .A2(n13620), .ZN(n16386) );
  NAND2_X2 U11188 ( .A1(n9795), .A2(n10437), .ZN(n10461) );
  NAND2_X2 U11189 ( .A1(n10330), .A2(n10329), .ZN(n10385) );
  NOR2_X2 U11190 ( .A1(n16084), .A2(n18232), .ZN(n16086) );
  INV_X2 U11191 ( .A(n10265), .ZN(n10345) );
  INV_X2 U11192 ( .A(n13019), .ZN(n13024) );
  AND2_X4 U11193 ( .A1(n9842), .A2(n12294), .ZN(n14419) );
  BUF_X4 U11194 ( .A(n13308), .Z(n9661) );
  AND2_X4 U11195 ( .A1(n10489), .A2(n10259), .ZN(n11666) );
  BUF_X2 U11196 ( .A(n11638), .Z(n9662) );
  BUF_X2 U11197 ( .A(n11638), .Z(n9663) );
  BUF_X4 U11198 ( .A(n11638), .Z(n9664) );
  NOR2_X2 U11199 ( .A1(n14525), .A2(n14488), .ZN(n14513) );
  AND2_X1 U11200 ( .A1(n15883), .A2(n10572), .ZN(n9665) );
  INV_X2 U11201 ( .A(n14037), .ZN(n9666) );
  AOI221_X2 U11202 ( .B1(n18380), .B2(n18560), .C1(n18372), .C2(n18560), .A(
        n18371), .ZN(n18379) );
  XNOR2_X1 U11203 ( .A(n11013), .B(n13235), .ZN(n11419) );
  AND2_X1 U11204 ( .A1(n11736), .A2(n9911), .ZN(n15238) );
  AND2_X2 U11205 ( .A1(n16269), .A2(n9767), .ZN(n14533) );
  AND2_X1 U11206 ( .A1(n10871), .A2(n15846), .ZN(n10872) );
  AND2_X1 U11207 ( .A1(n16138), .A2(n10079), .ZN(n16188) );
  OR2_X1 U11208 ( .A1(n15300), .A2(n11396), .ZN(n16552) );
  OR2_X1 U11209 ( .A1(n15435), .A2(n10802), .ZN(n9907) );
  NAND2_X1 U11210 ( .A1(n10072), .A2(n10070), .ZN(n15085) );
  INV_X1 U11211 ( .A(n15363), .ZN(n10072) );
  NAND2_X1 U11212 ( .A1(n9778), .A2(n11455), .ZN(n12562) );
  NOR4_X1 U11213 ( .A1(n15463), .A2(n15456), .A3(n15460), .A4(n15533), .ZN(
        n10769) );
  CLKBUF_X2 U11214 ( .A(n12616), .Z(n9680) );
  BUF_X1 U11215 ( .A(n10621), .Z(n19894) );
  BUF_X1 U11216 ( .A(n10619), .Z(n19836) );
  OR2_X1 U11217 ( .A1(n10793), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U11218 ( .A1(n12670), .A2(n12600), .ZN(n12616) );
  AND2_X1 U11219 ( .A1(n10442), .A2(n15894), .ZN(n10466) );
  NAND2_X1 U11220 ( .A1(n10463), .A2(n15894), .ZN(n19982) );
  OR2_X1 U11221 ( .A1(n10462), .A2(n10458), .ZN(n19865) );
  NOR2_X2 U11222 ( .A1(n10759), .A2(n10755), .ZN(n10770) );
  CLKBUF_X2 U11223 ( .A(n10451), .Z(n11439) );
  NAND2_X1 U11224 ( .A1(n18122), .A2(n16126), .ZN(n18497) );
  OR3_X1 U11225 ( .A1(n13025), .A2(n13024), .A3(n13023), .ZN(n16239) );
  INV_X2 U11226 ( .A(n18451), .ZN(n19037) );
  AOI21_X2 U11227 ( .B1(n13234), .B2(n20278), .A(n10048), .ZN(n13308) );
  AOI21_X2 U11228 ( .B1(n16212), .B2(n16211), .A(n19254), .ZN(n17631) );
  NOR2_X1 U11229 ( .A1(n17082), .A2(n17261), .ZN(n17075) );
  INV_X2 U11230 ( .A(n11301), .ZN(n10052) );
  INV_X1 U11231 ( .A(n10413), .ZN(n10890) );
  NAND2_X1 U11232 ( .A1(n18609), .A2(n17717), .ZN(n15955) );
  INV_X1 U11233 ( .A(n16081), .ZN(n17775) );
  INV_X1 U11234 ( .A(n16102), .ZN(n18633) );
  INV_X4 U11235 ( .A(n18639), .ZN(n17717) );
  NAND2_X2 U11236 ( .A1(n11979), .A2(n12539), .ZN(n12050) );
  INV_X2 U11237 ( .A(n10385), .ZN(n10582) );
  AOI211_X1 U11238 ( .C1(n9669), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n13930), .B(n13929), .ZN(n13931) );
  INV_X1 U11239 ( .A(n9658), .ZN(n9679) );
  INV_X2 U11240 ( .A(n9658), .ZN(n9669) );
  BUF_X2 U11241 ( .A(n11923), .Z(n14219) );
  CLKBUF_X2 U11242 ( .A(n13964), .Z(n17561) );
  BUF_X2 U11243 ( .A(n10483), .Z(n11793) );
  CLKBUF_X2 U11244 ( .A(n13986), .Z(n17471) );
  BUF_X2 U11245 ( .A(n12217), .Z(n9686) );
  CLKBUF_X2 U11246 ( .A(n12198), .Z(n12199) );
  CLKBUF_X2 U11247 ( .A(n12211), .Z(n14365) );
  AND2_X2 U11248 ( .A1(n12797), .A2(n11878), .ZN(n12198) );
  AND2_X2 U11249 ( .A1(n11880), .A2(n11878), .ZN(n12217) );
  INV_X1 U11250 ( .A(n9714), .ZN(n17501) );
  BUF_X4 U11252 ( .A(n14024), .Z(n9667) );
  CLKBUF_X2 U11253 ( .A(n12200), .Z(n14359) );
  CLKBUF_X2 U11254 ( .A(n10350), .Z(n11792) );
  AND3_X1 U11255 ( .A1(n12798), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n12376), .ZN(n11913) );
  AND2_X1 U11256 ( .A1(n12329), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11878) );
  NOR2_X1 U11257 ( .A1(n12329), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11879) );
  OR2_X1 U11258 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17321) );
  OR2_X1 U11259 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13879) );
  CLKBUF_X2 U11260 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15871) );
  OAI211_X1 U11261 ( .C1(n15618), .C2(n9895), .A(n9893), .B(n9894), .ZN(n11394) );
  OAI211_X1 U11262 ( .C1(n10134), .C2(n10128), .A(n10127), .B(n10242), .ZN(
        n11012) );
  OAI21_X1 U11263 ( .B1(n11404), .B2(n19532), .A(n10986), .ZN(n10987) );
  OAI21_X1 U11264 ( .B1(n11419), .B2(n16710), .A(n9695), .ZN(n11420) );
  OAI211_X1 U11265 ( .C1(n10991), .C2(n10130), .A(n10126), .B(n10124), .ZN(
        n10127) );
  OAI21_X1 U11266 ( .B1(n11419), .B2(n19532), .A(n11028), .ZN(n11029) );
  AND2_X1 U11267 ( .A1(n10141), .A2(n9746), .ZN(n15402) );
  NOR2_X1 U11268 ( .A1(n14758), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14749) );
  OR2_X1 U11269 ( .A1(n15390), .A2(n10167), .ZN(n11013) );
  NAND2_X1 U11270 ( .A1(n14781), .A2(n14440), .ZN(n14757) );
  OR2_X1 U11271 ( .A1(n14774), .A2(n14888), .ZN(n9843) );
  NOR2_X1 U11272 ( .A1(n15424), .A2(n10803), .ZN(n10806) );
  AOI21_X1 U11273 ( .B1(n14755), .B2(n20456), .A(n14754), .ZN(n14756) );
  NAND2_X1 U11274 ( .A1(n9844), .A2(n14511), .ZN(n14774) );
  AOI21_X1 U11275 ( .B1(n14767), .B2(n14949), .A(n20885), .ZN(n14779) );
  NAND2_X1 U11276 ( .A1(n9903), .A2(n9907), .ZN(n15424) );
  XNOR2_X1 U11277 ( .A(n9719), .B(n14447), .ZN(n14499) );
  OR2_X1 U11278 ( .A1(n14521), .A2(n10177), .ZN(n14511) );
  NAND2_X1 U11279 ( .A1(n9742), .A2(n9880), .ZN(n15560) );
  AND2_X1 U11280 ( .A1(n13588), .A2(n10871), .ZN(n10873) );
  AND2_X1 U11281 ( .A1(n14651), .A2(n14133), .ZN(n16269) );
  NAND2_X1 U11282 ( .A1(n9933), .A2(n9716), .ZN(n14880) );
  AOI21_X1 U11283 ( .B1(n9933), .B2(n9694), .A(n9740), .ZN(n9931) );
  XNOR2_X1 U11284 ( .A(n11713), .B(n11714), .ZN(n15246) );
  NAND2_X1 U11285 ( .A1(n9811), .A2(n13722), .ZN(n14424) );
  OAI21_X1 U11286 ( .B1(n16376), .B2(n9810), .A(n9808), .ZN(n9811) );
  AND2_X1 U11287 ( .A1(n13388), .A2(n10182), .ZN(n13822) );
  NAND2_X1 U11288 ( .A1(n10189), .A2(n10192), .ZN(n16376) );
  NOR2_X1 U11289 ( .A1(n15258), .A2(n11662), .ZN(n11690) );
  NAND2_X1 U11290 ( .A1(n13417), .A2(n13422), .ZN(n13416) );
  NOR2_X1 U11291 ( .A1(n9906), .A2(n9902), .ZN(n9901) );
  NOR2_X1 U11292 ( .A1(n15271), .A2(n11637), .ZN(n15260) );
  NOR2_X1 U11293 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  OR2_X1 U11294 ( .A1(n10202), .A2(n9935), .ZN(n9934) );
  OR2_X1 U11295 ( .A1(n10204), .A2(n10206), .ZN(n10201) );
  OAI21_X1 U11296 ( .B1(n12995), .B2(n9815), .A(n9812), .ZN(n20451) );
  AND2_X1 U11297 ( .A1(n16342), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10204) );
  NAND2_X1 U11298 ( .A1(n11009), .A2(n10816), .ZN(n10998) );
  AND2_X1 U11299 ( .A1(n15270), .A2(n15269), .ZN(n15271) );
  AND2_X1 U11300 ( .A1(n14435), .A2(n10203), .ZN(n10202) );
  XNOR2_X1 U11301 ( .A(n10861), .B(n10860), .ZN(n10862) );
  AND2_X1 U11302 ( .A1(n10814), .A2(n10815), .ZN(n16576) );
  NOR2_X2 U11303 ( .A1(n12970), .A2(n12969), .ZN(n12895) );
  NOR2_X1 U11304 ( .A1(n10195), .A2(n10191), .ZN(n10190) );
  NAND3_X1 U11305 ( .A1(n10617), .A2(n10616), .A3(n11126), .ZN(n10668) );
  NAND2_X1 U11306 ( .A1(n10617), .A2(n10616), .ZN(n10861) );
  AND2_X1 U11307 ( .A1(n12872), .A2(n12871), .ZN(n12969) );
  INV_X1 U11308 ( .A(n14877), .ZN(n10206) );
  OR2_X2 U11309 ( .A1(n15146), .A2(n15145), .ZN(n15363) );
  NAND2_X1 U11310 ( .A1(n10707), .A2(n10706), .ZN(n10850) );
  NAND2_X1 U11311 ( .A1(n12893), .A2(n12892), .ZN(n12894) );
  OR2_X1 U11312 ( .A1(n10693), .A2(n10692), .ZN(n10707) );
  AND2_X1 U11313 ( .A1(n13636), .A2(n13635), .ZN(n16379) );
  INV_X1 U11314 ( .A(n14877), .ZN(n9668) );
  AND2_X1 U11315 ( .A1(n10754), .A2(n10753), .ZN(n10776) );
  AND2_X1 U11316 ( .A1(n13723), .A2(n16453), .ZN(n14868) );
  OAI21_X1 U11317 ( .B1(n13164), .B2(n10172), .A(n10171), .ZN(n13648) );
  AND2_X1 U11318 ( .A1(n13723), .A2(n13659), .ZN(n13720) );
  AND3_X1 U11319 ( .A1(n10460), .A2(n10439), .A3(n10443), .ZN(n10010) );
  OAI22_X1 U11320 ( .A1(n10464), .A2(n11640), .B1(n19982), .B2(n11159), .ZN(
        n10465) );
  OAI21_X1 U11321 ( .B1(n13164), .B2(n13165), .A(n13171), .ZN(n10171) );
  NAND2_X1 U11322 ( .A1(n9926), .A2(n12671), .ZN(n15012) );
  AND2_X1 U11323 ( .A1(n19295), .A2(n10779), .ZN(n15479) );
  OR2_X1 U11324 ( .A1(n12884), .A2(n9943), .ZN(n13654) );
  NOR2_X1 U11325 ( .A1(n10461), .A2(n10441), .ZN(n10621) );
  AND2_X1 U11326 ( .A1(n10466), .A2(n10437), .ZN(n20026) );
  NAND2_X1 U11327 ( .A1(n12859), .A2(n12860), .ZN(n12884) );
  INV_X1 U11328 ( .A(n10684), .ZN(n19678) );
  NAND2_X1 U11329 ( .A1(n9891), .A2(n9892), .ZN(n10682) );
  OR2_X1 U11330 ( .A1(n10756), .A2(n10770), .ZN(n15157) );
  OR2_X1 U11331 ( .A1(n10445), .A2(n11439), .ZN(n10631) );
  NAND2_X1 U11332 ( .A1(n10468), .A2(n19414), .ZN(n10470) );
  NAND2_X1 U11333 ( .A1(n12232), .A2(n10198), .ZN(n13539) );
  AND2_X1 U11334 ( .A1(n13595), .A2(n13594), .ZN(n13597) );
  NAND2_X1 U11335 ( .A1(n12231), .A2(n9938), .ZN(n12232) );
  OAI21_X1 U11336 ( .B1(n12494), .B2(n12227), .A(n12493), .ZN(n10198) );
  NAND2_X1 U11337 ( .A1(n11086), .A2(n20122), .ZN(n11370) );
  NOR2_X1 U11338 ( .A1(n12911), .A2(n14498), .ZN(n20751) );
  NOR2_X1 U11339 ( .A1(n12911), .A2(n12905), .ZN(n20743) );
  NOR2_X1 U11340 ( .A1(n12911), .A2(n14478), .ZN(n20737) );
  OR2_X1 U11341 ( .A1(n19046), .A2(n19254), .ZN(n16946) );
  NOR2_X1 U11342 ( .A1(n12911), .A2(n12910), .ZN(n20731) );
  NAND3_X1 U11343 ( .A1(n9862), .A2(n9863), .A3(n10429), .ZN(n9796) );
  NOR2_X1 U11344 ( .A1(n16099), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10101) );
  NOR2_X1 U11345 ( .A1(n12911), .A2(n11978), .ZN(n20719) );
  NOR2_X1 U11346 ( .A1(n12911), .A2(n12059), .ZN(n20713) );
  CLKBUF_X1 U11347 ( .A(n12492), .Z(n20591) );
  OR2_X1 U11348 ( .A1(n12584), .A2(n12583), .ZN(n9824) );
  NOR2_X1 U11349 ( .A1(n19545), .A2(n19544), .ZN(n19583) );
  XNOR2_X1 U11350 ( .A(n9951), .B(n9950), .ZN(n18183) );
  NAND2_X1 U11351 ( .A1(n10434), .A2(n10435), .ZN(n10436) );
  INV_X2 U11352 ( .A(n15291), .ZN(n15279) );
  OR2_X1 U11353 ( .A1(n10394), .A2(n10393), .ZN(n10423) );
  XNOR2_X1 U11354 ( .A(n12270), .B(n12269), .ZN(n12678) );
  NAND2_X1 U11355 ( .A1(n10428), .A2(n10421), .ZN(n10429) );
  XNOR2_X1 U11356 ( .A(n10898), .B(n10897), .ZN(n10896) );
  CLKBUF_X1 U11357 ( .A(n10888), .Z(n10977) );
  NAND2_X1 U11358 ( .A1(n9841), .A2(n12181), .ZN(n12197) );
  OAI211_X1 U11359 ( .C1(n10902), .C2(n11372), .A(n10431), .B(n10430), .ZN(
        n10897) );
  NAND2_X1 U11360 ( .A1(n9898), .A2(n10395), .ZN(n10433) );
  NAND3_X1 U11361 ( .A1(n10414), .A2(n9826), .A3(n10415), .ZN(n10426) );
  INV_X1 U11362 ( .A(n10032), .ZN(n10031) );
  AND3_X1 U11363 ( .A1(n10090), .A2(n9743), .A3(n10088), .ZN(n16091) );
  NOR2_X1 U11364 ( .A1(n10403), .A2(n10245), .ZN(n10405) );
  OR2_X1 U11365 ( .A1(n11858), .A2(n11857), .ZN(n11860) );
  INV_X2 U11366 ( .A(n17292), .ZN(n17261) );
  OR2_X1 U11367 ( .A1(n10398), .A2(n10397), .ZN(n10403) );
  INV_X2 U11368 ( .A(n17863), .ZN(n17893) );
  XNOR2_X1 U11369 ( .A(n16086), .B(n16087), .ZN(n18226) );
  XNOR2_X1 U11370 ( .A(n16794), .B(n9963), .ZN(n17292) );
  AND2_X1 U11371 ( .A1(n11349), .A2(n10362), .ZN(n11336) );
  NAND2_X1 U11372 ( .A1(n10054), .A2(n10053), .ZN(n16699) );
  NAND2_X1 U11373 ( .A1(n19265), .A2(n16945), .ZN(n16960) );
  NAND2_X1 U11374 ( .A1(n12183), .A2(n9928), .ZN(n12283) );
  INV_X2 U11375 ( .A(n10890), .ZN(n9678) );
  AND4_X1 U11376 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12319), .ZN(
        n12191) );
  CLKBUF_X1 U11377 ( .A(n11338), .Z(n16728) );
  NOR2_X1 U11378 ( .A1(n12175), .A2(n9819), .ZN(n9818) );
  OR2_X1 U11379 ( .A1(n10722), .A2(n10030), .ZN(n10029) );
  INV_X2 U11380 ( .A(n11335), .ZN(n11328) );
  NAND2_X2 U11381 ( .A1(n12272), .A2(n12294), .ZN(n11946) );
  NAND2_X1 U11382 ( .A1(n11094), .A2(n9659), .ZN(n11301) );
  AND2_X1 U11383 ( .A1(n13014), .A2(n14454), .ZN(n12186) );
  AND2_X1 U11384 ( .A1(n11980), .A2(n12065), .ZN(n9817) );
  AND2_X1 U11385 ( .A1(n11077), .A2(n10406), .ZN(n10413) );
  NAND2_X1 U11386 ( .A1(n11918), .A2(n10255), .ZN(n12272) );
  NAND2_X1 U11387 ( .A1(n14454), .A2(n9988), .ZN(n14417) );
  NOR2_X1 U11388 ( .A1(n10331), .A2(n10332), .ZN(n11077) );
  INV_X1 U11389 ( .A(n20860), .ZN(n13657) );
  NAND2_X1 U11390 ( .A1(n10364), .A2(n10363), .ZN(n10381) );
  NAND2_X1 U11391 ( .A1(n12497), .A2(n12226), .ZN(n13167) );
  INV_X1 U11392 ( .A(n11802), .ZN(n11062) );
  AND2_X1 U11393 ( .A1(n12169), .A2(n12905), .ZN(n12065) );
  NAND2_X1 U11394 ( .A1(n10372), .A2(n10582), .ZN(n11096) );
  INV_X2 U11395 ( .A(n14419), .ZN(n14454) );
  NAND3_X1 U11396 ( .A1(n13923), .A2(n13922), .A3(n13921), .ZN(n16101) );
  AND2_X1 U11397 ( .A1(n10379), .A2(n10378), .ZN(n11065) );
  OR2_X1 U11398 ( .A1(n10614), .A2(n10613), .ZN(n11126) );
  AND2_X1 U11399 ( .A1(n10343), .A2(n19564), .ZN(n11802) );
  INV_X1 U11400 ( .A(n18625), .ZN(n16114) );
  NOR2_X2 U11402 ( .A1(n13970), .A2(n13969), .ZN(n18639) );
  NOR2_X1 U11403 ( .A1(n12286), .A2(n12294), .ZN(n12788) );
  NAND3_X1 U11404 ( .A1(n13933), .A2(n13932), .A3(n13931), .ZN(n16102) );
  NAND2_X1 U11405 ( .A1(n9800), .A2(n9797), .ZN(n10849) );
  NAND2_X1 U11406 ( .A1(n10306), .A2(n10305), .ZN(n19569) );
  NAND2_X1 U11407 ( .A1(n20279), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20277) );
  OR2_X2 U11408 ( .A1(n16895), .A2(n16849), .ZN(n16897) );
  OR2_X2 U11409 ( .A1(n11908), .A2(n11907), .ZN(n14477) );
  NAND2_X2 U11410 ( .A1(n10318), .A2(n10317), .ZN(n11352) );
  NAND3_X1 U11411 ( .A1(n10323), .A2(n10322), .A3(n10321), .ZN(n10330) );
  NAND2_X1 U11412 ( .A1(n10275), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10282) );
  NAND2_X1 U11413 ( .A1(n10253), .A2(n10263), .ZN(n10271) );
  NAND2_X1 U11414 ( .A1(n10287), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10294) );
  AND2_X2 U11415 ( .A1(n11760), .A2(n9802), .ZN(n11623) );
  AND2_X1 U11416 ( .A1(n10277), .A2(n10276), .ZN(n10280) );
  NOR2_X1 U11417 ( .A1(n9803), .A2(n9802), .ZN(n9801) );
  NOR2_X1 U11418 ( .A1(n9799), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9798) );
  AND4_X1 U11419 ( .A1(n10273), .A2(n10274), .A3(n9869), .A4(n10272), .ZN(
        n10275) );
  AND4_X1 U11420 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10311) );
  AND4_X1 U11421 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10287) );
  AND4_X1 U11422 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11887) );
  AND3_X1 U11423 ( .A1(n10320), .A2(n10319), .A3(n9802), .ZN(n10323) );
  AND2_X1 U11424 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  INV_X2 U11425 ( .A(n15903), .ZN(n11760) );
  AND2_X1 U11426 ( .A1(n11889), .A2(n11888), .ZN(n11890) );
  NAND2_X2 U11427 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20197), .ZN(n20203) );
  BUF_X4 U11429 ( .A(n12219), .Z(n14364) );
  AND2_X1 U11431 ( .A1(n10324), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10328) );
  BUF_X2 U11432 ( .A(n13949), .Z(n17556) );
  CLKBUF_X2 U11433 ( .A(n13949), .Z(n17540) );
  NAND2_X2 U11434 ( .A1(n19260), .A2(n19125), .ZN(n19183) );
  OR2_X1 U11435 ( .A1(n13884), .A2(n13880), .ZN(n17458) );
  AND2_X4 U11436 ( .A1(n11880), .A2(n12800), .ZN(n13337) );
  BUF_X2 U11437 ( .A(n11913), .Z(n9674) );
  INV_X2 U11438 ( .A(n16934), .ZN(n16936) );
  INV_X2 U11439 ( .A(n20289), .ZN(n20197) );
  AND3_X2 U11440 ( .A1(n10259), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n10162), .ZN(n11638) );
  AND2_X1 U11441 ( .A1(n12273), .A2(n11881), .ZN(n11947) );
  AND2_X2 U11442 ( .A1(n11872), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11880) );
  CLKBUF_X1 U11443 ( .A(n10489), .Z(n15907) );
  INV_X2 U11444 ( .A(n20126), .ZN(n9671) );
  NOR2_X1 U11445 ( .A1(n13879), .A2(n17321), .ZN(n17584) );
  INV_X1 U11446 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12376) );
  AND2_X1 U11447 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11882) );
  AND2_X2 U11448 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12800) );
  NAND2_X2 U11449 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19061) );
  NAND2_X1 U11450 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13880) );
  INV_X2 U11451 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19232) );
  INV_X1 U11452 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11872) );
  AND2_X1 U11453 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12798) );
  INV_X1 U11454 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10259) );
  INV_X1 U11455 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10572) );
  AND2_X1 U11456 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10489) );
  NOR2_X2 U11457 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15876) );
  NAND3_X2 U11458 ( .A1(n9948), .A2(n9947), .A3(n9946), .ZN(n18253) );
  INV_X2 U11459 ( .A(n12286), .ZN(n11978) );
  NAND2_X2 U11460 ( .A1(n15590), .A2(n10883), .ZN(n15550) );
  NOR2_X2 U11461 ( .A1(n10471), .A2(n10470), .ZN(n10618) );
  NOR2_X2 U11462 ( .A1(n14757), .A2(n14441), .ZN(n14748) );
  AND2_X1 U11463 ( .A1(n12273), .A2(n11882), .ZN(n9672) );
  AND2_X4 U11464 ( .A1(n12798), .A2(n11873), .ZN(n11984) );
  AND2_X1 U11465 ( .A1(n11881), .A2(n11879), .ZN(n9673) );
  AND2_X1 U11466 ( .A1(n11881), .A2(n11879), .ZN(n12218) );
  AND2_X4 U11467 ( .A1(n11091), .A2(n11090), .ZN(n11236) );
  NOR2_X1 U11468 ( .A1(n13879), .A2(n17321), .ZN(n9676) );
  AND2_X4 U11469 ( .A1(n11880), .A2(n12273), .ZN(n12219) );
  NAND2_X1 U11470 ( .A1(n11364), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9677) );
  INV_X4 U11471 ( .A(n10408), .ZN(n10889) );
  AOI21_X2 U11472 ( .B1(n15958), .B2(n18613), .A(n15957), .ZN(n19055) );
  AND2_X4 U11473 ( .A1(n12797), .A2(n12800), .ZN(n11989) );
  XNOR2_X2 U11474 ( .A(n10444), .B(n10420), .ZN(n10437) );
  NAND3_X2 U11475 ( .A1(n11945), .A2(n11946), .A3(n9696), .ZN(n12172) );
  NAND2_X2 U11476 ( .A1(n14816), .A2(n14777), .ZN(n14767) );
  AND2_X1 U11478 ( .A1(n11880), .A2(n11879), .ZN(n9683) );
  AND2_X1 U11479 ( .A1(n11878), .A2(n11882), .ZN(n9684) );
  XNOR2_X2 U11480 ( .A(n12657), .B(n12762), .ZN(n12677) );
  NAND2_X2 U11481 ( .A1(n12584), .A2(n12583), .ZN(n12657) );
  NAND3_X2 U11482 ( .A1(n19262), .A2(n19249), .A3(n19261), .ZN(n18476) );
  NAND2_X1 U11483 ( .A1(n12184), .A2(n12050), .ZN(n12183) );
  OAI211_X1 U11484 ( .C1(n12232), .C2(n12295), .A(n9984), .B(n9982), .ZN(
        n12545) );
  AOI21_X1 U11485 ( .B1(n12296), .B2(n13651), .A(n9985), .ZN(n9984) );
  NAND2_X1 U11486 ( .A1(n9983), .A2(n12296), .ZN(n9982) );
  INV_X1 U11487 ( .A(n10198), .ZN(n9983) );
  AOI22_X1 U11488 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11954) );
  AND3_X1 U11489 ( .A1(n16156), .A2(n12528), .A3(n12383), .ZN(n20457) );
  OR2_X1 U11490 ( .A1(n12009), .A2(n12059), .ZN(n12020) );
  NAND2_X1 U11491 ( .A1(n10381), .A2(n10343), .ZN(n10382) );
  NAND2_X1 U11492 ( .A1(n10358), .A2(n10343), .ZN(n10360) );
  NAND2_X1 U11493 ( .A1(n12283), .A2(n12052), .ZN(n12179) );
  OAI21_X1 U11494 ( .B1(n9986), .B2(n9988), .A(n9817), .ZN(n9816) );
  NOR2_X1 U11495 ( .A1(n13024), .A2(n9987), .ZN(n9986) );
  INV_X1 U11496 ( .A(n10426), .ZN(n10428) );
  AOI21_X1 U11497 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20236), .A(
        n10602), .ZN(n10836) );
  NOR2_X1 U11498 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  INV_X1 U11499 ( .A(n10599), .ZN(n10601) );
  NAND2_X1 U11500 ( .A1(n9668), .A2(n9783), .ZN(n10203) );
  INV_X1 U11501 ( .A(n14566), .ZN(n10008) );
  NAND2_X1 U11502 ( .A1(n9936), .A2(n9941), .ZN(n12494) );
  NAND2_X1 U11503 ( .A1(n9755), .A2(n13401), .ZN(n10065) );
  AND2_X2 U11504 ( .A1(n11793), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11573) );
  AND2_X1 U11505 ( .A1(n15907), .A2(n10490), .ZN(n11562) );
  NAND2_X1 U11506 ( .A1(n15251), .A2(n11691), .ZN(n11713) );
  OR2_X1 U11507 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  NOR2_X1 U11508 ( .A1(n15364), .A2(n10074), .ZN(n10073) );
  INV_X1 U11509 ( .A(n15133), .ZN(n10074) );
  NOR2_X1 U11510 ( .A1(n10230), .A2(n15276), .ZN(n10229) );
  NAND2_X1 U11511 ( .A1(n9701), .A2(n9922), .ZN(n9921) );
  NOR2_X1 U11512 ( .A1(n9924), .A2(n9923), .ZN(n9922) );
  AND2_X1 U11513 ( .A1(n13304), .A2(n16684), .ZN(n13324) );
  INV_X1 U11514 ( .A(n11732), .ZN(n11684) );
  AND3_X1 U11515 ( .A1(n15403), .A2(n10147), .A3(n10146), .ZN(n10145) );
  AND2_X1 U11516 ( .A1(n10149), .A2(n10150), .ZN(n9910) );
  INV_X1 U11517 ( .A(n10151), .ZN(n10150) );
  NAND2_X1 U11518 ( .A1(n10775), .A2(n10155), .ZN(n10149) );
  OAI21_X1 U11519 ( .B1(n10154), .B2(n15452), .A(n10152), .ZN(n10151) );
  AND2_X1 U11520 ( .A1(n15819), .A2(n15197), .ZN(n10062) );
  NAND2_X1 U11521 ( .A1(n10875), .A2(n11137), .ZN(n10881) );
  AND2_X1 U11522 ( .A1(n16723), .A2(n11821), .ZN(n11090) );
  NAND2_X1 U11523 ( .A1(n11336), .A2(n11802), .ZN(n15886) );
  NOR2_X1 U11524 ( .A1(n17758), .A2(n16090), .ZN(n16095) );
  NOR3_X1 U11525 ( .A1(n16136), .A2(n18316), .A3(n17963), .ZN(n17926) );
  INV_X1 U11526 ( .A(n9951), .ZN(n16097) );
  NOR2_X1 U11527 ( .A1(n18629), .A2(n16101), .ZN(n16110) );
  NOR2_X1 U11528 ( .A1(n13019), .A2(n9842), .ZN(n12787) );
  OAI21_X1 U11529 ( .B1(n9680), .B2(n13476), .A(n12604), .ZN(n12605) );
  INV_X1 U11530 ( .A(n20293), .ZN(n12534) );
  NAND2_X1 U11531 ( .A1(n9990), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9989) );
  INV_X1 U11532 ( .A(n16197), .ZN(n9990) );
  NAND3_X1 U11533 ( .A1(n12895), .A2(n12894), .A3(n13177), .ZN(n13181) );
  NAND2_X1 U11534 ( .A1(n13167), .A2(n11982), .ZN(n12028) );
  OAI21_X1 U11535 ( .B1(n12026), .B2(n9779), .A(n12027), .ZN(n9840) );
  AND2_X1 U11536 ( .A1(n12673), .A2(n15009), .ZN(n12949) );
  OR2_X1 U11537 ( .A1(n9680), .A2(n12708), .ZN(n20704) );
  AND3_X1 U11538 ( .A1(n12063), .A2(n12540), .A3(n12062), .ZN(n16156) );
  OR2_X1 U11539 ( .A1(n16725), .A2(n12243), .ZN(n11867) );
  INV_X1 U11540 ( .A(n15315), .ZN(n10067) );
  NAND2_X1 U11541 ( .A1(n13285), .A2(n11133), .ZN(n13595) );
  AND2_X1 U11542 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10013) );
  NAND2_X1 U11543 ( .A1(n10129), .A2(n10134), .ZN(n15377) );
  AOI21_X1 U11544 ( .B1(n10991), .B2(n10133), .A(n10130), .ZN(n10129) );
  NAND2_X1 U11545 ( .A1(n10062), .A2(n10059), .ZN(n10058) );
  INV_X1 U11546 ( .A(n13257), .ZN(n10059) );
  AND2_X1 U11547 ( .A1(n12102), .A2(n11435), .ZN(n12134) );
  OAI211_X1 U11548 ( .C1(n15894), .C2(n10220), .A(n10214), .B(n10212), .ZN(
        n12135) );
  AND2_X1 U11549 ( .A1(n10215), .A2(n10217), .ZN(n10214) );
  NAND2_X1 U11550 ( .A1(n10218), .A2(n11436), .ZN(n10217) );
  AND4_X1 U11551 ( .A1(n11803), .A2(n11802), .A3(n10385), .A4(n10355), .ZN(
        n10356) );
  INV_X2 U11552 ( .A(n9720), .ZN(n17575) );
  INV_X1 U11553 ( .A(n18613), .ZN(n19246) );
  NAND2_X1 U11554 ( .A1(n16125), .A2(n18168), .ZN(n16129) );
  NAND2_X1 U11555 ( .A1(n9954), .A2(n9762), .ZN(n16127) );
  NAND2_X1 U11556 ( .A1(n16128), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9954) );
  AND2_X1 U11557 ( .A1(n16333), .A2(n12548), .ZN(n16365) );
  AND3_X1 U11558 ( .A1(n10252), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n10824), .ZN(n15618) );
  NAND2_X1 U11559 ( .A1(n12000), .A2(n11999), .ZN(n12009) );
  NAND2_X1 U11560 ( .A1(n9842), .A2(n13167), .ZN(n12000) );
  NAND2_X1 U11561 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n9793) );
  NAND2_X1 U11562 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9794) );
  NAND2_X1 U11563 ( .A1(n9693), .A2(n9891), .ZN(n9889) );
  AND4_X1 U11564 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        n10700) );
  NOR2_X1 U11565 ( .A1(n9677), .A2(n10366), .ZN(n10369) );
  NAND2_X1 U11566 ( .A1(n20243), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10584) );
  NAND2_X1 U11567 ( .A1(n20252), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10570) );
  NAND2_X1 U11568 ( .A1(n10585), .A2(n10584), .ZN(n10599) );
  NAND2_X1 U11569 ( .A1(n11065), .A2(n11352), .ZN(n11063) );
  NAND2_X1 U11570 ( .A1(n11945), .A2(n11946), .ZN(n12182) );
  INV_X1 U11571 ( .A(n13656), .ZN(n13644) );
  NAND3_X1 U11572 ( .A1(n12049), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13019), 
        .ZN(n13169) );
  NAND2_X1 U11573 ( .A1(n9834), .A2(n9832), .ZN(n9831) );
  NAND2_X1 U11574 ( .A1(n12014), .A2(n9833), .ZN(n9832) );
  INV_X1 U11575 ( .A(n12015), .ZN(n9833) );
  AND2_X1 U11576 ( .A1(n12018), .A2(n12017), .ZN(n9830) );
  NAND2_X1 U11577 ( .A1(n12051), .A2(n20860), .ZN(n9928) );
  NAND2_X1 U11578 ( .A1(n10033), .A2(n10662), .ZN(n10032) );
  INV_X1 U11579 ( .A(n10658), .ZN(n10033) );
  NAND2_X1 U11580 ( .A1(n9899), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U11581 ( .A1(n10158), .A2(n10159), .ZN(n9899) );
  INV_X1 U11582 ( .A(n10400), .ZN(n10158) );
  INV_X1 U11583 ( .A(n10850), .ZN(n10708) );
  INV_X1 U11584 ( .A(n10709), .ZN(n10157) );
  OR2_X1 U11585 ( .A1(n10655), .A2(n10654), .ZN(n10660) );
  AOI22_X1 U11586 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11781), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U11587 ( .A1(n11342), .A2(n9825), .ZN(n9826) );
  AND2_X1 U11588 ( .A1(n10571), .A2(n10570), .ZN(n10574) );
  OR2_X1 U11589 ( .A1(n11038), .A2(n10842), .ZN(n10571) );
  NOR2_X1 U11590 ( .A1(n17765), .A2(n16085), .ZN(n16080) );
  AND2_X1 U11591 ( .A1(n9761), .A2(n14183), .ZN(n10180) );
  NAND2_X1 U11592 ( .A1(n14091), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14348) );
  INV_X1 U11593 ( .A(n14348), .ZN(n14375) );
  NOR2_X1 U11594 ( .A1(n10188), .A2(n13753), .ZN(n10186) );
  INV_X1 U11595 ( .A(n13832), .ZN(n10188) );
  NAND2_X1 U11596 ( .A1(n10184), .A2(n13753), .ZN(n13820) );
  INV_X1 U11597 ( .A(n13750), .ZN(n10184) );
  AND2_X1 U11598 ( .A1(n13480), .A2(n13389), .ZN(n10187) );
  OR2_X1 U11599 ( .A1(n14477), .A2(n20697), .ZN(n14285) );
  INV_X1 U11600 ( .A(n14615), .ZN(n9999) );
  AND2_X1 U11601 ( .A1(n14631), .A2(n10001), .ZN(n10000) );
  INV_X1 U11602 ( .A(n14622), .ZN(n10001) );
  INV_X1 U11603 ( .A(n16373), .ZN(n9810) );
  AOI21_X1 U11604 ( .B1(n16373), .B2(n9809), .A(n9738), .ZN(n9808) );
  INV_X1 U11605 ( .A(n16374), .ZN(n9809) );
  NAND2_X1 U11606 ( .A1(n9988), .A2(n14419), .ZN(n14410) );
  AND2_X1 U11607 ( .A1(n12540), .A2(n14477), .ZN(n11980) );
  NAND2_X1 U11608 ( .A1(n12910), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U11609 ( .A1(n12334), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9841) );
  OR2_X1 U11610 ( .A1(n13019), .A2(n16503), .ZN(n12497) );
  INV_X1 U11611 ( .A(n12226), .ZN(n12495) );
  OR2_X1 U11612 ( .A1(n12490), .A2(n12489), .ZN(n12618) );
  INV_X1 U11613 ( .A(n13169), .ZN(n13044) );
  INV_X1 U11614 ( .A(n12859), .ZN(n9926) );
  OR2_X1 U11615 ( .A1(n12268), .A2(n12331), .ZN(n12332) );
  NOR2_X1 U11616 ( .A1(n10197), .A2(n10196), .ZN(n11981) );
  OAI21_X1 U11617 ( .B1(n20861), .B2(n12819), .A(n15028), .ZN(n12680) );
  INV_X1 U11618 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20554) );
  INV_X1 U11619 ( .A(n9817), .ZN(n12301) );
  OAI21_X1 U11620 ( .B1(n13262), .B2(n10022), .A(n10019), .ZN(n10830) );
  NOR2_X1 U11621 ( .A1(n10799), .A2(n10798), .ZN(n10018) );
  NAND2_X1 U11622 ( .A1(n10770), .A2(n10951), .ZN(n10793) );
  INV_X1 U11623 ( .A(n11576), .ZN(n11612) );
  INV_X1 U11624 ( .A(n11575), .ZN(n11613) );
  INV_X1 U11625 ( .A(n11574), .ZN(n11609) );
  AND2_X1 U11626 ( .A1(n11661), .A2(n11660), .ZN(n11662) );
  INV_X1 U11627 ( .A(n11661), .ZN(n10227) );
  INV_X1 U11628 ( .A(n10229), .ZN(n10224) );
  NAND2_X1 U11629 ( .A1(n15286), .A2(n10231), .ZN(n10230) );
  INV_X1 U11630 ( .A(n15280), .ZN(n10231) );
  AND2_X1 U11631 ( .A1(n11457), .A2(n13395), .ZN(n10237) );
  INV_X1 U11632 ( .A(n15170), .ZN(n10066) );
  NOR2_X1 U11633 ( .A1(n15263), .A2(n10116), .ZN(n10115) );
  INV_X1 U11634 ( .A(n15080), .ZN(n10116) );
  NAND2_X1 U11635 ( .A1(n10131), .A2(n10994), .ZN(n10130) );
  NAND2_X1 U11636 ( .A1(n10992), .A2(n10132), .ZN(n10131) );
  NAND2_X1 U11637 ( .A1(n10995), .A2(n15626), .ZN(n10132) );
  AND2_X1 U11638 ( .A1(n10115), .A2(n10114), .ZN(n10113) );
  INV_X1 U11639 ( .A(n15254), .ZN(n10114) );
  INV_X1 U11640 ( .A(n15422), .ZN(n10143) );
  INV_X1 U11641 ( .A(n10806), .ZN(n10144) );
  OR2_X1 U11642 ( .A1(n10792), .A2(n15479), .ZN(n10156) );
  NAND2_X1 U11643 ( .A1(n15560), .A2(n15452), .ZN(n15530) );
  OAI21_X1 U11644 ( .B1(n10136), .B2(n10729), .A(n15454), .ZN(n9883) );
  NAND2_X1 U11645 ( .A1(n10716), .A2(n10135), .ZN(n9884) );
  NAND2_X1 U11646 ( .A1(n9888), .A2(n9886), .ZN(n10140) );
  NOR2_X1 U11647 ( .A1(n10716), .A2(n9887), .ZN(n9886) );
  NAND2_X1 U11648 ( .A1(n10107), .A2(n12556), .ZN(n10106) );
  INV_X1 U11649 ( .A(n12406), .ZN(n10107) );
  INV_X1 U11650 ( .A(n9763), .ZN(n9791) );
  NAND2_X1 U11651 ( .A1(n10015), .A2(n10160), .ZN(n10863) );
  NAND2_X1 U11652 ( .A1(n10859), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10160) );
  NOR2_X1 U11653 ( .A1(n13143), .A2(n11372), .ZN(n9878) );
  NAND2_X1 U11654 ( .A1(n13143), .A2(n11372), .ZN(n9877) );
  NAND2_X1 U11655 ( .A1(n13275), .A2(n11137), .ZN(n9872) );
  NOR2_X1 U11656 ( .A1(n9878), .A2(n9875), .ZN(n9874) );
  INV_X1 U11657 ( .A(n13275), .ZN(n9875) );
  NAND2_X1 U11658 ( .A1(n9866), .A2(n9864), .ZN(n10553) );
  INV_X1 U11659 ( .A(n10617), .ZN(n9866) );
  INV_X1 U11660 ( .A(n10616), .ZN(n9864) );
  OR2_X1 U11661 ( .A1(n10495), .A2(n10494), .ZN(n11095) );
  INV_X1 U11662 ( .A(n19564), .ZN(n11350) );
  NAND2_X1 U11663 ( .A1(n16699), .A2(n16698), .ZN(n11109) );
  NAND4_X1 U11664 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10329) );
  AND2_X1 U11665 ( .A1(n11056), .A2(n11054), .ZN(n11830) );
  INV_X1 U11666 ( .A(n10470), .ZN(n10438) );
  AOI21_X1 U11667 ( .B1(n17540), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n10086), .ZN(n10085) );
  INV_X1 U11668 ( .A(n16015), .ZN(n10083) );
  INV_X1 U11669 ( .A(n16014), .ZN(n10087) );
  NOR2_X1 U11670 ( .A1(n13884), .A2(n13879), .ZN(n14024) );
  NOR2_X1 U11671 ( .A1(n10240), .A2(n9957), .ZN(n9956) );
  NOR2_X1 U11672 ( .A1(n18639), .A2(n18621), .ZN(n15966) );
  NAND3_X1 U11673 ( .A1(n10093), .A2(n9952), .A3(n9730), .ZN(n9951) );
  OAI21_X1 U11674 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n21004), .A(
        n13981), .ZN(n15933) );
  INV_X1 U11675 ( .A(n18621), .ZN(n15953) );
  AOI211_X1 U11676 ( .C1(n17572), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n13920), .B(n13919), .ZN(n13921) );
  NAND2_X1 U11677 ( .A1(n10005), .A2(n10003), .ZN(n10002) );
  NOR2_X1 U11678 ( .A1(n10008), .A2(n14653), .ZN(n10003) );
  OR2_X1 U11679 ( .A1(n20855), .A2(n13011), .ZN(n16238) );
  OR2_X1 U11680 ( .A1(n12786), .A2(n12528), .ZN(n12291) );
  INV_X1 U11681 ( .A(n12280), .ZN(n12529) );
  INV_X1 U11682 ( .A(n10176), .ZN(n10174) );
  NAND2_X1 U11683 ( .A1(n14436), .A2(n10206), .ZN(n14816) );
  AND2_X1 U11684 ( .A1(n10202), .A2(n9787), .ZN(n10199) );
  NAND2_X1 U11685 ( .A1(n13822), .A2(n9846), .ZN(n14658) );
  NOR2_X1 U11686 ( .A1(n9847), .A2(n14561), .ZN(n9846) );
  INV_X1 U11687 ( .A(n9848), .ZN(n9847) );
  AND2_X1 U11688 ( .A1(n14738), .A2(n14739), .ZN(n14740) );
  INV_X1 U11689 ( .A(n13181), .ZN(n13178) );
  INV_X1 U11690 ( .A(n9934), .ZN(n9932) );
  AND2_X1 U11691 ( .A1(n10193), .A2(n13639), .ZN(n10192) );
  NAND2_X1 U11692 ( .A1(n16386), .A2(n16385), .ZN(n16384) );
  NAND2_X1 U11693 ( .A1(n12309), .A2(n12534), .ZN(n12323) );
  NAND2_X1 U11694 ( .A1(n9820), .A2(n14478), .ZN(n9819) );
  INV_X1 U11695 ( .A(n12494), .ZN(n12231) );
  NAND2_X1 U11696 ( .A1(n12342), .A2(n12341), .ZN(n12762) );
  NAND2_X1 U11697 ( .A1(n16503), .A2(n12680), .ZN(n13496) );
  NOR2_X1 U11698 ( .A1(n12301), .A2(n13024), .ZN(n16166) );
  INV_X2 U11699 ( .A(n9842), .ZN(n12059) );
  NAND2_X1 U11700 ( .A1(n10018), .A2(n10017), .ZN(n10807) );
  INV_X1 U11701 ( .A(n10018), .ZN(n10804) );
  NOR2_X1 U11702 ( .A1(n10037), .A2(n10763), .ZN(n10036) );
  INV_X1 U11703 ( .A(n10038), .ZN(n10037) );
  NOR2_X1 U11704 ( .A1(n10039), .A2(n10747), .ZN(n10038) );
  INV_X1 U11705 ( .A(n10743), .ZN(n10039) );
  NOR2_X1 U11706 ( .A1(n10026), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10025) );
  INV_X1 U11707 ( .A(n10419), .ZN(n10444) );
  AND2_X1 U11708 ( .A1(n9664), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11565) );
  OR2_X1 U11709 ( .A1(n11736), .A2(n9915), .ZN(n9914) );
  INV_X1 U11710 ( .A(n9916), .ZN(n9915) );
  INV_X1 U11711 ( .A(n11734), .ZN(n10209) );
  NAND2_X1 U11712 ( .A1(n11713), .A2(n10211), .ZN(n10210) );
  AND2_X1 U11713 ( .A1(n9727), .A2(n11661), .ZN(n11637) );
  AND2_X1 U11714 ( .A1(n10073), .A2(n10071), .ZN(n10070) );
  INV_X1 U11715 ( .A(n15118), .ZN(n10071) );
  NAND2_X1 U11716 ( .A1(n12398), .A2(n11452), .ZN(n12369) );
  AND2_X1 U11717 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12368) );
  XNOR2_X1 U11718 ( .A(n11025), .B(n11024), .ZN(n13234) );
  NAND2_X1 U11719 ( .A1(n9829), .A2(n9828), .ZN(n15380) );
  INV_X1 U11720 ( .A(n10169), .ZN(n9828) );
  INV_X1 U11721 ( .A(n15390), .ZN(n9829) );
  AOI21_X1 U11722 ( .B1(n9907), .B2(n9905), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9904) );
  INV_X1 U11723 ( .A(n9722), .ZN(n9905) );
  NOR2_X1 U11724 ( .A1(n15530), .A2(n10775), .ZN(n10153) );
  AND2_X1 U11725 ( .A1(n10886), .A2(n10170), .ZN(n15485) );
  NOR2_X1 U11726 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  INV_X1 U11727 ( .A(n15189), .ZN(n10057) );
  NOR2_X1 U11728 ( .A1(n10728), .A2(n10139), .ZN(n10138) );
  INV_X1 U11729 ( .A(n15829), .ZN(n10139) );
  XNOR2_X1 U11730 ( .A(n10881), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15591) );
  OAI21_X1 U11731 ( .B1(n15840), .B2(n9806), .A(n9804), .ZN(n15590) );
  INV_X1 U11732 ( .A(n10880), .ZN(n9806) );
  AOI21_X1 U11733 ( .B1(n10880), .B2(n16682), .A(n9805), .ZN(n9804) );
  INV_X1 U11734 ( .A(n15591), .ZN(n9805) );
  NAND2_X1 U11735 ( .A1(n13416), .A2(n10865), .ZN(n13448) );
  AND2_X1 U11736 ( .A1(n13424), .A2(n13281), .ZN(n10055) );
  INV_X1 U11737 ( .A(n9879), .ZN(n9876) );
  OAI21_X1 U11738 ( .B1(n10851), .B2(n11137), .A(n13275), .ZN(n9879) );
  OR2_X1 U11739 ( .A1(n20239), .A2(n20227), .ZN(n19802) );
  INV_X1 U11740 ( .A(n9661), .ZN(n19379) );
  NAND2_X1 U11741 ( .A1(n12133), .A2(n11438), .ZN(n12400) );
  NAND2_X1 U11742 ( .A1(n10222), .A2(n11427), .ZN(n11437) );
  NAND2_X1 U11743 ( .A1(n15894), .A2(n11440), .ZN(n10222) );
  AND2_X1 U11744 ( .A1(n11451), .A2(n11449), .ZN(n12399) );
  NOR2_X2 U11745 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20223) );
  AND2_X1 U11746 ( .A1(n19860), .A2(n20256), .ZN(n19767) );
  AND2_X1 U11747 ( .A1(n19860), .A2(n19827), .ZN(n19807) );
  AND2_X1 U11748 ( .A1(n20239), .A2(n20227), .ZN(n19828) );
  NOR2_X1 U11749 ( .A1(n19860), .A2(n19827), .ZN(n20019) );
  NOR2_X1 U11750 ( .A1(n19860), .A2(n20256), .ZN(n19927) );
  INV_X1 U11751 ( .A(n19802), .ZN(n20062) );
  NAND2_X2 U11752 ( .A1(n10282), .A2(n10281), .ZN(n19590) );
  NAND2_X1 U11753 ( .A1(n10280), .A2(n10238), .ZN(n10281) );
  INV_X1 U11754 ( .A(n20067), .ZN(n19775) );
  INV_X1 U11755 ( .A(n17919), .ZN(n9970) );
  INV_X1 U11756 ( .A(n9971), .ZN(n17008) );
  OAI21_X1 U11757 ( .B1(n17025), .B2(n17261), .A(n9968), .ZN(n9971) );
  NOR2_X1 U11758 ( .A1(n9969), .A2(n17908), .ZN(n9968) );
  NOR2_X1 U11759 ( .A1(n17261), .A2(n9970), .ZN(n9969) );
  INV_X1 U11760 ( .A(n17310), .ZN(n17326) );
  NOR3_X1 U11761 ( .A1(n17456), .A2(n13985), .A3(n17469), .ZN(n17342) );
  OR2_X1 U11762 ( .A1(n13983), .A2(n15947), .ZN(n9861) );
  NOR3_X1 U11763 ( .A1(n15954), .A2(n16114), .A3(n17717), .ZN(n13983) );
  INV_X1 U11764 ( .A(n15956), .ZN(n17827) );
  NOR2_X1 U11765 ( .A1(n21010), .A2(n16808), .ZN(n16794) );
  AND2_X1 U11766 ( .A1(n17928), .A2(n9972), .ZN(n16968) );
  AND2_X1 U11767 ( .A1(n9707), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9972) );
  NOR2_X1 U11768 ( .A1(n10081), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10079) );
  OR2_X1 U11769 ( .A1(n18052), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10081) );
  NAND2_X1 U11770 ( .A1(n16129), .A2(n18378), .ZN(n9953) );
  NOR2_X1 U11771 ( .A1(n15953), .A2(n16101), .ZN(n19052) );
  INV_X1 U11772 ( .A(n18122), .ZN(n18453) );
  NOR2_X1 U11773 ( .A1(n16091), .A2(n16092), .ZN(n16093) );
  OR2_X1 U11774 ( .A1(n18202), .A2(n10095), .ZN(n9952) );
  OR2_X1 U11775 ( .A1(n18189), .A2(n18526), .ZN(n10095) );
  NAND2_X1 U11776 ( .A1(n16093), .A2(n10094), .ZN(n10093) );
  INV_X1 U11777 ( .A(n18189), .ZN(n10094) );
  OR2_X1 U11778 ( .A1(n18202), .A2(n18526), .ZN(n10097) );
  NAND2_X1 U11779 ( .A1(n9739), .A2(n9962), .ZN(n10090) );
  INV_X1 U11780 ( .A(n18226), .ZN(n9962) );
  NAND2_X1 U11781 ( .A1(n16088), .A2(n10089), .ZN(n10088) );
  INV_X1 U11782 ( .A(n18216), .ZN(n10089) );
  OR2_X1 U11783 ( .A1(n18226), .A2(n18549), .ZN(n10092) );
  AOI211_X1 U11784 ( .C1(n15931), .C2(n16105), .A(n15934), .B(n15933), .ZN(
        n19038) );
  NOR2_X1 U11785 ( .A1(n13956), .A2(n13955), .ZN(n18625) );
  NOR2_X1 U11786 ( .A1(n19102), .A2(n19261), .ZN(n19090) );
  INV_X1 U11787 ( .A(n20372), .ZN(n20354) );
  OR2_X1 U11788 ( .A1(n14472), .A2(n14473), .ZN(n9844) );
  OR2_X1 U11789 ( .A1(n20457), .A2(n12385), .ZN(n16333) );
  INV_X1 U11790 ( .A(n20456), .ZN(n14888) );
  INV_X1 U11791 ( .A(n20457), .ZN(n20299) );
  INV_X1 U11792 ( .A(n20503), .ZN(n20481) );
  INV_X1 U11793 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20693) );
  NAND2_X1 U11794 ( .A1(n12502), .A2(n12575), .ZN(n15009) );
  CLKBUF_X1 U11795 ( .A(n20658), .Z(n20622) );
  INV_X1 U11796 ( .A(n12597), .ZN(n12598) );
  NAND2_X1 U11797 ( .A1(n9824), .A2(n12657), .ZN(n12940) );
  NOR2_X1 U11798 ( .A1(n11867), .A2(n11808), .ZN(n19272) );
  NAND2_X1 U11799 ( .A1(n16731), .A2(n20122), .ZN(n19275) );
  AND2_X1 U11800 ( .A1(n10742), .A2(n10036), .ZN(n15178) );
  AND2_X1 U11801 ( .A1(n15291), .A2(n10102), .ZN(n15281) );
  AND2_X1 U11802 ( .A1(n16666), .A2(n16203), .ZN(n19538) );
  OR2_X1 U11803 ( .A1(n19275), .A2(n9659), .ZN(n19534) );
  OR2_X1 U11804 ( .A1(n19275), .A2(n20281), .ZN(n19532) );
  INV_X1 U11805 ( .A(n19534), .ZN(n16662) );
  OR2_X1 U11806 ( .A1(n10168), .A2(n11416), .ZN(n10167) );
  XNOR2_X1 U11807 ( .A(n11035), .B(n11034), .ZN(n11385) );
  OAI21_X1 U11808 ( .B1(n11390), .B2(n16710), .A(n10110), .ZN(n10109) );
  INV_X1 U11809 ( .A(n11382), .ZN(n10110) );
  OR2_X1 U11810 ( .A1(n10077), .A2(n15609), .ZN(n10076) );
  OAI21_X1 U11811 ( .B1(n15612), .B2(n15611), .A(n15606), .ZN(n10077) );
  NAND2_X1 U11812 ( .A1(n15301), .A2(n15302), .ZN(n16541) );
  NAND2_X1 U11813 ( .A1(n10826), .A2(n9897), .ZN(n9894) );
  NAND2_X1 U11814 ( .A1(n9896), .A2(n10827), .ZN(n9895) );
  INV_X1 U11815 ( .A(n16702), .ZN(n16689) );
  INV_X1 U11816 ( .A(n16697), .ZN(n16673) );
  OR2_X1 U11817 ( .A1(n11370), .A2(n16711), .ZN(n16710) );
  OR2_X1 U11818 ( .A1(n11370), .A2(n11343), .ZN(n16702) );
  INV_X1 U11819 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20252) );
  INV_X1 U11820 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20236) );
  OR2_X1 U11821 ( .A1(n16993), .A2(n9979), .ZN(n9978) );
  NAND2_X1 U11822 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  NAND2_X1 U11823 ( .A1(n17267), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9980) );
  INV_X1 U11824 ( .A(n16995), .ZN(n9977) );
  NOR2_X1 U11825 ( .A1(n16996), .A2(n17261), .ZN(n16990) );
  NOR2_X1 U11826 ( .A1(n17083), .A2(n18013), .ZN(n17082) );
  AND2_X1 U11827 ( .A1(n9861), .A2(n9860), .ZN(n17621) );
  NOR3_X1 U11828 ( .A1(n18613), .A2(n18609), .A3(n19254), .ZN(n9860) );
  AND2_X1 U11829 ( .A1(n17621), .A2(n17717), .ZN(n17625) );
  OAI211_X1 U11830 ( .C1(n12011), .C2(n12012), .A(n12010), .B(n12020), .ZN(
        n9839) );
  NAND2_X1 U11831 ( .A1(n12008), .A2(n12011), .ZN(n9838) );
  NAND2_X1 U11832 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  INV_X1 U11833 ( .A(n12013), .ZN(n9836) );
  INV_X1 U11834 ( .A(n12173), .ZN(n9987) );
  INV_X1 U11835 ( .A(n13262), .ZN(n11037) );
  NAND2_X1 U11836 ( .A1(n11358), .A2(n10377), .ZN(n10400) );
  AND4_X1 U11837 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10539) );
  AND4_X1 U11838 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n20281), .ZN(
        n10538) );
  AND2_X1 U11839 ( .A1(n9744), .A2(n10475), .ZN(n9868) );
  NAND2_X1 U11840 ( .A1(n10466), .A2(n9734), .ZN(n9792) );
  NOR2_X1 U11841 ( .A1(n10011), .A2(n10465), .ZN(n10009) );
  NAND2_X1 U11842 ( .A1(n20058), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9890) );
  NAND2_X1 U11843 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10443) );
  OR2_X1 U11844 ( .A1(n10551), .A2(n10550), .ZN(n10586) );
  NOR2_X1 U11845 ( .A1(n11347), .A2(n20278), .ZN(n9825) );
  XNOR2_X1 U11846 ( .A(n9802), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10600) );
  OR2_X1 U11847 ( .A1(n12856), .A2(n12855), .ZN(n13622) );
  NAND2_X1 U11848 ( .A1(n9926), .A2(n12861), .ZN(n12862) );
  NAND2_X1 U11849 ( .A1(n13044), .A2(n13647), .ZN(n12003) );
  AND2_X1 U11850 ( .A1(n12340), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12328) );
  NAND2_X1 U11851 ( .A1(n13262), .A2(n11044), .ZN(n10019) );
  INV_X1 U11852 ( .A(n10713), .ZN(n10030) );
  INV_X1 U11853 ( .A(n11044), .ZN(n10021) );
  NOR2_X1 U11854 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11587) );
  INV_X1 U11855 ( .A(n15294), .ZN(n9923) );
  OR2_X1 U11856 ( .A1(n10705), .A2(n10704), .ZN(n10711) );
  AND2_X1 U11857 ( .A1(n19590), .A2(n11352), .ZN(n10363) );
  AND2_X1 U11858 ( .A1(n10164), .A2(n10868), .ZN(n10163) );
  NAND2_X1 U11859 ( .A1(n9763), .A2(n10869), .ZN(n10164) );
  NAND2_X1 U11860 ( .A1(n9725), .A2(n10023), .ZN(n10022) );
  NOR2_X1 U11861 ( .A1(n10520), .A2(n9737), .ZN(n10023) );
  INV_X1 U11862 ( .A(n10351), .ZN(n9803) );
  INV_X1 U11863 ( .A(n10348), .ZN(n9799) );
  OR2_X1 U11864 ( .A1(n10507), .A2(n10506), .ZN(n10581) );
  NAND2_X1 U11865 ( .A1(n12094), .A2(n20281), .ZN(n11732) );
  NAND2_X1 U11866 ( .A1(n10360), .A2(n10374), .ZN(n10361) );
  AND2_X1 U11867 ( .A1(n11067), .A2(n10102), .ZN(n10380) );
  NAND2_X1 U11868 ( .A1(n11352), .A2(n10372), .ZN(n10371) );
  NOR2_X1 U11869 ( .A1(n10447), .A2(n10449), .ZN(n10467) );
  NAND2_X1 U11870 ( .A1(n9795), .A2(n12104), .ZN(n10471) );
  AND2_X1 U11871 ( .A1(n10264), .A2(n9802), .ZN(n10269) );
  NAND2_X1 U11872 ( .A1(n10577), .A2(n10576), .ZN(n10585) );
  INV_X1 U11873 ( .A(n10574), .ZN(n10577) );
  NAND2_X1 U11874 ( .A1(n10570), .A2(n10569), .ZN(n11038) );
  NOR2_X1 U11875 ( .A1(n9714), .A2(n17618), .ZN(n10086) );
  AOI22_X1 U11876 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U11877 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11985) );
  NOR2_X1 U11878 ( .A1(n10177), .A2(n14512), .ZN(n10176) );
  NAND2_X1 U11879 ( .A1(n14473), .A2(n10178), .ZN(n10177) );
  INV_X1 U11880 ( .A(n14522), .ZN(n10178) );
  INV_X1 U11881 ( .A(n14548), .ZN(n9851) );
  AND2_X1 U11882 ( .A1(n9757), .A2(n9853), .ZN(n9852) );
  INV_X1 U11883 ( .A(n14614), .ZN(n9853) );
  NOR2_X1 U11884 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10205) );
  AND2_X1 U11885 ( .A1(n10180), .A2(n14629), .ZN(n10179) );
  INV_X1 U11886 ( .A(n16268), .ZN(n10181) );
  NOR2_X1 U11887 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  INV_X1 U11888 ( .A(n13800), .ZN(n9849) );
  INV_X1 U11889 ( .A(n13863), .ZN(n9850) );
  NAND2_X1 U11890 ( .A1(n10173), .A2(n13166), .ZN(n10172) );
  INV_X1 U11891 ( .A(n13171), .ZN(n10173) );
  AND2_X1 U11892 ( .A1(n9820), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12865) );
  NAND2_X1 U11893 ( .A1(n14779), .A2(n14797), .ZN(n14439) );
  INV_X1 U11894 ( .A(n14832), .ZN(n9935) );
  INV_X1 U11895 ( .A(n14660), .ZN(n10006) );
  NAND2_X1 U11896 ( .A1(n14855), .A2(n14429), .ZN(n14838) );
  INV_X1 U11897 ( .A(n13637), .ZN(n10195) );
  INV_X1 U11898 ( .A(n16385), .ZN(n10191) );
  NAND2_X1 U11899 ( .A1(n13637), .A2(n10194), .ZN(n10193) );
  INV_X1 U11900 ( .A(n13630), .ZN(n10194) );
  INV_X1 U11901 ( .A(n14417), .ZN(n14399) );
  NAND2_X1 U11902 ( .A1(n13166), .A2(n9944), .ZN(n9943) );
  INV_X1 U11903 ( .A(n12883), .ZN(n9944) );
  INV_X1 U11904 ( .A(n13651), .ZN(n13647) );
  INV_X1 U11905 ( .A(n12994), .ZN(n9814) );
  NAND2_X1 U11906 ( .A1(n12986), .A2(n12985), .ZN(n13610) );
  NAND2_X1 U11907 ( .A1(n12183), .A2(n9732), .ZN(n12192) );
  NAND2_X1 U11908 ( .A1(n9942), .A2(n12617), .ZN(n9941) );
  INV_X1 U11909 ( .A(n12501), .ZN(n9942) );
  OR2_X1 U11910 ( .A1(n12667), .A2(n12666), .ZN(n13623) );
  INV_X1 U11911 ( .A(n12265), .ZN(n12340) );
  OAI21_X1 U11912 ( .B1(n12179), .B2(n12178), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12180) );
  OR2_X1 U11913 ( .A1(n11970), .A2(n11967), .ZN(n11968) );
  AOI21_X1 U11914 ( .B1(n9831), .B2(n12016), .A(n9830), .ZN(n12025) );
  OR2_X1 U11915 ( .A1(n12003), .A2(n11996), .ZN(n12027) );
  AND2_X1 U11916 ( .A1(n12054), .A2(n12053), .ZN(n12063) );
  NAND2_X1 U11917 ( .A1(n10812), .A2(n10811), .ZN(n10817) );
  NAND2_X1 U11918 ( .A1(n12471), .A2(n19339), .ZN(n10026) );
  NAND2_X1 U11919 ( .A1(n10031), .A2(n10027), .ZN(n10724) );
  NOR2_X1 U11920 ( .A1(n10659), .A2(n10030), .ZN(n10027) );
  OAI21_X1 U11921 ( .B1(n10580), .B2(n11007), .A(n10579), .ZN(n10589) );
  NAND2_X1 U11922 ( .A1(n11007), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10579) );
  OAI21_X1 U11923 ( .B1(n11112), .B2(n13262), .A(n10020), .ZN(n10580) );
  NAND2_X1 U11924 ( .A1(n13262), .A2(n10021), .ZN(n10020) );
  INV_X1 U11925 ( .A(n11573), .ZN(n11608) );
  INV_X1 U11926 ( .A(n11563), .ZN(n11629) );
  INV_X1 U11927 ( .A(n11565), .ZN(n11625) );
  AND2_X1 U11928 ( .A1(n11666), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11575) );
  INV_X1 U11929 ( .A(n15326), .ZN(n10068) );
  AND2_X1 U11930 ( .A1(n15334), .A2(n15343), .ZN(n10069) );
  INV_X1 U11931 ( .A(n13578), .ZN(n10234) );
  AND2_X1 U11932 ( .A1(n10237), .A2(n10236), .ZN(n10235) );
  INV_X1 U11933 ( .A(n13431), .ZN(n10236) );
  INV_X1 U11934 ( .A(n15405), .ZN(n15391) );
  NOR2_X1 U11935 ( .A1(n15089), .A2(n10042), .ZN(n10041) );
  NOR2_X1 U11936 ( .A1(n13397), .A2(n10123), .ZN(n10122) );
  INV_X1 U11937 ( .A(n13299), .ZN(n10123) );
  AND2_X1 U11938 ( .A1(n10122), .A2(n10121), .ZN(n10120) );
  INV_X1 U11939 ( .A(n13440), .ZN(n10121) );
  NOR2_X1 U11940 ( .A1(n15563), .A2(n10051), .ZN(n10050) );
  INV_X1 U11941 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U11942 ( .A1(n16656), .A2(n10046), .ZN(n10045) );
  AOI21_X1 U11943 ( .B1(n10433), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10432), .ZN(n10898) );
  NAND2_X1 U11944 ( .A1(n10425), .A2(n10424), .ZN(n9863) );
  INV_X1 U11945 ( .A(n10815), .ZN(n11009) );
  NOR2_X1 U11946 ( .A1(n10995), .A2(n15626), .ZN(n10133) );
  NAND2_X1 U11947 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10169) );
  AND2_X1 U11948 ( .A1(n16551), .A2(n11137), .ZN(n10992) );
  OR2_X1 U11949 ( .A1(n16563), .A2(n10717), .ZN(n10825) );
  AND2_X1 U11950 ( .A1(n9687), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10014) );
  INV_X1 U11951 ( .A(n9910), .ZN(n9902) );
  INV_X1 U11952 ( .A(n9907), .ZN(n9906) );
  AND2_X1 U11953 ( .A1(n11318), .A2(n11317), .ZN(n15118) );
  NOR2_X1 U11954 ( .A1(n15694), .A2(n11366), .ZN(n10170) );
  OR2_X1 U11955 ( .A1(n19305), .A2(n10717), .ZN(n10789) );
  AND3_X1 U11956 ( .A1(n10908), .A2(n10907), .A3(n10906), .ZN(n12406) );
  INV_X1 U11957 ( .A(n10022), .ZN(n11112) );
  INV_X1 U11958 ( .A(n10581), .ZN(n11108) );
  NAND2_X1 U11959 ( .A1(n11430), .A2(n11429), .ZN(n11433) );
  OR2_X1 U11960 ( .A1(n11732), .A2(n11160), .ZN(n11434) );
  INV_X1 U11961 ( .A(n11427), .ZN(n10218) );
  NOR2_X1 U11962 ( .A1(n10221), .A2(n10216), .ZN(n10213) );
  NAND2_X1 U11963 ( .A1(n10219), .A2(n10216), .ZN(n10215) );
  INV_X1 U11964 ( .A(n11045), .ZN(n11803) );
  INV_X1 U11965 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U11966 ( .A1(n11439), .A2(n11440), .ZN(n11446) );
  AND2_X1 U11967 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11447) );
  NOR2_X1 U11968 ( .A1(n10471), .A2(n10441), .ZN(n10619) );
  AND2_X1 U11969 ( .A1(n10312), .A2(n9802), .ZN(n10316) );
  NAND3_X1 U11970 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20223), .A3(n20067), 
        .ZN(n19544) );
  AOI221_X1 U11971 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10836), 
        .C1(n20221), .C2(n10836), .A(n10835), .ZN(n11053) );
  NOR3_X1 U11972 ( .A1(n16101), .A2(n16102), .A3(n16114), .ZN(n15950) );
  OR2_X1 U11973 ( .A1(n17321), .A2(n13883), .ZN(n10251) );
  OR2_X1 U11974 ( .A1(n19061), .A2(n13883), .ZN(n9720) );
  INV_X1 U11975 ( .A(n17584), .ZN(n13962) );
  NOR2_X1 U11976 ( .A1(n16971), .A2(n9974), .ZN(n9973) );
  INV_X1 U11977 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9974) );
  AND2_X1 U11978 ( .A1(n10101), .A2(n18168), .ZN(n10100) );
  XNOR2_X1 U11979 ( .A(n17770), .B(n16081), .ZN(n16083) );
  NOR2_X1 U11980 ( .A1(n13982), .A2(n15965), .ZN(n15947) );
  AND2_X1 U11981 ( .A1(n13007), .A2(n16503), .ZN(n12384) );
  NAND2_X1 U11982 ( .A1(n16253), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16291) );
  NOR2_X1 U11983 ( .A1(n20803), .A2(n14563), .ZN(n16253) );
  NAND2_X1 U11984 ( .A1(n14589), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14563) );
  NAND2_X1 U11985 ( .A1(n20325), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14599) );
  AND2_X1 U11986 ( .A1(n13349), .A2(n13348), .ZN(n13351) );
  INV_X1 U11987 ( .A(n12609), .ZN(n12606) );
  NAND3_X1 U11988 ( .A1(n9994), .A2(n9736), .A3(n12474), .ZN(n9996) );
  OR2_X1 U11989 ( .A1(n14417), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n9994) );
  INV_X1 U11990 ( .A(n14405), .ZN(n14457) );
  AND2_X1 U11991 ( .A1(n14383), .A2(n14382), .ZN(n14566) );
  AND2_X1 U11992 ( .A1(n12140), .A2(n16165), .ZN(n20396) );
  AND2_X1 U11993 ( .A1(n20697), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14444) );
  NAND2_X1 U11994 ( .A1(n10176), .A2(n14443), .ZN(n10175) );
  NOR2_X1 U11995 ( .A1(n14270), .A2(n14791), .ZN(n14289) );
  AOI21_X1 U11996 ( .B1(n14795), .B2(n12477), .A(n14288), .ZN(n14534) );
  NAND2_X1 U11997 ( .A1(n13003), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14251) );
  INV_X1 U11998 ( .A(n14231), .ZN(n13003) );
  NOR2_X1 U11999 ( .A1(n14164), .A2(n16261), .ZN(n14167) );
  NAND2_X1 U12000 ( .A1(n14167), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14199) );
  NOR2_X1 U12001 ( .A1(n14116), .A2(n16280), .ZN(n14134) );
  NAND2_X1 U12002 ( .A1(n14134), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14164) );
  OR2_X1 U12003 ( .A1(n14100), .A2(n16289), .ZN(n14116) );
  OR2_X1 U12004 ( .A1(n14080), .A2(n14571), .ZN(n14100) );
  NAND2_X1 U12005 ( .A1(n13847), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14080) );
  NAND2_X1 U12006 ( .A1(n13001), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13754) );
  INV_X1 U12007 ( .A(n13779), .ZN(n13001) );
  NOR2_X1 U12008 ( .A1(n10185), .A2(n10183), .ZN(n10182) );
  OR2_X1 U12009 ( .A1(n13783), .A2(n10186), .ZN(n10185) );
  INV_X1 U12010 ( .A(n10187), .ZN(n10183) );
  AND2_X1 U12011 ( .A1(n13462), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13751) );
  NAND2_X1 U12012 ( .A1(n13751), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13779) );
  NOR2_X1 U12013 ( .A1(n13374), .A2(n20315), .ZN(n13462) );
  NAND2_X1 U12014 ( .A1(n13334), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13374) );
  INV_X1 U12015 ( .A(n13172), .ZN(n13334) );
  INV_X1 U12016 ( .A(n13045), .ZN(n13173) );
  NAND2_X1 U12017 ( .A1(n13173), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13172) );
  NAND2_X1 U12018 ( .A1(n13046), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13045) );
  INV_X1 U12019 ( .A(n12887), .ZN(n12888) );
  NAND2_X1 U12020 ( .A1(n12888), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13000) );
  NAND2_X1 U12021 ( .A1(n12886), .A2(n13859), .ZN(n12893) );
  NAND2_X1 U12022 ( .A1(n12864), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12887) );
  NAND2_X1 U12023 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12744) );
  NOR2_X1 U12024 ( .A1(n12744), .A2(n12743), .ZN(n12864) );
  INV_X1 U12025 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U12026 ( .A1(n12742), .A2(n12741), .ZN(n12752) );
  NAND2_X1 U12027 ( .A1(n12752), .A2(n12751), .ZN(n12970) );
  XNOR2_X1 U12028 ( .A(n12612), .B(n12545), .ZN(n12546) );
  AOI21_X1 U12029 ( .B1(n13539), .B2(n12905), .A(n20697), .ZN(n12238) );
  OR2_X1 U12030 ( .A1(n14537), .A2(n14523), .ZN(n14525) );
  INV_X1 U12031 ( .A(n14765), .ZN(n9930) );
  AND2_X1 U12032 ( .A1(n9704), .A2(n14549), .ZN(n9998) );
  NAND2_X1 U12033 ( .A1(n14638), .A2(n14631), .ZN(n14633) );
  NAND2_X1 U12034 ( .A1(n14638), .A2(n10000), .ZN(n14624) );
  NOR2_X1 U12035 ( .A1(n16272), .A2(n14396), .ZN(n14647) );
  NAND2_X1 U12036 ( .A1(n10200), .A2(n10202), .ZN(n14833) );
  AOI21_X1 U12037 ( .B1(n14838), .B2(n16341), .A(n9927), .ZN(n16342) );
  NAND2_X1 U12038 ( .A1(n14845), .A2(n14843), .ZN(n9927) );
  NOR3_X1 U12039 ( .A1(n13869), .A2(n10008), .A3(n13868), .ZN(n14661) );
  NOR2_X1 U12040 ( .A1(n13869), .A2(n13868), .ZN(n14567) );
  OR2_X1 U12041 ( .A1(n13826), .A2(n13816), .ZN(n13869) );
  NAND2_X1 U12042 ( .A1(n16295), .A2(n13825), .ZN(n13826) );
  NOR2_X1 U12043 ( .A1(n16296), .A2(n16297), .ZN(n16295) );
  NAND2_X1 U12044 ( .A1(n9993), .A2(n9992), .ZN(n16296) );
  INV_X1 U12045 ( .A(n13833), .ZN(n9992) );
  AND2_X1 U12046 ( .A1(n13358), .A2(n13357), .ZN(n13413) );
  OR2_X1 U12047 ( .A1(n20369), .A2(n12901), .ZN(n20370) );
  INV_X1 U12048 ( .A(n20498), .ZN(n20484) );
  NOR2_X1 U12049 ( .A1(n9996), .A2(n9995), .ZN(n12706) );
  NOR2_X1 U12050 ( .A1(n12475), .A2(n14456), .ZN(n9995) );
  AND2_X1 U12051 ( .A1(n20498), .A2(n16473), .ZN(n16476) );
  AND2_X1 U12052 ( .A1(n14454), .A2(n12753), .ZN(n14405) );
  NAND2_X1 U12053 ( .A1(n12496), .A2(n13652), .ZN(n12578) );
  AOI21_X1 U12054 ( .B1(n9939), .B2(n9940), .A(n9937), .ZN(n12496) );
  NOR2_X1 U12055 ( .A1(n9941), .A2(n9938), .ZN(n9937) );
  AND2_X1 U12056 ( .A1(n12271), .A2(n9729), .ZN(n9939) );
  AND3_X1 U12057 ( .A1(n12501), .A2(n12500), .A3(n12499), .ZN(n12575) );
  NAND2_X1 U12058 ( .A1(n9823), .A2(n12595), .ZN(n12597) );
  AND3_X1 U12059 ( .A1(n12321), .A2(n12060), .A3(n12172), .ZN(n12791) );
  OAI211_X1 U12060 ( .C1(n15073), .C2(n16512), .A(n20527), .B(n15039), .ZN(
        n15072) );
  NOR2_X1 U12061 ( .A1(n13675), .A2(n13496), .ZN(n20527) );
  OR2_X1 U12062 ( .A1(n15012), .A2(n12672), .ZN(n20655) );
  INV_X1 U12063 ( .A(n20655), .ZN(n15035) );
  NOR2_X1 U12064 ( .A1(n15009), .A2(n13539), .ZN(n13670) );
  INV_X1 U12065 ( .A(n20704), .ZN(n13491) );
  AND2_X1 U12066 ( .A1(n15009), .A2(n13539), .ZN(n12939) );
  AND2_X1 U12067 ( .A1(n16510), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12265) );
  NOR2_X1 U12068 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20270) );
  NAND2_X1 U12069 ( .A1(n10999), .A2(n11000), .ZN(n11004) );
  AND2_X1 U12070 ( .A1(n15391), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15393) );
  AND2_X1 U12071 ( .A1(n10813), .A2(n10817), .ZN(n10815) );
  NAND2_X1 U12072 ( .A1(n15119), .A2(n9661), .ZN(n15107) );
  NAND2_X1 U12073 ( .A1(n15107), .A2(n15436), .ZN(n16514) );
  NAND2_X1 U12074 ( .A1(n10795), .A2(n10794), .ZN(n10799) );
  NAND2_X1 U12075 ( .A1(n10072), .A2(n10073), .ZN(n15135) );
  AND2_X1 U12076 ( .A1(n11310), .A2(n11309), .ZN(n13580) );
  NOR2_X1 U12077 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  INV_X1 U12078 ( .A(n13432), .ZN(n10064) );
  NOR2_X1 U12079 ( .A1(n15781), .A2(n10065), .ZN(n13433) );
  NAND2_X1 U12080 ( .A1(n10742), .A2(n10743), .ZN(n10748) );
  AND2_X1 U12081 ( .A1(n10731), .A2(n10024), .ZN(n10736) );
  INV_X1 U12082 ( .A(n10026), .ZN(n10024) );
  NOR2_X1 U12083 ( .A1(n10659), .A2(n10658), .ZN(n10663) );
  INV_X1 U12084 ( .A(n19411), .ZN(n19352) );
  NOR2_X1 U12085 ( .A1(n9917), .A2(n11771), .ZN(n9916) );
  INV_X1 U12086 ( .A(n15226), .ZN(n9917) );
  AND2_X1 U12087 ( .A1(n11731), .A2(n11730), .ZN(n15230) );
  NAND2_X1 U12088 ( .A1(n15083), .A2(n9770), .ZN(n15324) );
  NAND2_X1 U12089 ( .A1(n15083), .A2(n10069), .ZN(n15336) );
  XNOR2_X1 U12090 ( .A(n11690), .B(n11686), .ZN(n15253) );
  NAND2_X1 U12091 ( .A1(n15253), .A2(n15252), .ZN(n15251) );
  AND2_X1 U12092 ( .A1(n15083), .A2(n15343), .ZN(n15345) );
  NOR2_X1 U12093 ( .A1(n15260), .A2(n15259), .ZN(n15258) );
  AND2_X1 U12094 ( .A1(n11320), .A2(n11319), .ZN(n15084) );
  NAND2_X1 U12095 ( .A1(n10224), .A2(n11661), .ZN(n10223) );
  OR2_X1 U12096 ( .A1(n15284), .A2(n10227), .ZN(n10226) );
  INV_X1 U12097 ( .A(n10230), .ZN(n10228) );
  AND2_X1 U12098 ( .A1(n11314), .A2(n11313), .ZN(n15364) );
  NOR2_X1 U12099 ( .A1(n15363), .A2(n15364), .ZN(n15362) );
  NAND2_X1 U12100 ( .A1(n15284), .A2(n15286), .ZN(n15285) );
  NOR2_X1 U12101 ( .A1(n9925), .A2(n9920), .ZN(n15295) );
  NAND2_X1 U12102 ( .A1(n9701), .A2(n12831), .ZN(n9920) );
  NAND2_X1 U12103 ( .A1(n12829), .A2(n10235), .ZN(n13577) );
  NAND2_X1 U12104 ( .A1(n11284), .A2(n10254), .ZN(n15782) );
  AND3_X1 U12105 ( .A1(n11235), .A2(n11234), .A3(n11233), .ZN(n13257) );
  AND2_X1 U12106 ( .A1(n11099), .A2(n11113), .ZN(n10053) );
  AND2_X1 U12107 ( .A1(n19463), .A2(n10355), .ZN(n19426) );
  INV_X1 U12108 ( .A(n20277), .ZN(n12245) );
  AND2_X1 U12109 ( .A1(n12244), .A2(n20280), .ZN(n19494) );
  OAI21_X1 U12110 ( .B1(n11820), .B2(n11819), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12447) );
  INV_X1 U12111 ( .A(n12447), .ZN(n19545) );
  NAND2_X1 U12112 ( .A1(n15391), .A2(n9706), .ZN(n15381) );
  NAND2_X1 U12113 ( .A1(n15092), .A2(n10040), .ZN(n15425) );
  AND2_X1 U12114 ( .A1(n9703), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10040) );
  NOR2_X1 U12115 ( .A1(n15425), .A2(n15415), .ZN(n15414) );
  NAND2_X1 U12116 ( .A1(n15117), .A2(n10115), .ZN(n15266) );
  NAND2_X1 U12117 ( .A1(n15117), .A2(n15080), .ZN(n15264) );
  INV_X1 U12118 ( .A(n15093), .ZN(n15092) );
  NAND2_X1 U12119 ( .A1(n15092), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15091) );
  NOR2_X1 U12120 ( .A1(n15105), .A2(n15494), .ZN(n15094) );
  AND2_X1 U12121 ( .A1(n13300), .A2(n10118), .ZN(n15151) );
  AND2_X1 U12122 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  INV_X1 U12123 ( .A(n13667), .ZN(n10119) );
  NOR2_X1 U12124 ( .A1(n15103), .A2(n15515), .ZN(n15106) );
  NAND2_X1 U12125 ( .A1(n15106), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15105) );
  NAND2_X1 U12126 ( .A1(n13300), .A2(n10122), .ZN(n13441) );
  NAND2_X1 U12127 ( .A1(n13300), .A2(n10120), .ZN(n13666) );
  AND2_X1 U12128 ( .A1(n13245), .A2(n10049), .ZN(n15104) );
  AND2_X1 U12129 ( .A1(n9689), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10049) );
  NAND2_X1 U12130 ( .A1(n15104), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15103) );
  AND2_X1 U12131 ( .A1(n13095), .A2(n12976), .ZN(n13300) );
  NAND2_X1 U12132 ( .A1(n13300), .A2(n13299), .ZN(n13398) );
  NAND2_X1 U12133 ( .A1(n13245), .A2(n9689), .ZN(n15102) );
  INV_X1 U12134 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15563) );
  NAND2_X1 U12135 ( .A1(n13245), .A2(n10050), .ZN(n15100) );
  NOR2_X2 U12136 ( .A1(n13094), .A2(n13093), .ZN(n13095) );
  NAND2_X1 U12137 ( .A1(n13245), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15099) );
  NOR2_X1 U12138 ( .A1(n13244), .A2(n16635), .ZN(n13245) );
  NAND2_X1 U12139 ( .A1(n13242), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13244) );
  AND2_X1 U12140 ( .A1(n13239), .A2(n10044), .ZN(n13242) );
  AND2_X1 U12141 ( .A1(n9690), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10044) );
  NAND2_X1 U12142 ( .A1(n13239), .A2(n9690), .ZN(n13240) );
  AND2_X1 U12143 ( .A1(n13239), .A2(n10045), .ZN(n13241) );
  NOR2_X1 U12144 ( .A1(n12407), .A2(n12406), .ZN(n12557) );
  NAND2_X1 U12145 ( .A1(n13239), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13238) );
  NOR2_X1 U12146 ( .A1(n16667), .A2(n13236), .ZN(n13239) );
  NAND2_X1 U12147 ( .A1(n13237), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13236) );
  AND3_X1 U12148 ( .A1(n10905), .A2(n10904), .A3(n10903), .ZN(n12370) );
  OR2_X1 U12149 ( .A1(n12371), .A2(n12370), .ZN(n12407) );
  NOR2_X1 U12150 ( .A1(n13157), .A2(n13273), .ZN(n13237) );
  INV_X1 U12151 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13273) );
  OR2_X1 U12152 ( .A1(n10169), .A2(n15611), .ZN(n10168) );
  NAND2_X1 U12153 ( .A1(n10993), .A2(n10992), .ZN(n10134) );
  INV_X1 U12154 ( .A(n10125), .ZN(n10124) );
  OAI21_X1 U12155 ( .B1(n10130), .B2(n10133), .A(n15375), .ZN(n10125) );
  NAND2_X1 U12156 ( .A1(n10126), .A2(n15375), .ZN(n10128) );
  AND2_X1 U12157 ( .A1(n10113), .A2(n15248), .ZN(n10112) );
  INV_X1 U12158 ( .A(n15411), .ZN(n10146) );
  NAND2_X1 U12159 ( .A1(n9909), .A2(n9722), .ZN(n9903) );
  INV_X1 U12160 ( .A(n9883), .ZN(n9882) );
  NAND2_X1 U12161 ( .A1(n13325), .A2(n10062), .ZN(n15198) );
  INV_X1 U12162 ( .A(n15819), .ZN(n10060) );
  INV_X1 U12163 ( .A(n12570), .ZN(n12835) );
  NAND2_X1 U12164 ( .A1(n10104), .A2(n10103), .ZN(n12570) );
  NOR2_X1 U12165 ( .A1(n10106), .A2(n10105), .ZN(n10103) );
  INV_X1 U12166 ( .A(n12407), .ZN(n10104) );
  INV_X1 U12167 ( .A(n12568), .ZN(n10105) );
  NOR2_X1 U12168 ( .A1(n12407), .A2(n10106), .ZN(n12569) );
  INV_X1 U12169 ( .A(n10716), .ZN(n9885) );
  AND2_X1 U12170 ( .A1(n11137), .A2(n10052), .ZN(n11138) );
  OAI21_X1 U12171 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n13589) );
  INV_X1 U12172 ( .A(n10868), .ZN(n9789) );
  NAND2_X1 U12173 ( .A1(n9790), .A2(n10870), .ZN(n9788) );
  NAND2_X1 U12174 ( .A1(n9873), .A2(n9870), .ZN(n13419) );
  INV_X1 U12175 ( .A(n9871), .ZN(n9870) );
  OAI21_X1 U12176 ( .B1(n9878), .B2(n9872), .A(n9877), .ZN(n9871) );
  OR2_X1 U12177 ( .A1(n11370), .A2(n16720), .ZN(n12110) );
  OR2_X1 U12178 ( .A1(n11370), .A2(n11365), .ZN(n15743) );
  NAND2_X1 U12179 ( .A1(n12109), .A2(n12108), .ZN(n12107) );
  NOR2_X1 U12180 ( .A1(n11423), .A2(n20278), .ZN(n12094) );
  AND2_X2 U12181 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15883) );
  AOI21_X1 U12182 ( .B1(n10437), .B2(n11440), .A(n11432), .ZN(n12100) );
  AND2_X1 U12183 ( .A1(n13235), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10048) );
  INV_X1 U12184 ( .A(n19990), .ZN(n19984) );
  INV_X1 U12185 ( .A(n19927), .ZN(n19991) );
  NAND2_X2 U12186 ( .A1(n10294), .A2(n10293), .ZN(n19564) );
  INV_X1 U12187 ( .A(n19583), .ZN(n19585) );
  NAND2_X1 U12189 ( .A1(n10208), .A2(n10207), .ZN(n11866) );
  NOR2_X1 U12190 ( .A1(n11070), .A2(n10332), .ZN(n10208) );
  AOI21_X1 U12191 ( .B1(n15935), .B2(n15934), .A(n15933), .ZN(n19041) );
  NOR2_X1 U12192 ( .A1(n16962), .A2(n16961), .ZN(n19040) );
  OR2_X1 U12193 ( .A1(n17004), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U12194 ( .A1(n17041), .A2(n9856), .ZN(n9855) );
  INV_X1 U12195 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U12196 ( .A1(n17509), .A2(n9712), .ZN(n17456) );
  NOR2_X1 U12197 ( .A1(n17148), .A2(n9858), .ZN(n9857) );
  INV_X1 U12198 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U12199 ( .A1(n10082), .A2(n9728), .ZN(n16078) );
  NOR3_X1 U12200 ( .A1(n10087), .A2(n10084), .A3(n10083), .ZN(n10082) );
  NOR2_X1 U12201 ( .A1(n16960), .A2(n19116), .ZN(n17784) );
  NAND2_X1 U12202 ( .A1(n17928), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17902) );
  NOR2_X1 U12203 ( .A1(n17947), .A2(n17948), .ZN(n17928) );
  NOR2_X1 U12204 ( .A1(n17983), .A2(n16977), .ZN(n17967) );
  NAND2_X1 U12205 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18011), .ZN(
        n17983) );
  NAND2_X1 U12206 ( .A1(n17162), .A2(n9702), .ZN(n18018) );
  NOR2_X1 U12207 ( .A1(n18056), .A2(n9967), .ZN(n9966) );
  NAND2_X1 U12208 ( .A1(n17162), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18055) );
  NOR2_X1 U12209 ( .A1(n18100), .A2(n18102), .ZN(n17162) );
  INV_X1 U12210 ( .A(n17899), .ZN(n18101) );
  NAND2_X1 U12211 ( .A1(n18161), .A2(n18078), .ZN(n18100) );
  NOR2_X1 U12212 ( .A1(n18192), .A2(n18193), .ZN(n18161) );
  NAND2_X1 U12213 ( .A1(n16779), .A2(n10080), .ZN(n16189) );
  NAND2_X1 U12214 ( .A1(n9960), .A2(n9958), .ZN(n17916) );
  NAND2_X1 U12215 ( .A1(n18260), .A2(n17945), .ZN(n18263) );
  NOR2_X1 U12216 ( .A1(n18294), .A2(n18302), .ZN(n17944) );
  OAI21_X1 U12217 ( .B1(n16133), .B2(n16132), .A(n10241), .ZN(n16134) );
  NOR2_X1 U12218 ( .A1(n18167), .A2(n18138), .ZN(n18095) );
  NOR2_X1 U12219 ( .A1(n21047), .A2(n18444), .ZN(n18411) );
  NAND2_X1 U12220 ( .A1(n18613), .A2(n18491), .ZN(n18451) );
  NOR2_X1 U12221 ( .A1(n18497), .A2(n18168), .ZN(n18167) );
  NAND2_X1 U12222 ( .A1(n10098), .A2(n10101), .ZN(n16126) );
  NAND2_X1 U12223 ( .A1(n9724), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18122) );
  INV_X1 U12224 ( .A(n18465), .ZN(n18434) );
  INV_X1 U12225 ( .A(n16098), .ZN(n9950) );
  INV_X1 U12226 ( .A(n18487), .ZN(n18560) );
  XNOR2_X1 U12227 ( .A(n16083), .B(n18562), .ZN(n18233) );
  NOR2_X1 U12228 ( .A1(n18234), .A2(n18233), .ZN(n18232) );
  NOR2_X1 U12229 ( .A1(n16104), .A2(n16103), .ZN(n18507) );
  NOR2_X1 U12230 ( .A1(n13902), .A2(n13901), .ZN(n18609) );
  NOR2_X1 U12231 ( .A1(n13912), .A2(n13911), .ZN(n18621) );
  NOR2_X1 U12232 ( .A1(n13943), .A2(n13942), .ZN(n18629) );
  AOI22_X1 U12233 ( .A1(n19038), .A2(n19037), .B1(n19042), .B2(n18507), .ZN(
        n19046) );
  NAND3_X1 U12234 ( .A1(n16166), .A2(n12534), .A3(n12528), .ZN(n12392) );
  OR2_X1 U12235 ( .A1(n14526), .A2(n14491), .ZN(n14517) );
  NOR2_X1 U12236 ( .A1(n20808), .A2(n16291), .ZN(n16283) );
  NOR2_X1 U12237 ( .A1(n16298), .A2(n20798), .ZN(n14589) );
  INV_X1 U12238 ( .A(n20348), .ZN(n16255) );
  NAND2_X1 U12239 ( .A1(n20381), .A2(n14465), .ZN(n13364) );
  INV_X1 U12240 ( .A(n16303), .ZN(n20329) );
  NOR2_X1 U12241 ( .A1(n13364), .A2(n20793), .ZN(n20325) );
  NOR2_X2 U12242 ( .A1(n14449), .A2(n13013), .ZN(n20348) );
  OR3_X1 U12243 ( .A1(n13025), .A2(n13022), .A3(n13021), .ZN(n20372) );
  AND2_X1 U12244 ( .A1(n16238), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20374) );
  XNOR2_X1 U12245 ( .A(n9996), .B(n12475), .ZN(n13074) );
  INV_X1 U12246 ( .A(n20376), .ZN(n20356) );
  AND2_X1 U12247 ( .A1(n14449), .A2(n13012), .ZN(n20322) );
  OR3_X1 U12248 ( .A1(n13025), .A2(n13017), .A3(n13020), .ZN(n20376) );
  INV_X1 U12249 ( .A(n14666), .ZN(n20387) );
  AND2_X2 U12250 ( .A1(n12171), .A2(n12534), .ZN(n20390) );
  AND2_X1 U12251 ( .A1(n14476), .A2(n14475), .ZN(n21062) );
  NAND2_X1 U12252 ( .A1(n12535), .A2(n12534), .ZN(n21063) );
  INV_X1 U12253 ( .A(n21063), .ZN(n14745) );
  OR2_X1 U12254 ( .A1(n21063), .A2(n12536), .ZN(n14744) );
  BUF_X1 U12255 ( .A(n20413), .Z(n20858) );
  NOR2_X2 U12256 ( .A1(n20442), .A2(n12059), .ZN(n20432) );
  AOI21_X1 U12257 ( .B1(n14742), .B2(n14741), .A(n14740), .ZN(n16363) );
  AND2_X1 U12258 ( .A1(n16504), .A2(n20622), .ZN(n20456) );
  INV_X1 U12259 ( .A(n16333), .ZN(n20450) );
  NOR3_X1 U12260 ( .A1(n16449), .A2(n16438), .A3(n16448), .ZN(n16427) );
  NAND2_X1 U12261 ( .A1(n9807), .A2(n16373), .ZN(n13719) );
  NAND2_X1 U12262 ( .A1(n16376), .A2(n16374), .ZN(n9807) );
  NOR2_X1 U12263 ( .A1(n13730), .A2(n20478), .ZN(n16491) );
  NAND2_X1 U12264 ( .A1(n16384), .A2(n13630), .ZN(n16381) );
  OR2_X1 U12265 ( .A1(n12786), .A2(n12323), .ZN(n20498) );
  INV_X1 U12266 ( .A(n16476), .ZN(n20499) );
  AND2_X1 U12267 ( .A1(n12313), .A2(n12312), .ZN(n20509) );
  AND2_X1 U12268 ( .A1(n12172), .A2(n12280), .ZN(n12311) );
  AND2_X1 U12269 ( .A1(n14902), .A2(n9985), .ZN(n20514) );
  OAI21_X1 U12270 ( .B1(n13539), .B2(n13651), .A(n12296), .ZN(n12297) );
  OR2_X1 U12271 ( .A1(n12323), .A2(n12804), .ZN(n14902) );
  OR2_X1 U12272 ( .A1(n12323), .A2(n12316), .ZN(n20503) );
  INV_X1 U12273 ( .A(n20509), .ZN(n16457) );
  INV_X1 U12274 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20516) );
  OAI21_X1 U12275 ( .B1(n12818), .B2(n16511), .A(n13496), .ZN(n20515) );
  NAND2_X1 U12276 ( .A1(n12528), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15028) );
  OAI22_X1 U12277 ( .A1(n20532), .A2(n20531), .B1(n20530), .B2(n20588), .ZN(
        n20549) );
  NOR2_X1 U12278 ( .A1(n20704), .A2(n12709), .ZN(n20548) );
  OAI21_X1 U12279 ( .B1(n20594), .B2(n20610), .A(n20593), .ZN(n20612) );
  AND2_X1 U12280 ( .A1(n20517), .A2(n12949), .ZN(n20611) );
  AOI22_X1 U12281 ( .A1(n13681), .A2(n13678), .B1(n13675), .B2(n13674), .ZN(
        n13718) );
  INV_X1 U12282 ( .A(n20678), .ZN(n20686) );
  INV_X1 U12283 ( .A(n20753), .ZN(n13572) );
  INV_X1 U12284 ( .A(n13543), .ZN(n13574) );
  NOR2_X1 U12285 ( .A1(n12760), .A2(n13496), .ZN(n20712) );
  NOR2_X1 U12286 ( .A1(n12758), .A2(n13496), .ZN(n20718) );
  NOR2_X1 U12287 ( .A1(n12757), .A2(n13496), .ZN(n20724) );
  NOR2_X1 U12288 ( .A1(n12974), .A2(n13496), .ZN(n20736) );
  NOR2_X1 U12289 ( .A1(n13100), .A2(n13496), .ZN(n20742) );
  NOR2_X1 U12290 ( .A1(n20704), .A2(n15034), .ZN(n20753) );
  NOR2_X1 U12291 ( .A1(n13183), .A2(n13496), .ZN(n20749) );
  NAND2_X1 U12292 ( .A1(n13491), .A2(n12939), .ZN(n13534) );
  NOR2_X1 U12293 ( .A1(n12696), .A2(n13496), .ZN(n20700) );
  OAI21_X1 U12294 ( .B1(n12714), .B2(n12715), .A(n20705), .ZN(n12921) );
  INV_X1 U12295 ( .A(n13534), .ZN(n13492) );
  NAND2_X1 U12296 ( .A1(n12265), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20293) );
  INV_X1 U12297 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16510) );
  NOR2_X1 U12298 ( .A1(n11867), .A2(n11866), .ZN(n13252) );
  NAND2_X1 U12299 ( .A1(n16555), .A2(n9661), .ZN(n16545) );
  NAND2_X1 U12300 ( .A1(n16545), .A2(n16546), .ZN(n16544) );
  NAND2_X1 U12301 ( .A1(n16580), .A2(n13308), .ZN(n16570) );
  NAND2_X1 U12302 ( .A1(n16570), .A2(n16571), .ZN(n16569) );
  NAND2_X1 U12303 ( .A1(n16604), .A2(n13308), .ZN(n16593) );
  NAND2_X1 U12304 ( .A1(n16593), .A2(n16594), .ZN(n16592) );
  NAND2_X1 U12305 ( .A1(n16514), .A2(n9661), .ZN(n16605) );
  NAND2_X1 U12306 ( .A1(n16605), .A2(n16606), .ZN(n16604) );
  AND2_X1 U12307 ( .A1(n9661), .A2(n10047), .ZN(n15142) );
  NAND2_X1 U12308 ( .A1(n19308), .A2(n19309), .ZN(n10047) );
  OR2_X1 U12309 ( .A1(n15142), .A2(n15496), .ZN(n15144) );
  OR2_X1 U12310 ( .A1(n19272), .A2(n13256), .ZN(n19405) );
  NOR2_X1 U12311 ( .A1(n10035), .A2(n9754), .ZN(n10034) );
  INV_X1 U12312 ( .A(n10036), .ZN(n10035) );
  INV_X1 U12313 ( .A(n19404), .ZN(n19294) );
  NAND2_X1 U12314 ( .A1(n10742), .A2(n10038), .ZN(n10764) );
  INV_X1 U12315 ( .A(n19405), .ZN(n19392) );
  NOR2_X1 U12316 ( .A1(n13308), .A2(n20126), .ZN(n19397) );
  AND2_X1 U12317 ( .A1(n19272), .A2(n13263), .ZN(n19396) );
  AND2_X1 U12318 ( .A1(n11300), .A2(n11299), .ZN(n13297) );
  AND3_X1 U12319 ( .A1(n11280), .A2(n11279), .A3(n11278), .ZN(n12978) );
  AND2_X1 U12320 ( .A1(n11454), .A2(n12368), .ZN(n10233) );
  AND2_X1 U12321 ( .A1(n11153), .A2(n11152), .ZN(n12843) );
  INV_X1 U12322 ( .A(n15281), .ZN(n15298) );
  XNOR2_X1 U12323 ( .A(n9919), .B(n11801), .ZN(n11832) );
  OAI211_X1 U12324 ( .C1(n15236), .C2(n9915), .A(n11777), .B(n9914), .ZN(n9919) );
  AND2_X1 U12325 ( .A1(n19426), .A2(n19543), .ZN(n19422) );
  AND2_X1 U12326 ( .A1(n19426), .A2(n19545), .ZN(n19420) );
  NAND2_X1 U12327 ( .A1(n19463), .A2(n11822), .ZN(n19427) );
  AND2_X1 U12328 ( .A1(n12829), .A2(n11457), .ZN(n13396) );
  NAND2_X1 U12329 ( .A1(n11810), .A2(n11809), .ZN(n19463) );
  INV_X1 U12330 ( .A(n20256), .ZN(n19827) );
  INV_X1 U12331 ( .A(n15314), .ZN(n19486) );
  AND2_X1 U12332 ( .A1(n11368), .A2(n10885), .ZN(n10166) );
  AND2_X1 U12333 ( .A1(n10140), .A2(n9691), .ZN(n16628) );
  INV_X1 U12334 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16656) );
  INV_X1 U12335 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16667) );
  INV_X1 U12336 ( .A(n16658), .ZN(n19542) );
  NAND2_X1 U12337 ( .A1(n19275), .A2(n10980), .ZN(n16666) );
  AND2_X1 U12338 ( .A1(n16666), .A2(n12040), .ZN(n16658) );
  INV_X1 U12339 ( .A(n16666), .ZN(n19530) );
  INV_X1 U12340 ( .A(n19538), .ZN(n16648) );
  INV_X1 U12341 ( .A(n11418), .ZN(n10117) );
  NAND2_X1 U12342 ( .A1(n16525), .A2(n16689), .ZN(n10016) );
  NAND2_X1 U12343 ( .A1(n10252), .A2(n10824), .ZN(n15389) );
  NAND2_X1 U12344 ( .A1(n10141), .A2(n10147), .ZN(n15412) );
  NAND2_X1 U12345 ( .A1(n9909), .A2(n15441), .ZN(n15434) );
  NOR2_X1 U12346 ( .A1(n10153), .A2(n10154), .ZN(n15445) );
  NOR2_X1 U12347 ( .A1(n10058), .A2(n10061), .ZN(n15190) );
  NAND2_X1 U12348 ( .A1(n10140), .A2(n10138), .ZN(n15582) );
  INV_X1 U12349 ( .A(n10728), .ZN(n10137) );
  NAND2_X1 U12350 ( .A1(n15841), .A2(n10880), .ZN(n15592) );
  NOR3_X1 U12351 ( .A1(n13422), .A2(n13455), .A3(n13423), .ZN(n15847) );
  NOR2_X1 U12352 ( .A1(n13446), .A2(n9763), .ZN(n13447) );
  NAND2_X1 U12353 ( .A1(n13425), .A2(n13424), .ZN(n13283) );
  NAND2_X1 U12354 ( .A1(n9879), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13141) );
  NAND2_X1 U12355 ( .A1(n9876), .A2(n11372), .ZN(n13142) );
  NAND2_X1 U12356 ( .A1(n12110), .A2(n15743), .ZN(n16705) );
  INV_X1 U12357 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20263) );
  INV_X1 U12358 ( .A(n20227), .ZN(n20248) );
  INV_X1 U12359 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20243) );
  INV_X1 U12360 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16209) );
  AND2_X1 U12361 ( .A1(n12103), .A2(n12102), .ZN(n20227) );
  OR2_X1 U12362 ( .A1(n12101), .A2(n12100), .ZN(n12103) );
  NAND2_X1 U12363 ( .A1(n12133), .A2(n12136), .ZN(n20239) );
  AOI21_X1 U12364 ( .B1(n11439), .B2(n15912), .A(n15911), .ZN(n16740) );
  NAND2_X1 U12365 ( .A1(n16721), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16761) );
  NAND2_X1 U12366 ( .A1(n12398), .A2(n12401), .ZN(n19860) );
  INV_X1 U12367 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20221) );
  OR2_X1 U12368 ( .A1(n19655), .A2(n19775), .ZN(n19673) );
  OAI21_X1 U12369 ( .B1(n19717), .B2(n19713), .A(n19712), .ZN(n19736) );
  INV_X1 U12370 ( .A(n19766), .ZN(n19758) );
  NAND2_X1 U12371 ( .A1(n19767), .A2(n19984), .ZN(n19766) );
  OR3_X1 U12372 ( .A1(n19776), .A2(n19775), .A3(n19774), .ZN(n19794) );
  OAI21_X1 U12373 ( .B1(n19898), .B2(n19913), .A(n20067), .ZN(n19916) );
  NOR2_X2 U12374 ( .A1(n19991), .A2(n19861), .ZN(n19915) );
  INV_X1 U12375 ( .A(n19953), .ZN(n19977) );
  NAND2_X1 U12376 ( .A1(n20019), .A2(n19984), .ZN(n20018) );
  OAI22_X1 U12377 ( .A1(n14691), .A2(n19584), .B1(n15339), .B2(n19585), .ZN(
        n20032) );
  OAI21_X1 U12378 ( .B1(n20029), .B2(n20028), .A(n20027), .ZN(n20052) );
  NOR2_X2 U12379 ( .A1(n19991), .A2(n19990), .ZN(n20051) );
  OAI22_X1 U12380 ( .A1(n14697), .A2(n19584), .B1(n15349), .B2(n19585), .ZN(
        n20069) );
  OAI22_X1 U12381 ( .A1(n14721), .A2(n19584), .B1(n19563), .B2(n19585), .ZN(
        n20081) );
  AND2_X1 U12382 ( .A1(n19569), .A2(n19568), .ZN(n20085) );
  INV_X1 U12383 ( .A(n20120), .ZN(n20106) );
  INV_X1 U12384 ( .A(n20013), .ZN(n20105) );
  AND2_X1 U12385 ( .A1(n13254), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20122) );
  NAND2_X1 U12386 ( .A1(n19090), .A2(n19041), .ZN(n17825) );
  XOR2_X1 U12387 ( .A(n18613), .B(n18609), .Z(n19265) );
  INV_X1 U12388 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19261) );
  NOR2_X1 U12389 ( .A1(n19040), .A2(n17825), .ZN(n19264) );
  AOI21_X1 U12390 ( .B1(n17025), .B2(n9970), .A(n17261), .ZN(n17009) );
  NOR2_X1 U12391 ( .A1(n17017), .A2(n17919), .ZN(n17016) );
  NOR2_X1 U12392 ( .A1(n17025), .A2(n17261), .ZN(n17017) );
  NOR2_X1 U12393 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17040), .ZN(n17024) );
  NOR2_X1 U12394 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17060), .ZN(n17045) );
  NOR2_X1 U12395 ( .A1(n16983), .A2(n17081), .ZN(n17054) );
  NOR2_X1 U12396 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17078), .ZN(n17065) );
  AND2_X1 U12397 ( .A1(n17292), .A2(n9745), .ZN(n17083) );
  NOR2_X1 U12398 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17117), .ZN(n17104) );
  NOR2_X2 U12399 ( .A1(n19092), .A2(n16966), .ZN(n17310) );
  CLKBUF_X1 U12400 ( .A(n17305), .Z(n17267) );
  NOR2_X1 U12401 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17272), .ZN(n17252) );
  INV_X1 U12402 ( .A(n17305), .ZN(n17322) );
  NAND2_X1 U12403 ( .A1(n17400), .A2(n9713), .ZN(n17385) );
  NAND2_X1 U12404 ( .A1(n17385), .A2(n17619), .ZN(n17383) );
  NOR2_X1 U12405 ( .A1(n17343), .A2(n17395), .ZN(n17400) );
  AND3_X1 U12406 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17453), .ZN(n17426) );
  AND2_X1 U12407 ( .A1(n18639), .A2(n17342), .ZN(n17453) );
  NOR2_X1 U12408 ( .A1(n17168), .A2(n17521), .ZN(n17509) );
  NAND2_X1 U12409 ( .A1(n17509), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n17508) );
  NAND2_X1 U12410 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17536), .ZN(n17521) );
  NOR2_X1 U12411 ( .A1(n17194), .A2(n17550), .ZN(n17536) );
  NAND2_X1 U12412 ( .A1(n17570), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17550) );
  NOR2_X1 U12413 ( .A1(n17591), .A2(n17220), .ZN(n17570) );
  NAND2_X1 U12414 ( .A1(n17593), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17591) );
  NOR3_X1 U12415 ( .A1(n17599), .A2(n20911), .A3(n17602), .ZN(n17593) );
  AND2_X1 U12416 ( .A1(n17621), .A2(n9859), .ZN(n17603) );
  NOR2_X1 U12417 ( .A1(n17594), .A2(n13984), .ZN(n9859) );
  INV_X2 U12418 ( .A(n17625), .ZN(n17619) );
  INV_X1 U12419 ( .A(n17640), .ZN(n17635) );
  NOR2_X1 U12420 ( .A1(n17852), .A2(n17651), .ZN(n17644) );
  NOR2_X1 U12421 ( .A1(n17848), .A2(n17660), .ZN(n17655) );
  INV_X1 U12422 ( .A(n17665), .ZN(n17661) );
  NOR2_X1 U12423 ( .A1(n17717), .A2(n17670), .ZN(n17666) );
  NOR4_X1 U12424 ( .A1(n20871), .A2(n17710), .A3(n17840), .A4(n17630), .ZN(
        n17671) );
  NOR2_X1 U12425 ( .A1(n17894), .A2(n17723), .ZN(n17711) );
  NAND2_X1 U12426 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17711), .ZN(n17710) );
  INV_X1 U12427 ( .A(n17707), .ZN(n17709) );
  INV_X1 U12428 ( .A(n16096), .ZN(n17755) );
  NOR2_X1 U12429 ( .A1(n15990), .A2(n15989), .ZN(n17758) );
  NOR2_X1 U12430 ( .A1(n16028), .A2(n16027), .ZN(n17765) );
  INV_X1 U12431 ( .A(n16078), .ZN(n17770) );
  NAND2_X1 U12432 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n9948) );
  NOR2_X1 U12433 ( .A1(n15998), .A2(n9945), .ZN(n9946) );
  AND3_X1 U12434 ( .A1(n15996), .A2(n15995), .A3(n9949), .ZN(n9947) );
  OR3_X1 U12435 ( .A1(n16210), .A2(n17786), .A3(n19246), .ZN(n16211) );
  INV_X1 U12436 ( .A(n9861), .ZN(n16210) );
  INV_X1 U12437 ( .A(n17771), .ZN(n17776) );
  NOR2_X1 U12438 ( .A1(n18613), .A2(n17890), .ZN(n17883) );
  INV_X1 U12439 ( .A(n17865), .ZN(n17890) );
  NAND2_X1 U12441 ( .A1(n17928), .A2(n9707), .ZN(n16813) );
  AND2_X1 U12442 ( .A1(n17162), .A2(n9964), .ZN(n18011) );
  AND2_X1 U12443 ( .A1(n9702), .A2(n9965), .ZN(n9964) );
  INV_X1 U12444 ( .A(n18019), .ZN(n9965) );
  NAND2_X1 U12445 ( .A1(n16786), .A2(n18255), .ZN(n18170) );
  NAND2_X1 U12446 ( .A1(n18203), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18192) );
  NOR2_X1 U12447 ( .A1(n18209), .A2(n18221), .ZN(n18203) );
  OAI21_X1 U12448 ( .B1(n18600), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n16946), 
        .ZN(n18242) );
  NAND2_X1 U12449 ( .A1(n18947), .A2(n18662), .ZN(n18843) );
  INV_X1 U12450 ( .A(n18254), .ZN(n18238) );
  NOR2_X1 U12451 ( .A1(n17932), .A2(n18093), .ZN(n18250) );
  INV_X1 U12452 ( .A(n18242), .ZN(n18251) );
  AND3_X1 U12453 ( .A1(n9960), .A2(n9958), .A3(n9955), .ZN(n16187) );
  INV_X1 U12454 ( .A(n10240), .ZN(n9955) );
  NOR2_X1 U12456 ( .A1(n10078), .A2(n16127), .ZN(n18042) );
  INV_X1 U12457 ( .A(n18480), .ZN(n18504) );
  NAND2_X1 U12458 ( .A1(n18476), .A2(n18498), .ZN(n18575) );
  INV_X1 U12459 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18514) );
  INV_X1 U12460 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18518) );
  INV_X1 U12461 ( .A(n16093), .ZN(n10096) );
  NAND2_X1 U12462 ( .A1(n10090), .A2(n10088), .ZN(n18215) );
  AOI21_X2 U12463 ( .B1(n16117), .B2(n16116), .A(n19254), .ZN(n18586) );
  AOI211_X1 U12464 ( .C1(n16113), .C2(n19042), .A(n16112), .B(n16111), .ZN(
        n16117) );
  INV_X1 U12465 ( .A(n18575), .ZN(n18584) );
  INV_X1 U12466 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19079) );
  INV_X1 U12467 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19082) );
  INV_X1 U12468 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21004) );
  INV_X1 U12469 ( .A(n17239), .ZN(n19105) );
  AND2_X2 U12470 ( .A1(n11849), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14482)
         );
  CLKBUF_X1 U12471 ( .A(n16928), .Z(n16932) );
  OAI211_X1 U12472 ( .C1(n14938), .C2(n20299), .A(n9845), .B(n9843), .ZN(
        P1_U2971) );
  AOI21_X1 U12473 ( .B1(n14776), .B2(n16365), .A(n14775), .ZN(n9845) );
  INV_X1 U12474 ( .A(n9925), .ZN(n12832) );
  AOI21_X1 U12475 ( .B1(n16525), .B2(n19538), .A(n11027), .ZN(n11028) );
  INV_X1 U12476 ( .A(n11391), .ZN(n11392) );
  INV_X1 U12477 ( .A(n10987), .ZN(n10988) );
  INV_X1 U12478 ( .A(n11383), .ZN(n10111) );
  INV_X1 U12479 ( .A(n10109), .ZN(n10108) );
  OAI21_X1 U12480 ( .B1(n16541), .B2(n16701), .A(n10075), .ZN(n15613) );
  AOI21_X1 U12481 ( .B1(n15610), .B2(n16689), .A(n10076), .ZN(n10075) );
  INV_X1 U12482 ( .A(n11405), .ZN(n11406) );
  OAI21_X1 U12483 ( .B1(n11404), .B2(n16710), .A(n11403), .ZN(n11405) );
  OAI21_X1 U12484 ( .B1(n16989), .B2(n9731), .A(n9976), .ZN(P3_U2641) );
  NOR2_X1 U12485 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  INV_X1 U12486 ( .A(n17621), .ZN(n17624) );
  CLKBUF_X3 U12487 ( .A(n13986), .Z(n17581) );
  NAND2_X1 U12488 ( .A1(n10886), .A2(n9710), .ZN(n15430) );
  AND2_X2 U12489 ( .A1(n10568), .A2(n10567), .ZN(n10717) );
  AND2_X1 U12490 ( .A1(n9711), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9687) );
  INV_X1 U12491 ( .A(n11097), .ZN(n11335) );
  CLKBUF_X3 U12492 ( .A(n13964), .Z(n17539) );
  AND2_X1 U12493 ( .A1(n9959), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9958) );
  NAND2_X1 U12494 ( .A1(n16269), .A2(n9757), .ZN(n14613) );
  NAND2_X1 U12495 ( .A1(n9940), .A2(n12271), .ZN(n12233) );
  NAND2_X1 U12496 ( .A1(n16269), .A2(n9761), .ZN(n9688) );
  NAND2_X1 U12497 ( .A1(n9691), .A2(n16626), .ZN(n10136) );
  INV_X1 U12498 ( .A(n11032), .ZN(n10126) );
  AND2_X1 U12499 ( .A1(n10050), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9689) );
  AND2_X1 U12500 ( .A1(n10045), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9690) );
  AND2_X1 U12501 ( .A1(n10138), .A2(n9776), .ZN(n9691) );
  AND2_X1 U12502 ( .A1(n14816), .A2(n14980), .ZN(n9692) );
  NAND2_X1 U12503 ( .A1(n13388), .A2(n10187), .ZN(n13750) );
  NAND2_X1 U12504 ( .A1(n10886), .A2(n9687), .ZN(n15418) );
  AND2_X1 U12505 ( .A1(n9892), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n9693)
         );
  AND2_X1 U12506 ( .A1(n9934), .A2(n9716), .ZN(n9694) );
  NAND2_X1 U12507 ( .A1(n16269), .A2(n9852), .ZN(n9854) );
  AND2_X1 U12508 ( .A1(n9741), .A2(n10016), .ZN(n9695) );
  AND2_X1 U12509 ( .A1(n11959), .A2(n12059), .ZN(n9696) );
  AND2_X1 U12510 ( .A1(n9897), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9697) );
  AND2_X1 U12511 ( .A1(n9692), .A2(n9930), .ZN(n9698) );
  INV_X1 U12512 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10162) );
  AND2_X1 U12513 ( .A1(n9918), .A2(n15232), .ZN(n9699) );
  OR2_X1 U12514 ( .A1(n10099), .A2(n18182), .ZN(n9700) );
  AND2_X1 U12515 ( .A1(n10235), .A2(n10234), .ZN(n9701) );
  AND2_X1 U12516 ( .A1(n9966), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9702) );
  OR2_X1 U12517 ( .A1(n11732), .A2(n11428), .ZN(n11436) );
  INV_X1 U12518 ( .A(n11436), .ZN(n10221) );
  NAND2_X1 U12519 ( .A1(n15284), .A2(n10228), .ZN(n10232) );
  AND2_X1 U12520 ( .A1(n10041), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9703) );
  AND2_X1 U12521 ( .A1(n10000), .A2(n9999), .ZN(n9704) );
  NOR2_X1 U12522 ( .A1(n13279), .A2(n9780), .ZN(n9705) );
  AND2_X1 U12523 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9706) );
  AND2_X1 U12524 ( .A1(n9973), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9707) );
  AND2_X1 U12525 ( .A1(n9706), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9708) );
  AND2_X1 U12526 ( .A1(n9708), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9709) );
  AND2_X1 U12527 ( .A1(n10170), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9710) );
  AND2_X1 U12528 ( .A1(n9710), .A2(n15654), .ZN(n9711) );
  AND2_X1 U12529 ( .A1(n9857), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n9712) );
  AND2_X1 U12530 ( .A1(n9855), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n9713) );
  OR2_X1 U12531 ( .A1(n13880), .A2(n19061), .ZN(n9714) );
  NOR2_X1 U12532 ( .A1(n17321), .A2(n13880), .ZN(n13891) );
  INV_X1 U12533 ( .A(n11464), .ZN(n11478) );
  NAND2_X1 U12534 ( .A1(n15550), .A2(n11368), .ZN(n15510) );
  NAND2_X1 U12535 ( .A1(n15876), .A2(n11587), .ZN(n9715) );
  NOR2_X1 U12536 ( .A1(n13880), .A2(n13881), .ZN(n13896) );
  OR2_X1 U12537 ( .A1(n14877), .A2(n14425), .ZN(n9716) );
  NAND2_X1 U12538 ( .A1(n9900), .A2(n9904), .ZN(n10147) );
  OAI21_X1 U12539 ( .B1(n10201), .B2(n9932), .A(n9931), .ZN(n14823) );
  NAND2_X1 U12540 ( .A1(n19590), .A2(n20268), .ZN(n9717) );
  INV_X1 U12541 ( .A(n12493), .ZN(n9938) );
  OR2_X1 U12542 ( .A1(n9961), .A2(n17926), .ZN(n9960) );
  NAND2_X1 U12543 ( .A1(n11587), .A2(n15883), .ZN(n9718) );
  OR2_X1 U12544 ( .A1(n14521), .A2(n10175), .ZN(n9719) );
  NAND2_X2 U12545 ( .A1(n16840), .A2(n16786), .ZN(n18168) );
  AND2_X1 U12546 ( .A1(n9888), .A2(n9885), .ZN(n15594) );
  NAND2_X1 U12547 ( .A1(n15840), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15841) );
  NAND2_X1 U12548 ( .A1(n10140), .A2(n10135), .ZN(n15451) );
  NAND2_X1 U12549 ( .A1(n10813), .A2(n10718), .ZN(n10731) );
  INV_X1 U12550 ( .A(n11736), .ZN(n15231) );
  AND2_X1 U12551 ( .A1(n9913), .A2(n9912), .ZN(n11736) );
  NAND2_X1 U12552 ( .A1(n9918), .A2(n9916), .ZN(n15227) );
  XOR2_X1 U12553 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14750), .Z(
        n9721) );
  NAND2_X1 U12554 ( .A1(n12180), .A2(n12268), .ZN(n12334) );
  INV_X1 U12555 ( .A(n11352), .ZN(n11069) );
  AND2_X1 U12556 ( .A1(n9908), .A2(n15441), .ZN(n9722) );
  AND2_X1 U12557 ( .A1(n10448), .A2(n10436), .ZN(n15857) );
  OR3_X1 U12558 ( .A1(n11417), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11416), .ZN(n9723) );
  AND2_X1 U12559 ( .A1(n16269), .A2(n10179), .ZN(n14618) );
  OR2_X1 U12560 ( .A1(n18182), .A2(n16099), .ZN(n9724) );
  OR2_X1 U12561 ( .A1(n12210), .A2(n12209), .ZN(n12617) );
  AND4_X1 U12562 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n9725) );
  AND2_X1 U12563 ( .A1(n15117), .A2(n10113), .ZN(n9726) );
  AND2_X1 U12564 ( .A1(n10874), .A2(n10710), .ZN(n10868) );
  NAND2_X1 U12565 ( .A1(n14880), .A2(n14426), .ZN(n14837) );
  NAND2_X1 U12566 ( .A1(n10886), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15483) );
  INV_X1 U12567 ( .A(n19955), .ZN(n10636) );
  AND2_X1 U12568 ( .A1(n15284), .A2(n10229), .ZN(n9727) );
  AND2_X1 U12569 ( .A1(n10886), .A2(n9711), .ZN(n15421) );
  AND3_X1 U12570 ( .A1(n16017), .A2(n16011), .A3(n16012), .ZN(n9728) );
  AND2_X1 U12572 ( .A1(n12493), .A2(n16503), .ZN(n9729) );
  NAND2_X1 U12573 ( .A1(n12196), .A2(n12197), .ZN(n12271) );
  OR2_X1 U12574 ( .A1(n18518), .A2(n16094), .ZN(n9730) );
  AND2_X1 U12575 ( .A1(n16990), .A2(n16991), .ZN(n9731) );
  AND2_X1 U12576 ( .A1(n12272), .A2(n9842), .ZN(n9732) );
  AND3_X1 U12577 ( .A1(n11917), .A2(n11914), .A3(n11915), .ZN(n9733) );
  AND3_X1 U12578 ( .A1(n19564), .A2(n19569), .A3(n11352), .ZN(n10384) );
  INV_X1 U12579 ( .A(n11981), .ZN(n12049) );
  BUF_X1 U12580 ( .A(n11981), .Z(n12910) );
  AOI21_X1 U12581 ( .B1(n10433), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10416), .ZN(n10421) );
  INV_X1 U12582 ( .A(n10155), .ZN(n10154) );
  NOR2_X1 U12583 ( .A1(n10156), .A2(n15466), .ZN(n10155) );
  AND2_X1 U12584 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9734) );
  NAND2_X1 U12585 ( .A1(n14832), .A2(n14426), .ZN(n9735) );
  NAND2_X1 U12586 ( .A1(n16269), .A2(n16268), .ZN(n14642) );
  OR2_X1 U12587 ( .A1(n14454), .A2(n9997), .ZN(n9736) );
  NAND3_X1 U12588 ( .A1(n10510), .A2(n10509), .A3(n10508), .ZN(n9737) );
  AND2_X1 U12589 ( .A1(n13720), .A2(n16468), .ZN(n9738) );
  INV_X1 U12590 ( .A(n10826), .ZN(n9896) );
  INV_X1 U12591 ( .A(n9929), .ZN(n12184) );
  NAND2_X1 U12592 ( .A1(n12054), .A2(n12910), .ZN(n9929) );
  NOR2_X1 U12593 ( .A1(n18216), .A2(n18549), .ZN(n9739) );
  INV_X1 U12594 ( .A(n10729), .ZN(n9887) );
  AND2_X1 U12595 ( .A1(n9934), .A2(n9735), .ZN(n9740) );
  AND2_X1 U12596 ( .A1(n16269), .A2(n10180), .ZN(n14628) );
  NOR2_X1 U12597 ( .A1(n12005), .A2(n11997), .ZN(n12014) );
  INV_X1 U12598 ( .A(n12014), .ZN(n9837) );
  AND2_X1 U12599 ( .A1(n10886), .A2(n10014), .ZN(n15401) );
  AND2_X1 U12600 ( .A1(n10117), .A2(n9723), .ZN(n9741) );
  AND2_X1 U12601 ( .A1(n9884), .A2(n9882), .ZN(n9742) );
  INV_X1 U12602 ( .A(n10802), .ZN(n9908) );
  OR2_X1 U12603 ( .A1(n18524), .A2(n16089), .ZN(n9743) );
  AND3_X1 U12604 ( .A1(n9794), .A2(n9793), .A3(n9792), .ZN(n9744) );
  OR2_X1 U12605 ( .A1(n17984), .A2(n17133), .ZN(n9745) );
  AND2_X1 U12606 ( .A1(n10147), .A2(n10146), .ZN(n9746) );
  NOR2_X1 U12607 ( .A1(n15390), .A2(n10168), .ZN(n15379) );
  INV_X1 U12608 ( .A(n10136), .ZN(n10135) );
  AND2_X1 U12609 ( .A1(n10140), .A2(n10137), .ZN(n9747) );
  NAND2_X1 U12610 ( .A1(n14777), .A2(n9692), .ZN(n9748) );
  OR2_X1 U12611 ( .A1(n12562), .A2(n12649), .ZN(n9925) );
  NOR2_X1 U12612 ( .A1(n9925), .A2(n9924), .ZN(n12829) );
  AND2_X1 U12613 ( .A1(n17509), .A2(n9857), .ZN(n9749) );
  AND2_X1 U12614 ( .A1(n12369), .A2(n12368), .ZN(n12367) );
  AND2_X1 U12615 ( .A1(n12895), .A2(n12894), .ZN(n9750) );
  NOR2_X1 U12616 ( .A1(n13350), .A2(n13351), .ZN(n13388) );
  NAND2_X1 U12617 ( .A1(n12829), .A2(n10237), .ZN(n13394) );
  AND2_X1 U12618 ( .A1(n11804), .A2(n10365), .ZN(n11364) );
  AND2_X1 U12619 ( .A1(n17400), .A2(n9855), .ZN(n9751) );
  AND2_X1 U12620 ( .A1(n17400), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n9752) );
  OR2_X1 U12621 ( .A1(n10061), .A2(n10060), .ZN(n9753) );
  AND2_X1 U12622 ( .A1(n11007), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n9754) );
  AND2_X1 U12623 ( .A1(n10066), .A2(n10254), .ZN(n9755) );
  AND2_X1 U12624 ( .A1(n13388), .A2(n13389), .ZN(n9756) );
  NAND2_X1 U12625 ( .A1(n13822), .A2(n9848), .ZN(n14099) );
  OAI22_X1 U12626 ( .A1(n13419), .A2(n13420), .B1(n19375), .B2(n13422), .ZN(
        n13449) );
  AND2_X1 U12627 ( .A1(n10179), .A2(n14230), .ZN(n9757) );
  AND2_X1 U12628 ( .A1(n13822), .A2(n13800), .ZN(n13862) );
  AND2_X1 U12629 ( .A1(n14638), .A2(n9704), .ZN(n9758) );
  NOR2_X1 U12630 ( .A1(n10032), .A2(n10659), .ZN(n10712) );
  INV_X1 U12631 ( .A(n14474), .ZN(n9820) );
  AND2_X1 U12632 ( .A1(n11284), .A2(n9755), .ZN(n9759) );
  OR3_X1 U12633 ( .A1(n13869), .A2(n10004), .A3(n10008), .ZN(n9760) );
  NOR2_X1 U12634 ( .A1(n14643), .A2(n10181), .ZN(n9761) );
  OR2_X1 U12635 ( .A1(n18168), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9762) );
  NOR2_X1 U12636 ( .A1(n13869), .A2(n10002), .ZN(n10007) );
  AND2_X1 U12637 ( .A1(n10867), .A2(n13455), .ZN(n9763) );
  INV_X1 U12638 ( .A(n15781), .ZN(n11284) );
  INV_X1 U12639 ( .A(n18182), .ZN(n10098) );
  AND2_X1 U12640 ( .A1(n13324), .A2(n13323), .ZN(n13325) );
  INV_X1 U12641 ( .A(n13325), .ZN(n10061) );
  OR2_X1 U12642 ( .A1(n9921), .A2(n12649), .ZN(n9764) );
  NOR2_X1 U12643 ( .A1(n14658), .A2(n14659), .ZN(n14651) );
  INV_X1 U12644 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n19328) );
  INV_X1 U12645 ( .A(n10232), .ZN(n15275) );
  INV_X1 U12646 ( .A(n10005), .ZN(n10004) );
  NOR2_X1 U12647 ( .A1(n13868), .A2(n10006), .ZN(n10005) );
  INV_X1 U12648 ( .A(n10220), .ZN(n10219) );
  NAND2_X1 U12649 ( .A1(n10221), .A2(n11427), .ZN(n10220) );
  OAI22_X1 U12650 ( .A1(n14801), .A2(n14351), .B1(n14269), .B2(n14268), .ZN(
        n14548) );
  AND2_X1 U12651 ( .A1(n10229), .A2(n10227), .ZN(n9765) );
  AND2_X1 U12652 ( .A1(n10206), .A2(n14931), .ZN(n9766) );
  NAND2_X1 U12653 ( .A1(n12787), .A2(n14478), .ZN(n9822) );
  AND2_X1 U12654 ( .A1(n9851), .A2(n9852), .ZN(n9767) );
  INV_X1 U12655 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16645) );
  INV_X1 U12656 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15538) );
  INV_X1 U12657 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n16503) );
  INV_X1 U12658 ( .A(n12477), .ZN(n14351) );
  NOR2_X1 U12659 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12477) );
  NAND2_X1 U12660 ( .A1(n9817), .A2(n9988), .ZN(n12280) );
  AND2_X1 U12661 ( .A1(n15391), .A2(n9708), .ZN(n9768) );
  NOR2_X1 U12662 ( .A1(n13305), .A2(n13306), .ZN(n13304) );
  AND2_X1 U12663 ( .A1(n17928), .A2(n9973), .ZN(n9769) );
  NAND2_X1 U12664 ( .A1(n12031), .A2(n12392), .ZN(n20855) );
  AND2_X1 U12665 ( .A1(n10069), .A2(n10068), .ZN(n9770) );
  AND2_X1 U12666 ( .A1(n15092), .A2(n10041), .ZN(n9771) );
  AND2_X1 U12667 ( .A1(n15092), .A2(n9703), .ZN(n9772) );
  INV_X1 U12668 ( .A(n11439), .ZN(n9891) );
  OR2_X1 U12669 ( .A1(n20442), .A2(n9842), .ZN(n9773) );
  AND2_X1 U12670 ( .A1(n11734), .A2(n10211), .ZN(n9774) );
  AND2_X1 U12671 ( .A1(n11734), .A2(n15245), .ZN(n9775) );
  OR2_X1 U12672 ( .A1(n10739), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9776) );
  OR2_X1 U12673 ( .A1(n16137), .A2(n18260), .ZN(n9777) );
  INV_X1 U12674 ( .A(n9993), .ZN(n13834) );
  NOR2_X1 U12675 ( .A1(n13488), .A2(n13489), .ZN(n9993) );
  AND2_X1 U12676 ( .A1(n12369), .A2(n10233), .ZN(n9778) );
  AND2_X1 U12677 ( .A1(n16503), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9779) );
  INV_X1 U12678 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17329) );
  AND2_X1 U12679 ( .A1(n11439), .A2(n19396), .ZN(n9780) );
  AND2_X1 U12680 ( .A1(n9770), .A2(n10067), .ZN(n9781) );
  AND2_X1 U12681 ( .A1(n10097), .A2(n10096), .ZN(n9782) );
  AND2_X2 U12682 ( .A1(n20622), .A2(n12314), .ZN(n16482) );
  INV_X1 U12683 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n9985) );
  INV_X1 U12684 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9991) );
  INV_X1 U12685 ( .A(n12831), .ZN(n9924) );
  NAND3_X1 U12686 ( .A1(n14431), .A2(n14381), .A3(n16413), .ZN(n9783) );
  INV_X1 U12687 ( .A(n9821), .ZN(n12315) );
  NAND2_X1 U12688 ( .A1(n9818), .A2(n12787), .ZN(n9821) );
  AND2_X1 U12689 ( .A1(n10092), .A2(n10091), .ZN(n9784) );
  INV_X1 U12690 ( .A(n13914), .ZN(n14037) );
  INV_X1 U12691 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10046) );
  AND2_X1 U12692 ( .A1(n17162), .A2(n9966), .ZN(n9785) );
  INV_X1 U12693 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9975) );
  AND2_X1 U12694 ( .A1(n20278), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11440) );
  INV_X1 U12695 ( .A(n11440), .ZN(n10216) );
  AND2_X1 U12696 ( .A1(n14991), .A2(n16180), .ZN(n9786) );
  INV_X1 U12697 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10017) );
  AND2_X1 U12698 ( .A1(n9786), .A2(n10205), .ZN(n9787) );
  INV_X1 U12699 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9957) );
  INV_X1 U12700 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9967) );
  INV_X1 U12701 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9963) );
  INV_X1 U12702 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10043) );
  INV_X1 U12703 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10042) );
  INV_X1 U12704 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n9997) );
  AOI22_X2 U12705 ( .A1(DATAI_19_), .A2(n9650), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9656), .ZN(n20729) );
  AOI22_X2 U12706 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9656), .B1(DATAI_23_), 
        .B2(n9650), .ZN(n20758) );
  AOI22_X2 U12707 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9656), .B1(DATAI_18_), 
        .B2(n9650), .ZN(n20723) );
  AOI22_X2 U12708 ( .A1(DATAI_16_), .A2(n9650), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n9656), .ZN(n20711) );
  AOI22_X2 U12709 ( .A1(DATAI_17_), .A2(n9650), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n9656), .ZN(n20717) );
  AOI22_X2 U12710 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n9656), .B1(DATAI_22_), 
        .B2(n9650), .ZN(n20747) );
  AOI22_X2 U12711 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9656), .B1(DATAI_20_), 
        .B2(n9650), .ZN(n20735) );
  AOI22_X2 U12712 ( .A1(DATAI_21_), .A2(n9650), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n9656), .ZN(n20741) );
  AND2_X1 U12713 ( .A1(n12463), .A2(n16755), .ZN(n19377) );
  AND2_X2 U12714 ( .A1(n13252), .A2(n9659), .ZN(n12463) );
  NAND3_X1 U12715 ( .A1(n10865), .A2(n9791), .A3(n13416), .ZN(n9790) );
  INV_X2 U12716 ( .A(n10265), .ZN(n11781) );
  NAND2_X2 U12717 ( .A1(n15883), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10265) );
  NAND2_X1 U12719 ( .A1(n9796), .A2(n10896), .ZN(n10901) );
  XNOR2_X2 U12720 ( .A(n9796), .B(n10896), .ZN(n10451) );
  NAND3_X1 U12721 ( .A1(n14439), .A2(n9766), .A3(n14789), .ZN(n14758) );
  INV_X4 U12722 ( .A(n10849), .ZN(n20281) );
  NAND4_X1 U12723 ( .A1(n9798), .A2(n10347), .A3(n10346), .A4(n10349), .ZN(
        n9797) );
  NAND4_X1 U12724 ( .A1(n10354), .A2(n9801), .A3(n10352), .A4(n10353), .ZN(
        n9800) );
  NAND2_X1 U12725 ( .A1(n13611), .A2(n9814), .ZN(n9813) );
  INV_X1 U12726 ( .A(n13611), .ZN(n9815) );
  NAND2_X1 U12727 ( .A1(n13612), .A2(n13611), .ZN(n20453) );
  NAND2_X1 U12728 ( .A1(n12995), .A2(n12994), .ZN(n13612) );
  XNOR2_X1 U12729 ( .A(n13610), .B(n12987), .ZN(n12995) );
  NAND3_X1 U12730 ( .A1(n9816), .A2(n9821), .A3(n12172), .ZN(n12174) );
  NAND3_X1 U12731 ( .A1(n11945), .A2(n11946), .A3(n11959), .ZN(n12058) );
  NAND3_X1 U12732 ( .A1(n9824), .A2(n12657), .A3(n16503), .ZN(n9823) );
  NAND2_X2 U12733 ( .A1(n11342), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10902) );
  NAND2_X2 U12734 ( .A1(n9827), .A2(n15886), .ZN(n11342) );
  NAND2_X1 U12735 ( .A1(n10390), .A2(n9659), .ZN(n9827) );
  INV_X2 U12736 ( .A(n15506), .ZN(n10886) );
  NAND2_X2 U12737 ( .A1(n14817), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14777) );
  OAI21_X2 U12738 ( .B1(n14823), .B2(n9989), .A(n14877), .ZN(n14817) );
  NAND3_X1 U12739 ( .A1(n9839), .A2(n9838), .A3(n9835), .ZN(n9834) );
  NOR2_X2 U12740 ( .A1(n13063), .A2(n20785), .ZN(n20381) );
  AND2_X2 U12741 ( .A1(n9840), .A2(n12028), .ZN(n12528) );
  OR2_X4 U12742 ( .A1(n11995), .A2(n11994), .ZN(n9842) );
  NAND2_X1 U12743 ( .A1(n9842), .A2(n12539), .ZN(n13651) );
  OAI21_X1 U12744 ( .B1(n9842), .B2(n16165), .A(n20857), .ZN(n13018) );
  AOI21_X1 U12745 ( .B1(n9842), .B2(n16195), .A(n20773), .ZN(n12298) );
  NAND2_X1 U12746 ( .A1(n13019), .A2(n9842), .ZN(n13184) );
  NAND2_X1 U12747 ( .A1(n13024), .A2(n9842), .ZN(n13016) );
  NAND2_X1 U12748 ( .A1(n14091), .A2(n9842), .ZN(n12305) );
  OAI22_X1 U12749 ( .A1(n12392), .A2(n9842), .B1(n12804), .B2(n12139), .ZN(
        n12140) );
  INV_X1 U12750 ( .A(n9854), .ZN(n14547) );
  NAND3_X1 U12751 ( .A1(n10436), .A2(n10422), .A3(n10424), .ZN(n9862) );
  INV_X1 U12752 ( .A(n10451), .ZN(n10468) );
  AND2_X2 U12753 ( .A1(n9865), .A2(n10552), .ZN(n10616) );
  NAND3_X1 U12754 ( .A1(n10537), .A2(n10539), .A3(n10538), .ZN(n9865) );
  AND2_X2 U12755 ( .A1(n9867), .A2(n10522), .ZN(n10617) );
  NAND3_X1 U12756 ( .A1(n10009), .A2(n10010), .A3(n9868), .ZN(n9867) );
  AOI22_X1 U12757 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10345), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U12758 ( .A1(n10851), .A2(n9874), .ZN(n9873) );
  NAND2_X1 U12759 ( .A1(n13593), .A2(n13592), .ZN(n9888) );
  NAND2_X1 U12760 ( .A1(n13593), .A2(n9881), .ZN(n9880) );
  NAND3_X1 U12761 ( .A1(n10459), .A2(n9890), .A3(n9889), .ZN(n10011) );
  NOR2_X1 U12762 ( .A1(n10458), .A2(n10457), .ZN(n9892) );
  NAND3_X1 U12763 ( .A1(n10252), .A2(n10824), .A3(n9697), .ZN(n9893) );
  INV_X1 U12764 ( .A(n10827), .ZN(n9897) );
  NAND2_X1 U12765 ( .A1(n10148), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U12766 ( .A1(n10148), .A2(n9901), .ZN(n9900) );
  NAND3_X1 U12767 ( .A1(n15244), .A2(n10210), .A3(n10209), .ZN(n9911) );
  NAND2_X1 U12768 ( .A1(n15246), .A2(n15245), .ZN(n15244) );
  NAND2_X1 U12769 ( .A1(n11713), .A2(n9774), .ZN(n9912) );
  NAND2_X1 U12770 ( .A1(n15246), .A2(n9775), .ZN(n9913) );
  NAND2_X1 U12771 ( .A1(n15236), .A2(n11736), .ZN(n9918) );
  NOR2_X2 U12772 ( .A1(n12562), .A2(n9764), .ZN(n15284) );
  AND3_X2 U12773 ( .A1(n12596), .A2(n12597), .A3(n12761), .ZN(n12859) );
  NAND2_X2 U12774 ( .A1(n12059), .A2(n13019), .ZN(n20860) );
  NAND2_X1 U12775 ( .A1(n14777), .A2(n9698), .ZN(n14438) );
  INV_X1 U12776 ( .A(n14424), .ZN(n9933) );
  NAND3_X1 U12777 ( .A1(n14880), .A2(n14426), .A3(n10201), .ZN(n10200) );
  NAND2_X1 U12778 ( .A1(n12195), .A2(n12194), .ZN(n9940) );
  NAND3_X1 U12779 ( .A1(n9940), .A2(n12271), .A3(n16503), .ZN(n9936) );
  OR2_X1 U12780 ( .A1(n12884), .A2(n12883), .ZN(n13164) );
  INV_X1 U12781 ( .A(n15997), .ZN(n9945) );
  NAND2_X1 U12782 ( .A1(n17583), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n9949) );
  INV_X1 U12783 ( .A(n18253), .ZN(n16056) );
  NOR2_X2 U12784 ( .A1(n18183), .A2(n18514), .ZN(n18182) );
  NAND2_X1 U12785 ( .A1(n10093), .A2(n9952), .ZN(n18188) );
  OR2_X2 U12786 ( .A1(n16127), .A2(n9953), .ZN(n18041) );
  OR2_X1 U12787 ( .A1(n17941), .A2(n9777), .ZN(n9959) );
  NAND3_X1 U12788 ( .A1(n9960), .A2(n9958), .A3(n9956), .ZN(n16779) );
  AOI21_X2 U12789 ( .B1(n17926), .B2(n18260), .A(n9961), .ZN(n16138) );
  OR2_X2 U12790 ( .A1(n17941), .A2(n16137), .ZN(n9961) );
  NAND2_X1 U12791 ( .A1(n12625), .A2(n12626), .ZN(n12986) );
  XNOR2_X1 U12792 ( .A(n12984), .B(n20870), .ZN(n12626) );
  NAND2_X1 U12793 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  NAND2_X1 U12794 ( .A1(n10190), .A2(n16386), .ZN(n10189) );
  INV_X2 U12795 ( .A(n13184), .ZN(n9988) );
  AND2_X2 U12796 ( .A1(n9991), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12797) );
  NAND2_X1 U12797 ( .A1(n14638), .A2(n9998), .ZN(n14551) );
  INV_X1 U12798 ( .A(n10007), .ZN(n16272) );
  AND2_X4 U12799 ( .A1(n15888), .A2(n10259), .ZN(n10478) );
  AND2_X2 U12800 ( .A1(n10162), .A2(n10012), .ZN(n15888) );
  NAND2_X4 U12801 ( .A1(n20279), .A2(n20281), .ZN(n13262) );
  NAND3_X1 U12802 ( .A1(n10553), .A2(n10861), .A3(n10161), .ZN(n10015) );
  NOR2_X2 U12803 ( .A1(n10807), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U12804 ( .A1(n10731), .A2(n10025), .ZN(n10741) );
  NAND2_X1 U12805 ( .A1(n10731), .A2(n12471), .ZN(n10734) );
  AND2_X2 U12806 ( .A1(n10031), .A2(n10028), .ZN(n10720) );
  NAND2_X1 U12807 ( .A1(n10742), .A2(n10034), .ZN(n10760) );
  NAND2_X1 U12808 ( .A1(n15094), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15093) );
  NAND2_X1 U12809 ( .A1(n15391), .A2(n9709), .ZN(n11025) );
  NAND2_X1 U12810 ( .A1(n11095), .A2(n10052), .ZN(n10054) );
  NAND2_X1 U12811 ( .A1(n13425), .A2(n10055), .ZN(n13285) );
  NAND2_X1 U12812 ( .A1(n13325), .A2(n10056), .ZN(n15781) );
  NAND2_X1 U12813 ( .A1(n11284), .A2(n10063), .ZN(n13581) );
  AND2_X2 U12814 ( .A1(n15083), .A2(n9781), .ZN(n15317) );
  INV_X1 U12815 ( .A(n16129), .ZN(n10078) );
  NAND2_X1 U12816 ( .A1(n16138), .A2(n18267), .ZN(n16777) );
  NAND2_X1 U12817 ( .A1(n16188), .A2(n9957), .ZN(n10080) );
  NAND3_X1 U12818 ( .A1(n16016), .A2(n16013), .A3(n10085), .ZN(n10084) );
  INV_X1 U12819 ( .A(n10092), .ZN(n18225) );
  INV_X1 U12820 ( .A(n16088), .ZN(n10091) );
  INV_X2 U12821 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19207) );
  INV_X2 U12822 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19219) );
  INV_X1 U12823 ( .A(n10097), .ZN(n18201) );
  NAND3_X1 U12824 ( .A1(n10100), .A2(n10098), .A3(n18148), .ZN(n18120) );
  INV_X1 U12825 ( .A(n10100), .ZN(n10099) );
  NAND2_X1 U12826 ( .A1(n10102), .A2(n10372), .ZN(n10332) );
  NAND2_X2 U12827 ( .A1(n10271), .A2(n10270), .ZN(n10372) );
  INV_X2 U12828 ( .A(n19590), .ZN(n10102) );
  NAND3_X1 U12829 ( .A1(n11384), .A2(n10111), .A3(n10108), .ZN(P2_U3016) );
  NAND2_X1 U12830 ( .A1(n15117), .A2(n10112), .ZN(n15247) );
  NAND2_X1 U12831 ( .A1(n15377), .A2(n15375), .ZN(n11031) );
  CLKBUF_X1 U12832 ( .A(n10142), .Z(n10141) );
  NAND2_X2 U12833 ( .A1(n10145), .A2(n10142), .ZN(n10990) );
  NAND2_X2 U12834 ( .A1(n10144), .A2(n10143), .ZN(n10142) );
  INV_X1 U12835 ( .A(n15443), .ZN(n10152) );
  OR2_X2 U12836 ( .A1(n15560), .A2(n10154), .ZN(n10148) );
  NAND3_X1 U12837 ( .A1(n10874), .A2(n10710), .A3(n10717), .ZN(n10714) );
  NAND2_X2 U12838 ( .A1(n10157), .A2(n10708), .ZN(n10874) );
  NAND2_X1 U12839 ( .A1(n10399), .A2(n11037), .ZN(n10159) );
  NAND2_X1 U12840 ( .A1(n10383), .A2(n10382), .ZN(n10399) );
  XNOR2_X1 U12841 ( .A(n10862), .B(n10863), .ZN(n13417) );
  NAND2_X1 U12842 ( .A1(n10861), .A2(n10553), .ZN(n10851) );
  INV_X1 U12843 ( .A(n13145), .ZN(n10161) );
  NAND2_X1 U12844 ( .A1(n10165), .A2(n10163), .ZN(n10871) );
  NAND2_X1 U12845 ( .A1(n13448), .A2(n10869), .ZN(n10165) );
  NAND2_X1 U12846 ( .A1(n15550), .A2(n10166), .ZN(n15506) );
  NOR2_X1 U12847 ( .A1(n15390), .A2(n15626), .ZN(n10887) );
  NAND2_X1 U12848 ( .A1(n12596), .A2(n12597), .ZN(n12670) );
  AOI21_X1 U12849 ( .B1(n13648), .B2(n13859), .A(n13176), .ZN(n13180) );
  NOR2_X1 U12850 ( .A1(n14521), .A2(n14522), .ZN(n14472) );
  NOR2_X1 U12851 ( .A1(n14521), .A2(n10174), .ZN(n14510) );
  NAND3_X1 U12852 ( .A1(n11910), .A2(n11912), .A3(n11911), .ZN(n10196) );
  NAND3_X1 U12853 ( .A1(n11909), .A2(n9733), .A3(n11916), .ZN(n10197) );
  NAND2_X1 U12854 ( .A1(n12539), .A2(n11981), .ZN(n12382) );
  NAND2_X1 U12855 ( .A1(n14438), .A2(n10206), .ZN(n14789) );
  NAND2_X1 U12856 ( .A1(n14789), .A2(n14439), .ZN(n14781) );
  NAND2_X1 U12857 ( .A1(n10200), .A2(n10199), .ZN(n14436) );
  INV_X1 U12858 ( .A(n10331), .ZN(n10207) );
  INV_X1 U12859 ( .A(n11714), .ZN(n10211) );
  NAND2_X1 U12860 ( .A1(n15894), .A2(n10213), .ZN(n10212) );
  NAND2_X1 U12861 ( .A1(n12134), .A2(n12135), .ZN(n12133) );
  NAND2_X1 U12862 ( .A1(n15284), .A2(n9765), .ZN(n10225) );
  NAND3_X1 U12863 ( .A1(n10226), .A2(n10225), .A3(n10223), .ZN(n15270) );
  NAND2_X1 U12864 ( .A1(n17962), .A2(n18000), .ZN(n18037) );
  NAND2_X1 U12865 ( .A1(n17962), .A2(n16134), .ZN(n17956) );
  INV_X1 U12866 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10260) );
  NOR2_X4 U12867 ( .A1(n15085), .A2(n15084), .ZN(n15083) );
  NAND2_X1 U12868 ( .A1(n12107), .A2(n11120), .ZN(n13150) );
  INV_X1 U12869 ( .A(n10874), .ZN(n10875) );
  INV_X1 U12870 ( .A(n12578), .ZN(n12579) );
  NAND2_X1 U12871 ( .A1(n15151), .A2(n15150), .ZN(n15289) );
  OAI22_X1 U12872 ( .A1(n10452), .A2(n19865), .B1(n10628), .B2(n11158), .ZN(
        n10453) );
  NAND2_X1 U12873 ( .A1(n12333), .A2(n20553), .ZN(n12492) );
  NAND2_X1 U12874 ( .A1(n10357), .A2(n10849), .ZN(n10358) );
  NAND2_X1 U12875 ( .A1(n11070), .A2(n10849), .ZN(n11045) );
  NAND2_X1 U12876 ( .A1(n14533), .A2(n14534), .ZN(n14521) );
  OAI21_X2 U12877 ( .B1(n12492), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12491), 
        .ZN(n12577) );
  NAND2_X1 U12878 ( .A1(n10250), .A2(n11070), .ZN(n11066) );
  AOI21_X1 U12879 ( .B1(n14499), .B2(n20456), .A(n14450), .ZN(n14451) );
  NAND2_X1 U12880 ( .A1(n11096), .A2(n19569), .ZN(n10374) );
  AOI22_X1 U12881 ( .A1(n16828), .A2(n18156), .B1(n16829), .B2(n18123), .ZN(
        n16789) );
  INV_X1 U12882 ( .A(n10902), .ZN(n10888) );
  OAI21_X1 U12883 ( .B1(n11834), .B2(n15279), .A(n11833), .ZN(n11835) );
  OR2_X1 U12884 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  AOI22_X1 U12885 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10312) );
  NOR2_X1 U12886 ( .A1(n13882), .A2(n17321), .ZN(n13963) );
  INV_X1 U12887 ( .A(n13891), .ZN(n13957) );
  NAND2_X1 U12888 ( .A1(n20390), .A2(n14498), .ZN(n20385) );
  OR2_X2 U12889 ( .A1(n12392), .A2(n12391), .ZN(n20442) );
  OR2_X1 U12890 ( .A1(n12463), .A2(n12128), .ZN(n12412) );
  INV_X1 U12891 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16261) );
  AND3_X1 U12892 ( .A1(n10279), .A2(n10278), .A3(n9802), .ZN(n10238) );
  NOR2_X1 U12893 ( .A1(n16283), .A2(n20329), .ZN(n10239) );
  OR2_X1 U12894 ( .A1(n18168), .A2(n17898), .ZN(n10240) );
  OR3_X1 U12895 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17979), .ZN(n10241) );
  INV_X1 U12896 ( .A(n13476), .ZN(n13859) );
  AND2_X1 U12897 ( .A1(n11033), .A2(n15376), .ZN(n10242) );
  AND2_X1 U12898 ( .A1(n10371), .A2(n10102), .ZN(n10243) );
  NAND2_X1 U12899 ( .A1(n10102), .A2(n11069), .ZN(n10244) );
  NOR2_X1 U12900 ( .A1(n10402), .A2(n20278), .ZN(n10245) );
  AND2_X1 U12901 ( .A1(n10468), .A2(n10467), .ZN(n10246) );
  OR2_X1 U12902 ( .A1(n11453), .A2(n12552), .ZN(n10247) );
  INV_X1 U12903 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14590) );
  NAND2_X2 U12904 ( .A1(n14745), .A2(n12536), .ZN(n14717) );
  INV_X2 U12905 ( .A(n9773), .ZN(n20447) );
  INV_X1 U12906 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16289) );
  INV_X1 U12907 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21015) );
  OR2_X1 U12908 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19110), .ZN(n19258) );
  INV_X1 U12909 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16280) );
  NOR2_X1 U12910 ( .A1(n20585), .A2(n20692), .ZN(n10248) );
  NAND2_X1 U12911 ( .A1(n17985), .A2(n18242), .ZN(n18012) );
  AND4_X1 U12912 ( .A1(n10355), .A2(n10344), .A3(n11352), .A4(n10343), .ZN(
        n10250) );
  AND2_X1 U12913 ( .A1(n11194), .A2(n11193), .ZN(n12561) );
  AND2_X1 U12914 ( .A1(n10823), .A2(n10994), .ZN(n10252) );
  AND3_X1 U12915 ( .A1(n10258), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10257), .ZN(n10253) );
  NOR2_X1 U12916 ( .A1(n19061), .A2(n13879), .ZN(n13914) );
  NAND3_X1 U12917 ( .A1(n11283), .A2(n11282), .A3(n11281), .ZN(n10254) );
  INV_X1 U12918 ( .A(n12367), .ZN(n12405) );
  AND2_X1 U12919 ( .A1(n14477), .A2(n12049), .ZN(n10255) );
  INV_X1 U12920 ( .A(n12050), .ZN(n11918) );
  AND4_X1 U12921 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n10256) );
  INV_X1 U12922 ( .A(n13167), .ZN(n12005) );
  INV_X1 U12923 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11964) );
  INV_X1 U12924 ( .A(n12020), .ZN(n12022) );
  AOI22_X1 U12925 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10618), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10523) );
  INV_X1 U12926 ( .A(n12001), .ZN(n11973) );
  OR2_X1 U12927 ( .A1(n12882), .A2(n12881), .ZN(n13640) );
  AND2_X1 U12928 ( .A1(n20516), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11967) );
  NOR2_X1 U12929 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11873) );
  OR2_X1 U12930 ( .A1(n12594), .A2(n12593), .ZN(n12619) );
  OR2_X1 U12931 ( .A1(n13043), .A2(n13042), .ZN(n13641) );
  INV_X1 U12932 ( .A(n12540), .ZN(n12056) );
  INV_X1 U12933 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12329) );
  NOR2_X1 U12934 ( .A1(n10361), .A2(n10244), .ZN(n10362) );
  NOR2_X1 U12935 ( .A1(n10369), .A2(n10368), .ZN(n10370) );
  INV_X1 U12936 ( .A(n13165), .ZN(n13166) );
  OR2_X1 U12937 ( .A1(n12225), .A2(n12224), .ZN(n13656) );
  NAND2_X1 U12938 ( .A1(n11968), .A2(n11969), .ZN(n11996) );
  INV_X1 U12939 ( .A(n12678), .ZN(n12679) );
  NOR2_X1 U12940 ( .A1(n13262), .A2(n11062), .ZN(n10365) );
  AND2_X1 U12941 ( .A1(n11606), .A2(n11605), .ZN(n11655) );
  NAND4_X1 U12943 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10317) );
  NAND2_X1 U12944 ( .A1(n15871), .A2(n20263), .ZN(n10842) );
  INV_X1 U12945 ( .A(n14635), .ZN(n14183) );
  INV_X1 U12946 ( .A(n14652), .ZN(n14133) );
  INV_X1 U12947 ( .A(n14351), .ZN(n14345) );
  INV_X1 U12948 ( .A(n14410), .ZN(n14412) );
  AND2_X1 U12949 ( .A1(n12057), .A2(n12318), .ZN(n12176) );
  INV_X1 U12950 ( .A(n12384), .ZN(n12337) );
  INV_X1 U12951 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11024) );
  AND2_X1 U12952 ( .A1(n11821), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U12953 ( .A1(n11424), .A2(n20268), .ZN(n11444) );
  AND2_X1 U12954 ( .A1(n11665), .A2(n11664), .ZN(n11685) );
  INV_X1 U12955 ( .A(n11562), .ZN(n11627) );
  INV_X1 U12956 ( .A(n10381), .ZN(n11804) );
  AND4_X1 U12957 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n9802), .ZN(
        n10292) );
  AND2_X1 U12958 ( .A1(n13004), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14327) );
  AND2_X1 U12959 ( .A1(n14345), .A2(n16235), .ZN(n14200) );
  AND2_X1 U12960 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  INV_X1 U12961 ( .A(n14285), .ZN(n14445) );
  AOI22_X1 U12962 ( .A1(n12217), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11993) );
  OR2_X1 U12963 ( .A1(n14352), .A2(n14753), .ZN(n13006) );
  NOR2_X1 U12964 ( .A1(n13754), .A2(n14590), .ZN(n13784) );
  INV_X1 U12965 ( .A(n13180), .ZN(n13179) );
  AND2_X1 U12966 ( .A1(n13809), .A2(n13808), .ZN(n13833) );
  INV_X1 U12967 ( .A(n20514), .ZN(n13729) );
  INV_X1 U12968 ( .A(n16473), .ZN(n20483) );
  INV_X1 U12969 ( .A(n12272), .ZN(n14091) );
  OAI211_X1 U12970 ( .C1(n13107), .C2(n12337), .A(n12336), .B(n12335), .ZN(
        n12583) );
  NAND2_X1 U12971 ( .A1(n12677), .A2(n16503), .ZN(n12669) );
  AND2_X1 U12972 ( .A1(n15037), .A2(n15036), .ZN(n15040) );
  AND2_X2 U12973 ( .A1(n10256), .A2(n11887), .ZN(n11979) );
  INV_X1 U12974 ( .A(n12814), .ZN(n16145) );
  INV_X1 U12975 ( .A(n12561), .ZN(n11455) );
  NAND2_X1 U12976 ( .A1(n15857), .A2(n11440), .ZN(n11430) );
  AND2_X1 U12977 ( .A1(n11312), .A2(n11311), .ZN(n15145) );
  AND3_X1 U12978 ( .A1(n11304), .A2(n11303), .A3(n11302), .ZN(n15170) );
  AND4_X1 U12979 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n13151) );
  NOR2_X1 U12980 ( .A1(n15721), .A2(n11376), .ZN(n15676) );
  NAND2_X1 U12981 ( .A1(n15597), .A2(n15842), .ZN(n10728) );
  BUF_X1 U12982 ( .A(n10618), .Z(n19554) );
  NOR2_X1 U12983 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19232), .ZN(
        n15932) );
  NAND2_X1 U12984 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16968), .ZN(
        n16808) );
  OAI21_X1 U12985 ( .B1(n16840), .B2(n16786), .A(n18168), .ZN(n16098) );
  NOR2_X1 U12986 ( .A1(n18302), .A2(n18293), .ZN(n17945) );
  NOR2_X1 U12987 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18052), .ZN(
        n18036) );
  INV_X1 U12988 ( .A(n18452), .ZN(n18432) );
  AOI21_X1 U12989 ( .B1(n15953), .B2(n15952), .A(n15951), .ZN(n15969) );
  NAND2_X1 U12990 ( .A1(n14327), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14352) );
  AND2_X1 U12991 ( .A1(n14404), .A2(n14403), .ZN(n14622) );
  INV_X1 U12992 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14571) );
  INV_X1 U12993 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20315) );
  OR2_X1 U12994 ( .A1(n12531), .A2(n14456), .ZN(n12170) );
  OR2_X1 U12995 ( .A1(n12533), .A2(n12532), .ZN(n12535) );
  XNOR2_X1 U12996 ( .A(n13006), .B(n13005), .ZN(n14449) );
  OR2_X1 U12997 ( .A1(n14251), .A2(n14250), .ZN(n14270) );
  NOR2_X1 U12998 ( .A1(n13002), .A2(n14199), .ZN(n14203) );
  AND2_X1 U12999 ( .A1(n13784), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13847) );
  NAND2_X1 U13000 ( .A1(n12905), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13476) );
  OR2_X1 U13001 ( .A1(n12323), .A2(n12322), .ZN(n13727) );
  AND2_X1 U13002 ( .A1(n13727), .A2(n14902), .ZN(n16473) );
  NAND2_X1 U13003 ( .A1(n20483), .A2(n13729), .ZN(n20493) );
  OR2_X1 U13004 ( .A1(n12058), .A2(n12059), .ZN(n12804) );
  AND2_X1 U13005 ( .A1(n12291), .A2(n12290), .ZN(n12814) );
  NAND2_X1 U13006 ( .A1(n20584), .A2(n12939), .ZN(n13714) );
  NOR2_X1 U13007 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20658) );
  NAND3_X1 U13008 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16503), .A3(n12680), 
        .ZN(n12911) );
  NOR2_X1 U13009 ( .A1(n20529), .A2(n13496), .ZN(n20593) );
  AOI21_X1 U13010 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20693), .A(n13496), 
        .ZN(n20705) );
  NOR2_X1 U13011 ( .A1(n11346), .A2(n11345), .ZN(n15882) );
  INV_X1 U13012 ( .A(n19417), .ZN(n19389) );
  AND2_X1 U13013 ( .A1(n11507), .A2(n11506), .ZN(n13578) );
  OR2_X1 U13014 ( .A1(n15818), .A2(n11377), .ZN(n15721) );
  NOR2_X1 U13015 ( .A1(n15845), .A2(n11375), .ZN(n15831) );
  OR2_X1 U13016 ( .A1(n19270), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15727) );
  OR2_X1 U13017 ( .A1(n16761), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16207) );
  INV_X1 U13018 ( .A(n19828), .ZN(n19861) );
  OR2_X1 U13019 ( .A1(n20239), .A2(n20248), .ZN(n19990) );
  NAND2_X1 U13020 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20067), .ZN(n19589) );
  NOR2_X1 U13021 ( .A1(n13978), .A2(n13977), .ZN(n15934) );
  NOR2_X1 U13022 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17147), .ZN(n17128) );
  NOR2_X1 U13023 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17193), .ZN(n17177) );
  NOR2_X1 U13024 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17246), .ZN(n17226) );
  NAND2_X1 U13025 ( .A1(n19264), .A2(n17786), .ZN(n16966) );
  NOR3_X1 U13026 ( .A1(n17779), .A2(n17629), .A3(n17628), .ZN(n17716) );
  OAI21_X1 U13027 ( .B1(n15970), .B2(n15962), .A(n15959), .ZN(n16961) );
  NAND2_X1 U13028 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17967), .ZN(
        n17947) );
  AOI21_X1 U13029 ( .B1(n19248), .B2(n18596), .A(n19228), .ZN(n18606) );
  INV_X1 U13030 ( .A(n17916), .ZN(n16839) );
  NOR2_X2 U13031 ( .A1(n17956), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16136) );
  NOR2_X1 U13032 ( .A1(n18410), .A2(n18082), .ZN(n18397) );
  NOR2_X1 U13033 ( .A1(n18077), .A2(n18410), .ZN(n18396) );
  NOR2_X1 U13034 ( .A1(n19066), .A2(n18585), .ZN(n18465) );
  AND2_X1 U13035 ( .A1(n16096), .A2(n16095), .ZN(n16840) );
  INV_X1 U13036 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18549) );
  INV_X1 U13037 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19074) );
  INV_X1 U13038 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19212) );
  NAND2_X1 U13039 ( .A1(n14289), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14310) );
  INV_X1 U13040 ( .A(n16239), .ZN(n20331) );
  INV_X1 U13041 ( .A(n20385), .ZN(n16315) );
  INV_X1 U13042 ( .A(n14477), .ZN(n14498) );
  INV_X1 U13043 ( .A(n14717), .ZN(n16319) );
  NOR2_X1 U13044 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16506), .ZN(n20413) );
  NAND2_X1 U13045 ( .A1(n14203), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14231) );
  INV_X1 U13046 ( .A(n13000), .ZN(n13046) );
  NOR2_X1 U13047 ( .A1(n16197), .A2(n16407), .ZN(n16390) );
  NOR2_X1 U13048 ( .A1(n20493), .A2(n20465), .ZN(n16475) );
  NAND2_X1 U13049 ( .A1(n12791), .A2(n12300), .ZN(n12786) );
  NOR2_X1 U13050 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13007) );
  OAI211_X1 U13051 ( .C1(n13197), .C2(n13196), .A(n20527), .B(n13195), .ZN(
        n13228) );
  AND2_X1 U13052 ( .A1(n20517), .A2(n13670), .ZN(n20578) );
  AND2_X1 U13053 ( .A1(n15012), .A2(n9680), .ZN(n20517) );
  NOR2_X1 U13054 ( .A1(n9680), .A2(n12761), .ZN(n20584) );
  NOR2_X2 U13055 ( .A1(n20619), .A2(n13671), .ZN(n20645) );
  INV_X1 U13056 ( .A(n13714), .ZN(n12934) );
  AND2_X1 U13057 ( .A1(n20584), .A2(n12949), .ZN(n15075) );
  INV_X1 U13058 ( .A(n20690), .ZN(n20675) );
  INV_X1 U13059 ( .A(n15034), .ZN(n20583) );
  OAI211_X1 U13060 ( .C1(n13113), .C2(n13112), .A(n20527), .B(n13111), .ZN(
        n13137) );
  NOR2_X1 U13061 ( .A1(n20655), .A2(n12674), .ZN(n13103) );
  INV_X1 U13062 ( .A(n20626), .ZN(n20708) );
  NOR2_X1 U13063 ( .A1(n12973), .A2(n13496), .ZN(n20730) );
  INV_X1 U13064 ( .A(n20664), .ZN(n20714) );
  INV_X1 U13065 ( .A(n20640), .ZN(n20738) );
  AND3_X1 U13066 ( .A1(n16503), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16504) );
  INV_X1 U13067 ( .A(n20866), .ZN(n20812) );
  INV_X1 U13068 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20763) );
  INV_X1 U13069 ( .A(n11830), .ZN(n16721) );
  NAND2_X1 U13070 ( .A1(n16521), .A2(n13253), .ZN(n19411) );
  AND3_X1 U13071 ( .A1(n11215), .A2(n11214), .A3(n11213), .ZN(n12649) );
  OR2_X1 U13072 ( .A1(n12553), .A2(n12552), .ZN(n12840) );
  OR2_X1 U13073 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  AND2_X1 U13074 ( .A1(n19463), .A2(n11811), .ZN(n19487) );
  INV_X1 U13075 ( .A(n20273), .ZN(n19521) );
  OAI21_X1 U13076 ( .B1(n11390), .B2(n19532), .A(n11389), .ZN(n11391) );
  INV_X1 U13077 ( .A(n19532), .ZN(n16660) );
  AND2_X1 U13078 ( .A1(n15550), .A2(n15778), .ZN(n16631) );
  NOR2_X1 U13079 ( .A1(n15581), .A2(n15836), .ZN(n16638) );
  INV_X1 U13080 ( .A(n16701), .ZN(n16669) );
  INV_X1 U13081 ( .A(n16710), .ZN(n16690) );
  OR2_X1 U13082 ( .A1(n11370), .A2(n11340), .ZN(n16701) );
  INV_X1 U13083 ( .A(n19529), .ZN(n19363) );
  NAND2_X1 U13084 ( .A1(n16207), .A2(n16206), .ZN(n20067) );
  OAI21_X1 U13085 ( .B1(n19557), .B2(n19556), .A(n19555), .ZN(n19593) );
  INV_X1 U13086 ( .A(n19650), .ZN(n19672) );
  OAI21_X1 U13087 ( .B1(n19717), .B2(n19716), .A(n19715), .ZN(n19735) );
  INV_X1 U13088 ( .A(n19732), .ZN(n19734) );
  AND2_X1 U13089 ( .A1(n19807), .A2(n19984), .ZN(n19793) );
  INV_X1 U13090 ( .A(n19851), .ZN(n19855) );
  AND2_X1 U13091 ( .A1(n20239), .A2(n20248), .ZN(n20224) );
  INV_X1 U13092 ( .A(n20090), .ZN(n19965) );
  AND2_X1 U13093 ( .A1(n19988), .A2(n19983), .ZN(n20014) );
  INV_X1 U13094 ( .A(n20084), .ZN(n20036) );
  AND2_X1 U13095 ( .A1(n19927), .A2(n20062), .ZN(n20116) );
  INV_X1 U13096 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20149) );
  NOR2_X1 U13097 ( .A1(n19175), .A2(n17029), .ZN(n17015) );
  INV_X1 U13098 ( .A(n17336), .ZN(n17325) );
  NOR2_X1 U13099 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17097), .ZN(n17084) );
  NOR2_X1 U13100 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17167), .ZN(n17155) );
  NOR2_X1 U13101 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17219), .ZN(n17198) );
  NOR2_X1 U13102 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17299), .ZN(n17283) );
  NOR2_X1 U13103 ( .A1(n17333), .A2(n19202), .ZN(n17305) );
  INV_X1 U13104 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20911) );
  NOR2_X2 U13105 ( .A1(n13890), .A2(n13889), .ZN(n18613) );
  NAND2_X1 U13106 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17661), .ZN(n17660) );
  NOR2_X1 U13107 ( .A1(n17833), .A2(n17703), .ZN(n17697) );
  INV_X1 U13108 ( .A(n17769), .ZN(n17696) );
  NOR2_X1 U13109 ( .A1(n16102), .A2(n18629), .ZN(n19069) );
  INV_X1 U13110 ( .A(n18609), .ZN(n17786) );
  INV_X1 U13111 ( .A(n17824), .ZN(n17817) );
  OAI211_X1 U13112 ( .C1(n18613), .C2(n19093), .A(n17827), .B(n17826), .ZN(
        n17882) );
  INV_X1 U13113 ( .A(n17751), .ZN(n16786) );
  INV_X1 U13114 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18193) );
  NOR2_X1 U13115 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18606), .ZN(n18947) );
  NOR2_X1 U13116 ( .A1(n19246), .A2(n16946), .ZN(n18254) );
  INV_X1 U13117 ( .A(n18168), .ZN(n18052) );
  NOR2_X1 U13118 ( .A1(n18399), .A2(n18410), .ZN(n18366) );
  NAND2_X1 U13119 ( .A1(n16100), .A2(n18450), .ZN(n18077) );
  INV_X1 U13120 ( .A(n18586), .ZN(n18498) );
  INV_X1 U13121 ( .A(n18582), .ZN(n18592) );
  INV_X1 U13122 ( .A(n18947), .ZN(n18842) );
  NOR2_X1 U13123 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19202), .ZN(
        n19228) );
  INV_X1 U13124 ( .A(n18739), .ZN(n18745) );
  INV_X1 U13125 ( .A(n18840), .ZN(n18833) );
  INV_X1 U13126 ( .A(n18925), .ZN(n18938) );
  NAND2_X1 U13127 ( .A1(n19212), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19102) );
  INV_X1 U13128 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19110) );
  INV_X1 U13129 ( .A(n19545), .ZN(n19543) );
  INV_X1 U13130 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20702) );
  INV_X1 U13131 ( .A(n20374), .ZN(n20316) );
  NOR2_X1 U13132 ( .A1(n14562), .A2(n14599), .ZN(n16312) );
  NAND2_X1 U13133 ( .A1(n20390), .A2(n14477), .ZN(n14666) );
  NAND2_X1 U13134 ( .A1(n14476), .A2(n14482), .ZN(n21068) );
  OR2_X1 U13135 ( .A1(n20396), .A2(n20858), .ZN(n20395) );
  INV_X1 U13136 ( .A(n20396), .ZN(n20418) );
  INV_X1 U13137 ( .A(n20442), .ZN(n12515) );
  OAI21_X1 U13138 ( .B1(n14740), .B2(n13824), .A(n13823), .ZN(n14875) );
  INV_X1 U13139 ( .A(n16365), .ZN(n20461) );
  AND2_X1 U13140 ( .A1(n16391), .A2(n14901), .ZN(n14981) );
  OAI21_X1 U13141 ( .B1(n20484), .B2(n16475), .A(n20497), .ZN(n20478) );
  INV_X1 U13142 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16151) );
  INV_X1 U13143 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12868) );
  NAND2_X1 U13144 ( .A1(n20517), .A2(n20583), .ZN(n20582) );
  AOI22_X1 U13145 ( .A1(n13194), .A2(n13196), .B1(n13674), .B2(n20529), .ZN(
        n13231) );
  NAND2_X1 U13146 ( .A1(n20517), .A2(n12939), .ZN(n13226) );
  NAND2_X1 U13147 ( .A1(n20584), .A2(n20583), .ZN(n20649) );
  INV_X1 U13148 ( .A(n15075), .ZN(n12938) );
  NAND2_X1 U13149 ( .A1(n15035), .A2(n20583), .ZN(n20690) );
  AOI22_X1 U13150 ( .A1(n13102), .A2(n13112), .B1(n13500), .B2(n20529), .ZN(
        n13140) );
  NAND2_X1 U13151 ( .A1(n15035), .A2(n12949), .ZN(n13543) );
  INV_X1 U13152 ( .A(n20700), .ZN(n13686) );
  AOI22_X1 U13153 ( .A1(n13547), .A2(n13544), .B1(n13675), .B2(n15041), .ZN(
        n13576) );
  NAND2_X1 U13154 ( .A1(n13491), .A2(n13670), .ZN(n20757) );
  INV_X1 U13155 ( .A(n20548), .ZN(n12927) );
  AND2_X1 U13156 ( .A1(n20778), .A2(n20867), .ZN(n20845) );
  CLKBUF_X1 U13157 ( .A(n20812), .Z(n20867) );
  INV_X1 U13158 ( .A(n10776), .ZN(n15141) );
  INV_X1 U13159 ( .A(n19396), .ZN(n19413) );
  INV_X1 U13160 ( .A(n19377), .ZN(n19408) );
  INV_X1 U13161 ( .A(n11835), .ZN(n11836) );
  AND2_X1 U13162 ( .A1(n11831), .A2(n20122), .ZN(n15291) );
  NAND2_X1 U13163 ( .A1(n12097), .A2(n12096), .ZN(n20256) );
  INV_X1 U13164 ( .A(n19487), .ZN(n19458) );
  NOR2_X1 U13165 ( .A1(n19486), .A2(n19487), .ZN(n19462) );
  AND2_X1 U13166 ( .A1(n19428), .A2(n19427), .ZN(n19492) );
  OR2_X1 U13167 ( .A1(n19494), .A2(n19521), .ZN(n19509) );
  INV_X1 U13168 ( .A(n19494), .ZN(n19527) );
  INV_X1 U13169 ( .A(n12463), .ZN(n12366) );
  INV_X1 U13170 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16635) );
  OR2_X1 U13171 ( .A1(n11370), .A2(n16716), .ZN(n16697) );
  NAND2_X1 U13172 ( .A1(n19828), .A2(n19767), .ZN(n19647) );
  NAND2_X1 U13173 ( .A1(n19767), .A2(n20224), .ZN(n19706) );
  NAND2_X1 U13174 ( .A1(n19807), .A2(n20224), .ZN(n19732) );
  INV_X1 U13175 ( .A(n19793), .ZN(n19770) );
  NAND2_X1 U13176 ( .A1(n20062), .A2(n19767), .ZN(n19826) );
  NAND2_X1 U13177 ( .A1(n20019), .A2(n19828), .ZN(n19882) );
  NAND2_X1 U13178 ( .A1(n20019), .A2(n20224), .ZN(n19942) );
  INV_X1 U13179 ( .A(n20069), .ZN(n19995) );
  INV_X1 U13180 ( .A(n20093), .ZN(n20005) );
  INV_X1 U13181 ( .A(n20081), .ZN(n20039) );
  INV_X1 U13182 ( .A(n20032), .ZN(n20078) );
  NAND2_X1 U13183 ( .A1(n20019), .A2(n20062), .ZN(n20120) );
  OR4_X1 U13184 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), 
        .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n15859), .ZN(n20126) );
  INV_X1 U13185 ( .A(n20217), .ZN(n20129) );
  INV_X1 U13186 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16967) );
  OR2_X1 U13187 ( .A1(n17326), .A2(n16982), .ZN(n17081) );
  INV_X1 U13188 ( .A(n17337), .ZN(n17275) );
  NOR2_X1 U13189 ( .A1(n17348), .A2(n17347), .ZN(n17373) );
  INV_X1 U13190 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17618) );
  NOR2_X1 U13191 ( .A1(n15980), .A2(n15979), .ZN(n17751) );
  NOR2_X1 U13192 ( .A1(n17717), .A2(n17747), .ZN(n17753) );
  NAND2_X1 U13193 ( .A1(n19069), .A2(n17631), .ZN(n17771) );
  NAND2_X1 U13194 ( .A1(n17817), .A2(n17786), .ZN(n17803) );
  OR2_X1 U13195 ( .A1(n19096), .A2(n17817), .ZN(n17811) );
  NAND2_X1 U13196 ( .A1(n17826), .A2(n17784), .ZN(n17824) );
  INV_X1 U13197 ( .A(n17882), .ZN(n17865) );
  NAND2_X1 U13198 ( .A1(n18366), .A2(n18125), .ZN(n18063) );
  INV_X1 U13199 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18221) );
  INV_X1 U13200 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21047) );
  INV_X1 U13201 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18484) );
  INV_X1 U13202 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18841) );
  INV_X1 U13203 ( .A(n18712), .ZN(n18727) );
  INV_X1 U13204 ( .A(n18892), .ZN(n18992) );
  INV_X1 U13205 ( .A(n19090), .ZN(n19254) );
  INV_X1 U13206 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19202) );
  INV_X1 U13207 ( .A(n19199), .ZN(n19196) );
  NOR2_X1 U13208 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n11852), .ZN(n16928)
         );
  AOI22_X1 U13209 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11781), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13210 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10257) );
  AND2_X4 U13211 ( .A1(n15888), .A2(n15871), .ZN(n10483) );
  AND2_X4 U13212 ( .A1(n15876), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11674) );
  AOI22_X1 U13213 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10262) );
  AND3_X4 U13214 ( .A1(n10260), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13215 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13216 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13217 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10345), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U13218 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13219 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10266) );
  NAND4_X1 U13220 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10270) );
  AOI22_X1 U13221 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U13222 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13223 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13224 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11781), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13225 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10484), .B1(
        n11666), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13226 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13227 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9663), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13228 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U13229 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13230 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11666), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13231 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13232 ( .A1(n10345), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11666), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13233 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13234 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13235 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U13236 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  AOI22_X1 U13237 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10478), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13238 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13239 ( .A1(n11674), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13240 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11666), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10295) );
  NAND4_X1 U13241 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10299) );
  NAND2_X1 U13242 ( .A1(n10299), .A2(n9802), .ZN(n10306) );
  AOI22_X1 U13243 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13244 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11666), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13245 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13246 ( .A1(n10345), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10300) );
  NAND4_X1 U13247 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10304) );
  NAND2_X1 U13248 ( .A1(n10304), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10305) );
  AOI22_X1 U13249 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13250 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13251 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13252 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10345), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U13253 ( .A1(n10311), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10318) );
  AOI22_X1 U13254 ( .A1(n10345), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11666), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13255 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13256 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13257 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13258 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13259 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13260 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10345), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13261 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13262 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13263 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13264 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11781), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10325) );
  NAND2_X1 U13265 ( .A1(n10384), .A2(n10385), .ZN(n10331) );
  AOI22_X1 U13266 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11781), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13267 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13268 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13269 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U13270 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10342) );
  AOI22_X1 U13271 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U13272 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13273 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10345), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13274 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10337) );
  NAND4_X1 U13275 ( .A1(n10340), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        n10341) );
  MUX2_X2 U13276 ( .A(n10342), .B(n10341), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n20279) );
  NOR2_X2 U13277 ( .A1(n19590), .A2(n10372), .ZN(n10355) );
  NOR2_X1 U13278 ( .A1(n19564), .A2(n10385), .ZN(n10344) );
  INV_X1 U13279 ( .A(n19569), .ZN(n10343) );
  NAND2_X1 U13280 ( .A1(n11866), .A2(n11066), .ZN(n11338) );
  AOI22_X1 U13281 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13282 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13283 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13284 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11674), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13285 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13286 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11781), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13287 ( .A1(n11666), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10484), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10353) );
  OR2_X2 U13288 ( .A1(n11338), .A2(n10356), .ZN(n10390) );
  NAND2_X1 U13289 ( .A1(n10385), .A2(n10372), .ZN(n10378) );
  INV_X1 U13290 ( .A(n10378), .ZN(n10357) );
  INV_X1 U13291 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10594) );
  AND2_X1 U13292 ( .A1(n10385), .A2(n11423), .ZN(n10364) );
  NAND2_X2 U13293 ( .A1(n11364), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10408) );
  INV_X1 U13294 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10366) );
  NOR2_X1 U13295 ( .A1(n20277), .A2(n16723), .ZN(n10406) );
  AOI22_X1 U13296 ( .A1(n10413), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10367) );
  INV_X1 U13297 ( .A(n10367), .ZN(n10368) );
  OAI21_X2 U13298 ( .B1(n10902), .B2(n10594), .A(n10370), .ZN(n10394) );
  NOR2_X1 U13299 ( .A1(n10250), .A2(n20279), .ZN(n10376) );
  OR2_X1 U13300 ( .A1(n10372), .A2(n10385), .ZN(n10379) );
  AND2_X1 U13301 ( .A1(n10379), .A2(n19564), .ZN(n10373) );
  NAND3_X1 U13302 ( .A1(n10243), .A2(n10374), .A3(n10373), .ZN(n10375) );
  NAND2_X1 U13303 ( .A1(n10376), .A2(n10375), .ZN(n11358) );
  AND2_X1 U13304 ( .A1(n11096), .A2(n10849), .ZN(n11354) );
  INV_X1 U13305 ( .A(n11354), .ZN(n10401) );
  NAND2_X1 U13306 ( .A1(n10401), .A2(n11070), .ZN(n10377) );
  NAND2_X1 U13307 ( .A1(n11096), .A2(n11069), .ZN(n11067) );
  NAND2_X1 U13308 ( .A1(n11063), .A2(n10380), .ZN(n11359) );
  NAND2_X1 U13309 ( .A1(n11359), .A2(n19569), .ZN(n10383) );
  INV_X1 U13310 ( .A(n10355), .ZN(n10386) );
  NOR2_X1 U13311 ( .A1(n10386), .A2(n11821), .ZN(n10387) );
  NAND2_X1 U13312 ( .A1(n10384), .A2(n10387), .ZN(n11089) );
  AND2_X1 U13313 ( .A1(n19564), .A2(n20281), .ZN(n10388) );
  NAND2_X1 U13314 ( .A1(n11089), .A2(n10388), .ZN(n11337) );
  INV_X1 U13315 ( .A(n11077), .ZN(n10389) );
  NAND3_X1 U13316 ( .A1(n11337), .A2(n12245), .A3(n10389), .ZN(n10395) );
  NAND2_X1 U13317 ( .A1(n10433), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10392) );
  AOI22_X1 U13318 ( .A1(n10390), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20270), .ZN(n10391) );
  NAND2_X1 U13319 ( .A1(n10392), .A2(n10391), .ZN(n10393) );
  NAND2_X1 U13320 ( .A1(n10394), .A2(n10393), .ZN(n10422) );
  AND2_X2 U13321 ( .A1(n10423), .A2(n10422), .ZN(n10419) );
  INV_X1 U13322 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12098) );
  OAI21_X1 U13323 ( .B1(n10408), .B2(n12098), .A(n10395), .ZN(n10398) );
  INV_X1 U13324 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19406) );
  INV_X1 U13325 ( .A(n20270), .ZN(n16756) );
  NAND2_X1 U13326 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10396) );
  OAI211_X1 U13327 ( .C1(n10890), .C2(n19406), .A(n16756), .B(n10396), .ZN(
        n10397) );
  AOI21_X1 U13328 ( .B1(n10399), .B2(n10401), .A(n10400), .ZN(n10402) );
  NAND2_X1 U13329 ( .A1(n10888), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13330 ( .A1(n10405), .A2(n10404), .ZN(n10434) );
  INV_X1 U13331 ( .A(n10406), .ZN(n10407) );
  NOR2_X1 U13332 ( .A1(n10407), .A2(n11062), .ZN(n10409) );
  OAI22_X1 U13333 ( .A1(n10433), .A2(n10409), .B1(n15871), .B2(n10889), .ZN(
        n10412) );
  INV_X1 U13334 ( .A(n15886), .ZN(n10410) );
  AOI22_X1 U13335 ( .A1(n10410), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n20270), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U13336 ( .A1(n10412), .A2(n10411), .ZN(n10435) );
  NAND2_X1 U13337 ( .A1(n10419), .A2(n10436), .ZN(n10447) );
  NAND2_X1 U13338 ( .A1(n10447), .A2(n10423), .ZN(n10418) );
  INV_X1 U13339 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U13340 ( .A1(n9678), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10415) );
  NAND2_X1 U13341 ( .A1(n10889), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10414) );
  INV_X1 U13342 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15859) );
  OAI21_X1 U13343 ( .B1(n20243), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15859), 
        .ZN(n10416) );
  XNOR2_X1 U13344 ( .A(n10426), .B(n10421), .ZN(n10417) );
  XNOR2_X2 U13345 ( .A(n10418), .B(n10417), .ZN(n10446) );
  BUF_X4 U13346 ( .A(n10446), .Z(n15894) );
  INV_X1 U13347 ( .A(n10436), .ZN(n10420) );
  INV_X1 U13348 ( .A(n10421), .ZN(n10427) );
  NAND2_X1 U13349 ( .A1(n10427), .A2(n10426), .ZN(n10424) );
  INV_X1 U13350 ( .A(n10423), .ZN(n10425) );
  INV_X1 U13351 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11372) );
  INV_X2 U13352 ( .A(n10890), .ZN(n10942) );
  AOI22_X1 U13353 ( .A1(n10942), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10431) );
  NAND2_X1 U13354 ( .A1(n10889), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10430) );
  AND2_X1 U13355 ( .A1(n20270), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10432) );
  OR2_X1 U13356 ( .A1(n10435), .A2(n10434), .ZN(n10448) );
  INV_X1 U13357 ( .A(n15857), .ZN(n19414) );
  NAND2_X1 U13358 ( .A1(n10451), .A2(n19414), .ZN(n10441) );
  AND2_X2 U13359 ( .A1(n15894), .A2(n10438), .ZN(n10440) );
  AND2_X2 U13360 ( .A1(n10440), .A2(n12104), .ZN(n19714) );
  NAND2_X1 U13361 ( .A1(n19714), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10439) );
  AND2_X2 U13362 ( .A1(n10440), .A2(n10437), .ZN(n10622) );
  INV_X1 U13363 ( .A(n10441), .ZN(n10442) );
  AND2_X1 U13364 ( .A1(n10444), .A2(n15857), .ZN(n10456) );
  NAND2_X1 U13365 ( .A1(n15894), .A2(n10456), .ZN(n10445) );
  INV_X1 U13366 ( .A(n10631), .ZN(n19742) );
  INV_X1 U13367 ( .A(n10448), .ZN(n10449) );
  INV_X1 U13368 ( .A(n10467), .ZN(n10450) );
  AOI22_X1 U13369 ( .A1(n19742), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n19678), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10460) );
  INV_X1 U13370 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U13371 ( .A1(n10456), .A2(n10451), .ZN(n10462) );
  NAND2_X1 U13372 ( .A1(n10451), .A2(n10467), .ZN(n10454) );
  INV_X1 U13373 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11158) );
  INV_X1 U13374 ( .A(n10453), .ZN(n10459) );
  INV_X1 U13375 ( .A(n10454), .ZN(n10455) );
  NAND2_X1 U13376 ( .A1(n10455), .A2(n10458), .ZN(n10676) );
  INV_X1 U13377 ( .A(n10676), .ZN(n20058) );
  INV_X1 U13378 ( .A(n10456), .ZN(n10457) );
  NOR2_X2 U13379 ( .A1(n10461), .A2(n10470), .ZN(n10620) );
  INV_X1 U13380 ( .A(n10620), .ZN(n10464) );
  INV_X1 U13381 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11640) );
  INV_X1 U13382 ( .A(n10462), .ZN(n10463) );
  INV_X1 U13383 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U13384 ( .A1(n10466), .A2(n12104), .ZN(n19955) );
  INV_X1 U13385 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11168) );
  NAND2_X2 U13386 ( .A1(n15894), .A2(n10246), .ZN(n19798) );
  INV_X1 U13387 ( .A(n19798), .ZN(n10469) );
  AOI21_X1 U13388 ( .B1(n10469), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(n9659), .ZN(n10473) );
  NAND2_X1 U13389 ( .A1(n10618), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10472) );
  OAI211_X1 U13390 ( .C1(n19955), .C2(n11168), .A(n10473), .B(n10472), .ZN(
        n10474) );
  INV_X1 U13391 ( .A(n10474), .ZN(n10475) );
  AND2_X1 U13392 ( .A1(n10260), .A2(n15871), .ZN(n10476) );
  AOI22_X1 U13393 ( .A1(n11617), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10482) );
  NOR2_X1 U13394 ( .A1(n10260), .A2(n15871), .ZN(n10477) );
  AOI22_X1 U13395 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U13396 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10480) );
  CLKBUF_X3 U13397 ( .A(n10478), .Z(n11794) );
  AND2_X2 U13398 ( .A1(n11794), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11258) );
  NAND2_X1 U13399 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10479) );
  AND4_X1 U13400 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10488) );
  AND2_X2 U13401 ( .A1(n11778), .A2(n9802), .ZN(n11574) );
  AOI22_X1 U13402 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10487) );
  INV_X1 U13403 ( .A(n10484), .ZN(n11585) );
  AND2_X2 U13404 ( .A1(n10485), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11576) );
  AOI22_X1 U13405 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11576), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10486) );
  NAND3_X1 U13406 ( .A1(n10488), .A2(n10487), .A3(n10486), .ZN(n10495) );
  INV_X1 U13407 ( .A(n11781), .ZN(n15903) );
  AOI22_X1 U13408 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10493) );
  AND2_X2 U13409 ( .A1(n11792), .A2(n9802), .ZN(n11563) );
  AND2_X1 U13410 ( .A1(n15871), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10490) );
  AOI22_X1 U13411 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11562), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10492) );
  INV_X1 U13412 ( .A(n9663), .ZN(n11586) );
  AOI22_X1 U13413 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10491) );
  NAND3_X1 U13414 ( .A1(n10493), .A2(n10492), .A3(n10491), .ZN(n10494) );
  AND2_X1 U13415 ( .A1(n9659), .A2(n11095), .ZN(n12035) );
  AOI22_X1 U13416 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11617), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13417 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10498) );
  NAND2_X1 U13418 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10497) );
  NAND2_X1 U13419 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10496) );
  AND4_X1 U13420 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10502) );
  AOI22_X1 U13421 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11574), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13422 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10500) );
  NAND3_X1 U13423 ( .A1(n10502), .A2(n10501), .A3(n10500), .ZN(n10507) );
  AOI22_X1 U13424 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11576), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13425 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n11562), .ZN(n10504) );
  AOI22_X1 U13426 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11563), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10503) );
  NAND3_X1 U13427 ( .A1(n10505), .A2(n10504), .A3(n10503), .ZN(n10506) );
  AND2_X1 U13428 ( .A1(n12035), .A2(n10581), .ZN(n10856) );
  INV_X1 U13429 ( .A(n10856), .ZN(n10521) );
  AOI22_X1 U13430 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11201), .B1(
        n11576), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13431 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n11562), .ZN(n10509) );
  AOI22_X1 U13432 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11563), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13433 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13434 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U13435 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10512) );
  NAND2_X1 U13436 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10511) );
  NAND4_X1 U13437 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10520) );
  NAND2_X1 U13438 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10519) );
  NAND2_X1 U13439 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10518) );
  NAND2_X1 U13440 ( .A1(n11623), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10517) );
  NAND2_X1 U13441 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10516) );
  NAND2_X1 U13442 ( .A1(n10521), .A2(n11112), .ZN(n10522) );
  AOI22_X1 U13443 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10619), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10526) );
  NAND2_X1 U13444 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10525) );
  NAND2_X1 U13445 ( .A1(n20026), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13446 ( .A1(n19714), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10532) );
  INV_X1 U13447 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11519) );
  INV_X1 U13448 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10527) );
  OAI22_X1 U13449 ( .A1(n11519), .A2(n19982), .B1(n10676), .B2(n10527), .ZN(
        n10529) );
  INV_X1 U13450 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11202) );
  INV_X1 U13451 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11197) );
  OAI22_X1 U13452 ( .A1(n11202), .A2(n19865), .B1(n10628), .B2(n11197), .ZN(
        n10528) );
  NOR2_X1 U13453 ( .A1(n10529), .A2(n10528), .ZN(n10531) );
  NAND2_X1 U13454 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10530) );
  INV_X1 U13455 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10533) );
  INV_X1 U13456 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11509) );
  OAI22_X1 U13457 ( .A1(n10533), .A2(n10631), .B1(n19798), .B2(n11509), .ZN(
        n10536) );
  INV_X1 U13458 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11511) );
  INV_X1 U13459 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10534) );
  OAI22_X1 U13460 ( .A1(n11511), .A2(n10682), .B1(n10684), .B2(n10534), .ZN(
        n10535) );
  NOR2_X1 U13461 ( .A1(n10536), .A2(n10535), .ZN(n10537) );
  AOI22_X1 U13462 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11617), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13463 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U13464 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10541) );
  NAND2_X1 U13465 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10540) );
  AND4_X1 U13466 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10546) );
  AOI22_X1 U13467 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11574), .B1(
        n11258), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13468 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11623), .B1(
        n11576), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10544) );
  NAND3_X1 U13469 ( .A1(n10546), .A2(n10545), .A3(n10544), .ZN(n10551) );
  AOI22_X1 U13470 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11201), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13471 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11562), .ZN(n10548) );
  AOI22_X1 U13472 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10547) );
  NAND3_X1 U13473 ( .A1(n10549), .A2(n10548), .A3(n10547), .ZN(n10550) );
  INV_X1 U13474 ( .A(n10586), .ZN(n11121) );
  NAND2_X1 U13475 ( .A1(n11121), .A2(n9659), .ZN(n10552) );
  AOI22_X1 U13476 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13477 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n11562), .ZN(n10555) );
  AOI22_X1 U13478 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10554) );
  AND3_X1 U13479 ( .A1(n10556), .A2(n10555), .A3(n10554), .ZN(n10568) );
  AOI22_X1 U13480 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11617), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13481 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10559) );
  NAND2_X1 U13482 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13483 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10557) );
  NAND4_X1 U13484 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10566) );
  NAND2_X1 U13485 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U13486 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U13487 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10562) );
  NAND2_X1 U13488 ( .A1(n11576), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10561) );
  NAND4_X1 U13489 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10565) );
  NOR2_X1 U13490 ( .A1(n10566), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U13491 ( .A1(n10260), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10569) );
  NAND2_X1 U13492 ( .A1(n10572), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10573) );
  NAND2_X1 U13493 ( .A1(n10584), .A2(n10573), .ZN(n10575) );
  NAND2_X1 U13494 ( .A1(n10574), .A2(n10575), .ZN(n10578) );
  INV_X1 U13495 ( .A(n10575), .ZN(n10576) );
  NAND2_X1 U13496 ( .A1(n10578), .A2(n10585), .ZN(n11044) );
  NAND2_X1 U13497 ( .A1(n10366), .A2(n12098), .ZN(n10583) );
  MUX2_X1 U13498 ( .A(n11108), .B(n10583), .S(n11821), .Z(n10592) );
  NOR2_X2 U13499 ( .A1(n10589), .A2(n10592), .ZN(n10588) );
  XNOR2_X1 U13500 ( .A(n10599), .B(n10600), .ZN(n10840) );
  MUX2_X1 U13501 ( .A(n10586), .B(n10840), .S(n13262), .Z(n10833) );
  INV_X1 U13502 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13274) );
  MUX2_X1 U13503 ( .A(n10833), .B(n13274), .S(n11821), .Z(n10587) );
  OAI21_X1 U13504 ( .B1(n10588), .B2(n10587), .A(n10659), .ZN(n13275) );
  XNOR2_X1 U13505 ( .A(n10589), .B(n10592), .ZN(n15217) );
  XNOR2_X1 U13506 ( .A(n15217), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12082) );
  OAI21_X1 U13507 ( .B1(n15871), .B2(n20263), .A(n10842), .ZN(n11039) );
  INV_X1 U13508 ( .A(n11039), .ZN(n11041) );
  MUX2_X1 U13509 ( .A(n11095), .B(n11041), .S(n13262), .Z(n10829) );
  MUX2_X1 U13510 ( .A(n10829), .B(P2_EBX_REG_0__SCAN_IN), .S(n11007), .Z(
        n19402) );
  NAND2_X1 U13511 ( .A1(n19402), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12034) );
  AND2_X1 U13512 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10590) );
  NAND2_X1 U13513 ( .A1(n11007), .A2(n10590), .ZN(n10591) );
  NAND2_X1 U13514 ( .A1(n10592), .A2(n10591), .ZN(n19390) );
  INV_X1 U13515 ( .A(n19390), .ZN(n10593) );
  NAND2_X1 U13516 ( .A1(n10593), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10596) );
  AND2_X1 U13517 ( .A1(n19390), .A2(n10594), .ZN(n10595) );
  AOI21_X1 U13518 ( .B1(n12034), .B2(n10596), .A(n10595), .ZN(n12081) );
  NAND2_X1 U13519 ( .A1(n12082), .A2(n12081), .ZN(n12080) );
  INV_X1 U13520 ( .A(n15217), .ZN(n10597) );
  NAND2_X1 U13521 ( .A1(n10597), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10598) );
  AND2_X1 U13522 ( .A1(n12080), .A2(n10598), .ZN(n13143) );
  NAND3_X1 U13523 ( .A1(n20221), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10836), .ZN(n10841) );
  AOI22_X1 U13524 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11617), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13525 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13526 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10604) );
  NAND2_X1 U13527 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10603) );
  AND4_X1 U13528 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n10609) );
  AOI22_X1 U13529 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11574), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13530 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11576), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10607) );
  NAND3_X1 U13531 ( .A1(n10609), .A2(n10608), .A3(n10607), .ZN(n10614) );
  AOI22_X1 U13532 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13533 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n11562), .ZN(n10611) );
  AOI22_X1 U13534 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10610) );
  NAND3_X1 U13535 ( .A1(n10612), .A2(n10611), .A3(n10610), .ZN(n10613) );
  MUX2_X1 U13536 ( .A(n10841), .B(n11126), .S(n11037), .Z(n10834) );
  INV_X1 U13537 ( .A(n10834), .ZN(n10615) );
  MUX2_X1 U13538 ( .A(n10615), .B(P2_EBX_REG_4__SCAN_IN), .S(n11821), .Z(
        n10658) );
  XNOR2_X1 U13539 ( .A(n10658), .B(n10659), .ZN(n19375) );
  INV_X1 U13540 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13422) );
  XNOR2_X1 U13541 ( .A(n19375), .B(n13422), .ZN(n13420) );
  AOI22_X1 U13542 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19554), .B1(
        n19836), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13543 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10620), .B1(
        n19894), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13544 ( .A1(n19714), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10624) );
  NAND2_X1 U13545 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10623) );
  NAND4_X1 U13546 ( .A1(n10626), .A2(n10625), .A3(n10624), .A4(n10623), .ZN(
        n10642) );
  INV_X1 U13547 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11246) );
  INV_X1 U13548 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10627) );
  OAI22_X1 U13549 ( .A1(n11246), .A2(n10676), .B1(n19865), .B2(n10627), .ZN(
        n10630) );
  INV_X1 U13550 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11239) );
  INV_X1 U13551 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11238) );
  OAI22_X1 U13552 ( .A1(n11239), .A2(n19982), .B1(n10628), .B2(n11238), .ZN(
        n10629) );
  NOR2_X1 U13553 ( .A1(n10630), .A2(n10629), .ZN(n10640) );
  INV_X1 U13554 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11249) );
  INV_X1 U13555 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11248) );
  OAI22_X1 U13556 ( .A1(n19798), .A2(n11249), .B1(n10682), .B2(n11248), .ZN(
        n10635) );
  INV_X1 U13557 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10633) );
  INV_X1 U13558 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10632) );
  OAI22_X1 U13559 ( .A1(n10631), .A2(n10633), .B1(n10684), .B2(n10632), .ZN(
        n10634) );
  NOR2_X1 U13560 ( .A1(n10635), .A2(n10634), .ZN(n10639) );
  NAND2_X1 U13561 ( .A1(n20026), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10638) );
  NAND2_X1 U13562 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10637) );
  NAND4_X1 U13563 ( .A1(n10640), .A2(n10639), .A3(n10638), .A4(n10637), .ZN(
        n10641) );
  NOR2_X1 U13564 ( .A1(n10642), .A2(n10641), .ZN(n10643) );
  INV_X1 U13565 ( .A(n10643), .ZN(n10657) );
  AOI22_X1 U13566 ( .A1(n11617), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13567 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U13568 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10645) );
  NAND2_X1 U13569 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10644) );
  AND4_X1 U13570 ( .A1(n10647), .A2(n10646), .A3(n10645), .A4(n10644), .ZN(
        n10650) );
  AOI22_X1 U13571 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13572 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11576), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10648) );
  NAND3_X1 U13573 ( .A1(n10650), .A2(n10649), .A3(n10648), .ZN(n10655) );
  AOI22_X1 U13574 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13575 ( .A1(n11564), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11562), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13576 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11563), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10651) );
  NAND3_X1 U13577 ( .A1(n10653), .A2(n10652), .A3(n10651), .ZN(n10654) );
  INV_X1 U13578 ( .A(n10660), .ZN(n11131) );
  NAND2_X1 U13579 ( .A1(n11131), .A2(n9659), .ZN(n10656) );
  XNOR2_X2 U13580 ( .A(n10668), .B(n10669), .ZN(n10866) );
  NAND2_X1 U13581 ( .A1(n10866), .A2(n10717), .ZN(n10664) );
  INV_X1 U13582 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12411) );
  MUX2_X1 U13583 ( .A(n10660), .B(n12411), .S(n11821), .Z(n10662) );
  INV_X1 U13584 ( .A(n10712), .ZN(n10661) );
  OAI21_X1 U13585 ( .B1(n10663), .B2(n10662), .A(n10661), .ZN(n13292) );
  NAND2_X1 U13586 ( .A1(n10664), .A2(n13292), .ZN(n10665) );
  INV_X1 U13587 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13455) );
  XNOR2_X1 U13588 ( .A(n10665), .B(n13455), .ZN(n13450) );
  NAND2_X1 U13589 ( .A1(n13449), .A2(n13450), .ZN(n10667) );
  NAND2_X1 U13590 ( .A1(n10665), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10666) );
  NAND2_X1 U13591 ( .A1(n10667), .A2(n10666), .ZN(n13593) );
  INV_X1 U13592 ( .A(n10668), .ZN(n10670) );
  NAND2_X1 U13593 ( .A1(n10670), .A2(n10669), .ZN(n10709) );
  AOI22_X1 U13594 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19554), .B1(
        n19894), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13595 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10620), .B1(
        n19836), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U13596 ( .A1(n19714), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10672) );
  NAND2_X1 U13597 ( .A1(n20026), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10671) );
  NAND4_X1 U13598 ( .A1(n10674), .A2(n10673), .A3(n10672), .A4(n10671), .ZN(
        n10693) );
  INV_X1 U13599 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11267) );
  INV_X1 U13600 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10675) );
  OAI22_X1 U13601 ( .A1(n11267), .A2(n19982), .B1(n10676), .B2(n10675), .ZN(
        n10679) );
  INV_X1 U13602 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10677) );
  INV_X1 U13603 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11265) );
  OAI22_X1 U13604 ( .A1(n10677), .A2(n10628), .B1(n19865), .B2(n11265), .ZN(
        n10678) );
  NOR2_X1 U13605 ( .A1(n10679), .A2(n10678), .ZN(n10691) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10681) );
  INV_X1 U13607 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10680) );
  OAI22_X1 U13608 ( .A1(n10681), .A2(n10631), .B1(n19798), .B2(n10680), .ZN(
        n10687) );
  INV_X1 U13609 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10685) );
  INV_X1 U13610 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10683) );
  OAI22_X1 U13611 ( .A1(n10685), .A2(n10684), .B1(n10682), .B2(n10683), .ZN(
        n10686) );
  NOR2_X1 U13612 ( .A1(n10687), .A2(n10686), .ZN(n10690) );
  NAND2_X1 U13613 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10689) );
  NAND2_X1 U13614 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10688) );
  NAND4_X1 U13615 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .ZN(
        n10692) );
  AOI22_X1 U13616 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13617 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11464), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10696) );
  NAND2_X1 U13618 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10695) );
  NAND2_X1 U13619 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10694) );
  AOI22_X1 U13620 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11574), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13621 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11576), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10698) );
  NAND3_X1 U13622 ( .A1(n10700), .A2(n10699), .A3(n10698), .ZN(n10705) );
  AOI22_X1 U13623 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13624 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n11562), .ZN(n10702) );
  AOI22_X1 U13625 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10701) );
  NAND3_X1 U13626 ( .A1(n10703), .A2(n10702), .A3(n10701), .ZN(n10704) );
  INV_X1 U13627 ( .A(n10711), .ZN(n11132) );
  NAND2_X1 U13628 ( .A1(n11132), .A2(n9659), .ZN(n10706) );
  NAND2_X1 U13629 ( .A1(n10709), .A2(n10850), .ZN(n10710) );
  INV_X1 U13630 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12560) );
  MUX2_X1 U13631 ( .A(n10711), .B(n12560), .S(n11821), .Z(n10713) );
  OAI21_X1 U13632 ( .B1(n10712), .B2(n10713), .A(n10724), .ZN(n19364) );
  NAND2_X1 U13633 ( .A1(n10714), .A2(n19364), .ZN(n10715) );
  INV_X1 U13634 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15846) );
  AND2_X1 U13635 ( .A1(n10715), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10716) );
  MUX2_X1 U13636 ( .A(n10717), .B(P2_EBX_REG_7__SCAN_IN), .S(n11821), .Z(
        n10722) );
  NAND2_X2 U13637 ( .A1(n10582), .A2(n10720), .ZN(n10813) );
  INV_X1 U13638 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n19353) );
  NAND2_X1 U13639 ( .A1(n10720), .A2(n19353), .ZN(n10718) );
  NAND2_X1 U13640 ( .A1(n11007), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10719) );
  NOR2_X1 U13641 ( .A1(n10720), .A2(n10719), .ZN(n10721) );
  OR2_X1 U13642 ( .A1(n10731), .A2(n10721), .ZN(n19354) );
  NOR2_X1 U13643 ( .A1(n19354), .A2(n10717), .ZN(n10725) );
  NAND2_X1 U13644 ( .A1(n10725), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15598) );
  INV_X1 U13645 ( .A(n10722), .ZN(n10723) );
  XNOR2_X1 U13646 ( .A(n10724), .B(n10723), .ZN(n13313) );
  NAND2_X1 U13647 ( .A1(n13313), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15843) );
  AND2_X1 U13648 ( .A1(n15598), .A2(n15843), .ZN(n10729) );
  INV_X1 U13649 ( .A(n10725), .ZN(n10726) );
  INV_X1 U13650 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16685) );
  NAND2_X1 U13651 ( .A1(n10726), .A2(n16685), .ZN(n15597) );
  INV_X1 U13652 ( .A(n13313), .ZN(n10727) );
  INV_X1 U13653 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16682) );
  NAND2_X1 U13654 ( .A1(n10727), .A2(n16682), .ZN(n15842) );
  NAND2_X1 U13655 ( .A1(n11007), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10730) );
  XNOR2_X1 U13656 ( .A(n10731), .B(n10730), .ZN(n13333) );
  INV_X1 U13657 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15836) );
  OAI21_X1 U13658 ( .B1(n13333), .B2(n10717), .A(n15836), .ZN(n15829) );
  NAND2_X1 U13659 ( .A1(n11007), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10732) );
  INV_X1 U13660 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12471) );
  MUX2_X1 U13661 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n10732), .S(n10734), .Z(
        n10733) );
  NAND2_X1 U13662 ( .A1(n10733), .A2(n10813), .ZN(n19340) );
  NOR2_X1 U13663 ( .A1(n19340), .A2(n10717), .ZN(n10739) );
  NAND2_X1 U13664 ( .A1(n11007), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10735) );
  OR2_X1 U13665 ( .A1(n10736), .A2(n10735), .ZN(n10738) );
  INV_X1 U13666 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n15201) );
  NAND2_X2 U13667 ( .A1(n10813), .A2(n10741), .ZN(n10742) );
  INV_X1 U13668 ( .A(n10742), .ZN(n10737) );
  NAND2_X1 U13669 ( .A1(n10738), .A2(n10737), .ZN(n15209) );
  INV_X1 U13670 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10921) );
  OAI21_X1 U13671 ( .B1(n15209), .B2(n10717), .A(n10921), .ZN(n16626) );
  OR3_X1 U13672 ( .A1(n15209), .A2(n10717), .A3(n10921), .ZN(n16625) );
  OR3_X1 U13673 ( .A1(n13333), .A2(n10717), .A3(n15836), .ZN(n15828) );
  NAND2_X1 U13674 ( .A1(n10739), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15583) );
  NAND2_X1 U13675 ( .A1(n15828), .A2(n15583), .ZN(n16627) );
  INV_X1 U13676 ( .A(n16627), .ZN(n10740) );
  NAND2_X1 U13677 ( .A1(n16625), .A2(n10740), .ZN(n15569) );
  INV_X1 U13678 ( .A(n10741), .ZN(n10744) );
  NAND2_X1 U13679 ( .A1(n11007), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10743) );
  OAI21_X1 U13680 ( .B1(n10744), .B2(n10743), .A(n10748), .ZN(n13268) );
  NOR2_X1 U13681 ( .A1(n13268), .A2(n10717), .ZN(n10745) );
  AND2_X1 U13682 ( .A1(n10745), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15573) );
  NOR2_X1 U13683 ( .A1(n15569), .A2(n15573), .ZN(n15454) );
  OR2_X1 U13684 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n10745), .ZN(
        n15571) );
  INV_X1 U13685 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10785) );
  INV_X1 U13686 ( .A(n10747), .ZN(n10746) );
  XNOR2_X1 U13687 ( .A(n10748), .B(n10746), .ZN(n15184) );
  NAND2_X1 U13688 ( .A1(n15184), .A2(n11137), .ZN(n10786) );
  NAND2_X1 U13689 ( .A1(n10785), .A2(n10786), .ZN(n15558) );
  AND2_X1 U13690 ( .A1(n15571), .A2(n15558), .ZN(n15452) );
  AND2_X1 U13691 ( .A1(n11821), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10763) );
  INV_X1 U13692 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10940) );
  INV_X1 U13693 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U13694 ( .A1(n10940), .A2(n10936), .ZN(n10749) );
  AND2_X1 U13695 ( .A1(n11821), .A2(n10749), .ZN(n10750) );
  OR2_X2 U13696 ( .A1(n10760), .A2(n10750), .ZN(n10761) );
  AND2_X1 U13697 ( .A1(n11821), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10757) );
  OR2_X2 U13698 ( .A1(n10761), .A2(n10757), .ZN(n10759) );
  AND2_X1 U13699 ( .A1(n11821), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10755) );
  INV_X1 U13700 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10951) );
  OR2_X1 U13701 ( .A1(n10793), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10754) );
  NAND2_X1 U13702 ( .A1(n10793), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10751) );
  OAI21_X1 U13703 ( .B1(n10751), .B2(n10582), .A(n10813), .ZN(n10752) );
  INV_X1 U13704 ( .A(n10752), .ZN(n10753) );
  INV_X1 U13705 ( .A(n10717), .ZN(n11137) );
  AOI21_X1 U13706 ( .B1(n10776), .B2(n11137), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15467) );
  AND2_X1 U13707 ( .A1(n10759), .A2(n10755), .ZN(n10756) );
  INV_X1 U13708 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15707) );
  OAI21_X2 U13709 ( .B1(n15157), .B2(n10717), .A(n15707), .ZN(n15489) );
  NAND2_X1 U13710 ( .A1(n10761), .A2(n10757), .ZN(n10758) );
  NAND2_X1 U13711 ( .A1(n10759), .A2(n10758), .ZN(n19305) );
  INV_X1 U13712 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11366) );
  NAND2_X1 U13713 ( .A1(n10789), .A2(n11366), .ZN(n15500) );
  NAND2_X1 U13714 ( .A1(n15489), .A2(n15500), .ZN(n15463) );
  AND2_X1 U13715 ( .A1(n10760), .A2(n11137), .ZN(n10783) );
  NOR2_X1 U13716 ( .A1(n10783), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15456) );
  OR2_X1 U13717 ( .A1(n10760), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10767) );
  NAND3_X1 U13718 ( .A1(n10767), .A2(P2_EBX_REG_17__SCAN_IN), .A3(n11821), 
        .ZN(n10762) );
  AND2_X1 U13719 ( .A1(n10762), .A2(n10761), .ZN(n10782) );
  AOI21_X1 U13720 ( .B1(n10782), .B2(n11137), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15460) );
  AND2_X1 U13721 ( .A1(n10764), .A2(n10763), .ZN(n10765) );
  OR2_X1 U13722 ( .A1(n15178), .A2(n10765), .ZN(n19332) );
  INV_X1 U13723 ( .A(n19332), .ZN(n10788) );
  AOI21_X1 U13724 ( .B1(n10788), .B2(n11137), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15533) );
  NAND3_X1 U13725 ( .A1(n10760), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n11821), 
        .ZN(n10766) );
  NAND3_X1 U13726 ( .A1(n10767), .A2(n10813), .A3(n10766), .ZN(n19316) );
  OR2_X1 U13727 ( .A1(n19316), .A2(n10717), .ZN(n10768) );
  XNOR2_X1 U13728 ( .A(n10768), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15523) );
  NAND2_X1 U13729 ( .A1(n10769), .A2(n15523), .ZN(n10773) );
  INV_X1 U13730 ( .A(n10770), .ZN(n10772) );
  NAND2_X1 U13731 ( .A1(n11007), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10771) );
  XNOR2_X1 U13732 ( .A(n10772), .B(n10771), .ZN(n19295) );
  AOI21_X1 U13733 ( .B1(n19295), .B2(n11137), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15477) );
  NOR3_X1 U13734 ( .A1(n15467), .A2(n10773), .A3(n15477), .ZN(n10774) );
  INV_X1 U13735 ( .A(n10774), .ZN(n10775) );
  INV_X1 U13736 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10777) );
  OR2_X1 U13737 ( .A1(n10717), .A2(n10777), .ZN(n10778) );
  NOR2_X1 U13738 ( .A1(n15141), .A2(n10778), .ZN(n15466) );
  INV_X1 U13739 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15708) );
  NOR2_X1 U13740 ( .A1(n10717), .A2(n15708), .ZN(n10779) );
  INV_X1 U13741 ( .A(n15157), .ZN(n10781) );
  NOR2_X1 U13742 ( .A1(n10717), .A2(n15707), .ZN(n10780) );
  NAND2_X1 U13743 ( .A1(n10781), .A2(n10780), .ZN(n15488) );
  INV_X1 U13744 ( .A(n10782), .ZN(n15167) );
  INV_X1 U13745 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15754) );
  OR3_X1 U13746 ( .A1(n15167), .A2(n10717), .A3(n15754), .ZN(n15461) );
  INV_X1 U13747 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15764) );
  OR3_X1 U13748 ( .A1(n19316), .A2(n10717), .A3(n15764), .ZN(n15458) );
  AND2_X1 U13749 ( .A1(n15461), .A2(n15458), .ZN(n10791) );
  INV_X1 U13750 ( .A(n10783), .ZN(n10784) );
  INV_X1 U13751 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15511) );
  OR2_X1 U13752 ( .A1(n10784), .A2(n15511), .ZN(n15534) );
  OR2_X1 U13753 ( .A1(n10786), .A2(n10785), .ZN(n15559) );
  INV_X1 U13754 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15552) );
  NOR2_X1 U13755 ( .A1(n10717), .A2(n15552), .ZN(n10787) );
  NAND2_X1 U13756 ( .A1(n10788), .A2(n10787), .ZN(n15531) );
  AND3_X1 U13757 ( .A1(n15534), .A2(n15559), .A3(n15531), .ZN(n15453) );
  INV_X1 U13758 ( .A(n10789), .ZN(n10790) );
  NAND2_X1 U13759 ( .A1(n10790), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15501) );
  NAND4_X1 U13760 ( .A1(n15488), .A2(n10791), .A3(n15453), .A4(n15501), .ZN(
        n10792) );
  NAND2_X1 U13761 ( .A1(n11007), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10794) );
  INV_X1 U13762 ( .A(n10794), .ZN(n10797) );
  NAND2_X1 U13763 ( .A1(n10813), .A2(n10249), .ZN(n10795) );
  INV_X1 U13764 ( .A(n10799), .ZN(n10796) );
  AOI21_X1 U13765 ( .B1(n10797), .B2(n10249), .A(n10796), .ZN(n15125) );
  AOI21_X1 U13766 ( .B1(n15125), .B2(n11137), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15443) );
  NAND3_X1 U13767 ( .A1(n15125), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11137), .ZN(n15441) );
  AND2_X1 U13768 ( .A1(n11821), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U13769 ( .A1(n10799), .A2(n10798), .ZN(n10800) );
  NAND2_X1 U13770 ( .A1(n10804), .A2(n10800), .ZN(n15114) );
  OR2_X1 U13771 ( .A1(n15114), .A2(n10717), .ZN(n10801) );
  XNOR2_X1 U13772 ( .A(n10801), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15435) );
  INV_X1 U13773 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15671) );
  NOR3_X1 U13774 ( .A1(n15114), .A2(n10717), .A3(n15671), .ZN(n10802) );
  INV_X1 U13775 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10803) );
  NAND3_X1 U13776 ( .A1(n10804), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n11007), 
        .ZN(n10805) );
  NAND3_X1 U13777 ( .A1(n10807), .A2(n10813), .A3(n10805), .ZN(n16599) );
  NOR2_X1 U13778 ( .A1(n16599), .A2(n10717), .ZN(n15422) );
  NAND3_X1 U13779 ( .A1(n10807), .A2(P2_EBX_REG_25__SCAN_IN), .A3(n11007), 
        .ZN(n10808) );
  NAND2_X1 U13780 ( .A1(n10808), .A2(n10813), .ZN(n10809) );
  NOR2_X1 U13781 ( .A1(n10812), .A2(n10809), .ZN(n16587) );
  AOI21_X1 U13782 ( .B1(n16587), .B2(n11137), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15411) );
  NAND2_X1 U13783 ( .A1(n11007), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10810) );
  OR2_X1 U13784 ( .A1(n10812), .A2(n10810), .ZN(n10814) );
  INV_X1 U13785 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10811) );
  NAND2_X1 U13786 ( .A1(n16576), .A2(n11137), .ZN(n10819) );
  XNOR2_X1 U13787 ( .A(n10819), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15403) );
  NAND2_X1 U13788 ( .A1(n11007), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10816) );
  NAND3_X1 U13789 ( .A1(n11821), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n10817), 
        .ZN(n10818) );
  NAND2_X1 U13790 ( .A1(n10998), .A2(n10818), .ZN(n16563) );
  NOR2_X2 U13791 ( .A1(n10990), .A2(n10825), .ZN(n10993) );
  INV_X1 U13792 ( .A(n10993), .ZN(n10824) );
  NAND2_X1 U13793 ( .A1(n10990), .A2(n10825), .ZN(n10823) );
  INV_X1 U13794 ( .A(n10819), .ZN(n10822) );
  INV_X1 U13795 ( .A(n16587), .ZN(n10821) );
  INV_X1 U13796 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15648) );
  OR2_X1 U13797 ( .A1(n10717), .A2(n15648), .ZN(n10820) );
  NOR2_X1 U13798 ( .A1(n10821), .A2(n10820), .ZN(n15410) );
  AOI21_X1 U13799 ( .B1(n10822), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15410), .ZN(n10994) );
  INV_X1 U13800 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15626) );
  AOI21_X1 U13801 ( .B1(n10990), .B2(n10994), .A(n10825), .ZN(n10826) );
  NAND2_X1 U13802 ( .A1(n11007), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10996) );
  XNOR2_X1 U13803 ( .A(n10998), .B(n10996), .ZN(n16551) );
  XOR2_X1 U13804 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n10992), .Z(
        n10827) );
  INV_X1 U13805 ( .A(n11038), .ZN(n10828) );
  NAND2_X1 U13806 ( .A1(n10829), .A2(n10828), .ZN(n10831) );
  NAND2_X1 U13807 ( .A1(n10831), .A2(n10830), .ZN(n10832) );
  AND3_X1 U13808 ( .A1(n10834), .A2(n10833), .A3(n10832), .ZN(n10837) );
  NOR2_X1 U13809 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16209), .ZN(
        n10835) );
  OR2_X1 U13810 ( .A1(n10837), .A2(n11053), .ZN(n16713) );
  AND2_X1 U13811 ( .A1(n9659), .A2(n20279), .ZN(n11064) );
  INV_X1 U13812 ( .A(n11064), .ZN(n11088) );
  NOR2_X1 U13813 ( .A1(n16713), .A2(n11088), .ZN(n11060) );
  INV_X1 U13814 ( .A(n11089), .ZN(n11081) );
  NAND2_X1 U13815 ( .A1(n11060), .A2(n11081), .ZN(n10848) );
  NOR2_X1 U13816 ( .A1(n11089), .A2(n13262), .ZN(n11087) );
  NAND2_X1 U13817 ( .A1(n15907), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10838) );
  NAND2_X1 U13818 ( .A1(n10838), .A2(n20221), .ZN(n16722) );
  OR2_X1 U13819 ( .A1(n11564), .A2(n16722), .ZN(n10839) );
  INV_X1 U13820 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19276) );
  NAND2_X1 U13821 ( .A1(n10839), .A2(n19276), .ZN(n20259) );
  NAND2_X1 U13822 ( .A1(n10841), .A2(n10840), .ZN(n11048) );
  NOR2_X1 U13823 ( .A1(n11048), .A2(n11044), .ZN(n10845) );
  INV_X1 U13824 ( .A(n10842), .ZN(n10843) );
  XNOR2_X1 U13825 ( .A(n11038), .B(n10843), .ZN(n11040) );
  AND2_X1 U13826 ( .A1(n11040), .A2(n10845), .ZN(n10844) );
  OR2_X1 U13827 ( .A1(n11053), .A2(n10844), .ZN(n16725) );
  AOI21_X1 U13828 ( .B1(n11041), .B2(n10845), .A(n16725), .ZN(n10846) );
  MUX2_X1 U13829 ( .A(n20259), .B(n10846), .S(n15859), .Z(n16753) );
  NAND2_X1 U13830 ( .A1(n11087), .A2(n16753), .ZN(n10847) );
  NAND2_X1 U13831 ( .A1(n10848), .A2(n10847), .ZN(n16731) );
  AND2_X1 U13832 ( .A1(n15859), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U13833 ( .A1(n11394), .A2(n16662), .ZN(n10989) );
  NAND2_X1 U13834 ( .A1(n10866), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10869) );
  INV_X1 U13835 ( .A(n10869), .ZN(n13446) );
  NAND2_X1 U13836 ( .A1(n13446), .A2(n10850), .ZN(n13588) );
  INV_X1 U13837 ( .A(n12035), .ZN(n10852) );
  NAND2_X1 U13838 ( .A1(n10852), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12037) );
  INV_X1 U13839 ( .A(n12037), .ZN(n10853) );
  XNOR2_X1 U13840 ( .A(n11095), .B(n11108), .ZN(n10854) );
  NAND2_X1 U13841 ( .A1(n10853), .A2(n10854), .ZN(n10855) );
  XNOR2_X1 U13842 ( .A(n12037), .B(n10854), .ZN(n11854) );
  NAND2_X1 U13843 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n11854), .ZN(
        n11855) );
  NAND2_X1 U13844 ( .A1(n10855), .A2(n11855), .ZN(n10857) );
  XOR2_X1 U13845 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10857), .Z(
        n12078) );
  XOR2_X1 U13846 ( .A(n11112), .B(n10856), .Z(n12077) );
  NAND2_X1 U13847 ( .A1(n12078), .A2(n12077), .ZN(n12076) );
  NAND2_X1 U13848 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10857), .ZN(
        n10858) );
  NAND2_X1 U13849 ( .A1(n12076), .A2(n10858), .ZN(n10859) );
  XNOR2_X1 U13850 ( .A(n10859), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13145) );
  INV_X1 U13851 ( .A(n11126), .ZN(n10860) );
  INV_X1 U13852 ( .A(n10862), .ZN(n10864) );
  OR2_X1 U13853 ( .A1(n10864), .A2(n10863), .ZN(n10865) );
  INV_X1 U13854 ( .A(n10866), .ZN(n10867) );
  NAND2_X1 U13855 ( .A1(n10868), .A2(n10869), .ZN(n10870) );
  AOI21_X2 U13856 ( .B1(n10873), .B2(n13589), .A(n10872), .ZN(n10879) );
  NAND2_X1 U13857 ( .A1(n10874), .A2(n10717), .ZN(n10876) );
  NAND2_X1 U13858 ( .A1(n10881), .A2(n10876), .ZN(n10877) );
  XNOR2_X1 U13859 ( .A(n10879), .B(n10877), .ZN(n15840) );
  INV_X1 U13860 ( .A(n10877), .ZN(n10878) );
  NAND2_X1 U13861 ( .A1(n10879), .A2(n10878), .ZN(n10880) );
  INV_X1 U13862 ( .A(n10881), .ZN(n10882) );
  NAND2_X1 U13863 ( .A1(n10882), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10883) );
  NAND2_X1 U13864 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15785) );
  NOR2_X1 U13865 ( .A1(n15785), .A2(n15552), .ZN(n10884) );
  AND3_X1 U13866 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15778) );
  NAND2_X1 U13867 ( .A1(n10884), .A2(n15778), .ZN(n15750) );
  INV_X1 U13868 ( .A(n15750), .ZN(n11368) );
  AND2_X1 U13869 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15751) );
  NAND2_X1 U13870 ( .A1(n15751), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15726) );
  INV_X1 U13871 ( .A(n15726), .ZN(n10885) );
  NAND2_X1 U13872 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15694) );
  NAND2_X1 U13873 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15665) );
  OAI21_X1 U13874 ( .B1(n10887), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15380), .ZN(n11404) );
  NAND2_X1 U13875 ( .A1(n10977), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10895) );
  NAND2_X1 U13876 ( .A1(n9678), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10892) );
  NAND2_X1 U13877 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10891) );
  OAI211_X1 U13878 ( .C1(n19353), .C2(n10408), .A(n10892), .B(n10891), .ZN(
        n10893) );
  INV_X1 U13879 ( .A(n10893), .ZN(n10894) );
  NAND2_X1 U13880 ( .A1(n10895), .A2(n10894), .ZN(n12836) );
  INV_X1 U13881 ( .A(n10897), .ZN(n10899) );
  NAND2_X1 U13882 ( .A1(n10899), .A2(n10898), .ZN(n10900) );
  NAND2_X1 U13883 ( .A1(n10901), .A2(n10900), .ZN(n12371) );
  OR2_X1 U13884 ( .A1(n11021), .A2(n13422), .ZN(n10905) );
  AOI22_X1 U13885 ( .A1(n10942), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10904) );
  NAND2_X1 U13886 ( .A1(n10889), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10903) );
  OR2_X1 U13887 ( .A1(n11021), .A2(n13455), .ZN(n10908) );
  AOI22_X1 U13888 ( .A1(n10942), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10907) );
  NAND2_X1 U13889 ( .A1(n10889), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13890 ( .A1(n10942), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10910) );
  NAND2_X1 U13891 ( .A1(n10889), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10909) );
  OAI211_X1 U13892 ( .C1(n11021), .C2(n15846), .A(n10910), .B(n10909), .ZN(
        n12556) );
  AOI22_X1 U13893 ( .A1(n10942), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10912) );
  NAND2_X1 U13894 ( .A1(n10889), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10911) );
  OAI211_X1 U13895 ( .C1(n11021), .C2(n16682), .A(n10912), .B(n10911), .ZN(
        n12568) );
  NAND2_X1 U13896 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  NAND2_X1 U13897 ( .A1(n10942), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U13898 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10913) );
  OAI211_X1 U13899 ( .C1(n12471), .C2(n10408), .A(n10914), .B(n10913), .ZN(
        n10915) );
  AOI21_X1 U13900 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10915), .ZN(n12469) );
  INV_X1 U13901 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19339) );
  NAND2_X1 U13902 ( .A1(n9678), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U13903 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10916) );
  OAI211_X1 U13904 ( .C1(n19339), .C2(n9677), .A(n10917), .B(n10916), .ZN(
        n10918) );
  AOI21_X1 U13905 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10918), .ZN(n12563) );
  NOR2_X2 U13906 ( .A1(n12564), .A2(n12563), .ZN(n12651) );
  AOI22_X1 U13907 ( .A1(n10942), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10920) );
  NAND2_X1 U13908 ( .A1(n10889), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10919) );
  OAI211_X1 U13909 ( .C1(n11021), .C2(n10921), .A(n10920), .B(n10919), .ZN(
        n12650) );
  NAND2_X1 U13910 ( .A1(n12651), .A2(n12650), .ZN(n12827) );
  INV_X1 U13911 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U13912 ( .A1(n9678), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U13913 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10922) );
  OAI211_X1 U13914 ( .C1(n10924), .C2(n10408), .A(n10923), .B(n10922), .ZN(
        n10925) );
  AOI21_X1 U13915 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10925), .ZN(n12826) );
  INV_X1 U13916 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10928) );
  NAND2_X1 U13917 ( .A1(n10942), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U13918 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10926) );
  OAI211_X1 U13919 ( .C1(n10928), .C2(n10408), .A(n10927), .B(n10926), .ZN(
        n10929) );
  AOI21_X1 U13920 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10929), .ZN(n13093) );
  AOI22_X1 U13921 ( .A1(n10942), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10931) );
  NAND2_X1 U13922 ( .A1(n10889), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10930) );
  OAI211_X1 U13923 ( .C1(n11021), .C2(n15552), .A(n10931), .B(n10930), .ZN(
        n12976) );
  AOI22_X1 U13924 ( .A1(n10942), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10933) );
  NAND2_X1 U13925 ( .A1(n10889), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10932) );
  OAI211_X1 U13926 ( .C1(n11021), .C2(n15511), .A(n10933), .B(n10932), .ZN(
        n13299) );
  NAND2_X1 U13927 ( .A1(n9678), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U13928 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10934) );
  OAI211_X1 U13929 ( .C1(n10936), .C2(n9677), .A(n10935), .B(n10934), .ZN(
        n10937) );
  AOI21_X1 U13930 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10937), .ZN(n13397) );
  NAND2_X1 U13931 ( .A1(n10942), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10939) );
  NAND2_X1 U13932 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10938) );
  OAI211_X1 U13933 ( .C1(n10940), .C2(n10408), .A(n10939), .B(n10938), .ZN(
        n10941) );
  AOI21_X1 U13934 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10941), .ZN(n13440) );
  INV_X1 U13935 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U13936 ( .A1(n9678), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U13937 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10943) );
  OAI211_X1 U13938 ( .C1(n10945), .C2(n9677), .A(n10944), .B(n10943), .ZN(
        n10946) );
  AOI21_X1 U13939 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10946), .ZN(n13667) );
  AOI22_X1 U13940 ( .A1(n9678), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10948) );
  NAND2_X1 U13941 ( .A1(n10889), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10947) );
  OAI211_X1 U13942 ( .C1(n11021), .C2(n15707), .A(n10948), .B(n10947), .ZN(
        n15150) );
  NAND2_X1 U13943 ( .A1(n10942), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U13944 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10949) );
  OAI211_X1 U13945 ( .C1(n10951), .C2(n10408), .A(n10950), .B(n10949), .ZN(
        n10952) );
  AOI21_X1 U13946 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10952), .ZN(n15290) );
  OR2_X2 U13947 ( .A1(n15289), .A2(n15290), .ZN(n15287) );
  INV_X1 U13948 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10955) );
  NAND2_X1 U13949 ( .A1(n9678), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U13950 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10953) );
  OAI211_X1 U13951 ( .C1(n10955), .C2(n10408), .A(n10954), .B(n10953), .ZN(
        n10956) );
  AOI21_X1 U13952 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10956), .ZN(n15130) );
  NOR2_X2 U13953 ( .A1(n15287), .A2(n15130), .ZN(n15132) );
  INV_X1 U13954 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U13955 ( .A1(n9678), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10958) );
  NAND2_X1 U13956 ( .A1(n10889), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10957) );
  OAI211_X1 U13957 ( .C1(n11021), .C2(n15431), .A(n10958), .B(n10957), .ZN(
        n15115) );
  AND2_X2 U13958 ( .A1(n15132), .A2(n15115), .ZN(n15117) );
  AOI22_X1 U13959 ( .A1(n9678), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10960) );
  NAND2_X1 U13960 ( .A1(n10889), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10959) );
  OAI211_X1 U13961 ( .C1(n11021), .C2(n15671), .A(n10960), .B(n10959), .ZN(
        n15080) );
  NAND2_X1 U13962 ( .A1(n9678), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U13963 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10961) );
  OAI211_X1 U13964 ( .C1(n10017), .C2(n9677), .A(n10962), .B(n10961), .ZN(
        n10963) );
  AOI21_X1 U13965 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10963), .ZN(n15263) );
  INV_X1 U13966 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U13967 ( .A1(n9678), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10965) );
  NAND2_X1 U13968 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10964) );
  OAI211_X1 U13969 ( .C1(n10966), .C2(n10408), .A(n10965), .B(n10964), .ZN(
        n10967) );
  AOI21_X1 U13970 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10967), .ZN(n15254) );
  INV_X1 U13971 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15633) );
  AOI22_X1 U13972 ( .A1(n10942), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10969) );
  NAND2_X1 U13973 ( .A1(n10889), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10968) );
  OAI211_X1 U13974 ( .C1(n11021), .C2(n15633), .A(n10969), .B(n10968), .ZN(
        n15248) );
  INV_X1 U13975 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16562) );
  NAND2_X1 U13976 ( .A1(n9678), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10971) );
  NAND2_X1 U13977 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10970) );
  OAI211_X1 U13978 ( .C1(n16562), .C2(n9677), .A(n10971), .B(n10970), .ZN(
        n10972) );
  AOI21_X1 U13979 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10972), .ZN(n15239) );
  OR2_X2 U13980 ( .A1(n15247), .A2(n15239), .ZN(n15241) );
  INV_X1 U13981 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U13982 ( .A1(n10942), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U13983 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10973) );
  OAI211_X1 U13984 ( .C1(n10975), .C2(n10408), .A(n10974), .B(n10973), .ZN(
        n10976) );
  AOI21_X1 U13985 ( .B1(n10977), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10976), .ZN(n10978) );
  NOR2_X2 U13986 ( .A1(n15241), .A2(n10978), .ZN(n15223) );
  AND2_X1 U13987 ( .A1(n15241), .A2(n10978), .ZN(n10979) );
  OR2_X1 U13988 ( .A1(n15223), .A2(n10979), .ZN(n16553) );
  INV_X1 U13989 ( .A(n16553), .ZN(n11402) );
  NOR2_X1 U13990 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20219) );
  OR2_X1 U13991 ( .A1(n20223), .A2(n20219), .ZN(n20254) );
  NAND2_X1 U13992 ( .A1(n20254), .A2(n20278), .ZN(n10980) );
  AND2_X1 U13993 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16203) );
  INV_X1 U13994 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10984) );
  INV_X1 U13995 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19952) );
  NAND2_X1 U13996 ( .A1(n19952), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10981) );
  NAND2_X1 U13997 ( .A1(n10216), .A2(n10981), .ZN(n12040) );
  INV_X1 U13998 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15515) );
  NAND2_X1 U13999 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13157) );
  INV_X1 U14000 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15494) );
  INV_X1 U14001 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15089) );
  INV_X1 U14002 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U14003 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n15414), .ZN(
        n15405) );
  OAI21_X1 U14004 ( .B1(n15393), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15381), .ZN(n16557) );
  INV_X1 U14005 ( .A(n16557), .ZN(n10982) );
  NAND2_X1 U14006 ( .A1(n16658), .A2(n10982), .ZN(n10983) );
  NAND2_X1 U14007 ( .A1(n20223), .A2(n15859), .ZN(n19270) );
  INV_X2 U14008 ( .A(n15727), .ZN(n19529) );
  INV_X1 U14009 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20199) );
  OR2_X1 U14010 ( .A1(n19363), .A2(n20199), .ZN(n11397) );
  OAI211_X1 U14011 ( .C1(n16666), .C2(n10984), .A(n10983), .B(n11397), .ZN(
        n10985) );
  AOI21_X1 U14012 ( .B1(n11402), .B2(n19538), .A(n10985), .ZN(n10986) );
  NAND2_X1 U14013 ( .A1(n10989), .A2(n10988), .ZN(P2_U2986) );
  INV_X1 U14014 ( .A(n10990), .ZN(n10991) );
  INV_X1 U14015 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10995) );
  INV_X1 U14016 ( .A(n10996), .ZN(n10997) );
  NAND2_X1 U14017 ( .A1(n11007), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11000) );
  XNOR2_X1 U14018 ( .A(n10999), .B(n11000), .ZN(n11003) );
  INV_X1 U14019 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15611) );
  OAI21_X1 U14020 ( .B1(n11003), .B2(n10717), .A(n15611), .ZN(n15375) );
  NAND2_X1 U14021 ( .A1(n11007), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11001) );
  XNOR2_X1 U14022 ( .A(n11004), .B(n11001), .ZN(n16529) );
  AOI21_X1 U14023 ( .B1(n16529), .B2(n11137), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11032) );
  INV_X1 U14024 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11416) );
  NOR2_X1 U14025 ( .A1(n10717), .A2(n11416), .ZN(n11002) );
  NAND2_X1 U14026 ( .A1(n16529), .A2(n11002), .ZN(n11033) );
  INV_X1 U14027 ( .A(n11003), .ZN(n16540) );
  NAND3_X1 U14028 ( .A1(n16540), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11137), .ZN(n15376) );
  INV_X1 U14029 ( .A(n11004), .ZN(n11006) );
  INV_X1 U14030 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11005) );
  NAND2_X1 U14031 ( .A1(n11006), .A2(n11005), .ZN(n11008) );
  MUX2_X1 U14032 ( .A(n11009), .B(n11008), .S(n11007), .Z(n16518) );
  NOR2_X1 U14033 ( .A1(n16518), .A2(n10717), .ZN(n11010) );
  XOR2_X1 U14034 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11010), .Z(
        n11011) );
  XNOR2_X1 U14035 ( .A(n11012), .B(n11011), .ZN(n11422) );
  AOI22_X1 U14036 ( .A1(n9678), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11015) );
  NAND2_X1 U14037 ( .A1(n10889), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11014) );
  OAI211_X1 U14038 ( .C1(n11021), .C2(n15611), .A(n11015), .B(n11014), .ZN(
        n15222) );
  NAND2_X1 U14039 ( .A1(n15223), .A2(n15222), .ZN(n15225) );
  INV_X1 U14040 ( .A(n15225), .ZN(n11018) );
  AOI22_X1 U14041 ( .A1(n10942), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11017) );
  NAND2_X1 U14042 ( .A1(n10889), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11016) );
  OAI211_X1 U14043 ( .C1(n11021), .C2(n11416), .A(n11017), .B(n11016), .ZN(
        n11341) );
  NAND2_X1 U14044 ( .A1(n11018), .A2(n11341), .ZN(n11023) );
  INV_X1 U14045 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U14046 ( .A1(n9678), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11020) );
  NAND2_X1 U14047 ( .A1(n10889), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11019) );
  OAI211_X1 U14048 ( .C1(n11021), .C2(n13235), .A(n11020), .B(n11019), .ZN(
        n11022) );
  INV_X1 U14049 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15384) );
  NAND2_X1 U14050 ( .A1(n19529), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11414) );
  NAND2_X1 U14051 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11026) );
  OAI211_X1 U14052 ( .C1(n19542), .C2(n13234), .A(n11414), .B(n11026), .ZN(
        n11027) );
  INV_X1 U14053 ( .A(n11029), .ZN(n11030) );
  OAI21_X1 U14054 ( .B1(n11422), .B2(n19534), .A(n11030), .ZN(P2_U2983) );
  NAND2_X1 U14055 ( .A1(n11031), .A2(n15376), .ZN(n11035) );
  NAND2_X1 U14056 ( .A1(n10126), .A2(n11033), .ZN(n11034) );
  INV_X1 U14057 ( .A(n11053), .ZN(n11051) );
  NAND2_X1 U14058 ( .A1(n20277), .A2(n20281), .ZN(n11036) );
  MUX2_X1 U14059 ( .A(n13262), .B(n11036), .S(n11044), .Z(n11047) );
  OAI21_X1 U14060 ( .B1(n11039), .B2(n11038), .A(n11037), .ZN(n11043) );
  OAI211_X1 U14061 ( .C1(n20281), .C2(n11041), .A(n11070), .B(n11040), .ZN(
        n11042) );
  OAI211_X1 U14062 ( .C1(n11045), .C2(n11044), .A(n11043), .B(n11042), .ZN(
        n11046) );
  NAND2_X1 U14063 ( .A1(n11047), .A2(n11046), .ZN(n11049) );
  MUX2_X1 U14064 ( .A(n11049), .B(n13262), .S(n11048), .Z(n11050) );
  NAND2_X1 U14065 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  MUX2_X1 U14066 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11052), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11056) );
  NAND2_X1 U14067 ( .A1(n11053), .A2(n12245), .ZN(n11054) );
  NOR2_X1 U14068 ( .A1(n11830), .A2(n9659), .ZN(n12242) );
  NAND2_X1 U14069 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20276) );
  INV_X1 U14070 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20130) );
  NOR2_X1 U14071 ( .A1(n20130), .A2(n20149), .ZN(n20141) );
  NOR2_X1 U14072 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20143) );
  NOR3_X1 U14073 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20141), .A3(n20143), 
        .ZN(n20280) );
  NAND2_X1 U14074 ( .A1(n20276), .A2(n20280), .ZN(n16729) );
  INV_X1 U14075 ( .A(n16729), .ZN(n11055) );
  NAND3_X1 U14076 ( .A1(n12242), .A2(n11350), .A3(n11055), .ZN(n11085) );
  INV_X1 U14077 ( .A(n12242), .ZN(n11058) );
  AOI21_X1 U14078 ( .B1(n11056), .B2(n11070), .A(n11352), .ZN(n11057) );
  NAND2_X1 U14079 ( .A1(n11058), .A2(n11057), .ZN(n11084) );
  INV_X1 U14080 ( .A(n16753), .ZN(n16208) );
  NOR2_X1 U14081 ( .A1(n16208), .A2(n9659), .ZN(n11059) );
  OR2_X1 U14082 ( .A1(n11060), .A2(n11059), .ZN(n11082) );
  MUX2_X1 U14083 ( .A(n11077), .B(n11350), .S(n9659), .Z(n11061) );
  NAND2_X1 U14084 ( .A1(n11061), .A2(n20276), .ZN(n11079) );
  AND2_X1 U14085 ( .A1(n11063), .A2(n11062), .ZN(n11075) );
  OAI21_X1 U14086 ( .B1(n11065), .B2(n19590), .A(n11064), .ZN(n11360) );
  NAND2_X1 U14087 ( .A1(n11067), .A2(n19564), .ZN(n11068) );
  NAND2_X1 U14088 ( .A1(n11066), .A2(n11068), .ZN(n11074) );
  NAND2_X1 U14089 ( .A1(n11069), .A2(n9659), .ZN(n11345) );
  NAND2_X1 U14090 ( .A1(n11345), .A2(n11070), .ZN(n11071) );
  NAND2_X1 U14091 ( .A1(n11071), .A2(n10102), .ZN(n11072) );
  NAND2_X1 U14092 ( .A1(n11072), .A2(n19564), .ZN(n11073) );
  NAND4_X1 U14093 ( .A1(n11075), .A2(n11360), .A3(n11074), .A4(n11073), .ZN(
        n11346) );
  NOR2_X1 U14094 ( .A1(n16725), .A2(n16729), .ZN(n11076) );
  AND2_X1 U14095 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  NOR2_X1 U14096 ( .A1(n11346), .A2(n11078), .ZN(n15864) );
  OAI21_X1 U14097 ( .B1(n16725), .B2(n11079), .A(n15864), .ZN(n11080) );
  AOI21_X1 U14098 ( .B1(n11082), .B2(n11081), .A(n11080), .ZN(n11083) );
  NAND3_X1 U14099 ( .A1(n11085), .A2(n11084), .A3(n11083), .ZN(n11086) );
  INV_X1 U14100 ( .A(n11087), .ZN(n16716) );
  NAND2_X1 U14101 ( .A1(n11385), .A2(n16673), .ZN(n11384) );
  XNOR2_X1 U14102 ( .A(n15379), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11390) );
  OR2_X1 U14103 ( .A1(n11089), .A2(n11088), .ZN(n16711) );
  NOR2_X1 U14104 ( .A1(n9659), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11097) );
  NOR2_X1 U14105 ( .A1(n19590), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U14106 ( .A1(n11236), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11093) );
  INV_X2 U14107 ( .A(n9717), .ZN(n11410) );
  NAND2_X1 U14108 ( .A1(n11410), .A2(P2_EAX_REG_30__SCAN_IN), .ZN(n11092) );
  OAI211_X1 U14109 ( .C1(n11416), .C2(n11335), .A(n11093), .B(n11092), .ZN(
        n11408) );
  AOI222_X1 U14110 ( .A1(n11236), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n11328), 
        .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n11410), .C2(
        P2_EAX_REG_7__SCAN_IN), .ZN(n13305) );
  NOR2_X1 U14111 ( .A1(n11821), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11094) );
  INV_X1 U14112 ( .A(n11096), .ZN(n11811) );
  NAND2_X1 U14113 ( .A1(n11097), .A2(n11811), .ZN(n11113) );
  AND2_X1 U14114 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11098) );
  NOR2_X1 U14115 ( .A1(n11410), .A2(n11098), .ZN(n11099) );
  NAND2_X1 U14116 ( .A1(n11236), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11103) );
  INV_X1 U14117 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16706) );
  NAND2_X1 U14118 ( .A1(n19590), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11100) );
  OAI211_X1 U14119 ( .C1(n9659), .C2(n16706), .A(n11100), .B(n20268), .ZN(
        n11101) );
  INV_X1 U14120 ( .A(n11101), .ZN(n11102) );
  NAND2_X1 U14121 ( .A1(n11103), .A2(n11102), .ZN(n16698) );
  AOI22_X1 U14122 ( .A1(n11097), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14123 ( .A1(n11236), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11104) );
  AND2_X1 U14124 ( .A1(n11105), .A2(n11104), .ZN(n11110) );
  XNOR2_X1 U14125 ( .A(n11109), .B(n11110), .ZN(n11858) );
  NAND2_X1 U14126 ( .A1(n11096), .A2(n10102), .ZN(n11106) );
  MUX2_X1 U14127 ( .A(n11106), .B(n20252), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11107) );
  OAI21_X1 U14128 ( .B1(n11108), .B2(n11301), .A(n11107), .ZN(n11857) );
  NAND2_X1 U14129 ( .A1(n11110), .A2(n11109), .ZN(n11111) );
  NAND2_X1 U14130 ( .A1(n11860), .A2(n11111), .ZN(n11118) );
  OR2_X1 U14131 ( .A1(n11301), .A2(n11112), .ZN(n11114) );
  OAI211_X1 U14132 ( .C1(n20268), .C2(n20243), .A(n11114), .B(n11113), .ZN(
        n11117) );
  XNOR2_X1 U14133 ( .A(n11118), .B(n11117), .ZN(n12109) );
  AOI22_X1 U14134 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n11116) );
  NAND2_X1 U14135 ( .A1(n11236), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11115) );
  AND2_X1 U14136 ( .A1(n11116), .A2(n11115), .ZN(n12108) );
  INV_X1 U14137 ( .A(n11117), .ZN(n11119) );
  NAND2_X1 U14138 ( .A1(n11119), .A2(n11118), .ZN(n11120) );
  AOI22_X1 U14139 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11125) );
  NAND2_X1 U14140 ( .A1(n11236), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U14141 ( .A1(n11410), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11123) );
  OR2_X1 U14142 ( .A1(n11301), .A2(n11121), .ZN(n11122) );
  NOR2_X2 U14143 ( .A1(n13150), .A2(n13151), .ZN(n13425) );
  AOI22_X1 U14144 ( .A1(n10052), .A2(n11126), .B1(n11236), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14145 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U14146 ( .A1(n11128), .A2(n11127), .ZN(n13424) );
  AOI22_X1 U14147 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U14148 ( .A1(n11236), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11129) );
  OAI211_X1 U14149 ( .C1(n11131), .C2(n11301), .A(n11130), .B(n11129), .ZN(
        n13281) );
  OR2_X1 U14150 ( .A1(n11301), .A2(n11132), .ZN(n11133) );
  INV_X1 U14151 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14152 ( .A1(n11236), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14153 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11134) );
  OAI211_X1 U14154 ( .C1(n9717), .C2(n11136), .A(n11135), .B(n11134), .ZN(
        n13594) );
  NOR2_X1 U14155 ( .A1(n13597), .A2(n11138), .ZN(n13306) );
  NAND2_X1 U14156 ( .A1(n11236), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14157 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14158 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11562), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U14159 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11139) );
  AND3_X1 U14160 ( .A1(n11141), .A2(n11140), .A3(n11139), .ZN(n11153) );
  AOI22_X1 U14161 ( .A1(n11617), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14162 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11144) );
  NAND2_X1 U14163 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U14164 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11142) );
  NAND4_X1 U14165 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n11151) );
  NAND2_X1 U14166 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11149) );
  NAND2_X1 U14167 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11148) );
  NAND2_X1 U14168 ( .A1(n11576), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14169 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11146) );
  NAND4_X1 U14170 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11150) );
  NOR2_X1 U14171 ( .A1(n11151), .A2(n11150), .ZN(n11152) );
  OR2_X1 U14172 ( .A1(n11301), .A2(n12843), .ZN(n11156) );
  NAND2_X1 U14173 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11155) );
  NAND2_X1 U14174 ( .A1(n11410), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n11154) );
  NAND4_X1 U14175 ( .A1(n11157), .A2(n11156), .A3(n11155), .A4(n11154), .ZN(
        n16684) );
  INV_X1 U14176 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11477) );
  OAI22_X1 U14177 ( .A1(n11477), .A2(n11609), .B1(n11608), .B2(n11158), .ZN(
        n11162) );
  INV_X1 U14178 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11160) );
  OAI22_X1 U14179 ( .A1(n11160), .A2(n11613), .B1(n11612), .B2(n11159), .ZN(
        n11161) );
  NOR2_X1 U14180 ( .A1(n11162), .A2(n11161), .ZN(n11176) );
  AOI22_X1 U14181 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14182 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U14183 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11164) );
  NAND2_X1 U14184 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11163) );
  AND4_X1 U14185 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(
        n11175) );
  AOI22_X1 U14186 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11623), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11174) );
  INV_X1 U14187 ( .A(n11564), .ZN(n11624) );
  INV_X1 U14188 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11167) );
  OAI22_X1 U14189 ( .A1(n11168), .A2(n11625), .B1(n11624), .B2(n11167), .ZN(
        n11172) );
  INV_X1 U14190 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11170) );
  INV_X1 U14191 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11169) );
  OAI22_X1 U14192 ( .A1(n11629), .A2(n11170), .B1(n11169), .B2(n11627), .ZN(
        n11171) );
  NOR2_X1 U14193 ( .A1(n11172), .A2(n11171), .ZN(n11173) );
  NAND4_X1 U14194 ( .A1(n11176), .A2(n11175), .A3(n11174), .A4(n11173), .ZN(
        n12468) );
  INV_X1 U14195 ( .A(n12468), .ZN(n11179) );
  AOI22_X1 U14196 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11178) );
  NAND2_X1 U14197 ( .A1(n11236), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11177) );
  OAI211_X1 U14198 ( .C1(n11179), .C2(n11301), .A(n11178), .B(n11177), .ZN(
        n13323) );
  AOI22_X1 U14199 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11623), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14200 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11562), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14201 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11563), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11180) );
  AND3_X1 U14202 ( .A1(n11182), .A2(n11181), .A3(n11180), .ZN(n11194) );
  AOI22_X1 U14203 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14204 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14205 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11184) );
  NAND2_X1 U14206 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11183) );
  NAND4_X1 U14207 ( .A1(n11186), .A2(n11185), .A3(n11184), .A4(n11183), .ZN(
        n11192) );
  NAND2_X1 U14208 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11190) );
  NAND2_X1 U14209 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11189) );
  NAND2_X1 U14210 ( .A1(n11576), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11188) );
  NAND2_X1 U14211 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11187) );
  NAND4_X1 U14212 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11191) );
  NOR2_X1 U14213 ( .A1(n11192), .A2(n11191), .ZN(n11193) );
  AOI22_X1 U14214 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U14215 ( .A1(n11236), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11195) );
  OAI211_X1 U14216 ( .C1(n12561), .C2(n11301), .A(n11196), .B(n11195), .ZN(
        n15819) );
  INV_X1 U14217 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11198) );
  OAI22_X1 U14218 ( .A1(n11198), .A2(n11609), .B1(n11608), .B2(n11197), .ZN(
        n11200) );
  INV_X1 U14219 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11518) );
  OAI22_X1 U14220 ( .A1(n11518), .A2(n11613), .B1(n11612), .B2(n11519), .ZN(
        n11199) );
  NOR2_X1 U14221 ( .A1(n11200), .A2(n11199), .ZN(n11215) );
  INV_X1 U14222 ( .A(n11623), .ZN(n11266) );
  INV_X1 U14223 ( .A(n11201), .ZN(n11262) );
  INV_X1 U14224 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11520) );
  OAI22_X1 U14225 ( .A1(n11202), .A2(n11266), .B1(n11262), .B2(n11520), .ZN(
        n11208) );
  NAND2_X1 U14226 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11206) );
  NAND2_X1 U14227 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11205) );
  NAND2_X1 U14228 ( .A1(n11564), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14229 ( .A1(n11562), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11203) );
  NAND4_X1 U14230 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n11207) );
  NOR2_X1 U14231 ( .A1(n11208), .A2(n11207), .ZN(n11214) );
  AOI22_X1 U14232 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14233 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U14234 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U14235 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11209) );
  AND4_X1 U14236 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11213) );
  AOI22_X1 U14237 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U14238 ( .A1(n11236), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11216) );
  OAI211_X1 U14239 ( .C1(n12649), .C2(n11301), .A(n11217), .B(n11216), .ZN(
        n15197) );
  AOI22_X1 U14240 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U14241 ( .A1(n11236), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11234) );
  INV_X1 U14242 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11219) );
  INV_X1 U14243 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11218) );
  OAI22_X1 U14244 ( .A1(n11219), .A2(n11609), .B1(n11608), .B2(n11218), .ZN(
        n11221) );
  INV_X1 U14245 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11537) );
  INV_X1 U14246 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11538) );
  OAI22_X1 U14247 ( .A1(n11537), .A2(n11613), .B1(n11612), .B2(n11538), .ZN(
        n11220) );
  NOR2_X1 U14248 ( .A1(n11221), .A2(n11220), .ZN(n11232) );
  AOI22_X1 U14249 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14250 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14251 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14252 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11222) );
  AND4_X1 U14253 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11231) );
  AOI22_X1 U14254 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11230) );
  INV_X1 U14255 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11528) );
  INV_X1 U14256 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11226) );
  OAI22_X1 U14257 ( .A1(n11528), .A2(n11629), .B1(n11624), .B2(n11226), .ZN(
        n11228) );
  INV_X1 U14258 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11527) );
  INV_X1 U14259 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11530) );
  OAI22_X1 U14260 ( .A1(n11625), .A2(n11527), .B1(n11530), .B2(n11627), .ZN(
        n11227) );
  NOR2_X1 U14261 ( .A1(n11228), .A2(n11227), .ZN(n11229) );
  NAND4_X1 U14262 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n12831) );
  NAND2_X1 U14263 ( .A1(n10052), .A2(n12831), .ZN(n11233) );
  INV_X1 U14264 ( .A(n11236), .ZN(n11323) );
  INV_X1 U14265 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20170) );
  AOI22_X1 U14266 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11257) );
  INV_X1 U14267 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11237) );
  OAI22_X1 U14268 ( .A1(n11608), .A2(n11238), .B1(n11609), .B2(n11237), .ZN(
        n11241) );
  OAI22_X1 U14269 ( .A1(n12404), .A2(n11613), .B1(n11612), .B2(n11239), .ZN(
        n11240) );
  NOR2_X1 U14270 ( .A1(n11241), .A2(n11240), .ZN(n11255) );
  AOI22_X1 U14271 ( .A1(n11617), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14272 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11244) );
  NAND2_X1 U14273 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11243) );
  NAND2_X1 U14274 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11242) );
  AND4_X1 U14275 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11254) );
  AOI22_X1 U14276 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11253) );
  INV_X1 U14277 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11247) );
  OAI22_X1 U14278 ( .A1(n11625), .A2(n11247), .B1(n11624), .B2(n11246), .ZN(
        n11251) );
  OAI22_X1 U14279 ( .A1(n11629), .A2(n11249), .B1(n11627), .B2(n11248), .ZN(
        n11250) );
  NOR2_X1 U14280 ( .A1(n11251), .A2(n11250), .ZN(n11252) );
  NAND4_X1 U14281 ( .A1(n11255), .A2(n11254), .A3(n11253), .A4(n11252), .ZN(
        n13092) );
  NAND2_X1 U14282 ( .A1(n10052), .A2(n13092), .ZN(n11256) );
  OAI211_X1 U14283 ( .C1(n11323), .C2(n20170), .A(n11257), .B(n11256), .ZN(
        n15189) );
  AOI22_X1 U14284 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11283) );
  NAND2_X1 U14285 ( .A1(n11236), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11282) );
  INV_X1 U14286 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11260) );
  INV_X1 U14287 ( .A(n11258), .ZN(n11259) );
  INV_X1 U14288 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11763) );
  OAI22_X1 U14289 ( .A1(n11260), .A2(n11609), .B1(n11259), .B2(n11763), .ZN(
        n11264) );
  INV_X1 U14290 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12552) );
  INV_X1 U14291 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11261) );
  OAI22_X1 U14292 ( .A1(n12552), .A2(n11613), .B1(n11262), .B2(n11261), .ZN(
        n11263) );
  NOR2_X1 U14293 ( .A1(n11264), .A2(n11263), .ZN(n11280) );
  OAI22_X1 U14294 ( .A1(n11267), .A2(n11612), .B1(n11266), .B2(n11265), .ZN(
        n11273) );
  NAND2_X1 U14295 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14296 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11270) );
  NAND2_X1 U14297 ( .A1(n11564), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11269) );
  NAND2_X1 U14298 ( .A1(n11562), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11268) );
  NAND4_X1 U14299 ( .A1(n11271), .A2(n11270), .A3(n11269), .A4(n11268), .ZN(
        n11272) );
  NOR2_X1 U14300 ( .A1(n11273), .A2(n11272), .ZN(n11279) );
  AOI22_X1 U14301 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11277) );
  AOI22_X1 U14302 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11276) );
  NAND2_X1 U14303 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11275) );
  NAND2_X1 U14304 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11274) );
  AND4_X1 U14305 ( .A1(n11277), .A2(n11276), .A3(n11275), .A4(n11274), .ZN(
        n11278) );
  OR2_X1 U14306 ( .A1(n11301), .A2(n12978), .ZN(n11281) );
  AOI22_X1 U14307 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11304) );
  NAND2_X1 U14308 ( .A1(n11236), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14309 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14310 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n11562), .ZN(n11286) );
  AOI22_X1 U14311 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11285) );
  AND3_X1 U14312 ( .A1(n11287), .A2(n11286), .A3(n11285), .ZN(n11300) );
  AOI22_X1 U14313 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14314 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11288), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U14315 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11290) );
  NAND2_X1 U14316 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11289) );
  NAND4_X1 U14317 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n11298) );
  NAND2_X1 U14318 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11296) );
  NAND2_X1 U14319 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11295) );
  NAND2_X1 U14320 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11294) );
  NAND2_X1 U14321 ( .A1(n11576), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11293) );
  NAND4_X1 U14322 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n11297) );
  NOR2_X1 U14323 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  OR2_X1 U14324 ( .A1(n11301), .A2(n13297), .ZN(n11302) );
  INV_X1 U14325 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13403) );
  NAND2_X1 U14326 ( .A1(n11236), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U14327 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11305) );
  OAI211_X1 U14328 ( .C1(n13403), .C2(n9717), .A(n11306), .B(n11305), .ZN(
        n13401) );
  INV_X1 U14329 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20178) );
  NAND2_X1 U14330 ( .A1(n11410), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n11308) );
  NAND2_X1 U14331 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11307) );
  OAI211_X1 U14332 ( .C1(n11323), .C2(n20178), .A(n11308), .B(n11307), .ZN(
        n13432) );
  AOI22_X1 U14333 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U14334 ( .A1(n11236), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11309) );
  OR2_X2 U14335 ( .A1(n13581), .A2(n13580), .ZN(n15146) );
  AOI22_X1 U14336 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11312) );
  NAND2_X1 U14337 ( .A1(n11236), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14338 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U14339 ( .A1(n11236), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11313) );
  INV_X1 U14340 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20185) );
  NAND2_X1 U14341 ( .A1(n11410), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n11316) );
  NAND2_X1 U14342 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11315) );
  OAI211_X1 U14343 ( .C1(n11323), .C2(n20185), .A(n11316), .B(n11315), .ZN(
        n15133) );
  AOI22_X1 U14344 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11318) );
  NAND2_X1 U14345 ( .A1(n11236), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14346 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U14347 ( .A1(n11236), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11319) );
  INV_X1 U14348 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20191) );
  NAND2_X1 U14349 ( .A1(n11410), .A2(P2_EAX_REG_24__SCAN_IN), .ZN(n11322) );
  NAND2_X1 U14350 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11321) );
  OAI211_X1 U14351 ( .C1(n11323), .C2(n20191), .A(n11322), .B(n11321), .ZN(
        n15343) );
  NAND2_X1 U14352 ( .A1(n11236), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U14353 ( .A1(n11410), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n11324) );
  OAI211_X1 U14354 ( .C1(n11335), .C2(n15648), .A(n11325), .B(n11324), .ZN(
        n15334) );
  AOI22_X1 U14355 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11327) );
  NAND2_X1 U14356 ( .A1(n11236), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11326) );
  AND2_X1 U14357 ( .A1(n11327), .A2(n11326), .ZN(n15326) );
  AOI22_X1 U14358 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n11410), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U14359 ( .A1(n11236), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11329) );
  AND2_X1 U14360 ( .A1(n11330), .A2(n11329), .ZN(n15315) );
  INV_X1 U14361 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n21039) );
  NAND2_X1 U14362 ( .A1(n11236), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14363 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11331) );
  OAI211_X1 U14364 ( .C1(n9717), .C2(n21039), .A(n11332), .B(n11331), .ZN(
        n11395) );
  AND2_X2 U14365 ( .A1(n15317), .A2(n11395), .ZN(n15300) );
  NAND2_X1 U14366 ( .A1(n11236), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11334) );
  NAND2_X1 U14367 ( .A1(n11410), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n11333) );
  OAI211_X1 U14368 ( .C1(n11335), .C2(n15611), .A(n11334), .B(n11333), .ZN(
        n15299) );
  XOR2_X1 U14369 ( .A(n11408), .B(n15302), .Z(n16530) );
  INV_X1 U14370 ( .A(n11336), .ZN(n15854) );
  NOR2_X1 U14371 ( .A1(n15854), .A2(n11337), .ZN(n16718) );
  AND2_X1 U14372 ( .A1(n16728), .A2(n20281), .ZN(n11339) );
  NOR2_X1 U14373 ( .A1(n16718), .A2(n11339), .ZN(n11340) );
  XOR2_X1 U14374 ( .A(n11341), .B(n15225), .Z(n11834) );
  INV_X1 U14375 ( .A(n11834), .ZN(n16532) );
  INV_X1 U14376 ( .A(n11342), .ZN(n11343) );
  NAND2_X1 U14377 ( .A1(n16532), .A2(n16689), .ZN(n11344) );
  NAND2_X1 U14378 ( .A1(n19529), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11387) );
  OAI211_X1 U14379 ( .C1(n16530), .C2(n16701), .A(n11344), .B(n11387), .ZN(
        n11383) );
  INV_X1 U14380 ( .A(n15882), .ZN(n16720) );
  INV_X1 U14381 ( .A(n12110), .ZN(n15740) );
  NAND2_X1 U14382 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U14383 ( .A1(n11347), .A2(n12127), .ZN(n12111) );
  INV_X1 U14384 ( .A(n12127), .ZN(n12106) );
  NAND2_X1 U14385 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12106), .ZN(
        n12112) );
  INV_X1 U14386 ( .A(n12112), .ZN(n11348) );
  AOI21_X1 U14387 ( .B1(n15740), .B2(n12111), .A(n11348), .ZN(n13147) );
  NOR2_X1 U14388 ( .A1(n13147), .A2(n11372), .ZN(n13452) );
  NAND2_X1 U14389 ( .A1(n11350), .A2(n20279), .ZN(n11351) );
  OAI21_X1 U14390 ( .B1(n11352), .B2(n11349), .A(n11351), .ZN(n11353) );
  INV_X1 U14391 ( .A(n11353), .ZN(n11357) );
  OAI21_X1 U14392 ( .B1(n11804), .B2(n11354), .A(n11349), .ZN(n11355) );
  NAND2_X1 U14393 ( .A1(n11355), .A2(n11802), .ZN(n11356) );
  AND3_X1 U14394 ( .A1(n11358), .A2(n11357), .A3(n11356), .ZN(n11363) );
  NAND2_X1 U14395 ( .A1(n11359), .A2(n20281), .ZN(n15853) );
  NAND2_X1 U14396 ( .A1(n15853), .A2(n11360), .ZN(n11361) );
  NAND2_X1 U14397 ( .A1(n11361), .A2(n19569), .ZN(n11362) );
  NAND2_X1 U14398 ( .A1(n11363), .A2(n11362), .ZN(n15912) );
  NOR2_X1 U14399 ( .A1(n15912), .A2(n11364), .ZN(n11365) );
  NAND2_X1 U14400 ( .A1(n13452), .A2(n16705), .ZN(n13423) );
  NOR3_X1 U14401 ( .A1(n15846), .A2(n16682), .A3(n16685), .ZN(n11373) );
  NAND2_X1 U14402 ( .A1(n15847), .A2(n11373), .ZN(n15818) );
  NOR2_X1 U14403 ( .A1(n15726), .A2(n11366), .ZN(n11367) );
  NAND2_X1 U14404 ( .A1(n11368), .A2(n11367), .ZN(n11377) );
  INV_X1 U14405 ( .A(n15694), .ZN(n15706) );
  NAND2_X1 U14406 ( .A1(n15706), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11376) );
  INV_X1 U14407 ( .A(n15665), .ZN(n15654) );
  NAND3_X1 U14408 ( .A1(n15676), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15654), .ZN(n15642) );
  NAND2_X1 U14409 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15631) );
  NOR2_X1 U14410 ( .A1(n15642), .A2(n15631), .ZN(n15627) );
  NAND2_X1 U14411 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15607) );
  NOR2_X1 U14412 ( .A1(n15607), .A2(n15611), .ZN(n11380) );
  NAND2_X1 U14413 ( .A1(n15627), .A2(n11380), .ZN(n11417) );
  INV_X1 U14414 ( .A(n16705), .ZN(n13146) );
  INV_X1 U14415 ( .A(n15743), .ZN(n11369) );
  NAND2_X1 U14416 ( .A1(n11369), .A2(n12112), .ZN(n12126) );
  NAND2_X1 U14417 ( .A1(n11370), .A2(n15727), .ZN(n16695) );
  OAI211_X1 U14418 ( .C1(n12110), .C2(n12111), .A(n12126), .B(n16695), .ZN(
        n13148) );
  INV_X1 U14419 ( .A(n13148), .ZN(n11371) );
  NAND2_X1 U14420 ( .A1(n13146), .A2(n11371), .ZN(n15816) );
  INV_X1 U14421 ( .A(n15816), .ZN(n15701) );
  OAI21_X1 U14422 ( .B1(n13148), .B2(n11372), .A(n15816), .ZN(n13456) );
  OAI21_X1 U14423 ( .B1(n13455), .B2(n13422), .A(n16705), .ZN(n13454) );
  NAND2_X1 U14424 ( .A1(n13456), .A2(n13454), .ZN(n15845) );
  INV_X1 U14425 ( .A(n11373), .ZN(n11374) );
  AND2_X1 U14426 ( .A1(n16705), .A2(n11374), .ZN(n11375) );
  INV_X1 U14427 ( .A(n11376), .ZN(n11378) );
  INV_X1 U14428 ( .A(n11377), .ZN(n15702) );
  NAND3_X1 U14429 ( .A1(n15831), .A2(n11378), .A3(n15702), .ZN(n11379) );
  NAND2_X1 U14430 ( .A1(n11379), .A2(n15816), .ZN(n15677) );
  OAI211_X1 U14431 ( .C1(n15654), .C2(n15701), .A(n15677), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15643) );
  OAI21_X1 U14432 ( .B1(n15643), .B2(n15631), .A(n15816), .ZN(n15621) );
  OAI211_X1 U14433 ( .C1(n11380), .C2(n13146), .A(n15621), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11413) );
  INV_X1 U14434 ( .A(n11413), .ZN(n11381) );
  AOI21_X1 U14435 ( .B1(n11417), .B2(n11416), .A(n11381), .ZN(n11382) );
  NAND2_X1 U14436 ( .A1(n11385), .A2(n16662), .ZN(n11393) );
  XNOR2_X1 U14437 ( .A(n9768), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16535) );
  NAND2_X1 U14438 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11386) );
  OAI211_X1 U14439 ( .C1(n19542), .C2(n16535), .A(n11387), .B(n11386), .ZN(
        n11388) );
  AOI21_X1 U14440 ( .B1(n16532), .B2(n19538), .A(n11388), .ZN(n11389) );
  NAND2_X1 U14441 ( .A1(n11393), .A2(n11392), .ZN(P2_U2984) );
  NAND2_X1 U14442 ( .A1(n11394), .A2(n16673), .ZN(n11407) );
  NOR2_X1 U14443 ( .A1(n15317), .A2(n11395), .ZN(n11396) );
  OAI21_X1 U14444 ( .B1(n16552), .B2(n16701), .A(n11397), .ZN(n11401) );
  INV_X1 U14445 ( .A(n15621), .ZN(n11398) );
  AOI21_X1 U14446 ( .B1(n15627), .B2(n15607), .A(n11398), .ZN(n15612) );
  AOI21_X1 U14447 ( .B1(n15627), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11399) );
  NOR2_X1 U14448 ( .A1(n15612), .A2(n11399), .ZN(n11400) );
  AOI211_X1 U14449 ( .C1(n16689), .C2(n11402), .A(n11401), .B(n11400), .ZN(
        n11403) );
  NAND2_X1 U14450 ( .A1(n11407), .A2(n11406), .ZN(P2_U3018) );
  INV_X1 U14451 ( .A(n15302), .ZN(n11409) );
  NAND2_X1 U14452 ( .A1(n11409), .A2(n11408), .ZN(n11412) );
  AOI222_X1 U14453 ( .A1(n11236), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11328), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n11410), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n11411) );
  XNOR2_X2 U14454 ( .A(n11412), .B(n11411), .ZN(n16524) );
  NAND3_X1 U14455 ( .A1(n11413), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15816), .ZN(n11415) );
  OAI211_X1 U14456 ( .C1(n16524), .C2(n16701), .A(n11415), .B(n11414), .ZN(
        n11418) );
  INV_X1 U14457 ( .A(n11420), .ZN(n11421) );
  OAI21_X1 U14458 ( .B1(n16697), .B2(n11422), .A(n11421), .ZN(P2_U3015) );
  NAND2_X1 U14459 ( .A1(n11423), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U14460 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19920) );
  NAND2_X1 U14461 ( .A1(n19920), .A2(n20243), .ZN(n11426) );
  NAND2_X1 U14462 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20057) );
  INV_X1 U14463 ( .A(n20057), .ZN(n11425) );
  NAND2_X1 U14464 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11425), .ZN(
        n19548) );
  AND2_X1 U14465 ( .A1(n11426), .A2(n19548), .ZN(n19709) );
  AOI22_X1 U14466 ( .A1(n11444), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20223), .B2(n19709), .ZN(n11427) );
  INV_X1 U14467 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14468 ( .A1(n11444), .A2(n15871), .B1(n20223), .B2(n20263), .ZN(
        n11429) );
  XNOR2_X1 U14469 ( .A(n11433), .B(n11434), .ZN(n12101) );
  NAND2_X1 U14470 ( .A1(n11444), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11431) );
  NAND2_X1 U14471 ( .A1(n20252), .A2(n20263), .ZN(n19829) );
  NAND2_X1 U14472 ( .A1(n19920), .A2(n19829), .ZN(n19708) );
  INV_X1 U14473 ( .A(n19708), .ZN(n19773) );
  NAND2_X1 U14474 ( .A1(n19773), .A2(n20223), .ZN(n19892) );
  NAND2_X1 U14475 ( .A1(n11431), .A2(n19892), .ZN(n11432) );
  NAND2_X1 U14476 ( .A1(n12101), .A2(n12100), .ZN(n12102) );
  INV_X1 U14477 ( .A(n11433), .ZN(n12097) );
  NAND2_X1 U14478 ( .A1(n12097), .A2(n11434), .ZN(n11435) );
  NAND2_X1 U14479 ( .A1(n11437), .A2(n10221), .ZN(n11438) );
  INV_X1 U14480 ( .A(n19920), .ZN(n11441) );
  NAND2_X1 U14481 ( .A1(n20236), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19769) );
  INV_X1 U14482 ( .A(n19769), .ZN(n19772) );
  NAND2_X1 U14483 ( .A1(n11441), .A2(n19772), .ZN(n19832) );
  NAND2_X1 U14484 ( .A1(n19548), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U14485 ( .A1(n19832), .A2(n11442), .ZN(n11443) );
  AOI22_X1 U14486 ( .A1(n11444), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20223), .B2(n11443), .ZN(n11445) );
  NAND2_X1 U14487 ( .A1(n11446), .A2(n11445), .ZN(n11448) );
  NAND2_X1 U14488 ( .A1(n11448), .A2(n11447), .ZN(n11451) );
  OR2_X1 U14489 ( .A1(n11448), .A2(n11447), .ZN(n11449) );
  NAND2_X1 U14490 ( .A1(n12400), .A2(n12399), .ZN(n12398) );
  NAND2_X1 U14491 ( .A1(n11423), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11450) );
  AND2_X1 U14492 ( .A1(n11451), .A2(n11450), .ZN(n11452) );
  INV_X1 U14493 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12839) );
  OR2_X1 U14494 ( .A1(n12843), .A2(n12839), .ZN(n11453) );
  INV_X1 U14495 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12404) );
  NOR2_X1 U14496 ( .A1(n10247), .A2(n12404), .ZN(n12467) );
  AND2_X1 U14497 ( .A1(n12468), .A2(n12467), .ZN(n11454) );
  NOR2_X1 U14498 ( .A1(n13297), .A2(n12978), .ZN(n11456) );
  AND2_X1 U14499 ( .A1(n11456), .A2(n13092), .ZN(n11457) );
  INV_X1 U14500 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11459) );
  INV_X1 U14501 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11458) );
  OAI22_X1 U14502 ( .A1(n11608), .A2(n11459), .B1(n11609), .B2(n11458), .ZN(
        n11463) );
  INV_X1 U14503 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11461) );
  INV_X1 U14504 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11460) );
  OAI22_X1 U14505 ( .A1(n11613), .A2(n11461), .B1(n11612), .B2(n11460), .ZN(
        n11462) );
  NOR2_X1 U14506 ( .A1(n11463), .A2(n11462), .ZN(n11476) );
  AOI22_X1 U14507 ( .A1(n11617), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14508 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U14509 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U14510 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11465) );
  AND4_X1 U14511 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(
        n11475) );
  AOI22_X1 U14512 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11474) );
  INV_X1 U14513 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11469) );
  INV_X1 U14514 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12095) );
  OAI22_X1 U14515 ( .A1(n11625), .A2(n11469), .B1(n11624), .B2(n12095), .ZN(
        n11472) );
  INV_X1 U14516 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11470) );
  INV_X1 U14517 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11591) );
  OAI22_X1 U14518 ( .A1(n11629), .A2(n11470), .B1(n11627), .B2(n11591), .ZN(
        n11471) );
  NOR2_X1 U14519 ( .A1(n11472), .A2(n11471), .ZN(n11473) );
  NAND4_X1 U14520 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(
        n13395) );
  AOI22_X1 U14521 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11258), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14522 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11574), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11486) );
  INV_X1 U14523 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11479) );
  OAI22_X1 U14524 ( .A1(n11479), .A2(n11478), .B1(n9718), .B2(n11477), .ZN(
        n11483) );
  INV_X1 U14525 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n20879) );
  INV_X1 U14526 ( .A(n11618), .ZN(n11481) );
  INV_X1 U14527 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11480) );
  OAI22_X1 U14528 ( .A1(n20879), .A2(n9715), .B1(n11481), .B2(n11480), .ZN(
        n11482) );
  NOR2_X1 U14529 ( .A1(n11483), .A2(n11482), .ZN(n11485) );
  AOI22_X1 U14530 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11575), .B1(
        n11576), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11484) );
  NAND4_X1 U14531 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n11492) );
  AOI22_X1 U14532 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14533 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n11562), .ZN(n11489) );
  AOI22_X1 U14534 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11488) );
  NAND3_X1 U14535 ( .A1(n11490), .A2(n11489), .A3(n11488), .ZN(n11491) );
  NOR2_X1 U14536 ( .A1(n11492), .A2(n11491), .ZN(n13431) );
  AOI22_X1 U14537 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14538 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n11562), .ZN(n11494) );
  AOI22_X1 U14539 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11493) );
  AND3_X1 U14540 ( .A1(n11495), .A2(n11494), .A3(n11493), .ZN(n11507) );
  AOI22_X1 U14541 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14542 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11464), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11498) );
  NAND2_X1 U14543 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11497) );
  NAND2_X1 U14544 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11496) );
  NAND4_X1 U14545 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11505) );
  NAND2_X1 U14546 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14547 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14548 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11501) );
  NAND2_X1 U14549 ( .A1(n11576), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11500) );
  NAND4_X1 U14550 ( .A1(n11503), .A2(n11502), .A3(n11501), .A4(n11500), .ZN(
        n11504) );
  NOR2_X1 U14551 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  INV_X1 U14552 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11508) );
  OAI22_X1 U14553 ( .A1(n11509), .A2(n11609), .B1(n11608), .B2(n11508), .ZN(
        n11513) );
  INV_X1 U14554 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11510) );
  OAI22_X1 U14555 ( .A1(n11511), .A2(n11613), .B1(n11612), .B2(n11510), .ZN(
        n11512) );
  NOR2_X1 U14556 ( .A1(n11513), .A2(n11512), .ZN(n11526) );
  AOI22_X1 U14557 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14558 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11464), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14559 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11515) );
  NAND2_X1 U14560 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11514) );
  AND4_X1 U14561 ( .A1(n11517), .A2(n11516), .A3(n11515), .A4(n11514), .ZN(
        n11525) );
  AOI22_X1 U14562 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11201), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11524) );
  OAI22_X1 U14563 ( .A1(n11519), .A2(n11625), .B1(n11624), .B2(n11518), .ZN(
        n11522) );
  INV_X1 U14564 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11693) );
  OAI22_X1 U14565 ( .A1(n11629), .A2(n11520), .B1(n11693), .B2(n11627), .ZN(
        n11521) );
  NOR2_X1 U14566 ( .A1(n11522), .A2(n11521), .ZN(n11523) );
  NAND4_X1 U14567 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n15294) );
  OAI22_X1 U14568 ( .A1(n11528), .A2(n11609), .B1(n11608), .B2(n11527), .ZN(
        n11532) );
  INV_X1 U14569 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11529) );
  OAI22_X1 U14570 ( .A1(n11530), .A2(n11613), .B1(n11612), .B2(n11529), .ZN(
        n11531) );
  NOR2_X1 U14571 ( .A1(n11532), .A2(n11531), .ZN(n11546) );
  AOI22_X1 U14572 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14573 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11464), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14574 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11534) );
  NAND2_X1 U14575 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11533) );
  AND4_X1 U14576 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11545) );
  AOI22_X1 U14577 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11623), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11544) );
  OAI22_X1 U14578 ( .A1(n11538), .A2(n11625), .B1(n11624), .B2(n11537), .ZN(
        n11542) );
  INV_X1 U14579 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11540) );
  INV_X1 U14580 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11539) );
  OAI22_X1 U14581 ( .A1(n11629), .A2(n11540), .B1(n11627), .B2(n11539), .ZN(
        n11541) );
  NOR2_X1 U14582 ( .A1(n11542), .A2(n11541), .ZN(n11543) );
  NAND4_X1 U14583 ( .A1(n11546), .A2(n11545), .A3(n11544), .A4(n11543), .ZN(
        n15286) );
  AOI22_X1 U14584 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11623), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14585 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11562), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14586 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11547) );
  AND3_X1 U14587 ( .A1(n11549), .A2(n11548), .A3(n11547), .ZN(n11561) );
  AOI22_X1 U14588 ( .A1(n11617), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14589 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11552) );
  NAND2_X1 U14590 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11551) );
  NAND2_X1 U14591 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11550) );
  NAND4_X1 U14592 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11559) );
  NAND2_X1 U14593 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11557) );
  NAND2_X1 U14594 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11556) );
  NAND2_X1 U14595 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11555) );
  NAND2_X1 U14596 ( .A1(n11576), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11554) );
  NAND4_X1 U14597 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n11558) );
  NOR2_X1 U14598 ( .A1(n11559), .A2(n11558), .ZN(n11560) );
  AND2_X1 U14599 ( .A1(n11561), .A2(n11560), .ZN(n15280) );
  AOI22_X1 U14600 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11623), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14601 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n11562), .ZN(n11567) );
  AOI22_X1 U14602 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11565), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11566) );
  AND3_X1 U14603 ( .A1(n11568), .A2(n11567), .A3(n11566), .ZN(n11584) );
  AOI22_X1 U14604 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11617), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14605 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11464), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11571) );
  NAND2_X1 U14606 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11570) );
  NAND2_X1 U14607 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11569) );
  NAND4_X1 U14608 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n11582) );
  NAND2_X1 U14609 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11580) );
  NAND2_X1 U14610 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11579) );
  NAND2_X1 U14611 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11578) );
  NAND2_X1 U14612 ( .A1(n11576), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11577) );
  NAND4_X1 U14613 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11581) );
  NOR2_X1 U14614 ( .A1(n11582), .A2(n11581), .ZN(n11583) );
  AND2_X1 U14615 ( .A1(n11584), .A2(n11583), .ZN(n15276) );
  AOI22_X1 U14616 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14617 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14618 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11594) );
  INV_X1 U14619 ( .A(n11666), .ZN(n11788) );
  INV_X1 U14620 ( .A(n11586), .ZN(n11597) );
  NAND2_X1 U14621 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11590) );
  INV_X1 U14622 ( .A(n11587), .ZN(n11589) );
  NAND2_X1 U14623 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U14624 ( .A1(n11589), .A2(n11588), .ZN(n11785) );
  OAI211_X1 U14625 ( .C1(n11788), .C2(n11591), .A(n11590), .B(n11785), .ZN(
        n11592) );
  INV_X1 U14626 ( .A(n11592), .ZN(n11593) );
  NAND4_X1 U14627 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11606) );
  AOI22_X1 U14628 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14629 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14630 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11602) );
  INV_X1 U14631 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U14632 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11598) );
  INV_X1 U14633 ( .A(n11785), .ZN(n11761) );
  OAI211_X1 U14634 ( .C1(n11788), .C2(n11599), .A(n11598), .B(n11761), .ZN(
        n11600) );
  INV_X1 U14635 ( .A(n11600), .ZN(n11601) );
  NAND4_X1 U14636 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .ZN(
        n11605) );
  NAND2_X1 U14637 ( .A1(n20281), .A2(n11655), .ZN(n11636) );
  INV_X1 U14638 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11610) );
  INV_X1 U14639 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11607) );
  OAI22_X1 U14640 ( .A1(n11610), .A2(n11609), .B1(n11608), .B2(n11607), .ZN(
        n11616) );
  INV_X1 U14641 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11614) );
  INV_X1 U14642 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11611) );
  OAI22_X1 U14643 ( .A1(n11614), .A2(n11613), .B1(n11612), .B2(n11611), .ZN(
        n11615) );
  NOR2_X1 U14644 ( .A1(n11616), .A2(n11615), .ZN(n11635) );
  AOI22_X1 U14645 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11618), .B1(
        n11617), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14646 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11464), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11621) );
  NAND2_X1 U14647 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U14648 ( .A1(n11258), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11619) );
  AND4_X1 U14649 ( .A1(n11622), .A2(n11621), .A3(n11620), .A4(n11619), .ZN(
        n11634) );
  AOI22_X1 U14650 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11623), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11633) );
  INV_X1 U14651 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11626) );
  OAI22_X1 U14652 ( .A1(n11626), .A2(n11625), .B1(n11624), .B2(n12839), .ZN(
        n11631) );
  INV_X1 U14653 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11628) );
  INV_X1 U14654 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11787) );
  OAI22_X1 U14655 ( .A1(n11629), .A2(n11628), .B1(n11787), .B2(n11627), .ZN(
        n11630) );
  NOR2_X1 U14656 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  NAND4_X1 U14657 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11656) );
  XNOR2_X1 U14658 ( .A(n11636), .B(n11656), .ZN(n11661) );
  INV_X1 U14659 ( .A(n11655), .ZN(n11659) );
  NOR2_X1 U14660 ( .A1(n20281), .A2(n11659), .ZN(n15269) );
  AOI22_X1 U14661 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14662 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14663 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11643) );
  NAND2_X1 U14664 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11639) );
  OAI211_X1 U14665 ( .C1(n11788), .C2(n11640), .A(n11639), .B(n11785), .ZN(
        n11641) );
  INV_X1 U14666 ( .A(n11641), .ZN(n11642) );
  NAND4_X1 U14667 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11654) );
  AOI22_X1 U14668 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14669 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14670 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11650) );
  INV_X1 U14671 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14672 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11646) );
  OAI211_X1 U14673 ( .C1(n11788), .C2(n11647), .A(n11646), .B(n11761), .ZN(
        n11648) );
  INV_X1 U14674 ( .A(n11648), .ZN(n11649) );
  NAND4_X1 U14675 ( .A1(n11652), .A2(n11651), .A3(n11650), .A4(n11649), .ZN(
        n11653) );
  NAND2_X1 U14676 ( .A1(n11654), .A2(n11653), .ZN(n11658) );
  NAND2_X1 U14677 ( .A1(n11656), .A2(n11655), .ZN(n11663) );
  XOR2_X1 U14678 ( .A(n11658), .B(n11663), .Z(n11657) );
  NAND2_X1 U14679 ( .A1(n11657), .A2(n11684), .ZN(n15259) );
  INV_X1 U14680 ( .A(n11658), .ZN(n11664) );
  NAND2_X1 U14681 ( .A1(n9659), .A2(n11664), .ZN(n15262) );
  NOR2_X1 U14682 ( .A1(n15262), .A2(n11659), .ZN(n11660) );
  INV_X1 U14683 ( .A(n11663), .ZN(n11665) );
  AOI22_X1 U14684 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14685 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14686 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11666), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11671) );
  INV_X1 U14687 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11668) );
  NAND2_X1 U14688 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11667) );
  OAI211_X1 U14689 ( .C1(n11585), .C2(n11668), .A(n11667), .B(n11785), .ZN(
        n11669) );
  INV_X1 U14690 ( .A(n11669), .ZN(n11670) );
  NAND4_X1 U14691 ( .A1(n11673), .A2(n11672), .A3(n11671), .A4(n11670), .ZN(
        n11683) );
  AOI22_X1 U14692 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14693 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14694 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11679) );
  INV_X1 U14695 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U14696 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11675) );
  OAI211_X1 U14697 ( .C1(n11788), .C2(n11676), .A(n11675), .B(n11761), .ZN(
        n11677) );
  INV_X1 U14698 ( .A(n11677), .ZN(n11678) );
  NAND4_X1 U14699 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n11682) );
  AND2_X1 U14700 ( .A1(n11683), .A2(n11682), .ZN(n11687) );
  NAND2_X1 U14701 ( .A1(n11685), .A2(n11687), .ZN(n11708) );
  OAI211_X1 U14702 ( .C1(n11685), .C2(n11687), .A(n11684), .B(n11708), .ZN(
        n11689) );
  INV_X1 U14703 ( .A(n11689), .ZN(n11686) );
  INV_X1 U14704 ( .A(n11687), .ZN(n11688) );
  NOR2_X1 U14705 ( .A1(n20281), .A2(n11688), .ZN(n15252) );
  AOI22_X1 U14706 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14707 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14708 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14709 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11692) );
  OAI211_X1 U14710 ( .C1(n11788), .C2(n11693), .A(n11692), .B(n11785), .ZN(
        n11694) );
  INV_X1 U14711 ( .A(n11694), .ZN(n11695) );
  NAND4_X1 U14712 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11707) );
  AOI22_X1 U14713 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14714 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14715 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11703) );
  INV_X1 U14716 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U14717 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11699) );
  OAI211_X1 U14718 ( .C1(n11788), .C2(n11700), .A(n11699), .B(n11761), .ZN(
        n11701) );
  INV_X1 U14719 ( .A(n11701), .ZN(n11702) );
  NAND4_X1 U14720 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  NAND2_X1 U14721 ( .A1(n11707), .A2(n11706), .ZN(n11712) );
  AOI21_X1 U14722 ( .B1(n11708), .B2(n11712), .A(n11732), .ZN(n11711) );
  INV_X1 U14723 ( .A(n11708), .ZN(n11710) );
  INV_X1 U14724 ( .A(n11712), .ZN(n11709) );
  NAND2_X1 U14725 ( .A1(n11710), .A2(n11709), .ZN(n11733) );
  NAND2_X1 U14726 ( .A1(n11711), .A2(n11733), .ZN(n11714) );
  NOR2_X1 U14727 ( .A1(n20281), .A2(n11712), .ZN(n15245) );
  AOI22_X1 U14728 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14729 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14730 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11718) );
  NAND2_X1 U14731 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11715) );
  OAI211_X1 U14732 ( .C1(n11539), .C2(n11788), .A(n11715), .B(n11785), .ZN(
        n11716) );
  INV_X1 U14733 ( .A(n11716), .ZN(n11717) );
  NAND4_X1 U14734 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11729) );
  AOI22_X1 U14735 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11794), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14736 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14737 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11725) );
  INV_X1 U14738 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U14739 ( .A1(n11792), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11721) );
  OAI211_X1 U14740 ( .C1(n11788), .C2(n11722), .A(n11721), .B(n11761), .ZN(
        n11723) );
  INV_X1 U14741 ( .A(n11723), .ZN(n11724) );
  NAND4_X1 U14742 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11728) );
  AND2_X1 U14743 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  INV_X1 U14744 ( .A(n11730), .ZN(n11735) );
  INV_X1 U14745 ( .A(n11733), .ZN(n11731) );
  AOI211_X1 U14746 ( .C1(n11735), .C2(n11733), .A(n11732), .B(n15230), .ZN(
        n11734) );
  NOR2_X1 U14747 ( .A1(n20281), .A2(n11735), .ZN(n15237) );
  AOI22_X1 U14748 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14749 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14750 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11741) );
  INV_X1 U14751 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11738) );
  NAND2_X1 U14752 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11737) );
  OAI211_X1 U14753 ( .C1(n11788), .C2(n11738), .A(n11737), .B(n11785), .ZN(
        n11739) );
  INV_X1 U14754 ( .A(n11739), .ZN(n11740) );
  NAND4_X1 U14755 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11752) );
  AOI22_X1 U14756 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14757 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14758 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11748) );
  INV_X1 U14759 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11745) );
  NAND2_X1 U14760 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11744) );
  OAI211_X1 U14761 ( .C1(n11788), .C2(n11745), .A(n11744), .B(n11761), .ZN(
        n11746) );
  INV_X1 U14762 ( .A(n11746), .ZN(n11747) );
  NAND4_X1 U14763 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  NAND2_X1 U14764 ( .A1(n11752), .A2(n11751), .ZN(n11771) );
  AOI22_X1 U14765 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14766 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14767 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11757) );
  INV_X1 U14768 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U14769 ( .A1(n11792), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11753) );
  OAI211_X1 U14770 ( .C1(n11788), .C2(n11754), .A(n11753), .B(n11785), .ZN(
        n11755) );
  INV_X1 U14771 ( .A(n11755), .ZN(n11756) );
  NAND4_X1 U14772 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11770) );
  AOI22_X1 U14773 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11794), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14774 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14775 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U14776 ( .A1(n11792), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11762) );
  OAI211_X1 U14777 ( .C1(n11788), .C2(n11763), .A(n11762), .B(n11761), .ZN(
        n11764) );
  INV_X1 U14778 ( .A(n11764), .ZN(n11765) );
  NAND4_X1 U14779 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11769) );
  NAND2_X1 U14780 ( .A1(n11770), .A2(n11769), .ZN(n11775) );
  INV_X1 U14781 ( .A(n15230), .ZN(n11773) );
  INV_X1 U14782 ( .A(n11771), .ZN(n15232) );
  NAND2_X1 U14783 ( .A1(n20281), .A2(n15232), .ZN(n11772) );
  OR2_X1 U14784 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  NOR2_X1 U14785 ( .A1(n11774), .A2(n11775), .ZN(n11776) );
  AOI21_X1 U14786 ( .B1(n11775), .B2(n11774), .A(n11776), .ZN(n15226) );
  INV_X1 U14787 ( .A(n11776), .ZN(n11777) );
  AOI22_X1 U14788 ( .A1(n11794), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14789 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11779) );
  NAND2_X1 U14790 ( .A1(n11780), .A2(n11779), .ZN(n11800) );
  INV_X1 U14791 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14792 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11783) );
  AOI21_X1 U14793 ( .B1(n11792), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n11785), .ZN(n11782) );
  OAI211_X1 U14794 ( .C1(n11788), .C2(n11784), .A(n11783), .B(n11782), .ZN(
        n11799) );
  INV_X1 U14795 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11786) );
  OAI21_X1 U14796 ( .B1(n11586), .B2(n11786), .A(n11785), .ZN(n11791) );
  INV_X1 U14797 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11789) );
  OAI22_X1 U14798 ( .A1(n15903), .A2(n11789), .B1(n11788), .B2(n11787), .ZN(
        n11790) );
  AOI211_X1 U14799 ( .C1(n10485), .C2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11791), .B(n11790), .ZN(n11797) );
  AOI22_X1 U14800 ( .A1(n11793), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11792), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14801 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11794), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11795) );
  NAND3_X1 U14802 ( .A1(n11797), .A2(n11796), .A3(n11795), .ZN(n11798) );
  OAI21_X1 U14803 ( .B1(n11800), .B2(n11799), .A(n11798), .ZN(n11801) );
  NAND2_X1 U14804 ( .A1(n16721), .A2(n15882), .ZN(n15865) );
  AND2_X1 U14805 ( .A1(n11803), .A2(n11802), .ZN(n11805) );
  NAND2_X1 U14806 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  NAND2_X1 U14807 ( .A1(n15865), .A2(n11806), .ZN(n11807) );
  NAND2_X1 U14808 ( .A1(n11807), .A2(n20122), .ZN(n11810) );
  INV_X1 U14809 ( .A(n20122), .ZN(n12243) );
  INV_X1 U14810 ( .A(n16728), .ZN(n11808) );
  AND2_X1 U14811 ( .A1(n11349), .A2(n20276), .ZN(n16726) );
  NAND2_X1 U14812 ( .A1(n19272), .A2(n16726), .ZN(n11809) );
  NAND2_X1 U14813 ( .A1(n11832), .A2(n19487), .ZN(n11829) );
  NAND2_X1 U14814 ( .A1(n19463), .A2(n19590), .ZN(n15314) );
  NOR4_X1 U14815 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n11815) );
  NOR4_X1 U14816 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n11814) );
  NOR4_X1 U14817 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11813) );
  NOR4_X1 U14818 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n11812) );
  NAND4_X1 U14819 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11820) );
  NOR4_X1 U14820 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n11818) );
  NOR4_X1 U14821 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n11817) );
  NOR4_X1 U14822 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n11816) );
  INV_X1 U14823 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20153) );
  NAND4_X1 U14824 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n20153), .ZN(
        n11819) );
  AND2_X1 U14825 ( .A1(n10102), .A2(n11821), .ZN(n11822) );
  AOI22_X1 U14826 ( .A1(n19545), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n12447), .ZN(n19431) );
  INV_X1 U14827 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12254) );
  OAI22_X1 U14828 ( .A1(n19427), .A2(n19431), .B1(n19463), .B2(n12254), .ZN(
        n11825) );
  INV_X1 U14829 ( .A(n19422), .ZN(n15350) );
  INV_X1 U14830 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n11823) );
  NOR2_X1 U14831 ( .A1(n15350), .A2(n11823), .ZN(n11824) );
  AOI211_X1 U14832 ( .C1(n19420), .C2(BUF1_REG_30__SCAN_IN), .A(n11825), .B(
        n11824), .ZN(n11826) );
  OAI21_X1 U14833 ( .B1(n16530), .B2(n15314), .A(n11826), .ZN(n11827) );
  INV_X1 U14834 ( .A(n11827), .ZN(n11828) );
  NAND2_X1 U14835 ( .A1(n11829), .A2(n11828), .ZN(P2_U2889) );
  NAND2_X1 U14836 ( .A1(n11830), .A2(n16718), .ZN(n15863) );
  INV_X1 U14837 ( .A(n11364), .ZN(n15885) );
  NAND2_X1 U14838 ( .A1(n15863), .A2(n15885), .ZN(n11831) );
  NAND2_X1 U14839 ( .A1(n11832), .A2(n15281), .ZN(n11837) );
  NAND2_X1 U14840 ( .A1(n15279), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11833) );
  NAND2_X1 U14841 ( .A1(n11837), .A2(n11836), .ZN(P2_U2857) );
  NOR2_X1 U14842 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n11839) );
  NOR4_X1 U14843 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n11838) );
  NAND4_X1 U14844 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n11839), .A4(n11838), .ZN(n11852) );
  NOR4_X1 U14845 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_16__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n11843) );
  NOR4_X1 U14846 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n11842) );
  NOR4_X1 U14847 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11841) );
  NOR4_X1 U14848 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_8__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n11840) );
  AND4_X1 U14849 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n11848) );
  NOR4_X1 U14850 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11846) );
  NOR4_X1 U14851 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11845) );
  NOR4_X1 U14852 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11844) );
  INV_X1 U14853 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20782) );
  AND4_X1 U14854 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n20782), .ZN(
        n11847) );
  NAND2_X1 U14855 ( .A1(n11848), .A2(n11847), .ZN(n11849) );
  INV_X1 U14856 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20854) );
  NOR3_X1 U14857 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20854), .ZN(n11851) );
  NOR4_X1 U14858 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n11850) );
  NAND4_X1 U14859 ( .A1(n14482), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n11851), .A4(
        n11850), .ZN(U214) );
  NOR2_X1 U14860 ( .A1(n19543), .A2(n11852), .ZN(n16849) );
  NAND2_X1 U14861 ( .A1(n16849), .A2(U214), .ZN(U212) );
  AOI211_X1 U14862 ( .C1(n16706), .C2(n10594), .A(n12106), .B(n13146), .ZN(
        n11864) );
  XNOR2_X1 U14863 ( .A(n19390), .B(n10594), .ZN(n11853) );
  XNOR2_X1 U14864 ( .A(n12034), .B(n11853), .ZN(n12088) );
  OR2_X1 U14865 ( .A1(n11854), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U14866 ( .A1(n11856), .A2(n11855), .ZN(n12089) );
  OAI22_X1 U14867 ( .A1(n12088), .A2(n16697), .B1(n16710), .B2(n12089), .ZN(
        n11863) );
  OAI22_X1 U14868 ( .A1(n12104), .A2(n16702), .B1(n16695), .B2(n10594), .ZN(
        n11862) );
  NAND2_X1 U14869 ( .A1(n11858), .A2(n11857), .ZN(n11859) );
  NAND2_X1 U14870 ( .A1(n11860), .A2(n11859), .ZN(n20250) );
  INV_X1 U14871 ( .A(n20250), .ZN(n19455) );
  NAND2_X1 U14872 ( .A1(n19529), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12087) );
  OAI21_X1 U14873 ( .B1(n16701), .B2(n19455), .A(n12087), .ZN(n11861) );
  OR4_X1 U14874 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .ZN(
        P2_U3045) );
  INV_X1 U14875 ( .A(n11867), .ZN(n11865) );
  INV_X1 U14876 ( .A(n11066), .ZN(n12241) );
  NAND2_X1 U14877 ( .A1(n11865), .A2(n12241), .ZN(n19382) );
  INV_X1 U14878 ( .A(n19382), .ZN(n19416) );
  INV_X1 U14879 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20291) );
  INV_X1 U14880 ( .A(n13252), .ZN(n11868) );
  OAI211_X1 U14881 ( .C1(n19416), .C2(n20291), .A(n19270), .B(n11868), .ZN(
        P2_U2814) );
  INV_X1 U14882 ( .A(n11349), .ZN(n11871) );
  INV_X1 U14883 ( .A(n19272), .ZN(n20272) );
  INV_X1 U14884 ( .A(n19270), .ZN(n11869) );
  OAI21_X1 U14885 ( .B1(n11869), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20272), 
        .ZN(n11870) );
  OAI21_X1 U14886 ( .B1(n11871), .B2(n20272), .A(n11870), .ZN(P2_U3612) );
  AOI22_X1 U14888 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14889 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11876) );
  NOR2_X4 U14890 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U14891 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11947), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14892 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14893 ( .A1(n12217), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11886) );
  AND2_X4 U14894 ( .A1(n12273), .A2(n11882), .ZN(n14337) );
  AOI22_X1 U14895 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11885) );
  AND2_X2 U14896 ( .A1(n12797), .A2(n12273), .ZN(n11923) );
  AND2_X4 U14897 ( .A1(n11881), .A2(n12800), .ZN(n14357) );
  AOI22_X1 U14898 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14899 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14900 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14901 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14902 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11989), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14903 ( .A1(n12217), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11888) );
  NAND3_X1 U14904 ( .A1(n11892), .A2(n11891), .A3(n11890), .ZN(n11898) );
  AOI22_X1 U14905 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14906 ( .A1(n9683), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11947), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14907 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14908 ( .A1(n14337), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11893) );
  NAND4_X1 U14909 ( .A1(n11896), .A2(n11895), .A3(n11894), .A4(n11893), .ZN(
        n11897) );
  OR2_X4 U14910 ( .A1(n11898), .A2(n11897), .ZN(n12539) );
  AOI22_X1 U14911 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12198), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14912 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14913 ( .A1(n12217), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14914 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11899) );
  NAND4_X1 U14915 ( .A1(n11902), .A2(n11901), .A3(n11900), .A4(n11899), .ZN(
        n11908) );
  AOI22_X1 U14916 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14917 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14918 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14919 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11903) );
  NAND4_X1 U14920 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11907) );
  AOI22_X1 U14921 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U14922 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14923 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14924 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14925 ( .A1(n12217), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U14926 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U14927 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14928 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14929 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12217), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U14930 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U14931 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U14932 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11919) );
  NAND4_X1 U14933 ( .A1(n11922), .A2(n11921), .A3(n11920), .A4(n11919), .ZN(
        n11929) );
  AOI22_X1 U14934 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U14935 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11926) );
  BUF_X4 U14936 ( .A(n11923), .Z(n14358) );
  AOI22_X1 U14937 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14938 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11924) );
  NAND4_X1 U14939 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11928) );
  OR2_X2 U14940 ( .A1(n11929), .A2(n11928), .ZN(n12294) );
  INV_X2 U14941 ( .A(n11979), .ZN(n12061) );
  AND2_X1 U14942 ( .A1(n12539), .A2(n12061), .ZN(n11940) );
  AOI22_X1 U14943 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14219), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14944 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14945 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14946 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11930) );
  NAND4_X1 U14947 ( .A1(n11933), .A2(n11932), .A3(n11931), .A4(n11930), .ZN(
        n11939) );
  AOI22_X1 U14948 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U14949 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U14950 ( .A1(n12217), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U14951 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11934) );
  NAND4_X1 U14952 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n11938) );
  OR2_X2 U14953 ( .A1(n11939), .A2(n11938), .ZN(n12286) );
  NAND2_X1 U14954 ( .A1(n11940), .A2(n11978), .ZN(n11944) );
  NAND2_X1 U14955 ( .A1(n12382), .A2(n12286), .ZN(n11943) );
  OAI21_X1 U14956 ( .B1(n12061), .B2(n12049), .A(n14477), .ZN(n11941) );
  INV_X1 U14957 ( .A(n11941), .ZN(n11942) );
  AOI22_X1 U14958 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14959 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U14960 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U14961 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11949) );
  NAND4_X1 U14962 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(
        n11958) );
  AOI22_X1 U14963 ( .A1(n12217), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11956) );
  BUF_X4 U14964 ( .A(n11989), .Z(n14293) );
  AOI22_X1 U14965 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11953) );
  NAND4_X1 U14966 ( .A1(n11956), .A2(n11955), .A3(n11954), .A4(n11953), .ZN(
        n11957) );
  NOR2_X1 U14967 ( .A1(n12382), .A2(n13019), .ZN(n11959) );
  XNOR2_X1 U14968 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11974) );
  NAND2_X1 U14969 ( .A1(n20693), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12001) );
  NAND2_X1 U14970 ( .A1(n11974), .A2(n11973), .ZN(n11961) );
  NAND2_X1 U14971 ( .A1(n20554), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11960) );
  NAND2_X1 U14972 ( .A1(n11961), .A2(n11960), .ZN(n11976) );
  XNOR2_X1 U14973 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11975) );
  NAND2_X1 U14974 ( .A1(n11976), .A2(n11975), .ZN(n11963) );
  NAND2_X1 U14975 ( .A1(n16151), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11962) );
  NAND2_X1 U14976 ( .A1(n11963), .A2(n11962), .ZN(n11972) );
  MUX2_X1 U14977 ( .A(n11964), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11971) );
  NAND2_X1 U14978 ( .A1(n11972), .A2(n11971), .ZN(n11966) );
  NAND2_X1 U14979 ( .A1(n11964), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11965) );
  NAND2_X1 U14980 ( .A1(n11966), .A2(n11965), .ZN(n11970) );
  NAND2_X1 U14981 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12868), .ZN(
        n11969) );
  NOR2_X1 U14982 ( .A1(n11970), .A2(n11969), .ZN(n12021) );
  XNOR2_X1 U14983 ( .A(n11972), .B(n11971), .ZN(n12017) );
  XNOR2_X1 U14984 ( .A(n11974), .B(n11973), .ZN(n12010) );
  XNOR2_X1 U14985 ( .A(n11976), .B(n11975), .ZN(n11997) );
  OR4_X1 U14986 ( .A1(n12021), .A2(n12017), .A3(n12010), .A4(n11997), .ZN(
        n11977) );
  AND2_X1 U14987 ( .A1(n11996), .A2(n11977), .ZN(n12299) );
  INV_X1 U14988 ( .A(n12299), .ZN(n12068) );
  NOR2_X1 U14989 ( .A1(n12058), .A2(n12068), .ZN(n12043) );
  NAND2_X1 U14990 ( .A1(n12043), .A2(n12534), .ZN(n12031) );
  AND2_X1 U14991 ( .A1(n20658), .A2(n16510), .ZN(n12032) );
  AND2_X2 U14992 ( .A1(n11978), .A2(n12294), .ZN(n12540) );
  NOR2_X1 U14993 ( .A1(n12049), .A2(n12539), .ZN(n12169) );
  INV_X1 U14994 ( .A(n11996), .ZN(n11982) );
  AOI22_X1 U14995 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U14996 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U14997 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U14998 ( .A1(n11988), .A2(n11987), .A3(n11986), .A4(n11985), .ZN(
        n11995) );
  AOI22_X1 U14999 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15000 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15001 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12200), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11990) );
  NAND4_X1 U15002 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11994) );
  INV_X1 U15003 ( .A(n12003), .ZN(n12018) );
  OAI21_X1 U15004 ( .B1(n13024), .B2(n12539), .A(n12059), .ZN(n12015) );
  INV_X1 U15005 ( .A(n11997), .ZN(n11998) );
  OAI21_X1 U15006 ( .B1(n11998), .B2(n13169), .A(n12015), .ZN(n12013) );
  INV_X2 U15007 ( .A(n12539), .ZN(n14478) );
  NAND2_X1 U15008 ( .A1(n14478), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11999) );
  NOR2_X1 U15009 ( .A1(n12010), .A2(n12009), .ZN(n12008) );
  OAI21_X1 U15010 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20693), .A(
        n12001), .ZN(n12004) );
  INV_X1 U15011 ( .A(n12004), .ZN(n12002) );
  OAI211_X1 U15012 ( .C1(n13024), .C2(n12382), .A(n12015), .B(n12002), .ZN(
        n12007) );
  OAI21_X1 U15013 ( .B1(n12005), .B2(n12004), .A(n12003), .ZN(n12006) );
  NAND2_X1 U15014 ( .A1(n12007), .A2(n12006), .ZN(n12011) );
  INV_X1 U15015 ( .A(n12009), .ZN(n12012) );
  NAND2_X1 U15016 ( .A1(n13169), .A2(n12017), .ZN(n12016) );
  INV_X1 U15017 ( .A(n12021), .ZN(n12019) );
  NOR2_X1 U15018 ( .A1(n13044), .A2(n12019), .ZN(n12024) );
  NAND3_X1 U15019 ( .A1(n13044), .A2(n12022), .A3(n12021), .ZN(n12023) );
  OAI21_X1 U15020 ( .B1(n12025), .B2(n12024), .A(n12023), .ZN(n12026) );
  INV_X1 U15021 ( .A(n12392), .ZN(n12029) );
  AOI211_X1 U15022 ( .C1(n12031), .C2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12032), 
        .B(n12029), .ZN(n12030) );
  INV_X1 U15023 ( .A(n12030), .ZN(P1_U2801) );
  INV_X1 U15024 ( .A(n12787), .ZN(n13014) );
  OAI21_X1 U15025 ( .B1(n12032), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13025), 
        .ZN(n12033) );
  OAI21_X1 U15026 ( .B1(n12186), .B2(n13025), .A(n12033), .ZN(P1_U3487) );
  OAI21_X1 U15027 ( .B1(n19402), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12034), .ZN(n16696) );
  INV_X1 U15028 ( .A(n16696), .ZN(n12039) );
  NAND2_X1 U15029 ( .A1(n12035), .A2(n16706), .ZN(n12036) );
  NAND2_X1 U15030 ( .A1(n12037), .A2(n12036), .ZN(n16709) );
  OR2_X1 U15031 ( .A1(n19363), .A2(n19406), .ZN(n16707) );
  OAI21_X1 U15032 ( .B1(n19532), .B2(n16709), .A(n16707), .ZN(n12038) );
  AOI21_X1 U15033 ( .B1(n16662), .B2(n12039), .A(n12038), .ZN(n12042) );
  OAI21_X1 U15034 ( .B1(n19530), .B2(n12040), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12041) );
  OAI211_X1 U15035 ( .C1(n16648), .C2(n19414), .A(n12042), .B(n12041), .ZN(
        P2_U3014) );
  OR2_X1 U15036 ( .A1(n12043), .A2(n16166), .ZN(n12045) );
  OR2_X1 U15037 ( .A1(n12528), .A2(n12787), .ZN(n12044) );
  NAND2_X1 U15038 ( .A1(n12045), .A2(n12044), .ZN(n20294) );
  XNOR2_X1 U15039 ( .A(n20763), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12173) );
  INV_X1 U15040 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U15041 ( .A1(n12173), .A2(n12046), .ZN(n16195) );
  NAND3_X1 U15042 ( .A1(n13014), .A2(n14456), .A3(n16195), .ZN(n12047) );
  NAND2_X1 U15043 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20857) );
  AND2_X1 U15044 ( .A1(n12047), .A2(n20857), .ZN(n20859) );
  NOR2_X1 U15045 ( .A1(n20294), .A2(n20859), .ZN(n16157) );
  OR2_X1 U15046 ( .A1(n16157), .A2(n20293), .ZN(n12072) );
  INV_X1 U15047 ( .A(n12072), .ZN(n20301) );
  INV_X1 U15048 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12074) );
  NAND2_X1 U15049 ( .A1(n14478), .A2(n12061), .ZN(n12048) );
  AND2_X2 U15050 ( .A1(n12048), .A2(n14477), .ZN(n12054) );
  NAND2_X1 U15051 ( .A1(n12050), .A2(n13019), .ZN(n12051) );
  NAND2_X1 U15052 ( .A1(n12182), .A2(n13024), .ZN(n12052) );
  NAND2_X1 U15053 ( .A1(n11918), .A2(n12910), .ZN(n12053) );
  INV_X1 U15054 ( .A(n12382), .ZN(n16155) );
  OAI22_X1 U15055 ( .A1(n12063), .A2(n14454), .B1(n16155), .B2(n13016), .ZN(
        n12055) );
  NOR2_X1 U15056 ( .A1(n12179), .A2(n12055), .ZN(n12321) );
  NAND2_X1 U15057 ( .A1(n16155), .A2(n14419), .ZN(n12057) );
  NAND2_X1 U15058 ( .A1(n12056), .A2(n13019), .ZN(n12318) );
  AND3_X1 U15059 ( .A1(n12176), .A2(n12301), .A3(n9822), .ZN(n12060) );
  NAND2_X1 U15060 ( .A1(n12061), .A2(n14477), .ZN(n14474) );
  AND2_X1 U15061 ( .A1(n14474), .A2(n13019), .ZN(n12300) );
  INV_X1 U15062 ( .A(n12528), .ZN(n12287) );
  INV_X1 U15063 ( .A(n12058), .ZN(n12069) );
  NAND2_X1 U15064 ( .A1(n12272), .A2(n13024), .ZN(n12062) );
  OR2_X1 U15065 ( .A1(n16155), .A2(n12787), .ZN(n12064) );
  NAND2_X1 U15066 ( .A1(n16156), .A2(n12064), .ZN(n12310) );
  NAND3_X1 U15067 ( .A1(n12065), .A2(n12540), .A3(n13019), .ZN(n12066) );
  AOI21_X1 U15068 ( .B1(n12310), .B2(n12066), .A(n12528), .ZN(n12067) );
  AOI21_X1 U15069 ( .B1(n12069), .B2(n12068), .A(n12067), .ZN(n12070) );
  OAI21_X1 U15070 ( .B1(n12786), .B2(n12287), .A(n12070), .ZN(n12071) );
  NAND2_X1 U15071 ( .A1(n12071), .A2(n14477), .ZN(n16159) );
  OR2_X1 U15072 ( .A1(n16159), .A2(n12072), .ZN(n12073) );
  OAI21_X1 U15073 ( .B1(n20301), .B2(n12074), .A(n12073), .ZN(P1_U3484) );
  INV_X1 U15074 ( .A(n15894), .ZN(n12075) );
  OAI21_X1 U15075 ( .B1(n12078), .B2(n12077), .A(n12076), .ZN(n12079) );
  INV_X1 U15076 ( .A(n12079), .ZN(n12123) );
  INV_X1 U15077 ( .A(n12080), .ZN(n12121) );
  NOR2_X1 U15078 ( .A1(n12082), .A2(n12081), .ZN(n12120) );
  NOR3_X1 U15079 ( .A1(n19534), .A2(n12121), .A3(n12120), .ZN(n12085) );
  OAI21_X1 U15080 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n13157), .ZN(n15212) );
  INV_X1 U15081 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20152) );
  OR2_X1 U15082 ( .A1(n19363), .A2(n20152), .ZN(n12114) );
  NAND2_X1 U15083 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12083) );
  OAI211_X1 U15084 ( .C1(n19542), .C2(n15212), .A(n12114), .B(n12083), .ZN(
        n12084) );
  AOI211_X1 U15085 ( .C1(n16660), .C2(n12123), .A(n12085), .B(n12084), .ZN(
        n12086) );
  OAI21_X1 U15086 ( .B1(n12075), .B2(n16648), .A(n12086), .ZN(P2_U3012) );
  INV_X1 U15087 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12092) );
  OAI21_X1 U15088 ( .B1(n19534), .B2(n12088), .A(n12087), .ZN(n12091) );
  OAI22_X1 U15089 ( .A1(n19532), .A2(n12089), .B1(n16666), .B2(n12092), .ZN(
        n12090) );
  AOI211_X1 U15090 ( .C1(n16658), .C2(n12092), .A(n12091), .B(n12090), .ZN(
        n12093) );
  OAI21_X1 U15091 ( .B1(n12104), .B2(n16648), .A(n12093), .ZN(P2_U3013) );
  OAI211_X1 U15092 ( .C1(n9659), .C2(n12095), .A(n12094), .B(n20268), .ZN(
        n12096) );
  MUX2_X1 U15093 ( .A(n12098), .B(n19414), .S(n15291), .Z(n12099) );
  OAI21_X1 U15094 ( .B1(n15298), .B2(n20256), .A(n12099), .ZN(P2_U2887) );
  MUX2_X1 U15095 ( .A(n10366), .B(n12104), .S(n15291), .Z(n12105) );
  OAI21_X1 U15096 ( .B1(n20227), .B2(n15298), .A(n12105), .ZN(P2_U2886) );
  OAI21_X1 U15097 ( .B1(n15743), .B2(n12106), .A(n16695), .ZN(n12119) );
  NOR2_X1 U15098 ( .A1(n12075), .A2(n16702), .ZN(n12118) );
  OAI21_X1 U15099 ( .B1(n12109), .B2(n12108), .A(n12107), .ZN(n20241) );
  INV_X1 U15100 ( .A(n20241), .ZN(n12116) );
  AOI21_X1 U15101 ( .B1(n12112), .B2(n12111), .A(n12110), .ZN(n12113) );
  INV_X1 U15102 ( .A(n12113), .ZN(n12115) );
  OAI211_X1 U15103 ( .C1(n16701), .C2(n12116), .A(n12115), .B(n12114), .ZN(
        n12117) );
  AOI211_X1 U15104 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n12119), .A(
        n12118), .B(n12117), .ZN(n12125) );
  NOR3_X1 U15105 ( .A1(n16697), .A2(n12121), .A3(n12120), .ZN(n12122) );
  AOI21_X1 U15106 ( .B1(n16690), .B2(n12123), .A(n12122), .ZN(n12124) );
  OAI211_X1 U15107 ( .C1(n12127), .C2(n12126), .A(n12125), .B(n12124), .ZN(
        P2_U3044) );
  INV_X1 U15108 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12132) );
  AND2_X1 U15109 ( .A1(n13252), .A2(n20276), .ZN(n12128) );
  INV_X1 U15110 ( .A(n12128), .ZN(n12129) );
  NOR2_X2 U15111 ( .A1(n12129), .A2(n9659), .ZN(n12449) );
  INV_X1 U15112 ( .A(n12449), .ZN(n12131) );
  AOI22_X1 U15113 ( .A1(n19545), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n12447), .ZN(n19429) );
  INV_X1 U15114 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12130) );
  OAI222_X1 U15115 ( .A1(n12132), .A2(n12412), .B1(n12131), .B2(n19429), .C1(
        n12130), .C2(n12366), .ZN(P2_U2982) );
  INV_X1 U15116 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12137) );
  MUX2_X1 U15117 ( .A(n12075), .B(n12137), .S(n15279), .Z(n12138) );
  OAI21_X1 U15118 ( .B1(n20239), .B2(n15298), .A(n12138), .ZN(P2_U2885) );
  INV_X1 U15119 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U15120 ( .A1(n12528), .A2(n12534), .ZN(n12139) );
  INV_X1 U15121 ( .A(n16195), .ZN(n16165) );
  NAND2_X1 U15122 ( .A1(n20396), .A2(n13019), .ZN(n20391) );
  NOR2_X1 U15123 ( .A1(n16510), .A2(n20697), .ZN(n12819) );
  INV_X1 U15124 ( .A(n12819), .ZN(n16506) );
  INV_X2 U15125 ( .A(n20395), .ZN(n20415) );
  AOI22_X1 U15126 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12141) );
  OAI21_X1 U15127 ( .B1(n12142), .B2(n20391), .A(n12141), .ZN(P1_U2918) );
  INV_X1 U15128 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15129 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12143) );
  OAI21_X1 U15130 ( .B1(n12144), .B2(n20391), .A(n12143), .ZN(P1_U2912) );
  INV_X1 U15131 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15132 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12145) );
  OAI21_X1 U15133 ( .B1(n12146), .B2(n20391), .A(n12145), .ZN(P1_U2914) );
  INV_X1 U15134 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15135 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12147) );
  OAI21_X1 U15136 ( .B1(n12148), .B2(n20391), .A(n12147), .ZN(P1_U2906) );
  INV_X1 U15137 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15138 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12149) );
  OAI21_X1 U15139 ( .B1(n12150), .B2(n20391), .A(n12149), .ZN(P1_U2907) );
  INV_X1 U15140 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15141 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12151) );
  OAI21_X1 U15142 ( .B1(n12152), .B2(n20391), .A(n12151), .ZN(P1_U2908) );
  INV_X1 U15143 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15144 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12153) );
  OAI21_X1 U15145 ( .B1(n12154), .B2(n20391), .A(n12153), .ZN(P1_U2916) );
  INV_X1 U15146 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15147 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12155) );
  OAI21_X1 U15148 ( .B1(n12156), .B2(n20391), .A(n12155), .ZN(P1_U2910) );
  INV_X1 U15149 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15150 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12157) );
  OAI21_X1 U15151 ( .B1(n12158), .B2(n20391), .A(n12157), .ZN(P1_U2915) );
  INV_X1 U15152 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15153 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12159) );
  OAI21_X1 U15154 ( .B1(n12160), .B2(n20391), .A(n12159), .ZN(P1_U2913) );
  INV_X1 U15155 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15156 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12161) );
  OAI21_X1 U15157 ( .B1(n12162), .B2(n20391), .A(n12161), .ZN(P1_U2909) );
  INV_X1 U15158 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15159 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12163) );
  OAI21_X1 U15160 ( .B1(n12164), .B2(n20391), .A(n12163), .ZN(P1_U2919) );
  INV_X1 U15161 ( .A(n12294), .ZN(n12675) );
  NAND2_X1 U15162 ( .A1(n12675), .A2(n13019), .ZN(n12753) );
  INV_X1 U15163 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U15164 ( .A1(n14419), .A2(n12166), .ZN(n12165) );
  OAI21_X1 U15165 ( .B1(n12753), .B2(n12166), .A(n12165), .ZN(n12475) );
  INV_X1 U15166 ( .A(n12475), .ZN(n12168) );
  NAND2_X1 U15167 ( .A1(n14405), .A2(n9985), .ZN(n12167) );
  NAND2_X1 U15168 ( .A1(n12168), .A2(n12167), .ZN(n13083) );
  NAND4_X1 U15169 ( .A1(n12788), .A2(n12169), .A3(n14498), .A4(n12061), .ZN(
        n12531) );
  NAND2_X1 U15170 ( .A1(n12291), .A2(n12170), .ZN(n12171) );
  INV_X1 U15171 ( .A(n12788), .ZN(n12175) );
  NAND2_X1 U15172 ( .A1(n12174), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12268) );
  NAND2_X1 U15173 ( .A1(n12183), .A2(n12272), .ZN(n12177) );
  NAND4_X1 U15174 ( .A1(n12177), .A2(n12176), .A3(n13016), .A4(n12175), .ZN(
        n12178) );
  MUX2_X1 U15175 ( .A(n12337), .B(n12265), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12181) );
  INV_X1 U15176 ( .A(n12197), .ZN(n12195) );
  OAI21_X1 U15177 ( .B1(n13024), .B2(n12286), .A(n12182), .ZN(n12193) );
  NAND2_X1 U15178 ( .A1(n9929), .A2(n13657), .ZN(n12190) );
  NAND2_X1 U15179 ( .A1(n12050), .A2(n12294), .ZN(n12185) );
  NAND2_X1 U15180 ( .A1(n12186), .A2(n12185), .ZN(n12189) );
  NAND2_X1 U15181 ( .A1(n13007), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20296) );
  INV_X1 U15182 ( .A(n20296), .ZN(n12187) );
  AND2_X1 U15183 ( .A1(n13016), .A2(n12187), .ZN(n12188) );
  NAND2_X1 U15184 ( .A1(n12788), .A2(n12905), .ZN(n12319) );
  NAND3_X1 U15185 ( .A1(n12193), .A2(n12192), .A3(n12191), .ZN(n12196) );
  INV_X1 U15186 ( .A(n12196), .ZN(n12194) );
  AOI22_X1 U15187 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15188 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15189 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15190 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12201) );
  NAND4_X1 U15191 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12210) );
  AOI22_X1 U15192 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15193 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15194 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15195 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12205) );
  NAND4_X1 U15196 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12209) );
  AOI22_X1 U15197 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15198 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15199 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15200 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12213) );
  NAND4_X1 U15201 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12225) );
  AOI22_X1 U15202 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15203 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15204 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15205 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12220) );
  NAND4_X1 U15206 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12224) );
  NAND2_X1 U15207 ( .A1(n12495), .A2(n13644), .ZN(n12501) );
  NOR2_X1 U15208 ( .A1(n12226), .A2(n12617), .ZN(n12227) );
  INV_X1 U15209 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12230) );
  AOI21_X1 U15210 ( .B1(n12910), .B2(n13656), .A(n16503), .ZN(n12229) );
  NAND2_X1 U15211 ( .A1(n13024), .A2(n12617), .ZN(n12228) );
  OAI211_X1 U15212 ( .C1(n13169), .C2(n12230), .A(n12229), .B(n12228), .ZN(
        n12493) );
  INV_X1 U15213 ( .A(n12233), .ZN(n13088) );
  NAND2_X1 U15214 ( .A1(n13088), .A2(n13859), .ZN(n12237) );
  INV_X1 U15215 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n12234) );
  INV_X1 U15216 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13084) );
  OAI22_X1 U15217 ( .A1(n14285), .A2(n12234), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13084), .ZN(n12235) );
  AOI21_X1 U15218 ( .B1(n12865), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12235), .ZN(n12236) );
  NAND2_X1 U15219 ( .A1(n12237), .A2(n12236), .ZN(n12476) );
  NAND2_X1 U15220 ( .A1(n12238), .A2(n12476), .ZN(n12480) );
  OAI21_X1 U15221 ( .B1(n12238), .B2(n12476), .A(n12480), .ZN(n13090) );
  OAI222_X1 U15222 ( .A1(n13083), .A2(n20385), .B1(n12166), .B2(n20390), .C1(
        n13090), .C2(n14666), .ZN(P1_U2872) );
  INV_X1 U15223 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15224 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12239) );
  OAI21_X1 U15225 ( .B1(n12240), .B2(n20391), .A(n12239), .ZN(P1_U2920) );
  NAND2_X1 U15226 ( .A1(n12242), .A2(n12241), .ZN(n15860) );
  OAI21_X1 U15227 ( .B1(n15860), .B2(n12243), .A(n12366), .ZN(n12244) );
  NAND2_X1 U15228 ( .A1(n19494), .A2(n12245), .ZN(n12263) );
  NAND2_X1 U15229 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20253) );
  NOR2_X1 U15230 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20253), .ZN(n19525) );
  INV_X1 U15231 ( .A(n19525), .ZN(n20273) );
  INV_X2 U15232 ( .A(n19509), .ZN(n19524) );
  AOI22_X1 U15233 ( .A1(n19521), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12246) );
  OAI21_X1 U15234 ( .B1(n21039), .B2(n12263), .A(n12246), .ZN(P2_U2923) );
  AOI22_X1 U15235 ( .A1(n19521), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12247) );
  OAI21_X1 U15236 ( .B1(n13403), .B2(n12263), .A(n12247), .ZN(P2_U2935) );
  INV_X1 U15237 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U15238 ( .A1(n19521), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12248) );
  OAI21_X1 U15239 ( .B1(n15346), .B2(n12263), .A(n12248), .ZN(P2_U2927) );
  INV_X1 U15240 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U15241 ( .A1(n19521), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12249) );
  OAI21_X1 U15242 ( .B1(n15365), .B2(n12263), .A(n12249), .ZN(P2_U2931) );
  INV_X1 U15243 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15356) );
  AOI22_X1 U15244 ( .A1(n19521), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12250) );
  OAI21_X1 U15245 ( .B1(n15356), .B2(n12263), .A(n12250), .ZN(P2_U2930) );
  INV_X1 U15246 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U15247 ( .A1(n19525), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12251) );
  OAI21_X1 U15248 ( .B1(n15370), .B2(n12263), .A(n12251), .ZN(P2_U2932) );
  INV_X1 U15249 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15250 ( .A1(n19521), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12252) );
  OAI21_X1 U15251 ( .B1(n12358), .B2(n12263), .A(n12252), .ZN(P2_U2922) );
  AOI22_X1 U15252 ( .A1(n19521), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12253) );
  OAI21_X1 U15253 ( .B1(n12254), .B2(n12263), .A(n12253), .ZN(P2_U2921) );
  INV_X1 U15254 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15255 ( .A1(n19521), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12255) );
  OAI21_X1 U15256 ( .B1(n12363), .B2(n12263), .A(n12255), .ZN(P2_U2926) );
  INV_X1 U15257 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15327) );
  AOI22_X1 U15258 ( .A1(n19521), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12256) );
  OAI21_X1 U15259 ( .B1(n15327), .B2(n12263), .A(n12256), .ZN(P2_U2925) );
  INV_X1 U15260 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15261 ( .A1(n19521), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12257) );
  OAI21_X1 U15262 ( .B1(n12354), .B2(n12263), .A(n12257), .ZN(P2_U2924) );
  INV_X1 U15263 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15264 ( .A1(n19521), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12258) );
  OAI21_X1 U15265 ( .B1(n12259), .B2(n12263), .A(n12258), .ZN(P2_U2929) );
  INV_X1 U15266 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U15267 ( .A1(n19525), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12260) );
  OAI21_X1 U15268 ( .B1(n13583), .B2(n12263), .A(n12260), .ZN(P2_U2933) );
  INV_X1 U15269 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U15270 ( .A1(n19525), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12261) );
  OAI21_X1 U15271 ( .B1(n13434), .B2(n12263), .A(n12261), .ZN(P2_U2934) );
  INV_X1 U15272 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15273 ( .A1(n19521), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12262) );
  OAI21_X1 U15274 ( .B1(n12264), .B2(n12263), .A(n12262), .ZN(P2_U2928) );
  NAND2_X1 U15275 ( .A1(n12334), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12267) );
  NAND2_X1 U15276 ( .A1(n20554), .A2(n20693), .ZN(n20585) );
  NAND2_X1 U15277 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12942) );
  AND2_X1 U15278 ( .A1(n20585), .A2(n12942), .ZN(n20523) );
  AOI21_X1 U15279 ( .B1(n20523), .B2(n12384), .A(n12328), .ZN(n12266) );
  NAND2_X1 U15280 ( .A1(n12267), .A2(n12266), .ZN(n12270) );
  INV_X1 U15281 ( .A(n12268), .ZN(n12269) );
  OR2_X2 U15282 ( .A1(n12678), .A2(n12271), .ZN(n12333) );
  NAND2_X1 U15283 ( .A1(n12678), .A2(n12271), .ZN(n20553) );
  INV_X1 U15284 ( .A(n20591), .ZN(n20521) );
  INV_X1 U15285 ( .A(n12791), .ZN(n12809) );
  NAND2_X1 U15286 ( .A1(n20521), .A2(n12809), .ZN(n12276) );
  INV_X1 U15287 ( .A(n12273), .ZN(n12813) );
  INV_X1 U15288 ( .A(n12800), .ZN(n12274) );
  NAND3_X1 U15289 ( .A1(n14091), .A2(n12813), .A3(n12274), .ZN(n12275) );
  OAI211_X1 U15290 ( .C1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n12804), .A(
        n12276), .B(n12275), .ZN(n16146) );
  INV_X1 U15291 ( .A(n15028), .ZN(n16172) );
  NAND2_X1 U15292 ( .A1(n12813), .A2(n16172), .ZN(n12278) );
  INV_X1 U15293 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20500) );
  INV_X1 U15294 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15295 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20500), .B2(n12277), .ZN(
        n15022) );
  NAND2_X1 U15296 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15021) );
  OAI22_X1 U15297 ( .A1(n12278), .A2(n12800), .B1(n15022), .B2(n15021), .ZN(
        n12279) );
  AOI21_X1 U15298 ( .B1(n16146), .B2(n13007), .A(n12279), .ZN(n12293) );
  NAND2_X1 U15299 ( .A1(n12804), .A2(n12301), .ZN(n12282) );
  INV_X1 U15300 ( .A(n20857), .ZN(n20773) );
  AOI21_X1 U15301 ( .B1(n12280), .B2(n16195), .A(n20773), .ZN(n12281) );
  NAND3_X1 U15302 ( .A1(n12282), .A2(n12528), .A3(n12281), .ZN(n12285) );
  NAND2_X1 U15303 ( .A1(n16156), .A2(n12283), .ZN(n12284) );
  NAND2_X1 U15304 ( .A1(n12058), .A2(n12284), .ZN(n12308) );
  OAI211_X1 U15305 ( .C1(n13016), .C2(n12286), .A(n12285), .B(n12308), .ZN(
        n12289) );
  NAND2_X1 U15306 ( .A1(n12299), .A2(n20857), .ZN(n12288) );
  NAND2_X1 U15307 ( .A1(n16156), .A2(n12787), .ZN(n12785) );
  OAI22_X1 U15308 ( .A1(n12172), .A2(n12288), .B1(n12287), .B2(n12785), .ZN(
        n12533) );
  NOR2_X1 U15309 ( .A1(n12289), .A2(n12533), .ZN(n12290) );
  INV_X1 U15310 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20300) );
  NAND2_X1 U15311 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12819), .ZN(n16511) );
  OAI22_X1 U15312 ( .A1(n12814), .A2(n20293), .B1(n20300), .B2(n16511), .ZN(
        n12344) );
  AOI21_X1 U15313 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n16503), .A(n12344), 
        .ZN(n15032) );
  NAND2_X1 U15314 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n15032), .ZN(
        n12292) );
  OAI21_X1 U15315 ( .B1(n12293), .B2(n15032), .A(n12292), .ZN(P1_U3473) );
  NAND2_X1 U15316 ( .A1(n13024), .A2(n12294), .ZN(n12620) );
  OAI21_X1 U15317 ( .B1(n20860), .B2(n12617), .A(n12620), .ZN(n12295) );
  INV_X1 U15318 ( .A(n12295), .ZN(n12296) );
  OAI21_X1 U15319 ( .B1(n12297), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12545), .ZN(n12386) );
  NAND2_X1 U15320 ( .A1(n12299), .A2(n12298), .ZN(n12304) );
  OAI21_X1 U15321 ( .B1(n12301), .B2(n13018), .A(n12300), .ZN(n12302) );
  NAND2_X1 U15322 ( .A1(n12302), .A2(n12528), .ZN(n12303) );
  MUX2_X1 U15323 ( .A(n12304), .B(n12303), .S(n11978), .Z(n12307) );
  OR2_X1 U15324 ( .A1(n12305), .A2(n12528), .ZN(n12306) );
  NAND3_X1 U15325 ( .A1(n12308), .A2(n12307), .A3(n12306), .ZN(n12309) );
  INV_X1 U15326 ( .A(n12323), .ZN(n12313) );
  OAI211_X1 U15327 ( .C1(n12910), .C2(n9821), .A(n12311), .B(n12310), .ZN(
        n12312) );
  NOR2_X1 U15328 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12314) );
  INV_X1 U15329 ( .A(n16482), .ZN(n16489) );
  NAND2_X1 U15330 ( .A1(n16489), .A2(n12323), .ZN(n20506) );
  AOI21_X1 U15331 ( .B1(n14902), .B2(n20506), .A(n9985), .ZN(n12326) );
  AOI22_X1 U15332 ( .A1(n16166), .A2(n12059), .B1(n12910), .B2(n12315), .ZN(
        n12316) );
  NOR2_X1 U15333 ( .A1(n20503), .A2(n13083), .ZN(n12325) );
  INV_X1 U15334 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n12317) );
  NOR2_X1 U15335 ( .A1(n16489), .A2(n12317), .ZN(n12388) );
  AND2_X1 U15336 ( .A1(n12319), .A2(n12318), .ZN(n12320) );
  AND2_X1 U15337 ( .A1(n12321), .A2(n12320), .ZN(n12322) );
  AND2_X1 U15338 ( .A1(n20498), .A2(n13727), .ZN(n20507) );
  NOR2_X1 U15339 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20507), .ZN(
        n12324) );
  NOR4_X1 U15340 ( .A1(n12326), .A2(n12325), .A3(n12388), .A4(n12324), .ZN(
        n12327) );
  OAI21_X1 U15341 ( .B1(n12386), .B2(n16457), .A(n12327), .ZN(P1_U3031) );
  INV_X1 U15342 ( .A(n12328), .ZN(n12330) );
  AND2_X1 U15343 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  NAND2_X2 U15344 ( .A1(n12333), .A2(n12332), .ZN(n12584) );
  XNOR2_X1 U15345 ( .A(n12942), .B(n16151), .ZN(n13107) );
  NAND2_X1 U15346 ( .A1(n12334), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12336) );
  NAND2_X1 U15347 ( .A1(n12340), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12335) );
  NAND2_X1 U15348 ( .A1(n12334), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12342) );
  OAI21_X1 U15349 ( .B1(n12942), .B2(n16151), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12339) );
  INV_X1 U15350 ( .A(n12942), .ZN(n12712) );
  NAND2_X1 U15351 ( .A1(n11964), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20615) );
  INV_X1 U15352 ( .A(n20615), .ZN(n12338) );
  NAND2_X1 U15353 ( .A1(n12712), .A2(n12338), .ZN(n12932) );
  NAND2_X1 U15354 ( .A1(n12339), .A2(n12932), .ZN(n20524) );
  AOI22_X1 U15355 ( .A1(n20524), .A2(n12384), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12340), .ZN(n12341) );
  INV_X1 U15356 ( .A(n12762), .ZN(n12710) );
  NOR2_X1 U15357 ( .A1(n12657), .A2(n12710), .ZN(n12343) );
  XNOR2_X1 U15358 ( .A(n12343), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20365) );
  INV_X1 U15359 ( .A(n12172), .ZN(n12345) );
  NAND3_X1 U15360 ( .A1(n12345), .A2(n13007), .A3(n12344), .ZN(n12347) );
  INV_X1 U15361 ( .A(n15032), .ZN(n12346) );
  OAI22_X1 U15362 ( .A1(n20365), .A2(n12347), .B1(n12868), .B2(n12346), .ZN(
        P1_U3468) );
  INV_X1 U15363 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19507) );
  NAND2_X1 U15364 ( .A1(n12464), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12350) );
  NAND2_X1 U15365 ( .A1(n19543), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12349) );
  INV_X1 U15366 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16879) );
  OR2_X1 U15367 ( .A1(n19543), .A2(n16879), .ZN(n12348) );
  NAND2_X1 U15368 ( .A1(n12349), .A2(n12348), .ZN(n19447) );
  NAND2_X1 U15369 ( .A1(n12449), .A2(n19447), .ZN(n12361) );
  OAI211_X1 U15370 ( .C1(n19507), .C2(n12366), .A(n12350), .B(n12361), .ZN(
        P2_U2976) );
  NAND2_X1 U15371 ( .A1(n12464), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12353) );
  NAND2_X1 U15372 ( .A1(n19543), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12352) );
  INV_X1 U15373 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16876) );
  OR2_X1 U15374 ( .A1(n19543), .A2(n16876), .ZN(n12351) );
  NAND2_X1 U15375 ( .A1(n12352), .A2(n12351), .ZN(n19440) );
  NAND2_X1 U15376 ( .A1(n12449), .A2(n19440), .ZN(n12359) );
  OAI211_X1 U15377 ( .C1(n12354), .C2(n12366), .A(n12353), .B(n12359), .ZN(
        P2_U2963) );
  NAND2_X1 U15378 ( .A1(n12464), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12357) );
  NAND2_X1 U15379 ( .A1(n19543), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12356) );
  INV_X1 U15380 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16872) );
  OR2_X1 U15381 ( .A1(n19543), .A2(n16872), .ZN(n12355) );
  NAND2_X1 U15382 ( .A1(n12356), .A2(n12355), .ZN(n19433) );
  NAND2_X1 U15383 ( .A1(n12449), .A2(n19433), .ZN(n12364) );
  OAI211_X1 U15384 ( .C1(n12358), .C2(n12366), .A(n12357), .B(n12364), .ZN(
        P2_U2965) );
  INV_X1 U15385 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19503) );
  NAND2_X1 U15386 ( .A1(n12464), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12360) );
  OAI211_X1 U15387 ( .C1(n19503), .C2(n12366), .A(n12360), .B(n12359), .ZN(
        P2_U2978) );
  NAND2_X1 U15388 ( .A1(n12464), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12362) );
  OAI211_X1 U15389 ( .C1(n12363), .C2(n12366), .A(n12362), .B(n12361), .ZN(
        P2_U2961) );
  INV_X1 U15390 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19499) );
  NAND2_X1 U15391 ( .A1(n12464), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n12365) );
  OAI211_X1 U15392 ( .C1(n19499), .C2(n12366), .A(n12365), .B(n12364), .ZN(
        P2_U2980) );
  OAI21_X1 U15393 ( .B1(n12369), .B2(n12368), .A(n12405), .ZN(n19466) );
  NAND2_X1 U15394 ( .A1(n12371), .A2(n12370), .ZN(n12372) );
  AND2_X1 U15395 ( .A1(n12407), .A2(n12372), .ZN(n19537) );
  INV_X1 U15396 ( .A(n19537), .ZN(n19381) );
  INV_X1 U15397 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12373) );
  MUX2_X1 U15398 ( .A(n19381), .B(n12373), .S(n15279), .Z(n12374) );
  OAI21_X1 U15399 ( .B1(n19466), .B2(n15298), .A(n12374), .ZN(P2_U2883) );
  AOI22_X1 U15400 ( .A1(n13088), .A2(n12809), .B1(n14091), .B2(n12376), .ZN(
        n16142) );
  OAI21_X1 U15401 ( .B1(n16142), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n16510), 
        .ZN(n12375) );
  AOI22_X1 U15402 ( .A1(n12375), .A2(n15021), .B1(n12376), .B2(n16172), .ZN(
        n12378) );
  NOR2_X1 U15403 ( .A1(n12804), .A2(n12376), .ZN(n16143) );
  AOI22_X1 U15404 ( .A1(n16143), .A2(n13007), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15032), .ZN(n12377) );
  OAI21_X1 U15405 ( .B1(n12378), .B2(n15032), .A(n12377), .ZN(P1_U3474) );
  AOI22_X1 U15406 ( .A1(n12464), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n12463), .ZN(n12380) );
  AOI22_X1 U15407 ( .A1(n19545), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19543), .ZN(n19437) );
  INV_X1 U15408 ( .A(n19437), .ZN(n12379) );
  NAND2_X1 U15409 ( .A1(n12449), .A2(n12379), .ZN(n12457) );
  NAND2_X1 U15410 ( .A1(n12380), .A2(n12457), .ZN(P2_U2979) );
  NAND2_X1 U15411 ( .A1(n20702), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13008) );
  NAND2_X1 U15412 ( .A1(n16503), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12381) );
  AND2_X1 U15413 ( .A1(n13008), .A2(n12381), .ZN(n12547) );
  NOR2_X1 U15414 ( .A1(n12382), .A2(n20293), .ZN(n12383) );
  OR2_X1 U15415 ( .A1(n12384), .A2(n20622), .ZN(n20856) );
  AND2_X1 U15416 ( .A1(n20856), .A2(n16503), .ZN(n12385) );
  NAND2_X1 U15417 ( .A1(n12547), .A2(n16333), .ZN(n12389) );
  NOR2_X1 U15418 ( .A1(n12386), .A2(n20299), .ZN(n12387) );
  AOI211_X1 U15419 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n12389), .A(
        n12388), .B(n12387), .ZN(n12390) );
  OAI21_X1 U15420 ( .B1(n14888), .B2(n13090), .A(n12390), .ZN(P1_U2999) );
  AND2_X1 U15421 ( .A1(n20860), .A2(n20773), .ZN(n12391) );
  INV_X1 U15422 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12397) );
  INV_X1 U15423 ( .A(n20432), .ZN(n12396) );
  INV_X1 U15424 ( .A(n14482), .ZN(n14475) );
  INV_X1 U15425 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12393) );
  NOR2_X1 U15426 ( .A1(n14475), .A2(n12393), .ZN(n12394) );
  AOI21_X1 U15427 ( .B1(DATAI_15_), .B2(n14475), .A(n12394), .ZN(n14736) );
  INV_X1 U15428 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12395) );
  OAI222_X1 U15429 ( .A1(n9773), .A2(n12397), .B1(n12396), .B2(n14736), .C1(
        n12395), .C2(n12515), .ZN(P1_U2967) );
  NOR2_X1 U15430 ( .A1(n9891), .A2(n15279), .ZN(n12402) );
  AOI21_X1 U15431 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n15279), .A(n12402), .ZN(
        n12403) );
  OAI21_X1 U15432 ( .B1(n19860), .B2(n15298), .A(n12403), .ZN(P2_U2884) );
  OR2_X1 U15433 ( .A1(n12405), .A2(n12404), .ZN(n12553) );
  OAI211_X1 U15434 ( .C1(n12367), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15281), .B(n12553), .ZN(n12410) );
  AND2_X1 U15435 ( .A1(n12407), .A2(n12406), .ZN(n12408) );
  OR2_X1 U15436 ( .A1(n12408), .A2(n12557), .ZN(n13451) );
  INV_X1 U15437 ( .A(n13451), .ZN(n16659) );
  NAND2_X1 U15438 ( .A1(n16659), .A2(n15291), .ZN(n12409) );
  OAI211_X1 U15439 ( .C1(n15291), .C2(n12411), .A(n12410), .B(n12409), .ZN(
        P2_U2882) );
  INV_X2 U15440 ( .A(n12412), .ZN(n12464) );
  AOI22_X1 U15441 ( .A1(n12464), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n12463), .ZN(n12413) );
  OAI22_X1 U15442 ( .A1(n19543), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19545), .ZN(n19580) );
  INV_X1 U15443 ( .A(n19580), .ZN(n16617) );
  NAND2_X1 U15444 ( .A1(n12449), .A2(n16617), .ZN(n12437) );
  NAND2_X1 U15445 ( .A1(n12413), .A2(n12437), .ZN(P2_U2958) );
  AOI22_X1 U15446 ( .A1(n12464), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n12463), .ZN(n12415) );
  AOI22_X1 U15447 ( .A1(n19545), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n12447), .ZN(n19570) );
  INV_X1 U15448 ( .A(n19570), .ZN(n12414) );
  NAND2_X1 U15449 ( .A1(n12449), .A2(n12414), .ZN(n12445) );
  NAND2_X1 U15450 ( .A1(n12415), .A2(n12445), .ZN(P2_U2955) );
  AOI22_X1 U15451 ( .A1(n12464), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15452 ( .A1(n19545), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n12447), .ZN(n19574) );
  INV_X1 U15453 ( .A(n19574), .ZN(n12416) );
  NAND2_X1 U15454 ( .A1(n12449), .A2(n12416), .ZN(n12443) );
  NAND2_X1 U15455 ( .A1(n12417), .A2(n12443), .ZN(P2_U2956) );
  AOI22_X1 U15456 ( .A1(n12464), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n12463), .ZN(n12419) );
  AOI22_X1 U15457 ( .A1(n19545), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n12447), .ZN(n19560) );
  INV_X1 U15458 ( .A(n19560), .ZN(n12418) );
  NAND2_X1 U15459 ( .A1(n12449), .A2(n12418), .ZN(n12465) );
  NAND2_X1 U15460 ( .A1(n12419), .A2(n12465), .ZN(P2_U2953) );
  AOI22_X1 U15461 ( .A1(n12464), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15462 ( .A1(n19545), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19543), .ZN(n19553) );
  INV_X1 U15463 ( .A(n19553), .ZN(n12420) );
  NAND2_X1 U15464 ( .A1(n12449), .A2(n12420), .ZN(n12453) );
  NAND2_X1 U15465 ( .A1(n12421), .A2(n12453), .ZN(P2_U2952) );
  AOI22_X1 U15466 ( .A1(n12464), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n12463), .ZN(n12426) );
  INV_X1 U15467 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n12422) );
  OR2_X1 U15468 ( .A1(n19543), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U15469 ( .A1(n19543), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12423) );
  AND2_X1 U15470 ( .A1(n12424), .A2(n12423), .ZN(n19443) );
  INV_X1 U15471 ( .A(n19443), .ZN(n12425) );
  NAND2_X1 U15472 ( .A1(n12449), .A2(n12425), .ZN(n12459) );
  NAND2_X1 U15473 ( .A1(n12426), .A2(n12459), .ZN(P2_U2977) );
  AOI22_X1 U15474 ( .A1(n12464), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n12463), .ZN(n12431) );
  INV_X1 U15475 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n12427) );
  OR2_X1 U15476 ( .A1(n19543), .A2(n12427), .ZN(n12429) );
  NAND2_X1 U15477 ( .A1(n19543), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12428) );
  AND2_X1 U15478 ( .A1(n12429), .A2(n12428), .ZN(n19450) );
  INV_X1 U15479 ( .A(n19450), .ZN(n12430) );
  NAND2_X1 U15480 ( .A1(n12449), .A2(n12430), .ZN(n12455) );
  NAND2_X1 U15481 ( .A1(n12431), .A2(n12455), .ZN(P2_U2975) );
  AOI22_X1 U15482 ( .A1(n12464), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n12463), .ZN(n12433) );
  AOI22_X1 U15483 ( .A1(n19545), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n12447), .ZN(n19577) );
  INV_X1 U15484 ( .A(n19577), .ZN(n12432) );
  NAND2_X1 U15485 ( .A1(n12449), .A2(n12432), .ZN(n12439) );
  NAND2_X1 U15486 ( .A1(n12433), .A2(n12439), .ZN(P2_U2957) );
  AOI22_X1 U15487 ( .A1(n12464), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n12463), .ZN(n12434) );
  OAI22_X1 U15488 ( .A1(n19543), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19545), .ZN(n19592) );
  INV_X1 U15489 ( .A(n19592), .ZN(n16611) );
  NAND2_X1 U15490 ( .A1(n12449), .A2(n16611), .ZN(n12435) );
  NAND2_X1 U15491 ( .A1(n12434), .A2(n12435), .ZN(P2_U2959) );
  AOI22_X1 U15492 ( .A1(n12464), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n12463), .ZN(n12436) );
  NAND2_X1 U15493 ( .A1(n12436), .A2(n12435), .ZN(P2_U2974) );
  AOI22_X1 U15494 ( .A1(n12464), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n12463), .ZN(n12438) );
  NAND2_X1 U15495 ( .A1(n12438), .A2(n12437), .ZN(P2_U2973) );
  AOI22_X1 U15496 ( .A1(n12464), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n12463), .ZN(n12440) );
  NAND2_X1 U15497 ( .A1(n12440), .A2(n12439), .ZN(P2_U2972) );
  AOI22_X1 U15498 ( .A1(n12464), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n12463), .ZN(n12442) );
  INV_X1 U15499 ( .A(n19431), .ZN(n12441) );
  NAND2_X1 U15500 ( .A1(n12449), .A2(n12441), .ZN(n12451) );
  NAND2_X1 U15501 ( .A1(n12442), .A2(n12451), .ZN(P2_U2966) );
  AOI22_X1 U15502 ( .A1(n12464), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12444) );
  NAND2_X1 U15503 ( .A1(n12444), .A2(n12443), .ZN(P2_U2971) );
  AOI22_X1 U15504 ( .A1(n12464), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12446) );
  NAND2_X1 U15505 ( .A1(n12446), .A2(n12445), .ZN(P2_U2970) );
  AOI22_X1 U15506 ( .A1(n12464), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15507 ( .A1(n19545), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n12447), .ZN(n19565) );
  INV_X1 U15508 ( .A(n19565), .ZN(n12448) );
  NAND2_X1 U15509 ( .A1(n12449), .A2(n12448), .ZN(n12461) );
  NAND2_X1 U15510 ( .A1(n12450), .A2(n12461), .ZN(P2_U2969) );
  AOI22_X1 U15511 ( .A1(n12464), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n12463), .ZN(n12452) );
  NAND2_X1 U15512 ( .A1(n12452), .A2(n12451), .ZN(P2_U2981) );
  AOI22_X1 U15513 ( .A1(n12464), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n12454) );
  NAND2_X1 U15514 ( .A1(n12454), .A2(n12453), .ZN(P2_U2967) );
  AOI22_X1 U15515 ( .A1(n12464), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n12463), .ZN(n12456) );
  NAND2_X1 U15516 ( .A1(n12456), .A2(n12455), .ZN(P2_U2960) );
  AOI22_X1 U15517 ( .A1(n12464), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n12463), .ZN(n12458) );
  NAND2_X1 U15518 ( .A1(n12458), .A2(n12457), .ZN(P2_U2964) );
  AOI22_X1 U15519 ( .A1(n12464), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n12463), .ZN(n12460) );
  NAND2_X1 U15520 ( .A1(n12460), .A2(n12459), .ZN(P2_U2962) );
  AOI22_X1 U15521 ( .A1(n12464), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U15522 ( .A1(n12462), .A2(n12461), .ZN(P2_U2954) );
  AOI22_X1 U15523 ( .A1(n12464), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n12463), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U15524 ( .A1(n12466), .A2(n12465), .ZN(P2_U2968) );
  AND2_X1 U15525 ( .A1(n12367), .A2(n12467), .ZN(n12841) );
  XNOR2_X1 U15526 ( .A(n12841), .B(n12468), .ZN(n12473) );
  NAND2_X1 U15527 ( .A1(n12837), .A2(n12469), .ZN(n12470) );
  NAND2_X1 U15528 ( .A1(n12564), .A2(n12470), .ZN(n16639) );
  MUX2_X1 U15529 ( .A(n12471), .B(n16639), .S(n15291), .Z(n12472) );
  OAI21_X1 U15530 ( .B1(n12473), .B2(n15298), .A(n12472), .ZN(P2_U2878) );
  NAND2_X1 U15531 ( .A1(n14405), .A2(n20500), .ZN(n12474) );
  XNOR2_X1 U15532 ( .A(n13074), .B(n14456), .ZN(n20502) );
  INV_X1 U15533 ( .A(n12476), .ZN(n12478) );
  NAND2_X1 U15534 ( .A1(n12478), .A2(n14345), .ZN(n12479) );
  NAND2_X1 U15535 ( .A1(n12480), .A2(n12479), .ZN(n12508) );
  AOI22_X1 U15536 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15537 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11948), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15538 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15539 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12481) );
  NAND4_X1 U15540 ( .A1(n12484), .A2(n12483), .A3(n12482), .A4(n12481), .ZN(
        n12490) );
  AOI22_X1 U15541 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15542 ( .A1(n14338), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15543 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15544 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12485) );
  NAND4_X1 U15545 ( .A1(n12488), .A2(n12487), .A3(n12486), .A4(n12485), .ZN(
        n12489) );
  NAND2_X1 U15546 ( .A1(n12495), .A2(n12618), .ZN(n12491) );
  NAND2_X1 U15547 ( .A1(n12495), .A2(n13656), .ZN(n13652) );
  XNOR2_X1 U15548 ( .A(n12577), .B(n12578), .ZN(n12502) );
  NAND2_X1 U15549 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12500) );
  INV_X1 U15550 ( .A(n12497), .ZN(n12498) );
  NAND2_X1 U15551 ( .A1(n12498), .A2(n12618), .ZN(n12499) );
  NAND2_X1 U15552 ( .A1(n15009), .A2(n13859), .ZN(n12506) );
  INV_X1 U15553 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12503) );
  INV_X1 U15554 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13078) );
  OAI22_X1 U15555 ( .A1(n14285), .A2(n12503), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13078), .ZN(n12504) );
  AOI21_X1 U15556 ( .B1(n12865), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12504), .ZN(n12505) );
  NAND2_X1 U15557 ( .A1(n12506), .A2(n12505), .ZN(n12507) );
  NAND2_X1 U15558 ( .A1(n12508), .A2(n12507), .ZN(n12609) );
  OAI21_X1 U15559 ( .B1(n12508), .B2(n12507), .A(n12609), .ZN(n13080) );
  OAI222_X1 U15560 ( .A1(n20502), .A2(n20385), .B1(n9997), .B2(n20390), .C1(
        n13080), .C2(n14666), .ZN(P1_U2871) );
  AOI22_X1 U15561 ( .A1(n20447), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20442), .ZN(n12511) );
  NAND2_X1 U15562 ( .A1(n14475), .A2(DATAI_5_), .ZN(n12510) );
  NAND2_X1 U15563 ( .A1(n14482), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12509) );
  AND2_X1 U15564 ( .A1(n12510), .A2(n12509), .ZN(n12974) );
  INV_X1 U15565 ( .A(n12974), .ZN(n14706) );
  NAND2_X1 U15566 ( .A1(n20432), .A2(n14706), .ZN(n12647) );
  NAND2_X1 U15567 ( .A1(n12511), .A2(n12647), .ZN(P1_U2957) );
  AOI22_X1 U15568 ( .A1(n20447), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20442), .ZN(n12514) );
  NAND2_X1 U15569 ( .A1(n14475), .A2(DATAI_4_), .ZN(n12513) );
  NAND2_X1 U15570 ( .A1(n14482), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12512) );
  AND2_X1 U15571 ( .A1(n12513), .A2(n12512), .ZN(n12973) );
  INV_X1 U15572 ( .A(n12973), .ZN(n14711) );
  NAND2_X1 U15573 ( .A1(n20432), .A2(n14711), .ZN(n12639) );
  NAND2_X1 U15574 ( .A1(n12514), .A2(n12639), .ZN(P1_U2956) );
  AOI22_X1 U15575 ( .A1(n20447), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20442), .ZN(n12518) );
  NAND2_X1 U15576 ( .A1(n14475), .A2(DATAI_7_), .ZN(n12517) );
  NAND2_X1 U15577 ( .A1(n14482), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12516) );
  AND2_X1 U15578 ( .A1(n12517), .A2(n12516), .ZN(n13183) );
  INV_X1 U15579 ( .A(n13183), .ZN(n14700) );
  NAND2_X1 U15580 ( .A1(n20432), .A2(n14700), .ZN(n12631) );
  NAND2_X1 U15581 ( .A1(n12518), .A2(n12631), .ZN(P1_U2959) );
  AOI22_X1 U15582 ( .A1(n20447), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20442), .ZN(n12521) );
  NAND2_X1 U15583 ( .A1(n14475), .A2(DATAI_6_), .ZN(n12520) );
  NAND2_X1 U15584 ( .A1(n14482), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12519) );
  AND2_X1 U15585 ( .A1(n12520), .A2(n12519), .ZN(n13100) );
  INV_X1 U15586 ( .A(n13100), .ZN(n21064) );
  NAND2_X1 U15587 ( .A1(n20432), .A2(n21064), .ZN(n12629) );
  NAND2_X1 U15588 ( .A1(n12521), .A2(n12629), .ZN(P1_U2958) );
  AOI22_X1 U15589 ( .A1(n20447), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20442), .ZN(n12524) );
  NAND2_X1 U15590 ( .A1(n14475), .A2(DATAI_2_), .ZN(n12523) );
  NAND2_X1 U15591 ( .A1(n14482), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12522) );
  AND2_X1 U15592 ( .A1(n12523), .A2(n12522), .ZN(n12758) );
  INV_X1 U15593 ( .A(n12758), .ZN(n14718) );
  NAND2_X1 U15594 ( .A1(n20432), .A2(n14718), .ZN(n12633) );
  NAND2_X1 U15595 ( .A1(n12524), .A2(n12633), .ZN(P1_U2954) );
  AOI22_X1 U15596 ( .A1(n20447), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20442), .ZN(n12527) );
  NAND2_X1 U15597 ( .A1(n14475), .A2(DATAI_3_), .ZN(n12526) );
  NAND2_X1 U15598 ( .A1(n14482), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12525) );
  AND2_X1 U15599 ( .A1(n12526), .A2(n12525), .ZN(n12757) );
  INV_X1 U15600 ( .A(n12757), .ZN(n16318) );
  NAND2_X1 U15601 ( .A1(n20432), .A2(n16318), .ZN(n12643) );
  NAND2_X1 U15602 ( .A1(n12527), .A2(n12643), .ZN(P1_U2955) );
  NAND3_X1 U15603 ( .A1(n12529), .A2(n12528), .A3(n20857), .ZN(n12530) );
  OAI21_X1 U15604 ( .B1(n12531), .B2(n13014), .A(n12530), .ZN(n12532) );
  NAND2_X1 U15605 ( .A1(n12050), .A2(n14477), .ZN(n12536) );
  NAND2_X1 U15606 ( .A1(n14475), .A2(DATAI_0_), .ZN(n12538) );
  NAND2_X1 U15607 ( .A1(n14482), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12537) );
  AND2_X1 U15608 ( .A1(n12538), .A2(n12537), .ZN(n12696) );
  OAI222_X1 U15609 ( .A1(n14717), .A2(n13090), .B1(n14745), .B2(n12234), .C1(
        n14744), .C2(n12696), .ZN(P1_U2904) );
  OR2_X1 U15610 ( .A1(n12577), .A2(n12059), .ZN(n12544) );
  XNOR2_X1 U15611 ( .A(n12618), .B(n12617), .ZN(n12541) );
  OAI211_X1 U15612 ( .C1(n12541), .C2(n20860), .A(n12540), .B(n12539), .ZN(
        n12542) );
  INV_X1 U15613 ( .A(n12542), .ZN(n12543) );
  NAND2_X1 U15614 ( .A1(n12544), .A2(n12543), .ZN(n12612) );
  NAND2_X1 U15615 ( .A1(n12546), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12615) );
  OAI21_X1 U15616 ( .B1(n12546), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12615), .ZN(n20505) );
  INV_X1 U15617 ( .A(n12547), .ZN(n12548) );
  NAND2_X1 U15618 ( .A1(n16482), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20501) );
  OAI21_X1 U15619 ( .B1(n16333), .B2(n13078), .A(n20501), .ZN(n12550) );
  NOR2_X1 U15620 ( .A1(n13080), .A2(n14888), .ZN(n12549) );
  AOI211_X1 U15621 ( .C1(n16365), .C2(n13078), .A(n12550), .B(n12549), .ZN(
        n12551) );
  OAI21_X1 U15622 ( .B1(n20299), .B2(n20505), .A(n12551), .ZN(P1_U2998) );
  INV_X1 U15623 ( .A(n12553), .ZN(n12554) );
  OAI211_X1 U15624 ( .C1(n12554), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15281), .B(n12840), .ZN(n12559) );
  INV_X1 U15625 ( .A(n12569), .ZN(n12555) );
  OAI21_X1 U15626 ( .B1(n12557), .B2(n12556), .A(n12555), .ZN(n13604) );
  INV_X1 U15627 ( .A(n13604), .ZN(n19370) );
  NAND2_X1 U15628 ( .A1(n19370), .A2(n15291), .ZN(n12558) );
  OAI211_X1 U15629 ( .C1(n15291), .C2(n12560), .A(n12559), .B(n12558), .ZN(
        P2_U2881) );
  OAI211_X1 U15630 ( .C1(n9778), .C2(n11455), .A(n15281), .B(n12562), .ZN(
        n12567) );
  AND2_X1 U15631 ( .A1(n12564), .A2(n12563), .ZN(n12565) );
  NOR2_X1 U15632 ( .A1(n12651), .A2(n12565), .ZN(n19347) );
  NAND2_X1 U15633 ( .A1(n19347), .A2(n15291), .ZN(n12566) );
  OAI211_X1 U15634 ( .C1(n15291), .C2(n19339), .A(n12567), .B(n12566), .ZN(
        P2_U2877) );
  XOR2_X1 U15635 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n12840), .Z(n12574)
         );
  OR2_X1 U15636 ( .A1(n12569), .A2(n12568), .ZN(n12571) );
  NAND2_X1 U15637 ( .A1(n12571), .A2(n12570), .ZN(n16649) );
  INV_X1 U15638 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12572) );
  MUX2_X1 U15639 ( .A(n16649), .B(n12572), .S(n15279), .Z(n12573) );
  OAI21_X1 U15640 ( .B1(n12574), .B2(n15298), .A(n12573), .ZN(P2_U2880) );
  NAND2_X1 U15641 ( .A1(n12577), .A2(n12578), .ZN(n12576) );
  NAND2_X1 U15642 ( .A1(n12576), .A2(n12575), .ZN(n12582) );
  INV_X1 U15643 ( .A(n12577), .ZN(n12580) );
  NAND2_X1 U15644 ( .A1(n12580), .A2(n12579), .ZN(n12581) );
  NAND2_X1 U15645 ( .A1(n12582), .A2(n12581), .ZN(n12599) );
  INV_X1 U15646 ( .A(n12599), .ZN(n12596) );
  AOI22_X1 U15647 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15648 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15649 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15650 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12585) );
  NAND4_X1 U15651 ( .A1(n12588), .A2(n12587), .A3(n12586), .A4(n12585), .ZN(
        n12594) );
  AOI22_X1 U15652 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15653 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15654 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15655 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U15656 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12593) );
  AOI22_X1 U15657 ( .A1(n13167), .A2(n12619), .B1(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n13044), .ZN(n12595) );
  NAND2_X1 U15658 ( .A1(n12599), .A2(n12598), .ZN(n12600) );
  INV_X1 U15659 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12602) );
  XNOR2_X1 U15660 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13033) );
  AOI21_X1 U15661 ( .B1(n14345), .B2(n13033), .A(n14444), .ZN(n12601) );
  OAI21_X1 U15662 ( .B1(n14285), .B2(n12602), .A(n12601), .ZN(n12603) );
  AOI21_X1 U15663 ( .B1(n12865), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12603), .ZN(n12604) );
  NAND2_X1 U15664 ( .A1(n14444), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12741) );
  NAND2_X1 U15665 ( .A1(n12605), .A2(n12741), .ZN(n12610) );
  INV_X1 U15666 ( .A(n12610), .ZN(n12607) );
  NAND2_X1 U15667 ( .A1(n12607), .A2(n12606), .ZN(n12742) );
  INV_X1 U15668 ( .A(n12742), .ZN(n12608) );
  AOI21_X1 U15669 ( .B1(n12610), .B2(n12609), .A(n12608), .ZN(n13015) );
  INV_X1 U15670 ( .A(n13015), .ZN(n12759) );
  AND2_X1 U15671 ( .A1(n16482), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20480) );
  NOR2_X1 U15672 ( .A1(n20461), .A2(n13033), .ZN(n12611) );
  AOI211_X1 U15673 ( .C1(n20450), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20480), .B(n12611), .ZN(n12628) );
  INV_X1 U15674 ( .A(n12545), .ZN(n12613) );
  NAND2_X1 U15675 ( .A1(n12613), .A2(n12612), .ZN(n12614) );
  NAND2_X1 U15676 ( .A1(n12615), .A2(n12614), .ZN(n12984) );
  INV_X1 U15677 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20870) );
  OR2_X1 U15678 ( .A1(n12616), .A2(n13651), .ZN(n12624) );
  NAND2_X1 U15679 ( .A1(n12618), .A2(n12617), .ZN(n12989) );
  INV_X1 U15680 ( .A(n12619), .ZN(n12988) );
  XNOR2_X1 U15681 ( .A(n12989), .B(n12988), .ZN(n12622) );
  INV_X1 U15682 ( .A(n12620), .ZN(n12621) );
  AOI21_X1 U15683 ( .B1(n12622), .B2(n13657), .A(n12621), .ZN(n12623) );
  OR2_X1 U15684 ( .A1(n12626), .A2(n12625), .ZN(n20489) );
  NAND3_X1 U15685 ( .A1(n20489), .A2(n12986), .A3(n20457), .ZN(n12627) );
  OAI211_X1 U15686 ( .C1(n12759), .C2(n14888), .A(n12628), .B(n12627), .ZN(
        P1_U2997) );
  AOI22_X1 U15687 ( .A1(n20447), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20442), .ZN(n12630) );
  NAND2_X1 U15688 ( .A1(n12630), .A2(n12629), .ZN(P1_U2943) );
  AOI22_X1 U15689 ( .A1(n20447), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20442), .ZN(n12632) );
  NAND2_X1 U15690 ( .A1(n12632), .A2(n12631), .ZN(P1_U2944) );
  AOI22_X1 U15691 ( .A1(n20447), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20442), .ZN(n12634) );
  NAND2_X1 U15692 ( .A1(n12634), .A2(n12633), .ZN(P1_U2939) );
  AOI22_X1 U15693 ( .A1(n20447), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20442), .ZN(n12635) );
  INV_X1 U15694 ( .A(n12696), .ZN(n14730) );
  NAND2_X1 U15695 ( .A1(n20432), .A2(n14730), .ZN(n12645) );
  NAND2_X1 U15696 ( .A1(n12635), .A2(n12645), .ZN(P1_U2952) );
  AOI22_X1 U15697 ( .A1(n20447), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20442), .ZN(n12638) );
  NAND2_X1 U15698 ( .A1(n14475), .A2(DATAI_1_), .ZN(n12637) );
  NAND2_X1 U15699 ( .A1(n14482), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12636) );
  AND2_X1 U15700 ( .A1(n12637), .A2(n12636), .ZN(n12760) );
  INV_X1 U15701 ( .A(n12760), .ZN(n14724) );
  NAND2_X1 U15702 ( .A1(n20432), .A2(n14724), .ZN(n12641) );
  NAND2_X1 U15703 ( .A1(n12638), .A2(n12641), .ZN(P1_U2953) );
  AOI22_X1 U15704 ( .A1(n20447), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20442), .ZN(n12640) );
  NAND2_X1 U15705 ( .A1(n12640), .A2(n12639), .ZN(P1_U2941) );
  AOI22_X1 U15706 ( .A1(n20447), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20442), .ZN(n12642) );
  NAND2_X1 U15707 ( .A1(n12642), .A2(n12641), .ZN(P1_U2938) );
  AOI22_X1 U15708 ( .A1(n20447), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20442), .ZN(n12644) );
  NAND2_X1 U15709 ( .A1(n12644), .A2(n12643), .ZN(P1_U2940) );
  AOI22_X1 U15710 ( .A1(n20447), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20442), .ZN(n12646) );
  NAND2_X1 U15711 ( .A1(n12646), .A2(n12645), .ZN(P1_U2937) );
  AOI22_X1 U15712 ( .A1(n20447), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20442), .ZN(n12648) );
  NAND2_X1 U15713 ( .A1(n12648), .A2(n12647), .ZN(P1_U2942) );
  XNOR2_X1 U15714 ( .A(n12562), .B(n12649), .ZN(n12655) );
  OR2_X1 U15715 ( .A1(n12651), .A2(n12650), .ZN(n12652) );
  AND2_X1 U15716 ( .A1(n12827), .A2(n12652), .ZN(n16672) );
  NOR2_X1 U15717 ( .A1(n15291), .A2(n15201), .ZN(n12653) );
  AOI21_X1 U15718 ( .B1(n16672), .B2(n15291), .A(n12653), .ZN(n12654) );
  OAI21_X1 U15719 ( .B1(n12655), .B2(n15298), .A(n12654), .ZN(P2_U2876) );
  AOI22_X1 U15720 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15721 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15722 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U15723 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12658) );
  NAND4_X1 U15724 ( .A1(n12661), .A2(n12660), .A3(n12659), .A4(n12658), .ZN(
        n12667) );
  AOI22_X1 U15725 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15726 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15727 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15728 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12662) );
  NAND4_X1 U15729 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12666) );
  AOI22_X1 U15730 ( .A1(n13167), .A2(n13623), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13044), .ZN(n12668) );
  NAND2_X2 U15731 ( .A1(n12669), .A2(n12668), .ZN(n12761) );
  INV_X1 U15732 ( .A(n12761), .ZN(n12708) );
  NAND2_X1 U15733 ( .A1(n12670), .A2(n12708), .ZN(n12671) );
  INV_X1 U15734 ( .A(n9680), .ZN(n12672) );
  INV_X1 U15735 ( .A(n13539), .ZN(n12673) );
  INV_X1 U15736 ( .A(n12939), .ZN(n12674) );
  AOI22_X1 U15737 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9656), .B1(DATAI_27_), 
        .B2(n9650), .ZN(n20672) );
  INV_X1 U15738 ( .A(n20672), .ZN(n20726) );
  NOR2_X1 U15739 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20861) );
  NOR2_X1 U15740 ( .A1(n12911), .A2(n12675), .ZN(n20725) );
  INV_X1 U15741 ( .A(n20725), .ZN(n13200) );
  NAND2_X1 U15742 ( .A1(n16151), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20651) );
  INV_X1 U15743 ( .A(n20651), .ZN(n12676) );
  NAND2_X1 U15744 ( .A1(n12712), .A2(n12676), .ZN(n12913) );
  NAND2_X1 U15745 ( .A1(n12677), .A2(n12940), .ZN(n20650) );
  NAND2_X1 U15746 ( .A1(n12679), .A2(n13088), .ZN(n12941) );
  OAI21_X1 U15747 ( .B1(n20650), .B2(n12941), .A(n12913), .ZN(n12682) );
  NOR2_X1 U15748 ( .A1(n20554), .A2(n20651), .ZN(n13104) );
  AOI22_X1 U15749 ( .A1(n12682), .A2(n20658), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13104), .ZN(n12912) );
  INV_X1 U15750 ( .A(n20724), .ZN(n13694) );
  OAI22_X1 U15751 ( .A1(n13200), .A2(n12913), .B1(n12912), .B2(n13694), .ZN(
        n12681) );
  AOI21_X1 U15752 ( .B1(n13103), .B2(n20726), .A(n12681), .ZN(n12686) );
  NAND2_X1 U15753 ( .A1(n15009), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15008) );
  INV_X1 U15754 ( .A(n12682), .ZN(n12683) );
  OAI211_X1 U15755 ( .C1(n20655), .C2(n15008), .A(n20622), .B(n12683), .ZN(
        n12684) );
  OAI211_X1 U15756 ( .C1(n20622), .C2(n13104), .A(n12684), .B(n20705), .ZN(
        n12915) );
  NAND2_X1 U15757 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12685) );
  OAI211_X1 U15758 ( .C1(n20729), .C2(n13543), .A(n12686), .B(n12685), .ZN(
        P1_U3124) );
  AOI22_X1 U15759 ( .A1(DATAI_31_), .A2(n9650), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9656), .ZN(n20691) );
  INV_X1 U15760 ( .A(n20691), .ZN(n20752) );
  INV_X1 U15761 ( .A(n20751), .ZN(n13216) );
  INV_X1 U15762 ( .A(n20749), .ZN(n13702) );
  OAI22_X1 U15763 ( .A1(n13216), .A2(n12913), .B1(n12912), .B2(n13702), .ZN(
        n12687) );
  AOI21_X1 U15764 ( .B1(n13103), .B2(n20752), .A(n12687), .ZN(n12689) );
  NAND2_X1 U15765 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12688) );
  OAI211_X1 U15766 ( .C1(n20758), .C2(n13543), .A(n12689), .B(n12688), .ZN(
        P1_U3128) );
  AOI22_X1 U15767 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9656), .B1(DATAI_26_), 
        .B2(n9650), .ZN(n20668) );
  INV_X1 U15768 ( .A(n20668), .ZN(n20720) );
  INV_X1 U15769 ( .A(n20719), .ZN(n13212) );
  INV_X1 U15770 ( .A(n20718), .ZN(n13706) );
  OAI22_X1 U15771 ( .A1(n13212), .A2(n12913), .B1(n12912), .B2(n13706), .ZN(
        n12690) );
  AOI21_X1 U15772 ( .B1(n13103), .B2(n20720), .A(n12690), .ZN(n12692) );
  NAND2_X1 U15773 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12691) );
  OAI211_X1 U15774 ( .C1(n20723), .C2(n13543), .A(n12692), .B(n12691), .ZN(
        P1_U3123) );
  AOI22_X1 U15775 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9656), .B1(DATAI_29_), 
        .B2(n9650), .ZN(n20640) );
  INV_X1 U15776 ( .A(n20737), .ZN(n13208) );
  INV_X1 U15777 ( .A(n20736), .ZN(n13710) );
  OAI22_X1 U15778 ( .A1(n13208), .A2(n12913), .B1(n12912), .B2(n13710), .ZN(
        n12693) );
  AOI21_X1 U15779 ( .B1(n13103), .B2(n20738), .A(n12693), .ZN(n12695) );
  NAND2_X1 U15780 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12694) );
  OAI211_X1 U15781 ( .C1(n20741), .C2(n13543), .A(n12695), .B(n12694), .ZN(
        P1_U3126) );
  AOI22_X1 U15782 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9656), .B1(DATAI_24_), 
        .B2(n9650), .ZN(n20626) );
  NOR2_X2 U15783 ( .A1(n12911), .A2(n13024), .ZN(n20701) );
  INV_X1 U15784 ( .A(n20701), .ZN(n13220) );
  OAI22_X1 U15785 ( .A1(n13220), .A2(n12913), .B1(n12912), .B2(n13686), .ZN(
        n12697) );
  AOI21_X1 U15786 ( .B1(n13103), .B2(n20708), .A(n12697), .ZN(n12699) );
  NAND2_X1 U15787 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12698) );
  OAI211_X1 U15788 ( .C1(n20711), .C2(n13543), .A(n12699), .B(n12698), .ZN(
        P1_U3121) );
  AOI22_X1 U15789 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9656), .B1(DATAI_25_), 
        .B2(n9650), .ZN(n20664) );
  INV_X1 U15790 ( .A(n20713), .ZN(n13192) );
  INV_X1 U15791 ( .A(n20712), .ZN(n13690) );
  OAI22_X1 U15792 ( .A1(n13192), .A2(n12913), .B1(n12912), .B2(n13690), .ZN(
        n12700) );
  AOI21_X1 U15793 ( .B1(n13103), .B2(n20714), .A(n12700), .ZN(n12702) );
  NAND2_X1 U15794 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12701) );
  OAI211_X1 U15795 ( .C1(n20717), .C2(n13543), .A(n12702), .B(n12701), .ZN(
        P1_U3122) );
  MUX2_X1 U15796 ( .A(n14417), .B(n14454), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12704) );
  NAND2_X1 U15797 ( .A1(n14405), .A2(n20870), .ZN(n12703) );
  AND2_X1 U15798 ( .A1(n12704), .A2(n12703), .ZN(n12705) );
  NAND2_X1 U15799 ( .A1(n12706), .A2(n12705), .ZN(n20369) );
  OAI21_X1 U15800 ( .B1(n12706), .B2(n12705), .A(n20369), .ZN(n20479) );
  INV_X1 U15801 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12707) );
  OAI222_X1 U15802 ( .A1(n20479), .A2(n20385), .B1(n12707), .B2(n20390), .C1(
        n12759), .C2(n14666), .ZN(P1_U2870) );
  INV_X1 U15803 ( .A(n12949), .ZN(n12709) );
  NAND2_X1 U15804 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20692) );
  OR2_X1 U15805 ( .A1(n20554), .A2(n20692), .ZN(n12716) );
  INV_X1 U15806 ( .A(n20658), .ZN(n20703) );
  NOR2_X1 U15807 ( .A1(n9680), .A2(n15008), .ZN(n15014) );
  AOI21_X1 U15808 ( .B1(n15014), .B2(n12761), .A(n20703), .ZN(n15013) );
  AOI21_X1 U15809 ( .B1(n12716), .B2(n20703), .A(n15013), .ZN(n12714) );
  OR2_X1 U15810 ( .A1(n12940), .A2(n12710), .ZN(n20694) );
  INV_X1 U15811 ( .A(n20692), .ZN(n12711) );
  NAND2_X1 U15812 ( .A1(n12712), .A2(n12711), .ZN(n12923) );
  OAI21_X1 U15813 ( .B1(n20694), .B2(n12941), .A(n12923), .ZN(n12713) );
  AND2_X1 U15814 ( .A1(n12713), .A2(n20658), .ZN(n12715) );
  NAND2_X1 U15815 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12722) );
  INV_X1 U15816 ( .A(n12715), .ZN(n12719) );
  INV_X1 U15817 ( .A(n12716), .ZN(n12717) );
  NAND2_X1 U15818 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n12717), .ZN(n12718) );
  AND2_X1 U15819 ( .A1(n12719), .A2(n12718), .ZN(n12922) );
  OAI22_X1 U15820 ( .A1(n13216), .A2(n12923), .B1(n12922), .B2(n13702), .ZN(
        n12720) );
  AOI21_X1 U15821 ( .B1(n13492), .B2(n20752), .A(n12720), .ZN(n12721) );
  OAI211_X1 U15822 ( .C1(n20758), .C2(n12927), .A(n12722), .B(n12721), .ZN(
        P1_U3160) );
  NAND2_X1 U15823 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12725) );
  OAI22_X1 U15824 ( .A1(n13192), .A2(n12923), .B1(n12922), .B2(n13690), .ZN(
        n12723) );
  AOI21_X1 U15825 ( .B1(n13492), .B2(n20714), .A(n12723), .ZN(n12724) );
  OAI211_X1 U15826 ( .C1(n20717), .C2(n12927), .A(n12725), .B(n12724), .ZN(
        P1_U3154) );
  NAND2_X1 U15827 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12728) );
  OAI22_X1 U15828 ( .A1(n13208), .A2(n12923), .B1(n12922), .B2(n13710), .ZN(
        n12726) );
  AOI21_X1 U15829 ( .B1(n13492), .B2(n20738), .A(n12726), .ZN(n12727) );
  OAI211_X1 U15830 ( .C1(n20741), .C2(n12927), .A(n12728), .B(n12727), .ZN(
        P1_U3158) );
  NAND2_X1 U15831 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12731) );
  OAI22_X1 U15832 ( .A1(n13212), .A2(n12923), .B1(n12922), .B2(n13706), .ZN(
        n12729) );
  AOI21_X1 U15833 ( .B1(n13492), .B2(n20720), .A(n12729), .ZN(n12730) );
  OAI211_X1 U15834 ( .C1(n20723), .C2(n12927), .A(n12731), .B(n12730), .ZN(
        P1_U3155) );
  NAND2_X1 U15835 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12734) );
  OAI22_X1 U15836 ( .A1(n13200), .A2(n12923), .B1(n12922), .B2(n13694), .ZN(
        n12732) );
  AOI21_X1 U15837 ( .B1(n13492), .B2(n20726), .A(n12732), .ZN(n12733) );
  OAI211_X1 U15838 ( .C1(n20729), .C2(n12927), .A(n12734), .B(n12733), .ZN(
        P1_U3156) );
  INV_X1 U15839 ( .A(n12923), .ZN(n12736) );
  INV_X1 U15840 ( .A(n12922), .ZN(n12735) );
  AOI22_X1 U15841 ( .A1(n20701), .A2(n12736), .B1(n20700), .B2(n12735), .ZN(
        n12738) );
  INV_X1 U15842 ( .A(n20711), .ZN(n20623) );
  NAND2_X1 U15843 ( .A1(n20548), .A2(n20623), .ZN(n12737) );
  OAI211_X1 U15844 ( .C1(n20626), .C2(n13534), .A(n12738), .B(n12737), .ZN(
        n12739) );
  AOI21_X1 U15845 ( .B1(n12921), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12739), .ZN(n12740) );
  INV_X1 U15846 ( .A(n12740), .ZN(P1_U3153) );
  INV_X1 U15847 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12748) );
  INV_X1 U15848 ( .A(n12744), .ZN(n12746) );
  INV_X1 U15849 ( .A(n12864), .ZN(n12745) );
  OAI21_X1 U15850 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12746), .A(
        n12745), .ZN(n13068) );
  AOI22_X1 U15851 ( .A1(n14345), .A2(n13068), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12747) );
  OAI21_X1 U15852 ( .B1(n14285), .B2(n12748), .A(n12747), .ZN(n12749) );
  AOI21_X1 U15853 ( .B1(n12865), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12749), .ZN(n12750) );
  OAI21_X1 U15854 ( .B1(n15012), .B2(n13476), .A(n12750), .ZN(n12751) );
  OAI21_X1 U15855 ( .B1(n12752), .B2(n12751), .A(n12970), .ZN(n13072) );
  INV_X1 U15856 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12756) );
  INV_X1 U15857 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U15858 ( .A1(n12753), .A2(n12987), .ZN(n12754) );
  OAI211_X1 U15859 ( .C1(P1_EBX_REG_3__SCAN_IN), .C2(n14456), .A(n12754), .B(
        n14454), .ZN(n12755) );
  OAI21_X1 U15860 ( .B1(n14410), .B2(P1_EBX_REG_3__SCAN_IN), .A(n12755), .ZN(
        n12900) );
  INV_X1 U15861 ( .A(n12900), .ZN(n20368) );
  XNOR2_X1 U15862 ( .A(n20369), .B(n20368), .ZN(n20471) );
  OAI222_X1 U15863 ( .A1(n14666), .A2(n13072), .B1(n12756), .B2(n20390), .C1(
        n20385), .C2(n20471), .ZN(P1_U2869) );
  OAI222_X1 U15864 ( .A1(n14717), .A2(n13072), .B1(n14745), .B2(n12748), .C1(
        n14744), .C2(n12757), .ZN(P1_U2901) );
  OAI222_X1 U15865 ( .A1(n14717), .A2(n12759), .B1(n14745), .B2(n12602), .C1(
        n14744), .C2(n12758), .ZN(P1_U2902) );
  OAI222_X1 U15866 ( .A1(n14717), .A2(n13080), .B1(n14745), .B2(n12503), .C1(
        n14744), .C2(n12760), .ZN(P1_U2903) );
  NOR2_X1 U15867 ( .A1(n12940), .A2(n12762), .ZN(n20616) );
  INV_X1 U15868 ( .A(n20616), .ZN(n12763) );
  OAI21_X1 U15869 ( .B1(n12763), .B2(n12941), .A(n12932), .ZN(n12765) );
  NOR2_X1 U15870 ( .A1(n20554), .A2(n20615), .ZN(n13676) );
  AOI22_X1 U15871 ( .A1(n12765), .A2(n20622), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13676), .ZN(n12931) );
  OAI22_X1 U15872 ( .A1(n12932), .A2(n13216), .B1(n12931), .B2(n13702), .ZN(
        n12764) );
  AOI21_X1 U15873 ( .B1(n12934), .B2(n20752), .A(n12764), .ZN(n12769) );
  INV_X1 U15874 ( .A(n20584), .ZN(n20619) );
  INV_X1 U15875 ( .A(n12765), .ZN(n12766) );
  OAI211_X1 U15876 ( .C1(n20619), .C2(n15008), .A(n20622), .B(n12766), .ZN(
        n12767) );
  OAI211_X1 U15877 ( .C1(n20622), .C2(n13676), .A(n12767), .B(n20705), .ZN(
        n12935) );
  NAND2_X1 U15878 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12768) );
  OAI211_X1 U15879 ( .C1(n20758), .C2(n12938), .A(n12769), .B(n12768), .ZN(
        P1_U3096) );
  OAI22_X1 U15880 ( .A1(n12932), .A2(n13200), .B1(n12931), .B2(n13694), .ZN(
        n12770) );
  AOI21_X1 U15881 ( .B1(n12934), .B2(n20726), .A(n12770), .ZN(n12772) );
  NAND2_X1 U15882 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12771) );
  OAI211_X1 U15883 ( .C1(n20729), .C2(n12938), .A(n12772), .B(n12771), .ZN(
        P1_U3092) );
  OAI22_X1 U15884 ( .A1(n12932), .A2(n13212), .B1(n12931), .B2(n13706), .ZN(
        n12773) );
  AOI21_X1 U15885 ( .B1(n12934), .B2(n20720), .A(n12773), .ZN(n12775) );
  NAND2_X1 U15886 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12774) );
  OAI211_X1 U15887 ( .C1(n20723), .C2(n12938), .A(n12775), .B(n12774), .ZN(
        P1_U3091) );
  OAI22_X1 U15888 ( .A1(n12932), .A2(n13220), .B1(n12931), .B2(n13686), .ZN(
        n12776) );
  AOI21_X1 U15889 ( .B1(n12934), .B2(n20708), .A(n12776), .ZN(n12778) );
  NAND2_X1 U15890 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12777) );
  OAI211_X1 U15891 ( .C1(n20711), .C2(n12938), .A(n12778), .B(n12777), .ZN(
        P1_U3089) );
  OAI22_X1 U15892 ( .A1(n12932), .A2(n13208), .B1(n12931), .B2(n13710), .ZN(
        n12779) );
  AOI21_X1 U15893 ( .B1(n12934), .B2(n20738), .A(n12779), .ZN(n12781) );
  NAND2_X1 U15894 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12780) );
  OAI211_X1 U15895 ( .C1(n20741), .C2(n12938), .A(n12781), .B(n12780), .ZN(
        P1_U3094) );
  OAI22_X1 U15896 ( .A1(n12932), .A2(n13192), .B1(n12931), .B2(n13690), .ZN(
        n12782) );
  AOI21_X1 U15897 ( .B1(n12934), .B2(n20714), .A(n12782), .ZN(n12784) );
  NAND2_X1 U15898 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12783) );
  OAI211_X1 U15899 ( .C1(n20717), .C2(n12938), .A(n12784), .B(n12783), .ZN(
        P1_U3090) );
  NOR2_X1 U15900 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16510), .ZN(n12815) );
  NAND2_X1 U15901 ( .A1(n12786), .A2(n12785), .ZN(n12795) );
  XNOR2_X1 U15902 ( .A(n12800), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15020) );
  XNOR2_X1 U15903 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12790) );
  AND2_X1 U15904 ( .A1(n12788), .A2(n12787), .ZN(n12789) );
  NAND2_X1 U15905 ( .A1(n14091), .A2(n12789), .ZN(n12802) );
  OAI22_X1 U15906 ( .A1(n12804), .A2(n12790), .B1(n12802), .B2(n15020), .ZN(
        n12793) );
  NOR2_X1 U15907 ( .A1(n12940), .A2(n12791), .ZN(n12792) );
  AOI211_X1 U15908 ( .C1(n12795), .C2(n15020), .A(n12793), .B(n12792), .ZN(
        n15026) );
  INV_X1 U15909 ( .A(n15026), .ZN(n12794) );
  MUX2_X1 U15910 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n12794), .S(
        n16145), .Z(n16152) );
  AOI22_X1 U15911 ( .A1(n12815), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16152), .B2(n16510), .ZN(n12812) );
  MUX2_X1 U15912 ( .A(n11880), .B(n9991), .S(n12800), .Z(n12796) );
  OAI21_X1 U15913 ( .B1(n12797), .B2(n12796), .A(n12795), .ZN(n12807) );
  XNOR2_X1 U15914 ( .A(n12798), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12803) );
  INV_X1 U15915 ( .A(n11880), .ZN(n12799) );
  OAI21_X1 U15916 ( .B1(n12800), .B2(n9991), .A(n12799), .ZN(n12801) );
  NOR2_X1 U15917 ( .A1(n12801), .A2(n14293), .ZN(n15029) );
  OAI22_X1 U15918 ( .A1(n12804), .A2(n12803), .B1(n15029), .B2(n12802), .ZN(
        n12805) );
  INV_X1 U15919 ( .A(n12805), .ZN(n12806) );
  NAND2_X1 U15920 ( .A1(n12807), .A2(n12806), .ZN(n12808) );
  AOI21_X1 U15921 ( .B1(n12677), .B2(n12809), .A(n12808), .ZN(n15031) );
  MUX2_X1 U15922 ( .A(n9991), .B(n15031), .S(n16145), .Z(n16154) );
  INV_X1 U15923 ( .A(n16154), .ZN(n12810) );
  AOI22_X1 U15924 ( .A1(n12815), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16510), .B2(n12810), .ZN(n12811) );
  NOR2_X1 U15925 ( .A1(n12812), .A2(n12811), .ZN(n16163) );
  NAND2_X1 U15926 ( .A1(n16163), .A2(n12813), .ZN(n12820) );
  OAI21_X1 U15927 ( .B1(n20365), .B2(n12172), .A(n16145), .ZN(n12817) );
  AOI21_X1 U15928 ( .B1(n12814), .B2(n12868), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n12816) );
  AOI22_X1 U15929 ( .A1(n12817), .A2(n12816), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n12815), .ZN(n16161) );
  AND3_X1 U15930 ( .A1(n12820), .A2(n16161), .A3(n20300), .ZN(n12818) );
  AND3_X1 U15931 ( .A1(n12820), .A2(n16161), .A3(n12819), .ZN(n16174) );
  INV_X1 U15932 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n16512) );
  AND2_X1 U15933 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n16512), .ZN(n15017) );
  OAI22_X1 U15934 ( .A1(n13539), .A2(n20703), .B1(n12233), .B2(n15017), .ZN(
        n12821) );
  OAI21_X1 U15935 ( .B1(n16174), .B2(n12821), .A(n20515), .ZN(n12822) );
  OAI21_X1 U15936 ( .B1(n20515), .B2(n20693), .A(n12822), .ZN(P1_U3478) );
  AOI211_X1 U15937 ( .C1(n9680), .C2(n15008), .A(n20703), .B(n15014), .ZN(
        n12824) );
  NOR2_X1 U15938 ( .A1(n12940), .A2(n15017), .ZN(n12823) );
  OAI21_X1 U15939 ( .B1(n12824), .B2(n12823), .A(n20515), .ZN(n12825) );
  OAI21_X1 U15940 ( .B1(n20515), .B2(n16151), .A(n12825), .ZN(P1_U3476) );
  NAND2_X1 U15941 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  NAND2_X1 U15942 ( .A1(n13094), .A2(n12828), .ZN(n15807) );
  INV_X1 U15943 ( .A(n12829), .ZN(n12830) );
  OAI211_X1 U15944 ( .C1(n12832), .C2(n12831), .A(n12830), .B(n15281), .ZN(
        n12834) );
  NAND2_X1 U15945 ( .A1(n15279), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12833) );
  OAI211_X1 U15946 ( .C1(n15807), .C2(n15279), .A(n12834), .B(n12833), .ZN(
        P2_U2875) );
  OR2_X1 U15947 ( .A1(n12836), .A2(n12835), .ZN(n12838) );
  AND2_X1 U15948 ( .A1(n12838), .A2(n12837), .ZN(n19359) );
  NOR2_X1 U15949 ( .A1(n15291), .A2(n19353), .ZN(n12845) );
  OR2_X1 U15950 ( .A1(n12840), .A2(n12839), .ZN(n12842) );
  AOI211_X1 U15951 ( .C1(n12843), .C2(n12842), .A(n15298), .B(n12841), .ZN(
        n12844) );
  AOI211_X1 U15952 ( .C1(n19359), .C2(n15291), .A(n12845), .B(n12844), .ZN(
        n12846) );
  INV_X1 U15953 ( .A(n12846), .ZN(P2_U2879) );
  AOI22_X1 U15954 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9681), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U15955 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12199), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U15956 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U15957 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12847) );
  NAND4_X1 U15958 ( .A1(n12850), .A2(n12849), .A3(n12848), .A4(n12847), .ZN(
        n12856) );
  AOI22_X1 U15959 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U15960 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U15961 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15962 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12851) );
  NAND4_X1 U15963 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12855) );
  NAND2_X1 U15964 ( .A1(n13167), .A2(n13622), .ZN(n12858) );
  NAND2_X1 U15965 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12857) );
  NAND2_X1 U15966 ( .A1(n12858), .A2(n12857), .ZN(n12860) );
  INV_X1 U15967 ( .A(n12860), .ZN(n12861) );
  NAND2_X1 U15968 ( .A1(n12884), .A2(n12862), .ZN(n13613) );
  INV_X1 U15969 ( .A(n13613), .ZN(n12863) );
  NAND2_X1 U15970 ( .A1(n12863), .A2(n13859), .ZN(n12872) );
  OAI21_X1 U15971 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12864), .A(
        n12887), .ZN(n20460) );
  INV_X1 U15972 ( .A(n12865), .ZN(n12869) );
  OAI21_X1 U15973 ( .B1(n20702), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20697), .ZN(n12867) );
  NAND2_X1 U15974 ( .A1(n14445), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12866) );
  OAI211_X1 U15975 ( .C1(n12869), .C2(n12868), .A(n12867), .B(n12866), .ZN(
        n12870) );
  OAI21_X1 U15976 ( .B1(n14351), .B2(n20460), .A(n12870), .ZN(n12871) );
  AOI22_X1 U15977 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U15978 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U15979 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U15980 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12873) );
  NAND4_X1 U15981 ( .A1(n12876), .A2(n12875), .A3(n12874), .A4(n12873), .ZN(
        n12882) );
  AOI22_X1 U15982 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U15983 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U15984 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U15985 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12877) );
  NAND4_X1 U15986 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n12881) );
  AOI22_X1 U15987 ( .A1(n13167), .A2(n13640), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n13044), .ZN(n12883) );
  NAND2_X1 U15988 ( .A1(n12884), .A2(n12883), .ZN(n12885) );
  NAND2_X1 U15989 ( .A1(n13164), .A2(n12885), .ZN(n13621) );
  INV_X1 U15990 ( .A(n13621), .ZN(n12886) );
  INV_X1 U15991 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12890) );
  OAI21_X1 U15992 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12888), .A(
        n13000), .ZN(n20358) );
  AOI22_X1 U15993 ( .A1(n14345), .A2(n20358), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12889) );
  OAI21_X1 U15994 ( .B1(n14285), .B2(n12890), .A(n12889), .ZN(n12891) );
  INV_X1 U15995 ( .A(n12891), .ZN(n12892) );
  NOR2_X1 U15996 ( .A1(n12895), .A2(n12894), .ZN(n12896) );
  NOR2_X1 U15997 ( .A1(n12896), .A2(n9750), .ZN(n20360) );
  INV_X1 U15998 ( .A(n20360), .ZN(n12975) );
  INV_X1 U15999 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20389) );
  NAND2_X1 U16000 ( .A1(n14399), .A2(n20389), .ZN(n12899) );
  INV_X1 U16001 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13618) );
  NAND2_X1 U16002 ( .A1(n9988), .A2(n20389), .ZN(n12897) );
  OAI211_X1 U16003 ( .C1(n14419), .C2(n13618), .A(n12897), .B(n12753), .ZN(
        n12898) );
  AND2_X1 U16004 ( .A1(n12899), .A2(n12898), .ZN(n20366) );
  NAND2_X1 U16005 ( .A1(n20366), .A2(n12900), .ZN(n12901) );
  INV_X1 U16006 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13725) );
  OAI21_X1 U16007 ( .B1(n14419), .B2(n13725), .A(n12753), .ZN(n12902) );
  OAI21_X1 U16008 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n14456), .A(n12902), .ZN(
        n12903) );
  OAI21_X1 U16009 ( .B1(n14410), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12903), .ZN(
        n13057) );
  XNOR2_X1 U16010 ( .A(n20370), .B(n13057), .ZN(n20355) );
  INV_X1 U16011 ( .A(n20390), .ZN(n14649) );
  AOI22_X1 U16012 ( .A1(n16315), .A2(n20355), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14649), .ZN(n12904) );
  OAI21_X1 U16013 ( .B1(n12975), .B2(n14666), .A(n12904), .ZN(P1_U2867) );
  AOI22_X1 U16014 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9656), .B1(DATAI_30_), 
        .B2(n9650), .ZN(n20682) );
  INV_X1 U16015 ( .A(n20682), .ZN(n20744) );
  INV_X1 U16016 ( .A(n20743), .ZN(n13204) );
  INV_X1 U16017 ( .A(n20742), .ZN(n13698) );
  OAI22_X1 U16018 ( .A1(n13204), .A2(n12913), .B1(n12912), .B2(n13698), .ZN(
        n12906) );
  AOI21_X1 U16019 ( .B1(n13103), .B2(n20744), .A(n12906), .ZN(n12908) );
  NAND2_X1 U16020 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12907) );
  OAI211_X1 U16021 ( .C1(n20747), .C2(n13543), .A(n12908), .B(n12907), .ZN(
        P1_U3127) );
  AOI22_X1 U16022 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9656), .B1(DATAI_28_), 
        .B2(n9650), .ZN(n20636) );
  INV_X1 U16023 ( .A(n20636), .ZN(n20732) );
  INV_X1 U16024 ( .A(n20731), .ZN(n13224) );
  INV_X1 U16025 ( .A(n20730), .ZN(n13717) );
  OAI22_X1 U16026 ( .A1(n13224), .A2(n12913), .B1(n12912), .B2(n13717), .ZN(
        n12914) );
  AOI21_X1 U16027 ( .B1(n13103), .B2(n20732), .A(n12914), .ZN(n12917) );
  NAND2_X1 U16028 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12916) );
  OAI211_X1 U16029 ( .C1(n20735), .C2(n13543), .A(n12917), .B(n12916), .ZN(
        P1_U3125) );
  NAND2_X1 U16030 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12920) );
  OAI22_X1 U16031 ( .A1(n13204), .A2(n12923), .B1(n12922), .B2(n13698), .ZN(
        n12918) );
  AOI21_X1 U16032 ( .B1(n13492), .B2(n20744), .A(n12918), .ZN(n12919) );
  OAI211_X1 U16033 ( .C1(n20747), .C2(n12927), .A(n12920), .B(n12919), .ZN(
        P1_U3159) );
  NAND2_X1 U16034 ( .A1(n12921), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12926) );
  OAI22_X1 U16035 ( .A1(n13224), .A2(n12923), .B1(n12922), .B2(n13717), .ZN(
        n12924) );
  AOI21_X1 U16036 ( .B1(n13492), .B2(n20732), .A(n12924), .ZN(n12925) );
  OAI211_X1 U16037 ( .C1(n20735), .C2(n12927), .A(n12926), .B(n12925), .ZN(
        P1_U3157) );
  OAI22_X1 U16038 ( .A1(n12932), .A2(n13204), .B1(n12931), .B2(n13698), .ZN(
        n12928) );
  AOI21_X1 U16039 ( .B1(n12934), .B2(n20744), .A(n12928), .ZN(n12930) );
  NAND2_X1 U16040 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12929) );
  OAI211_X1 U16041 ( .C1(n20747), .C2(n12938), .A(n12930), .B(n12929), .ZN(
        P1_U3095) );
  OAI22_X1 U16042 ( .A1(n12932), .A2(n13224), .B1(n12931), .B2(n13717), .ZN(
        n12933) );
  AOI21_X1 U16043 ( .B1(n12934), .B2(n20732), .A(n12933), .ZN(n12937) );
  NAND2_X1 U16044 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12936) );
  OAI211_X1 U16045 ( .C1(n20735), .C2(n12938), .A(n12937), .B(n12936), .ZN(
        P1_U3093) );
  INV_X1 U16046 ( .A(n12940), .ZN(n13030) );
  OR2_X1 U16047 ( .A1(n12677), .A2(n13030), .ZN(n20522) );
  INV_X1 U16048 ( .A(n20522), .ZN(n20556) );
  INV_X1 U16049 ( .A(n12941), .ZN(n12944) );
  NOR2_X1 U16050 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20555) );
  INV_X1 U16051 ( .A(n20555), .ZN(n12943) );
  NOR2_X1 U16052 ( .A1(n12943), .A2(n12942), .ZN(n12966) );
  AOI21_X1 U16053 ( .B1(n20556), .B2(n12944), .A(n12966), .ZN(n12948) );
  INV_X1 U16054 ( .A(n12948), .ZN(n12946) );
  INV_X1 U16055 ( .A(n20517), .ZN(n20559) );
  OAI21_X1 U16056 ( .B1(n20559), .B2(n15008), .A(n20658), .ZN(n12947) );
  NAND2_X1 U16057 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20555), .ZN(
        n13191) );
  NAND2_X1 U16058 ( .A1(n20703), .A2(n13191), .ZN(n12945) );
  OAI211_X1 U16059 ( .C1(n12946), .C2(n12947), .A(n20705), .B(n12945), .ZN(
        n12965) );
  OAI22_X1 U16060 ( .A1(n12948), .A2(n12947), .B1(n20697), .B2(n13191), .ZN(
        n12964) );
  AOI22_X1 U16061 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12965), .B1(
        n20700), .B2(n12964), .ZN(n12951) );
  AOI22_X1 U16062 ( .A1(n20611), .A2(n20623), .B1(n12966), .B2(n20701), .ZN(
        n12950) );
  OAI211_X1 U16063 ( .C1(n20626), .C2(n13226), .A(n12951), .B(n12950), .ZN(
        P1_U3057) );
  AOI22_X1 U16064 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n12965), .B1(
        n20736), .B2(n12964), .ZN(n12953) );
  INV_X1 U16065 ( .A(n20741), .ZN(n20637) );
  AOI22_X1 U16066 ( .A1(n20611), .A2(n20637), .B1(n12966), .B2(n20737), .ZN(
        n12952) );
  OAI211_X1 U16067 ( .C1(n20640), .C2(n13226), .A(n12953), .B(n12952), .ZN(
        P1_U3062) );
  AOI22_X1 U16068 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12965), .B1(
        n20724), .B2(n12964), .ZN(n12955) );
  INV_X1 U16069 ( .A(n20729), .ZN(n20669) );
  AOI22_X1 U16070 ( .A1(n20611), .A2(n20669), .B1(n12966), .B2(n20725), .ZN(
        n12954) );
  OAI211_X1 U16071 ( .C1(n20672), .C2(n13226), .A(n12955), .B(n12954), .ZN(
        P1_U3060) );
  AOI22_X1 U16072 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12965), .B1(
        n20730), .B2(n12964), .ZN(n12957) );
  INV_X1 U16073 ( .A(n20735), .ZN(n20633) );
  AOI22_X1 U16074 ( .A1(n20611), .A2(n20633), .B1(n12966), .B2(n20731), .ZN(
        n12956) );
  OAI211_X1 U16075 ( .C1(n20636), .C2(n13226), .A(n12957), .B(n12956), .ZN(
        P1_U3061) );
  AOI22_X1 U16076 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12965), .B1(
        n20749), .B2(n12964), .ZN(n12959) );
  INV_X1 U16077 ( .A(n20758), .ZN(n20685) );
  AOI22_X1 U16078 ( .A1(n20611), .A2(n20685), .B1(n12966), .B2(n20751), .ZN(
        n12958) );
  OAI211_X1 U16079 ( .C1(n20691), .C2(n13226), .A(n12959), .B(n12958), .ZN(
        P1_U3064) );
  AOI22_X1 U16080 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12965), .B1(
        n20712), .B2(n12964), .ZN(n12961) );
  INV_X1 U16081 ( .A(n20717), .ZN(n20661) );
  AOI22_X1 U16082 ( .A1(n20611), .A2(n20661), .B1(n12966), .B2(n20713), .ZN(
        n12960) );
  OAI211_X1 U16083 ( .C1(n20664), .C2(n13226), .A(n12961), .B(n12960), .ZN(
        P1_U3058) );
  AOI22_X1 U16084 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12965), .B1(
        n20718), .B2(n12964), .ZN(n12963) );
  INV_X1 U16085 ( .A(n20723), .ZN(n20665) );
  AOI22_X1 U16086 ( .A1(n20611), .A2(n20665), .B1(n12966), .B2(n20719), .ZN(
        n12962) );
  OAI211_X1 U16087 ( .C1(n20668), .C2(n13226), .A(n12963), .B(n12962), .ZN(
        P1_U3059) );
  AOI22_X1 U16088 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12965), .B1(
        n20742), .B2(n12964), .ZN(n12968) );
  INV_X1 U16089 ( .A(n20747), .ZN(n20679) );
  AOI22_X1 U16090 ( .A1(n20611), .A2(n20679), .B1(n12966), .B2(n21074), .ZN(
        n12967) );
  OAI211_X1 U16091 ( .C1(n20682), .C2(n13226), .A(n12968), .B(n12967), .ZN(
        P1_U3063) );
  INV_X1 U16092 ( .A(n12969), .ZN(n12971) );
  XNOR2_X1 U16093 ( .A(n12971), .B(n12970), .ZN(n20455) );
  INV_X1 U16094 ( .A(n20455), .ZN(n12972) );
  INV_X1 U16095 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20411) );
  OAI222_X1 U16096 ( .A1(n14744), .A2(n12973), .B1(n14717), .B2(n12972), .C1(
        n20411), .C2(n14745), .ZN(P1_U2900) );
  OAI222_X1 U16097 ( .A1(n14717), .A2(n12975), .B1(n14745), .B2(n12890), .C1(
        n14744), .C2(n12974), .ZN(P1_U2899) );
  NOR2_X1 U16098 ( .A1(n13095), .A2(n12976), .ZN(n12977) );
  OR2_X1 U16099 ( .A1(n13300), .A2(n12977), .ZN(n15547) );
  NAND2_X1 U16100 ( .A1(n12829), .A2(n13092), .ZN(n12979) );
  INV_X1 U16101 ( .A(n12979), .ZN(n12981) );
  INV_X1 U16102 ( .A(n12978), .ZN(n12980) );
  OR2_X1 U16103 ( .A1(n12979), .A2(n12978), .ZN(n13298) );
  OAI211_X1 U16104 ( .C1(n12981), .C2(n12980), .A(n15281), .B(n13298), .ZN(
        n12983) );
  NAND2_X1 U16105 ( .A1(n15279), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12982) );
  OAI211_X1 U16106 ( .C1(n15547), .C2(n15279), .A(n12983), .B(n12982), .ZN(
        P2_U2873) );
  NAND2_X1 U16107 ( .A1(n12984), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12985) );
  OR2_X1 U16108 ( .A1(n15012), .A2(n13651), .ZN(n12993) );
  NAND2_X1 U16109 ( .A1(n12989), .A2(n12988), .ZN(n13625) );
  INV_X1 U16110 ( .A(n13623), .ZN(n12990) );
  XNOR2_X1 U16111 ( .A(n13625), .B(n12990), .ZN(n12991) );
  NAND2_X1 U16112 ( .A1(n12991), .A2(n13657), .ZN(n12992) );
  NAND2_X1 U16113 ( .A1(n12993), .A2(n12992), .ZN(n12994) );
  OAI21_X1 U16114 ( .B1(n12995), .B2(n12994), .A(n13612), .ZN(n12996) );
  INV_X1 U16115 ( .A(n12996), .ZN(n20475) );
  NAND2_X1 U16116 ( .A1(n20475), .A2(n20457), .ZN(n12999) );
  AND2_X1 U16117 ( .A1(n16482), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20472) );
  NOR2_X1 U16118 ( .A1(n20461), .A2(n13068), .ZN(n12997) );
  AOI211_X1 U16119 ( .C1(n20450), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20472), .B(n12997), .ZN(n12998) );
  OAI211_X1 U16120 ( .C1(n14888), .C2(n13072), .A(n12999), .B(n12998), .ZN(
        P1_U2996) );
  INV_X1 U16121 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13002) );
  INV_X1 U16122 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14250) );
  INV_X1 U16123 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14791) );
  INV_X1 U16124 ( .A(n14310), .ZN(n13004) );
  INV_X1 U16125 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14753) );
  INV_X1 U16126 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13005) );
  INV_X1 U16127 ( .A(n13007), .ZN(n15030) );
  AND2_X1 U16128 ( .A1(n13008), .A2(n16503), .ZN(n13010) );
  AOI22_X1 U16129 ( .A1(n20861), .A2(P1_STATE2_REG_3__SCAN_IN), .B1(n16503), 
        .B2(n20697), .ZN(n13009) );
  AOI21_X1 U16130 ( .B1(n15030), .B2(n13010), .A(n13009), .ZN(n13011) );
  NAND2_X1 U16131 ( .A1(n16238), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13013) );
  INV_X1 U16132 ( .A(n13013), .ZN(n13012) );
  INV_X1 U16133 ( .A(n20855), .ZN(n13025) );
  OAI21_X1 U16134 ( .B1(n13014), .B2(n13025), .A(n16255), .ZN(n20379) );
  NAND2_X1 U16135 ( .A1(n20379), .A2(n13015), .ZN(n13032) );
  OR2_X1 U16136 ( .A1(n13025), .A2(n13016), .ZN(n20364) );
  INV_X1 U16137 ( .A(n20364), .ZN(n13087) );
  AND2_X1 U16138 ( .A1(n20857), .A2(n20702), .ZN(n13017) );
  NAND2_X1 U16139 ( .A1(n9988), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13020) );
  OR2_X1 U16140 ( .A1(n13018), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13023) );
  INV_X1 U16141 ( .A(n13023), .ZN(n13022) );
  NAND2_X1 U16142 ( .A1(n13020), .A2(n13019), .ZN(n13021) );
  AOI22_X1 U16143 ( .A1(n20354), .A2(P1_EBX_REG_2__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20374), .ZN(n13028) );
  INV_X1 U16144 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20846) );
  NOR2_X1 U16145 ( .A1(n16239), .A2(n20846), .ZN(n13026) );
  NAND2_X1 U16146 ( .A1(n16239), .A2(n16238), .ZN(n16303) );
  NAND3_X1 U16147 ( .A1(n20331), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13063) );
  OAI211_X1 U16148 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n13026), .A(n16303), .B(
        n13063), .ZN(n13027) );
  OAI211_X1 U16149 ( .C1(n20479), .C2(n20376), .A(n13028), .B(n13027), .ZN(
        n13029) );
  AOI21_X1 U16150 ( .B1(n13030), .B2(n13087), .A(n13029), .ZN(n13031) );
  OAI211_X1 U16151 ( .C1(n20384), .C2(n13033), .A(n13032), .B(n13031), .ZN(
        P1_U2838) );
  AOI22_X1 U16152 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16153 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16154 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U16155 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13034) );
  NAND4_X1 U16156 ( .A1(n13037), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        n13043) );
  AOI22_X1 U16157 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14219), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16158 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U16159 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16160 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13038) );
  NAND4_X1 U16161 ( .A1(n13041), .A2(n13040), .A3(n13039), .A4(n13038), .ZN(
        n13042) );
  AOI22_X1 U16162 ( .A1(n13167), .A2(n13641), .B1(n13044), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13165) );
  NAND2_X1 U16163 ( .A1(n13164), .A2(n13165), .ZN(n13631) );
  NAND2_X1 U16164 ( .A1(n13631), .A2(n13859), .ZN(n13051) );
  INV_X1 U16165 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13048) );
  OAI21_X1 U16166 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13046), .A(
        n13045), .ZN(n20353) );
  AOI22_X1 U16167 ( .A1(n14345), .A2(n20353), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13047) );
  OAI21_X1 U16168 ( .B1(n14285), .B2(n13048), .A(n13047), .ZN(n13049) );
  INV_X1 U16169 ( .A(n13049), .ZN(n13050) );
  NAND2_X1 U16170 ( .A1(n13051), .A2(n13050), .ZN(n13177) );
  INV_X1 U16171 ( .A(n13177), .ZN(n13052) );
  XNOR2_X1 U16172 ( .A(n9750), .B(n13052), .ZN(n20347) );
  INV_X1 U16173 ( .A(n20370), .ZN(n13056) );
  INV_X1 U16174 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20341) );
  NAND2_X1 U16175 ( .A1(n14399), .A2(n20341), .ZN(n13055) );
  INV_X1 U16176 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20999) );
  NAND2_X1 U16177 ( .A1(n9988), .A2(n20341), .ZN(n13053) );
  OAI211_X1 U16178 ( .C1(n14419), .C2(n20999), .A(n13053), .B(n12753), .ZN(
        n13054) );
  AND2_X1 U16179 ( .A1(n13055), .A2(n13054), .ZN(n13058) );
  AOI21_X1 U16180 ( .B1(n13056), .B2(n13057), .A(n13058), .ZN(n13060) );
  NAND2_X1 U16181 ( .A1(n13058), .A2(n13057), .ZN(n13059) );
  OR2_X1 U16182 ( .A1(n13060), .A2(n13358), .ZN(n20342) );
  OAI22_X1 U16183 ( .A1(n20385), .A2(n20342), .B1(n20341), .B2(n20390), .ZN(
        n13061) );
  AOI21_X1 U16184 ( .B1(n20347), .B2(n20387), .A(n13061), .ZN(n13062) );
  INV_X1 U16185 ( .A(n13062), .ZN(P1_U2866) );
  INV_X1 U16186 ( .A(n20379), .ZN(n13091) );
  INV_X1 U16187 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20785) );
  OAI21_X1 U16188 ( .B1(n20329), .B2(n20785), .A(n13063), .ZN(n13065) );
  INV_X1 U16189 ( .A(n20381), .ZN(n13064) );
  NAND2_X1 U16190 ( .A1(n13065), .A2(n13064), .ZN(n13067) );
  AOI22_X1 U16191 ( .A1(n20354), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20374), .ZN(n13066) );
  OAI211_X1 U16192 ( .C1(n20471), .C2(n20376), .A(n13067), .B(n13066), .ZN(
        n13070) );
  NOR2_X1 U16193 ( .A1(n20384), .A2(n13068), .ZN(n13069) );
  AOI211_X1 U16194 ( .C1(n13087), .C2(n12677), .A(n13070), .B(n13069), .ZN(
        n13071) );
  OAI21_X1 U16195 ( .B1(n13091), .B2(n13072), .A(n13071), .ZN(P1_U2837) );
  OAI22_X1 U16196 ( .A1(n20316), .A2(n13078), .B1(n20846), .B2(n16238), .ZN(
        n13073) );
  AOI21_X1 U16197 ( .B1(n20354), .B2(P1_EBX_REG_1__SCAN_IN), .A(n13073), .ZN(
        n13076) );
  AOI22_X1 U16198 ( .A1(n20331), .A2(n20846), .B1(n20356), .B2(n13074), .ZN(
        n13075) );
  OAI211_X1 U16199 ( .C1(n20591), .C2(n20364), .A(n13076), .B(n13075), .ZN(
        n13077) );
  AOI21_X1 U16200 ( .B1(n20322), .B2(n13078), .A(n13077), .ZN(n13079) );
  OAI21_X1 U16201 ( .B1(n13091), .B2(n13080), .A(n13079), .ZN(P1_U2839) );
  NAND2_X1 U16202 ( .A1(n16303), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13082) );
  NAND2_X1 U16203 ( .A1(n20354), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13081) );
  OAI211_X1 U16204 ( .C1(n20376), .C2(n13083), .A(n13082), .B(n13081), .ZN(
        n13086) );
  AOI21_X1 U16205 ( .B1(n20384), .B2(n20316), .A(n13084), .ZN(n13085) );
  AOI211_X1 U16206 ( .C1(n13088), .C2(n13087), .A(n13086), .B(n13085), .ZN(
        n13089) );
  OAI21_X1 U16207 ( .B1(n13091), .B2(n13090), .A(n13089), .ZN(P1_U2840) );
  XNOR2_X1 U16208 ( .A(n12829), .B(n13092), .ZN(n13098) );
  AND2_X1 U16209 ( .A1(n13094), .A2(n13093), .ZN(n13096) );
  OR2_X1 U16210 ( .A1(n13096), .A2(n13095), .ZN(n15795) );
  MUX2_X1 U16211 ( .A(n15795), .B(n10928), .S(n15279), .Z(n13097) );
  OAI21_X1 U16212 ( .B1(n13098), .B2(n15298), .A(n13097), .ZN(P2_U2874) );
  INV_X1 U16213 ( .A(n20347), .ZN(n13099) );
  OAI222_X1 U16214 ( .A1(n14744), .A2(n13100), .B1(n14717), .B2(n13099), .C1(
        n13048), .C2(n14745), .ZN(P1_U2898) );
  NAND2_X1 U16215 ( .A1(n15035), .A2(n13670), .ZN(n20678) );
  OAI21_X1 U16216 ( .B1(n20686), .B2(n13103), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13101) );
  NAND2_X1 U16217 ( .A1(n13101), .A2(n20658), .ZN(n13113) );
  INV_X1 U16218 ( .A(n13113), .ZN(n13102) );
  NOR2_X1 U16219 ( .A1(n20650), .A2(n20591), .ZN(n13112) );
  NAND2_X1 U16220 ( .A1(n20523), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13108) );
  INV_X1 U16221 ( .A(n13108), .ZN(n13500) );
  AND2_X1 U16222 ( .A1(n13107), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20529) );
  INV_X1 U16223 ( .A(n13103), .ZN(n13135) );
  INV_X1 U16224 ( .A(n13104), .ZN(n13105) );
  NOR2_X1 U16225 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13105), .ZN(
        n13109) );
  INV_X1 U16226 ( .A(n13109), .ZN(n13134) );
  OAI22_X1 U16227 ( .A1(n13135), .A2(n20735), .B1(n13134), .B2(n13224), .ZN(
        n13106) );
  AOI21_X1 U16228 ( .B1(n20686), .B2(n20732), .A(n13106), .ZN(n13115) );
  OR2_X1 U16229 ( .A1(n13107), .A2(n20697), .ZN(n20587) );
  INV_X1 U16230 ( .A(n20587), .ZN(n13675) );
  NAND2_X1 U16231 ( .A1(n13108), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13497) );
  OAI21_X1 U16232 ( .B1(n16512), .B2(n13109), .A(n13497), .ZN(n13110) );
  INV_X1 U16233 ( .A(n13110), .ZN(n13111) );
  NAND2_X1 U16234 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13114) );
  OAI211_X1 U16235 ( .C1(n13140), .C2(n13717), .A(n13115), .B(n13114), .ZN(
        P1_U3117) );
  OAI22_X1 U16236 ( .A1(n13135), .A2(n20717), .B1(n13134), .B2(n13192), .ZN(
        n13116) );
  AOI21_X1 U16237 ( .B1(n20686), .B2(n20714), .A(n13116), .ZN(n13118) );
  NAND2_X1 U16238 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13117) );
  OAI211_X1 U16239 ( .C1(n13140), .C2(n13690), .A(n13118), .B(n13117), .ZN(
        P1_U3114) );
  OAI22_X1 U16240 ( .A1(n13135), .A2(n20741), .B1(n13134), .B2(n13208), .ZN(
        n13119) );
  AOI21_X1 U16241 ( .B1(n20686), .B2(n20738), .A(n13119), .ZN(n13121) );
  NAND2_X1 U16242 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13120) );
  OAI211_X1 U16243 ( .C1(n13140), .C2(n13710), .A(n13121), .B(n13120), .ZN(
        P1_U3118) );
  OAI22_X1 U16244 ( .A1(n13135), .A2(n20711), .B1(n13134), .B2(n13220), .ZN(
        n13122) );
  AOI21_X1 U16245 ( .B1(n20686), .B2(n20708), .A(n13122), .ZN(n13124) );
  NAND2_X1 U16246 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13123) );
  OAI211_X1 U16247 ( .C1(n13140), .C2(n13686), .A(n13124), .B(n13123), .ZN(
        P1_U3113) );
  OAI22_X1 U16248 ( .A1(n13135), .A2(n20729), .B1(n13134), .B2(n13200), .ZN(
        n13125) );
  AOI21_X1 U16249 ( .B1(n20686), .B2(n20726), .A(n13125), .ZN(n13127) );
  NAND2_X1 U16250 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13126) );
  OAI211_X1 U16251 ( .C1(n13140), .C2(n13694), .A(n13127), .B(n13126), .ZN(
        P1_U3116) );
  OAI22_X1 U16252 ( .A1(n13135), .A2(n20758), .B1(n13134), .B2(n13216), .ZN(
        n13128) );
  AOI21_X1 U16253 ( .B1(n20686), .B2(n20752), .A(n13128), .ZN(n13130) );
  NAND2_X1 U16254 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13129) );
  OAI211_X1 U16255 ( .C1(n13140), .C2(n13702), .A(n13130), .B(n13129), .ZN(
        P1_U3120) );
  OAI22_X1 U16256 ( .A1(n13135), .A2(n20747), .B1(n13134), .B2(n13204), .ZN(
        n13131) );
  AOI21_X1 U16257 ( .B1(n20686), .B2(n20744), .A(n13131), .ZN(n13133) );
  NAND2_X1 U16258 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13132) );
  OAI211_X1 U16259 ( .C1(n13140), .C2(n13698), .A(n13133), .B(n13132), .ZN(
        P1_U3119) );
  OAI22_X1 U16260 ( .A1(n13135), .A2(n20723), .B1(n13134), .B2(n13212), .ZN(
        n13136) );
  AOI21_X1 U16261 ( .B1(n20686), .B2(n20720), .A(n13136), .ZN(n13139) );
  NAND2_X1 U16262 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13138) );
  OAI211_X1 U16263 ( .C1(n13140), .C2(n13706), .A(n13139), .B(n13138), .ZN(
        P1_U3115) );
  NAND2_X1 U16264 ( .A1(n13142), .A2(n13141), .ZN(n13144) );
  XNOR2_X1 U16265 ( .A(n13144), .B(n13143), .ZN(n13163) );
  XOR2_X1 U16266 ( .A(n10851), .B(n13145), .Z(n13161) );
  NOR2_X1 U16267 ( .A1(n13147), .A2(n13146), .ZN(n13149) );
  MUX2_X1 U16268 ( .A(n13149), .B(n13148), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13155) );
  XNOR2_X1 U16269 ( .A(n13151), .B(n13150), .ZN(n19454) );
  INV_X1 U16270 ( .A(n19454), .ZN(n20228) );
  INV_X1 U16271 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20154) );
  NOR2_X1 U16272 ( .A1(n20154), .A2(n15727), .ZN(n13152) );
  AOI21_X1 U16273 ( .B1(n16669), .B2(n20228), .A(n13152), .ZN(n13153) );
  OAI21_X1 U16274 ( .B1(n9891), .B2(n16702), .A(n13153), .ZN(n13154) );
  AOI211_X1 U16275 ( .C1(n13161), .C2(n16690), .A(n13155), .B(n13154), .ZN(
        n13156) );
  OAI21_X1 U16276 ( .B1(n13163), .B2(n16697), .A(n13156), .ZN(P2_U3043) );
  AOI22_X1 U16277 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n19529), .ZN(n13159) );
  AOI21_X1 U16278 ( .B1(n13273), .B2(n13157), .A(n13237), .ZN(n13271) );
  NAND2_X1 U16279 ( .A1(n16658), .A2(n13271), .ZN(n13158) );
  OAI211_X1 U16280 ( .C1(n9891), .C2(n16648), .A(n13159), .B(n13158), .ZN(
        n13160) );
  AOI21_X1 U16281 ( .B1(n13161), .B2(n16660), .A(n13160), .ZN(n13162) );
  OAI21_X1 U16282 ( .B1(n13163), .B2(n19534), .A(n13162), .ZN(P2_U3011) );
  INV_X1 U16283 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13170) );
  NAND2_X1 U16284 ( .A1(n13167), .A2(n13656), .ZN(n13168) );
  OAI21_X1 U16285 ( .B1(n13170), .B2(n13169), .A(n13168), .ZN(n13171) );
  INV_X1 U16286 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13175) );
  OAI21_X1 U16287 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13173), .A(
        n13172), .ZN(n20334) );
  AOI22_X1 U16288 ( .A1(n14345), .A2(n20334), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13174) );
  OAI21_X1 U16289 ( .B1(n14285), .B2(n13175), .A(n13174), .ZN(n13176) );
  NAND2_X1 U16290 ( .A1(n13179), .A2(n13178), .ZN(n13350) );
  NAND2_X1 U16291 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  AND2_X1 U16292 ( .A1(n13350), .A2(n13182), .ZN(n20338) );
  INV_X1 U16293 ( .A(n20338), .ZN(n13188) );
  OAI222_X1 U16294 ( .A1(n14717), .A2(n13188), .B1(n14745), .B2(n13175), .C1(
        n14744), .C2(n13183), .ZN(P1_U2897) );
  INV_X1 U16295 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13187) );
  INV_X1 U16296 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16469) );
  OAI21_X1 U16297 ( .B1(n14419), .B2(n16469), .A(n12753), .ZN(n13185) );
  OAI21_X1 U16298 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n14456), .A(n13185), .ZN(
        n13186) );
  OAI21_X1 U16299 ( .B1(n14410), .B2(P1_EBX_REG_7__SCAN_IN), .A(n13186), .ZN(
        n13355) );
  XNOR2_X1 U16300 ( .A(n13358), .B(n13355), .ZN(n16481) );
  OAI222_X1 U16301 ( .A1(n14666), .A2(n13188), .B1(n13187), .B2(n20390), .C1(
        n20385), .C2(n16481), .ZN(P1_U2865) );
  INV_X1 U16302 ( .A(n20578), .ZN(n13189) );
  AOI21_X1 U16303 ( .B1(n13189), .B2(n13226), .A(n20702), .ZN(n13190) );
  NOR2_X1 U16304 ( .A1(n13190), .A2(n20703), .ZN(n13194) );
  NOR2_X1 U16305 ( .A1(n20522), .A2(n20591), .ZN(n13196) );
  INV_X1 U16306 ( .A(n20523), .ZN(n13542) );
  NOR2_X1 U16307 ( .A1(n13542), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13674) );
  OR2_X1 U16308 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13191), .ZN(
        n13225) );
  OAI22_X1 U16309 ( .A1(n13226), .A2(n20717), .B1(n13225), .B2(n13192), .ZN(
        n13193) );
  AOI21_X1 U16310 ( .B1(n20578), .B2(n20714), .A(n13193), .ZN(n13199) );
  INV_X1 U16311 ( .A(n13194), .ZN(n13197) );
  NOR2_X1 U16312 ( .A1(n13674), .A2(n20697), .ZN(n13679) );
  AOI21_X1 U16313 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n13225), .A(n13679), 
        .ZN(n13195) );
  NAND2_X1 U16314 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13198) );
  OAI211_X1 U16315 ( .C1(n13231), .C2(n13690), .A(n13199), .B(n13198), .ZN(
        P1_U3050) );
  OAI22_X1 U16316 ( .A1(n13226), .A2(n20729), .B1(n13225), .B2(n13200), .ZN(
        n13201) );
  AOI21_X1 U16317 ( .B1(n20578), .B2(n20726), .A(n13201), .ZN(n13203) );
  NAND2_X1 U16318 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13202) );
  OAI211_X1 U16319 ( .C1(n13231), .C2(n13694), .A(n13203), .B(n13202), .ZN(
        P1_U3052) );
  OAI22_X1 U16320 ( .A1(n13226), .A2(n20747), .B1(n13225), .B2(n13204), .ZN(
        n13205) );
  AOI21_X1 U16321 ( .B1(n20578), .B2(n20744), .A(n13205), .ZN(n13207) );
  NAND2_X1 U16322 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13206) );
  OAI211_X1 U16323 ( .C1(n13231), .C2(n13698), .A(n13207), .B(n13206), .ZN(
        P1_U3055) );
  OAI22_X1 U16324 ( .A1(n13226), .A2(n20741), .B1(n13225), .B2(n13208), .ZN(
        n13209) );
  AOI21_X1 U16325 ( .B1(n20578), .B2(n20738), .A(n13209), .ZN(n13211) );
  NAND2_X1 U16326 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13210) );
  OAI211_X1 U16327 ( .C1(n13231), .C2(n13710), .A(n13211), .B(n13210), .ZN(
        P1_U3054) );
  OAI22_X1 U16328 ( .A1(n13226), .A2(n20723), .B1(n13225), .B2(n13212), .ZN(
        n13213) );
  AOI21_X1 U16329 ( .B1(n20578), .B2(n20720), .A(n13213), .ZN(n13215) );
  NAND2_X1 U16330 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13214) );
  OAI211_X1 U16331 ( .C1(n13231), .C2(n13706), .A(n13215), .B(n13214), .ZN(
        P1_U3051) );
  OAI22_X1 U16332 ( .A1(n13226), .A2(n20758), .B1(n13225), .B2(n13216), .ZN(
        n13217) );
  AOI21_X1 U16333 ( .B1(n20578), .B2(n20752), .A(n13217), .ZN(n13219) );
  NAND2_X1 U16334 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13218) );
  OAI211_X1 U16335 ( .C1(n13231), .C2(n13702), .A(n13219), .B(n13218), .ZN(
        P1_U3056) );
  OAI22_X1 U16336 ( .A1(n13226), .A2(n20711), .B1(n13225), .B2(n13220), .ZN(
        n13221) );
  AOI21_X1 U16337 ( .B1(n20578), .B2(n20708), .A(n13221), .ZN(n13223) );
  NAND2_X1 U16338 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13222) );
  OAI211_X1 U16339 ( .C1(n13231), .C2(n13686), .A(n13223), .B(n13222), .ZN(
        P1_U3049) );
  OAI22_X1 U16340 ( .A1(n13226), .A2(n20735), .B1(n13225), .B2(n13224), .ZN(
        n13227) );
  AOI21_X1 U16341 ( .B1(n20578), .B2(n20732), .A(n13227), .ZN(n13230) );
  NAND2_X1 U16342 ( .A1(n13228), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13229) );
  OAI211_X1 U16343 ( .C1(n13231), .C2(n13717), .A(n13230), .B(n13229), .ZN(
        P1_U3053) );
  INV_X1 U16344 ( .A(n20276), .ZN(n20274) );
  NOR2_X1 U16345 ( .A1(n20274), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13250) );
  INV_X1 U16346 ( .A(n13250), .ZN(n13261) );
  NAND2_X1 U16347 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13261), .ZN(n13232) );
  NOR2_X1 U16348 ( .A1(n13262), .A2(n13232), .ZN(n13233) );
  NAND2_X1 U16349 ( .A1(n19272), .A2(n13233), .ZN(n19404) );
  INV_X1 U16350 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20278) );
  AOI21_X1 U16351 ( .B1(n16635), .B2(n13244), .A(n13245), .ZN(n16624) );
  AOI21_X1 U16352 ( .B1(n16645), .B2(n13240), .A(n13242), .ZN(n16636) );
  AOI21_X1 U16353 ( .B1(n16656), .B2(n13238), .A(n13241), .ZN(n16646) );
  AOI21_X1 U16354 ( .B1(n16667), .B2(n13236), .A(n13239), .ZN(n16657) );
  OAI22_X1 U16355 ( .A1(n20278), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15875) );
  OAI22_X1 U16356 ( .A1(n20278), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n12092), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15874) );
  AND2_X1 U16357 ( .A1(n15875), .A2(n15874), .ZN(n15210) );
  NAND2_X1 U16358 ( .A1(n15210), .A2(n15212), .ZN(n13269) );
  NOR2_X1 U16359 ( .A1(n13271), .A2(n13269), .ZN(n19378) );
  OAI21_X1 U16360 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13237), .A(
        n13236), .ZN(n19541) );
  NAND2_X1 U16361 ( .A1(n19378), .A2(n19541), .ZN(n13286) );
  NOR2_X1 U16362 ( .A1(n16657), .A2(n13286), .ZN(n19367) );
  OAI21_X1 U16363 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13239), .A(
        n13238), .ZN(n19368) );
  NAND2_X1 U16364 ( .A1(n19367), .A2(n19368), .ZN(n13309) );
  NOR2_X1 U16365 ( .A1(n16646), .A2(n13309), .ZN(n19356) );
  OAI21_X1 U16366 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13241), .A(
        n13240), .ZN(n19357) );
  NAND2_X1 U16367 ( .A1(n19356), .A2(n19357), .ZN(n13320) );
  NOR2_X1 U16368 ( .A1(n16636), .A2(n13320), .ZN(n19344) );
  OR2_X1 U16369 ( .A1(n13242), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13243) );
  NAND2_X1 U16370 ( .A1(n13244), .A2(n13243), .ZN(n19345) );
  NAND2_X1 U16371 ( .A1(n19344), .A2(n19345), .ZN(n15195) );
  NOR2_X1 U16372 ( .A1(n16624), .A2(n15195), .ZN(n15194) );
  NOR2_X1 U16373 ( .A1(n19379), .A2(n15194), .ZN(n13247) );
  OR2_X1 U16374 ( .A1(n13245), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13246) );
  NAND2_X1 U16375 ( .A1(n15099), .A2(n13246), .ZN(n15577) );
  XNOR2_X1 U16376 ( .A(n13247), .B(n15577), .ZN(n13248) );
  NAND2_X1 U16377 ( .A1(n13248), .A2(n9671), .ZN(n13267) );
  NOR2_X1 U16378 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n16729), .ZN(n16755) );
  INV_X1 U16379 ( .A(n16755), .ZN(n13249) );
  NAND2_X1 U16380 ( .A1(n12463), .A2(n13249), .ZN(n16521) );
  NOR2_X1 U16381 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13250), .ZN(n13251) );
  NAND2_X1 U16382 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NOR2_X1 U16383 ( .A1(n20268), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19800) );
  AND2_X1 U16384 ( .A1(n13254), .A2(n19800), .ZN(n16765) );
  NOR2_X1 U16385 ( .A1(n9671), .A2(n16765), .ZN(n13255) );
  NAND2_X1 U16386 ( .A1(n15727), .A2(n13255), .ZN(n13256) );
  INV_X1 U16387 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13260) );
  XOR2_X1 U16388 ( .A(n13257), .B(n15198), .Z(n19436) );
  NAND2_X1 U16389 ( .A1(n19377), .A2(n19436), .ZN(n13259) );
  NOR2_X2 U16390 ( .A1(n19392), .A2(n20268), .ZN(n19417) );
  AOI21_X1 U16391 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19417), .A(
        n19529), .ZN(n13258) );
  OAI211_X1 U16392 ( .C1(n19405), .C2(n13260), .A(n13259), .B(n13258), .ZN(
        n13265) );
  NOR2_X1 U16393 ( .A1(n13262), .A2(n13261), .ZN(n13263) );
  NOR2_X1 U16394 ( .A1(n15807), .A2(n19413), .ZN(n13264) );
  AOI211_X1 U16395 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19411), .A(n13265), .B(
        n13264), .ZN(n13266) );
  OAI211_X1 U16396 ( .C1(n19404), .C2(n13268), .A(n13267), .B(n13266), .ZN(
        P2_U2843) );
  NAND2_X1 U16397 ( .A1(n9661), .A2(n13269), .ZN(n13270) );
  XNOR2_X1 U16398 ( .A(n13271), .B(n13270), .ZN(n13272) );
  NAND2_X1 U16399 ( .A1(n13272), .A2(n9671), .ZN(n13280) );
  OAI22_X1 U16400 ( .A1(n19352), .A2(n13274), .B1(n13273), .B2(n19389), .ZN(
        n13277) );
  NOR2_X1 U16401 ( .A1(n19404), .A2(n13275), .ZN(n13276) );
  AOI211_X1 U16402 ( .C1(n19392), .C2(P2_REIP_REG_3__SCAN_IN), .A(n13277), .B(
        n13276), .ZN(n13278) );
  OAI21_X1 U16403 ( .B1(n19408), .B2(n19454), .A(n13278), .ZN(n13279) );
  OAI211_X1 U16404 ( .C1(n19860), .C2(n19382), .A(n13280), .B(n9705), .ZN(
        P2_U2852) );
  INV_X1 U16405 ( .A(n13281), .ZN(n13282) );
  NAND2_X1 U16406 ( .A1(n13283), .A2(n13282), .ZN(n13284) );
  AND2_X1 U16407 ( .A1(n13285), .A2(n13284), .ZN(n19459) );
  INV_X1 U16408 ( .A(n19459), .ZN(n13296) );
  NAND2_X1 U16409 ( .A1(n9661), .A2(n13286), .ZN(n13287) );
  XNOR2_X1 U16410 ( .A(n16657), .B(n13287), .ZN(n13288) );
  NAND2_X1 U16411 ( .A1(n13288), .A2(n9671), .ZN(n13295) );
  NAND2_X1 U16412 ( .A1(n19411), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13291) );
  INV_X1 U16413 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20157) );
  OAI21_X1 U16414 ( .B1(n20157), .B2(n19405), .A(n15727), .ZN(n13289) );
  AOI21_X1 U16415 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19417), .A(
        n13289), .ZN(n13290) );
  OAI211_X1 U16416 ( .C1(n19404), .C2(n13292), .A(n13291), .B(n13290), .ZN(
        n13293) );
  AOI21_X1 U16417 ( .B1(n16659), .B2(n19396), .A(n13293), .ZN(n13294) );
  OAI211_X1 U16418 ( .C1(n19408), .C2(n13296), .A(n13295), .B(n13294), .ZN(
        P2_U2850) );
  XNOR2_X1 U16419 ( .A(n13298), .B(n13297), .ZN(n13303) );
  OR2_X1 U16420 ( .A1(n13300), .A2(n13299), .ZN(n13301) );
  NAND2_X1 U16421 ( .A1(n13398), .A2(n13301), .ZN(n15769) );
  INV_X1 U16422 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n15177) );
  MUX2_X1 U16423 ( .A(n15769), .B(n15177), .S(n15279), .Z(n13302) );
  OAI21_X1 U16424 ( .B1(n13303), .B2(n15298), .A(n13302), .ZN(P2_U2872) );
  AOI21_X1 U16425 ( .B1(n13306), .B2(n13305), .A(n13304), .ZN(n13307) );
  INV_X1 U16426 ( .A(n13307), .ZN(n19452) );
  NAND2_X1 U16427 ( .A1(n13308), .A2(n13309), .ZN(n13310) );
  XNOR2_X1 U16428 ( .A(n16646), .B(n13310), .ZN(n13311) );
  NAND2_X1 U16429 ( .A1(n13311), .A2(n9671), .ZN(n13319) );
  INV_X1 U16430 ( .A(n16649), .ZN(n13317) );
  INV_X1 U16431 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n13312) );
  OAI21_X1 U16432 ( .B1(n19405), .B2(n13312), .A(n15727), .ZN(n13316) );
  AOI22_X1 U16433 ( .A1(n19411), .A2(P2_EBX_REG_7__SCAN_IN), .B1(n13313), .B2(
        n19294), .ZN(n13314) );
  OAI21_X1 U16434 ( .B1(n16656), .B2(n19389), .A(n13314), .ZN(n13315) );
  AOI211_X1 U16435 ( .C1(n13317), .C2(n19396), .A(n13316), .B(n13315), .ZN(
        n13318) );
  OAI211_X1 U16436 ( .C1(n19408), .C2(n19452), .A(n13319), .B(n13318), .ZN(
        P2_U2848) );
  NAND2_X1 U16437 ( .A1(n13308), .A2(n13320), .ZN(n13321) );
  XNOR2_X1 U16438 ( .A(n16636), .B(n13321), .ZN(n13322) );
  NAND2_X1 U16439 ( .A1(n13322), .A2(n9671), .ZN(n13332) );
  INV_X1 U16440 ( .A(n13323), .ZN(n13326) );
  INV_X1 U16441 ( .A(n13324), .ZN(n16683) );
  AOI21_X1 U16442 ( .B1(n13326), .B2(n16683), .A(n13325), .ZN(n19445) );
  NAND2_X1 U16443 ( .A1(n19392), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n13327) );
  OAI211_X1 U16444 ( .C1(n16645), .C2(n19389), .A(n13327), .B(n15727), .ZN(
        n13328) );
  AOI21_X1 U16445 ( .B1(n19445), .B2(n19377), .A(n13328), .ZN(n13329) );
  OAI21_X1 U16446 ( .B1(n16639), .B2(n19413), .A(n13329), .ZN(n13330) );
  AOI21_X1 U16447 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(n19411), .A(n13330), .ZN(
        n13331) );
  OAI211_X1 U16448 ( .C1(n19404), .C2(n13333), .A(n13332), .B(n13331), .ZN(
        P2_U2846) );
  INV_X1 U16449 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13373) );
  XNOR2_X1 U16450 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13334), .ZN(
        n13661) );
  AOI22_X1 U16451 ( .A1(n14345), .A2(n13661), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13335) );
  OAI21_X1 U16452 ( .B1(n14285), .B2(n13373), .A(n13335), .ZN(n13336) );
  INV_X1 U16453 ( .A(n13336), .ZN(n13349) );
  AOI22_X1 U16454 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U16455 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13340) );
  AOI22_X1 U16456 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13339) );
  AOI22_X1 U16457 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13338) );
  NAND4_X1 U16458 ( .A1(n13341), .A2(n13340), .A3(n13339), .A4(n13338), .ZN(
        n13347) );
  AOI22_X1 U16459 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U16460 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14219), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U16461 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U16462 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13342) );
  NAND4_X1 U16463 ( .A1(n13345), .A2(n13344), .A3(n13343), .A4(n13342), .ZN(
        n13346) );
  OAI21_X1 U16464 ( .B1(n13347), .B2(n13346), .A(n13859), .ZN(n13348) );
  AOI21_X1 U16465 ( .B1(n13351), .B2(n13350), .A(n13388), .ZN(n13368) );
  INV_X1 U16466 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13361) );
  NAND2_X1 U16467 ( .A1(n14399), .A2(n13361), .ZN(n13354) );
  INV_X1 U16468 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16468) );
  NAND2_X1 U16469 ( .A1(n9988), .A2(n13361), .ZN(n13352) );
  OAI211_X1 U16470 ( .C1(n14419), .C2(n16468), .A(n13352), .B(n12753), .ZN(
        n13353) );
  AND2_X1 U16471 ( .A1(n13354), .A2(n13353), .ZN(n13356) );
  AOI21_X1 U16472 ( .B1(n13358), .B2(n13355), .A(n13356), .ZN(n13359) );
  AND2_X1 U16473 ( .A1(n13356), .A2(n13355), .ZN(n13357) );
  NOR2_X1 U16474 ( .A1(n13359), .A2(n13413), .ZN(n16471) );
  AOI21_X1 U16475 ( .B1(n20374), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16482), .ZN(n13360) );
  OAI21_X1 U16476 ( .B1(n13361), .B2(n20372), .A(n13360), .ZN(n13362) );
  AOI21_X1 U16477 ( .B1(n16471), .B2(n20356), .A(n13362), .ZN(n13363) );
  OAI21_X1 U16478 ( .B1(n20384), .B2(n13661), .A(n13363), .ZN(n13366) );
  INV_X1 U16479 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20790) );
  NAND3_X1 U16480 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n20336) );
  NOR2_X1 U16481 ( .A1(n20790), .A2(n20336), .ZN(n14465) );
  INV_X1 U16482 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20793) );
  AOI211_X1 U16483 ( .C1(n13364), .C2(n20793), .A(n20329), .B(n20325), .ZN(
        n13365) );
  AOI211_X1 U16484 ( .C1(n13368), .C2(n20348), .A(n13366), .B(n13365), .ZN(
        n13367) );
  INV_X1 U16485 ( .A(n13367), .ZN(P1_U2832) );
  INV_X1 U16486 ( .A(n13368), .ZN(n13665) );
  AOI22_X1 U16487 ( .A1(n16471), .A2(n16315), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14649), .ZN(n13369) );
  OAI21_X1 U16488 ( .B1(n13665), .B2(n14666), .A(n13369), .ZN(P1_U2864) );
  INV_X1 U16489 ( .A(DATAI_8_), .ZN(n13371) );
  NAND2_X1 U16490 ( .A1(n14482), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13370) );
  OAI21_X1 U16491 ( .B1(n14482), .B2(n13371), .A(n13370), .ZN(n20419) );
  INV_X1 U16492 ( .A(n20419), .ZN(n13372) );
  OAI222_X1 U16493 ( .A1(n13665), .A2(n14717), .B1(n13373), .B2(n14745), .C1(
        n14744), .C2(n13372), .ZN(P1_U2896) );
  XNOR2_X1 U16494 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13374), .ZN(
        n20321) );
  AOI22_X1 U16495 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U16496 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13377) );
  AOI22_X1 U16497 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U16498 ( .A1(n14337), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13375) );
  NAND4_X1 U16499 ( .A1(n13378), .A2(n13377), .A3(n13376), .A4(n13375), .ZN(
        n13384) );
  AOI22_X1 U16500 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11989), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13382) );
  AOI22_X1 U16501 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13381) );
  AOI22_X1 U16502 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U16503 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13379) );
  NAND4_X1 U16504 ( .A1(n13382), .A2(n13381), .A3(n13380), .A4(n13379), .ZN(
        n13383) );
  OR2_X1 U16505 ( .A1(n13384), .A2(n13383), .ZN(n13385) );
  AOI22_X1 U16506 ( .A1(n13859), .A2(n13385), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U16507 ( .A1(n14445), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13386) );
  OAI211_X1 U16508 ( .C1(n20321), .C2(n14351), .A(n13387), .B(n13386), .ZN(
        n13389) );
  NOR2_X1 U16509 ( .A1(n13388), .A2(n13389), .ZN(n13390) );
  OR2_X1 U16510 ( .A1(n9756), .A2(n13390), .ZN(n20320) );
  INV_X1 U16511 ( .A(n14744), .ZN(n13483) );
  INV_X1 U16512 ( .A(DATAI_9_), .ZN(n13392) );
  NAND2_X1 U16513 ( .A1(n14482), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13391) );
  OAI21_X1 U16514 ( .B1(n14482), .B2(n13392), .A(n13391), .ZN(n20421) );
  AOI22_X1 U16515 ( .A1(n13483), .A2(n20421), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n21063), .ZN(n13393) );
  OAI21_X1 U16516 ( .B1(n20320), .B2(n14717), .A(n13393), .ZN(P1_U2895) );
  OAI21_X1 U16517 ( .B1(n13396), .B2(n13395), .A(n13394), .ZN(n13409) );
  NAND2_X1 U16518 ( .A1(n13398), .A2(n13397), .ZN(n13399) );
  NAND2_X1 U16519 ( .A1(n13441), .A2(n13399), .ZN(n19319) );
  MUX2_X1 U16520 ( .A(n19319), .B(n10936), .S(n15279), .Z(n13400) );
  OAI21_X1 U16521 ( .B1(n13409), .B2(n15298), .A(n13400), .ZN(P2_U2871) );
  NOR2_X1 U16522 ( .A1(n9759), .A2(n13401), .ZN(n13402) );
  OR2_X1 U16523 ( .A1(n13433), .A2(n13402), .ZN(n19326) );
  INV_X1 U16524 ( .A(n19326), .ZN(n13407) );
  OAI22_X1 U16525 ( .A1(n19427), .A2(n19553), .B1(n13403), .B2(n19463), .ZN(
        n13406) );
  INV_X1 U16526 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n13404) );
  INV_X1 U16527 ( .A(n19420), .ZN(n15305) );
  INV_X1 U16528 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14733) );
  OAI22_X1 U16529 ( .A1(n15350), .A2(n13404), .B1(n15305), .B2(n14733), .ZN(
        n13405) );
  AOI211_X1 U16530 ( .C1(n19486), .C2(n13407), .A(n13406), .B(n13405), .ZN(
        n13408) );
  OAI21_X1 U16531 ( .B1(n13409), .B2(n19458), .A(n13408), .ZN(P2_U2903) );
  INV_X1 U16532 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13415) );
  INV_X1 U16533 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14425) );
  OAI21_X1 U16534 ( .B1(n14419), .B2(n14425), .A(n12753), .ZN(n13410) );
  OAI21_X1 U16535 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n14456), .A(n13410), .ZN(
        n13411) );
  OAI21_X1 U16536 ( .B1(n14410), .B2(P1_EBX_REG_9__SCAN_IN), .A(n13411), .ZN(
        n13412) );
  NAND2_X1 U16537 ( .A1(n13413), .A2(n13412), .ZN(n13488) );
  OR2_X1 U16538 ( .A1(n13413), .A2(n13412), .ZN(n13414) );
  NAND2_X1 U16539 ( .A1(n13488), .A2(n13414), .ZN(n20317) );
  OAI222_X1 U16540 ( .A1(n20320), .A2(n14666), .B1(n13415), .B2(n20390), .C1(
        n20317), .C2(n20385), .ZN(P1_U2863) );
  OAI21_X1 U16541 ( .B1(n13417), .B2(n13422), .A(n13416), .ZN(n13418) );
  INV_X1 U16542 ( .A(n13418), .ZN(n19533) );
  XOR2_X1 U16543 ( .A(n13419), .B(n13420), .Z(n19531) );
  NAND2_X1 U16544 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19529), .ZN(n13421) );
  OAI221_X1 U16545 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13423), .C1(
        n13422), .C2(n13456), .A(n13421), .ZN(n13428) );
  XOR2_X1 U16546 ( .A(n13425), .B(n13424), .Z(n19464) );
  INV_X1 U16547 ( .A(n19464), .ZN(n13426) );
  OAI22_X1 U16548 ( .A1(n13426), .A2(n16701), .B1(n16702), .B2(n19381), .ZN(
        n13427) );
  AOI211_X1 U16549 ( .C1(n19531), .C2(n16673), .A(n13428), .B(n13427), .ZN(
        n13429) );
  OAI21_X1 U16550 ( .B1(n19533), .B2(n16710), .A(n13429), .ZN(P2_U3042) );
  INV_X1 U16551 ( .A(n13577), .ZN(n13430) );
  AOI21_X1 U16552 ( .B1(n13431), .B2(n13394), .A(n13430), .ZN(n13443) );
  INV_X1 U16553 ( .A(n13443), .ZN(n13439) );
  OAI21_X1 U16554 ( .B1(n13433), .B2(n13432), .A(n13581), .ZN(n15746) );
  INV_X1 U16555 ( .A(n15746), .ZN(n13436) );
  OAI22_X1 U16556 ( .A1(n19427), .A2(n19560), .B1(n13434), .B2(n19463), .ZN(
        n13435) );
  AOI21_X1 U16557 ( .B1(n19486), .B2(n13436), .A(n13435), .ZN(n13438) );
  AOI22_X1 U16558 ( .A1(n19422), .A2(BUF2_REG_17__SCAN_IN), .B1(n19420), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13437) );
  OAI211_X1 U16559 ( .C1(n13439), .C2(n19458), .A(n13438), .B(n13437), .ZN(
        P2_U2902) );
  NAND2_X1 U16560 ( .A1(n13441), .A2(n13440), .ZN(n13442) );
  NAND2_X1 U16561 ( .A1(n13666), .A2(n13442), .ZN(n15744) );
  NAND2_X1 U16562 ( .A1(n13443), .A2(n15281), .ZN(n13445) );
  NAND2_X1 U16563 ( .A1(n15279), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13444) );
  OAI211_X1 U16564 ( .C1(n15744), .C2(n15279), .A(n13445), .B(n13444), .ZN(
        P2_U2870) );
  XNOR2_X1 U16565 ( .A(n13448), .B(n13447), .ZN(n16661) );
  INV_X1 U16566 ( .A(n16661), .ZN(n13461) );
  XOR2_X1 U16567 ( .A(n13450), .B(n13449), .Z(n16663) );
  NAND2_X1 U16568 ( .A1(n16663), .A2(n16673), .ZN(n13460) );
  OAI22_X1 U16569 ( .A1(n13451), .A2(n16702), .B1(n20157), .B2(n15727), .ZN(
        n13458) );
  OAI21_X1 U16570 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n13452), .ZN(n13453) );
  OAI22_X1 U16571 ( .A1(n13456), .A2(n13455), .B1(n13454), .B2(n13453), .ZN(
        n13457) );
  AOI211_X1 U16572 ( .C1(n16669), .C2(n19459), .A(n13458), .B(n13457), .ZN(
        n13459) );
  OAI211_X1 U16573 ( .C1(n13461), .C2(n16710), .A(n13460), .B(n13459), .ZN(
        P2_U3041) );
  XNOR2_X1 U16574 ( .A(n13462), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14883) );
  NAND2_X1 U16575 ( .A1(n14883), .A2(n12477), .ZN(n13479) );
  AOI22_X1 U16576 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11948), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U16577 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U16578 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13464) );
  AOI22_X1 U16579 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13463) );
  NAND4_X1 U16580 ( .A1(n13466), .A2(n13465), .A3(n13464), .A4(n13463), .ZN(
        n13472) );
  AOI22_X1 U16581 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U16582 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U16583 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U16584 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13467) );
  NAND4_X1 U16585 ( .A1(n13470), .A2(n13469), .A3(n13468), .A4(n13467), .ZN(
        n13471) );
  NOR2_X1 U16586 ( .A1(n13472), .A2(n13471), .ZN(n13475) );
  NAND2_X1 U16587 ( .A1(n14445), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U16588 ( .A1(n14444), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13473) );
  OAI211_X1 U16589 ( .C1(n13476), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13477) );
  INV_X1 U16590 ( .A(n13477), .ZN(n13478) );
  NAND2_X1 U16591 ( .A1(n13479), .A2(n13478), .ZN(n13480) );
  OAI21_X1 U16592 ( .B1(n9756), .B2(n13480), .A(n13750), .ZN(n14887) );
  INV_X1 U16593 ( .A(DATAI_10_), .ZN(n13482) );
  NAND2_X1 U16594 ( .A1(n14482), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13481) );
  OAI21_X1 U16595 ( .B1(n14482), .B2(n13482), .A(n13481), .ZN(n20423) );
  AOI22_X1 U16596 ( .A1(n13483), .A2(n20423), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n21063), .ZN(n13484) );
  OAI21_X1 U16597 ( .B1(n14887), .B2(n14717), .A(n13484), .ZN(P1_U2894) );
  INV_X1 U16598 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14602) );
  NAND2_X1 U16599 ( .A1(n14399), .A2(n14602), .ZN(n13487) );
  INV_X1 U16600 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14995) );
  NAND2_X1 U16601 ( .A1(n9988), .A2(n14602), .ZN(n13485) );
  OAI211_X1 U16602 ( .C1(n14419), .C2(n14995), .A(n13485), .B(n12753), .ZN(
        n13486) );
  NAND2_X1 U16603 ( .A1(n13487), .A2(n13486), .ZN(n13489) );
  AOI21_X1 U16604 ( .B1(n13489), .B2(n13488), .A(n9993), .ZN(n16461) );
  AOI22_X1 U16605 ( .A1(n16461), .A2(n16315), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14649), .ZN(n13490) );
  OAI21_X1 U16606 ( .B1(n14887), .B2(n14666), .A(n13490), .ZN(P1_U2862) );
  NOR3_X2 U16607 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20554), .A3(
        n20692), .ZN(n13532) );
  INV_X1 U16608 ( .A(n20757), .ZN(n13493) );
  OAI21_X1 U16609 ( .B1(n13493), .B2(n13492), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13495) );
  NOR2_X1 U16610 ( .A1(n20694), .A2(n20591), .ZN(n13499) );
  INV_X1 U16611 ( .A(n13499), .ZN(n13494) );
  AOI21_X1 U16612 ( .B1(n13495), .B2(n13494), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n13498) );
  OAI211_X1 U16613 ( .C1(n13532), .C2(n13498), .A(n20593), .B(n13497), .ZN(
        n13537) );
  NOR2_X1 U16614 ( .A1(n20757), .A2(n20668), .ZN(n13505) );
  NAND2_X1 U16615 ( .A1(n13499), .A2(n20658), .ZN(n13502) );
  NAND2_X1 U16616 ( .A1(n13675), .A2(n13500), .ZN(n13501) );
  NAND2_X1 U16617 ( .A1(n13502), .A2(n13501), .ZN(n13531) );
  AOI22_X1 U16618 ( .A1(n20719), .A2(n13532), .B1(n20718), .B2(n13531), .ZN(
        n13503) );
  OAI21_X1 U16619 ( .B1(n20723), .B2(n13534), .A(n13503), .ZN(n13504) );
  AOI211_X1 U16620 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n13505), .B(n13504), .ZN(n13506) );
  INV_X1 U16621 ( .A(n13506), .ZN(P1_U3147) );
  NOR2_X1 U16622 ( .A1(n20757), .A2(n20672), .ZN(n13509) );
  AOI22_X1 U16623 ( .A1(n20725), .A2(n13532), .B1(n20724), .B2(n13531), .ZN(
        n13507) );
  OAI21_X1 U16624 ( .B1(n20729), .B2(n13534), .A(n13507), .ZN(n13508) );
  AOI211_X1 U16625 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n13509), .B(n13508), .ZN(n13510) );
  INV_X1 U16626 ( .A(n13510), .ZN(P1_U3148) );
  NOR2_X1 U16627 ( .A1(n20757), .A2(n20636), .ZN(n13513) );
  AOI22_X1 U16628 ( .A1(n20731), .A2(n13532), .B1(n20730), .B2(n13531), .ZN(
        n13511) );
  OAI21_X1 U16629 ( .B1(n20735), .B2(n13534), .A(n13511), .ZN(n13512) );
  AOI211_X1 U16630 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n13513), .B(n13512), .ZN(n13514) );
  INV_X1 U16631 ( .A(n13514), .ZN(P1_U3149) );
  NOR2_X1 U16632 ( .A1(n20757), .A2(n20640), .ZN(n13517) );
  AOI22_X1 U16633 ( .A1(n20737), .A2(n13532), .B1(n20736), .B2(n13531), .ZN(
        n13515) );
  OAI21_X1 U16634 ( .B1(n20741), .B2(n13534), .A(n13515), .ZN(n13516) );
  AOI211_X1 U16635 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n13517), .B(n13516), .ZN(n13518) );
  INV_X1 U16636 ( .A(n13518), .ZN(P1_U3150) );
  NOR2_X1 U16637 ( .A1(n20757), .A2(n20664), .ZN(n13521) );
  AOI22_X1 U16638 ( .A1(n20713), .A2(n13532), .B1(n20712), .B2(n13531), .ZN(
        n13519) );
  OAI21_X1 U16639 ( .B1(n20717), .B2(n13534), .A(n13519), .ZN(n13520) );
  AOI211_X1 U16640 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n13521), .B(n13520), .ZN(n13522) );
  INV_X1 U16641 ( .A(n13522), .ZN(P1_U3146) );
  NOR2_X1 U16642 ( .A1(n20757), .A2(n20691), .ZN(n13525) );
  AOI22_X1 U16643 ( .A1(n20751), .A2(n13532), .B1(n20749), .B2(n13531), .ZN(
        n13523) );
  OAI21_X1 U16644 ( .B1(n20758), .B2(n13534), .A(n13523), .ZN(n13524) );
  AOI211_X1 U16645 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n13525), .B(n13524), .ZN(n13526) );
  INV_X1 U16646 ( .A(n13526), .ZN(P1_U3152) );
  NOR2_X1 U16647 ( .A1(n20757), .A2(n20626), .ZN(n13529) );
  AOI22_X1 U16648 ( .A1(n20701), .A2(n13532), .B1(n20700), .B2(n13531), .ZN(
        n13527) );
  OAI21_X1 U16649 ( .B1(n20711), .B2(n13534), .A(n13527), .ZN(n13528) );
  AOI211_X1 U16650 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n13529), .B(n13528), .ZN(n13530) );
  INV_X1 U16651 ( .A(n13530), .ZN(P1_U3145) );
  NOR2_X1 U16652 ( .A1(n20757), .A2(n20682), .ZN(n13536) );
  AOI22_X1 U16653 ( .A1(n20743), .A2(n13532), .B1(n20742), .B2(n13531), .ZN(
        n13533) );
  OAI21_X1 U16654 ( .B1(n20747), .B2(n13534), .A(n13533), .ZN(n13535) );
  AOI211_X1 U16655 ( .C1(n13537), .C2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n13536), .B(n13535), .ZN(n13538) );
  INV_X1 U16656 ( .A(n13538), .ZN(P1_U3151) );
  INV_X1 U16657 ( .A(n15009), .ZN(n13540) );
  NAND2_X1 U16658 ( .A1(n13540), .A2(n13539), .ZN(n15034) );
  NAND2_X1 U16659 ( .A1(n13543), .A2(n13572), .ZN(n13541) );
  AOI21_X1 U16660 ( .B1(n13541), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20703), 
        .ZN(n13547) );
  NOR2_X1 U16661 ( .A1(n20694), .A2(n20521), .ZN(n13544) );
  AND2_X1 U16662 ( .A1(n13542), .A2(n20524), .ZN(n15041) );
  INV_X1 U16663 ( .A(n13544), .ZN(n13546) );
  NOR2_X1 U16664 ( .A1(n15041), .A2(n20697), .ZN(n13545) );
  AOI21_X1 U16665 ( .B1(n13547), .B2(n13546), .A(n13545), .ZN(n13548) );
  OAI211_X1 U16666 ( .C1(n10248), .C2(n16512), .A(n20593), .B(n13548), .ZN(
        n13570) );
  AOI22_X1 U16667 ( .A1(n20701), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n13570), .ZN(n13549) );
  OAI21_X1 U16668 ( .B1(n13572), .B2(n20711), .A(n13549), .ZN(n13550) );
  AOI21_X1 U16669 ( .B1(n13574), .B2(n20708), .A(n13550), .ZN(n13551) );
  OAI21_X1 U16670 ( .B1(n13576), .B2(n13686), .A(n13551), .ZN(P1_U3129) );
  AOI22_X1 U16671 ( .A1(n20713), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n13570), .ZN(n13552) );
  OAI21_X1 U16672 ( .B1(n13572), .B2(n20717), .A(n13552), .ZN(n13553) );
  AOI21_X1 U16673 ( .B1(n13574), .B2(n20714), .A(n13553), .ZN(n13554) );
  OAI21_X1 U16674 ( .B1(n13576), .B2(n13690), .A(n13554), .ZN(P1_U3130) );
  AOI22_X1 U16675 ( .A1(n20725), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n13570), .ZN(n13555) );
  OAI21_X1 U16676 ( .B1(n13572), .B2(n20729), .A(n13555), .ZN(n13556) );
  AOI21_X1 U16677 ( .B1(n13574), .B2(n20726), .A(n13556), .ZN(n13557) );
  OAI21_X1 U16678 ( .B1(n13576), .B2(n13694), .A(n13557), .ZN(P1_U3132) );
  AOI22_X1 U16679 ( .A1(n20719), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n13570), .ZN(n13558) );
  OAI21_X1 U16680 ( .B1(n13572), .B2(n20723), .A(n13558), .ZN(n13559) );
  AOI21_X1 U16681 ( .B1(n13574), .B2(n20720), .A(n13559), .ZN(n13560) );
  OAI21_X1 U16682 ( .B1(n13576), .B2(n13706), .A(n13560), .ZN(P1_U3131) );
  AOI22_X1 U16683 ( .A1(n20751), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n13570), .ZN(n13561) );
  OAI21_X1 U16684 ( .B1(n13572), .B2(n20758), .A(n13561), .ZN(n13562) );
  AOI21_X1 U16685 ( .B1(n13574), .B2(n20752), .A(n13562), .ZN(n13563) );
  OAI21_X1 U16686 ( .B1(n13576), .B2(n13702), .A(n13563), .ZN(P1_U3136) );
  AOI22_X1 U16687 ( .A1(n20743), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n13570), .ZN(n13564) );
  OAI21_X1 U16688 ( .B1(n13572), .B2(n20747), .A(n13564), .ZN(n13565) );
  AOI21_X1 U16689 ( .B1(n13574), .B2(n20744), .A(n13565), .ZN(n13566) );
  OAI21_X1 U16690 ( .B1(n13576), .B2(n13698), .A(n13566), .ZN(P1_U3135) );
  AOI22_X1 U16691 ( .A1(n20737), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n13570), .ZN(n13567) );
  OAI21_X1 U16692 ( .B1(n13572), .B2(n20741), .A(n13567), .ZN(n13568) );
  AOI21_X1 U16693 ( .B1(n13574), .B2(n20738), .A(n13568), .ZN(n13569) );
  OAI21_X1 U16694 ( .B1(n13576), .B2(n13710), .A(n13569), .ZN(P1_U3134) );
  AOI22_X1 U16695 ( .A1(n20731), .A2(n10248), .B1(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n13570), .ZN(n13571) );
  OAI21_X1 U16696 ( .B1(n13572), .B2(n20735), .A(n13571), .ZN(n13573) );
  AOI21_X1 U16697 ( .B1(n13574), .B2(n20732), .A(n13573), .ZN(n13575) );
  OAI21_X1 U16698 ( .B1(n13576), .B2(n13717), .A(n13575), .ZN(P1_U3133) );
  AOI21_X1 U16699 ( .B1(n13578), .B2(n13577), .A(n15295), .ZN(n13579) );
  INV_X1 U16700 ( .A(n13579), .ZN(n13669) );
  NAND2_X1 U16701 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  NAND2_X1 U16702 ( .A1(n15146), .A2(n13582), .ZN(n19315) );
  INV_X1 U16703 ( .A(n19315), .ZN(n13585) );
  OAI22_X1 U16704 ( .A1(n19427), .A2(n19565), .B1(n13583), .B2(n19463), .ZN(
        n13584) );
  AOI21_X1 U16705 ( .B1(n13585), .B2(n19486), .A(n13584), .ZN(n13587) );
  AOI22_X1 U16706 ( .A1(n19422), .A2(BUF2_REG_18__SCAN_IN), .B1(n19420), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n13586) );
  OAI211_X1 U16707 ( .C1(n13669), .C2(n19458), .A(n13587), .B(n13586), .ZN(
        P2_U2901) );
  NAND2_X1 U16708 ( .A1(n13589), .A2(n13588), .ZN(n13591) );
  NAND2_X1 U16709 ( .A1(n13591), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13590) );
  OAI21_X1 U16710 ( .B1(n13591), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13590), .ZN(n13609) );
  XOR2_X1 U16711 ( .A(n13592), .B(n13593), .Z(n13607) );
  INV_X1 U16712 ( .A(n15847), .ZN(n13601) );
  NOR2_X1 U16713 ( .A1(n13595), .A2(n13594), .ZN(n13596) );
  OR2_X1 U16714 ( .A1(n13597), .A2(n13596), .ZN(n19453) );
  NOR2_X1 U16715 ( .A1(n19453), .A2(n16701), .ZN(n13599) );
  INV_X1 U16716 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20159) );
  OAI22_X1 U16717 ( .A1(n13604), .A2(n16702), .B1(n20159), .B2(n15727), .ZN(
        n13598) );
  AOI211_X1 U16718 ( .C1(n15845), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13599), .B(n13598), .ZN(n13600) );
  OAI21_X1 U16719 ( .B1(n13601), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13600), .ZN(n13602) );
  AOI21_X1 U16720 ( .B1(n13607), .B2(n16673), .A(n13602), .ZN(n13603) );
  OAI21_X1 U16721 ( .B1(n13609), .B2(n16710), .A(n13603), .ZN(P2_U3040) );
  OAI22_X1 U16722 ( .A1(n10046), .A2(n16666), .B1(n19542), .B2(n19368), .ZN(
        n13606) );
  OAI22_X1 U16723 ( .A1(n13604), .A2(n16648), .B1(n15727), .B2(n20159), .ZN(
        n13605) );
  AOI211_X1 U16724 ( .C1(n13607), .C2(n16662), .A(n13606), .B(n13605), .ZN(
        n13608) );
  OAI21_X1 U16725 ( .B1(n19532), .B2(n13609), .A(n13608), .ZN(P2_U3008) );
  NAND2_X1 U16726 ( .A1(n13610), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13611) );
  OR2_X1 U16727 ( .A1(n13613), .A2(n13651), .ZN(n13617) );
  NAND2_X1 U16728 ( .A1(n13625), .A2(n13623), .ZN(n13614) );
  XNOR2_X1 U16729 ( .A(n13614), .B(n13622), .ZN(n13615) );
  NAND2_X1 U16730 ( .A1(n13615), .A2(n13657), .ZN(n13616) );
  XNOR2_X1 U16731 ( .A(n13619), .B(n13618), .ZN(n20452) );
  NAND2_X1 U16732 ( .A1(n13619), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13620) );
  OR2_X1 U16733 ( .A1(n13621), .A2(n13651), .ZN(n13628) );
  AND2_X1 U16734 ( .A1(n13623), .A2(n13622), .ZN(n13624) );
  NAND2_X1 U16735 ( .A1(n13625), .A2(n13624), .ZN(n13643) );
  XNOR2_X1 U16736 ( .A(n13643), .B(n13640), .ZN(n13626) );
  NAND2_X1 U16737 ( .A1(n13626), .A2(n13657), .ZN(n13627) );
  NAND2_X1 U16738 ( .A1(n13628), .A2(n13627), .ZN(n13629) );
  NAND2_X1 U16739 ( .A1(n13629), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13630) );
  NAND3_X1 U16740 ( .A1(n13654), .A2(n13647), .A3(n13631), .ZN(n13636) );
  INV_X1 U16741 ( .A(n13643), .ZN(n13632) );
  NAND2_X1 U16742 ( .A1(n13632), .A2(n13640), .ZN(n13633) );
  XNOR2_X1 U16743 ( .A(n13633), .B(n13641), .ZN(n13634) );
  NAND2_X1 U16744 ( .A1(n13634), .A2(n13657), .ZN(n13635) );
  NAND2_X1 U16745 ( .A1(n16379), .A2(n20999), .ZN(n13637) );
  INV_X1 U16746 ( .A(n16379), .ZN(n13638) );
  NAND2_X1 U16747 ( .A1(n13638), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13639) );
  NAND2_X1 U16748 ( .A1(n13641), .A2(n13640), .ZN(n13642) );
  OR2_X1 U16749 ( .A1(n13643), .A2(n13642), .ZN(n13655) );
  XNOR2_X1 U16750 ( .A(n13655), .B(n13644), .ZN(n13645) );
  NOR2_X1 U16751 ( .A1(n13645), .A2(n20860), .ZN(n13646) );
  AOI21_X1 U16752 ( .B1(n13648), .B2(n13647), .A(n13646), .ZN(n13649) );
  NAND2_X1 U16753 ( .A1(n13649), .A2(n16469), .ZN(n16374) );
  INV_X1 U16754 ( .A(n13649), .ZN(n13650) );
  NAND2_X1 U16755 ( .A1(n13650), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16373) );
  NOR2_X1 U16756 ( .A1(n13652), .A2(n13651), .ZN(n13653) );
  INV_X1 U16757 ( .A(n13655), .ZN(n13658) );
  NAND3_X1 U16758 ( .A1(n13658), .A2(n13657), .A3(n13656), .ZN(n13659) );
  XNOR2_X1 U16759 ( .A(n13720), .B(n16468), .ZN(n13660) );
  XNOR2_X1 U16760 ( .A(n13719), .B(n13660), .ZN(n16477) );
  NAND2_X1 U16761 ( .A1(n16477), .A2(n20457), .ZN(n13664) );
  AND2_X1 U16762 ( .A1(n16482), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n16470) );
  NOR2_X1 U16763 ( .A1(n20461), .A2(n13661), .ZN(n13662) );
  AOI211_X1 U16764 ( .C1(n20450), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16470), .B(n13662), .ZN(n13663) );
  OAI211_X1 U16765 ( .C1(n14888), .C2(n13665), .A(n13664), .B(n13663), .ZN(
        P1_U2991) );
  AOI21_X1 U16766 ( .B1(n13667), .B2(n13666), .A(n15151), .ZN(n19311) );
  INV_X1 U16767 ( .A(n19311), .ZN(n15732) );
  MUX2_X1 U16768 ( .A(n10945), .B(n15732), .S(n15291), .Z(n13668) );
  OAI21_X1 U16769 ( .B1(n13669), .B2(n15298), .A(n13668), .ZN(P2_U2869) );
  INV_X1 U16770 ( .A(n13670), .ZN(n13671) );
  INV_X1 U16771 ( .A(n20645), .ZN(n13672) );
  AOI21_X1 U16772 ( .B1(n13672), .B2(n13714), .A(n20702), .ZN(n13673) );
  NOR2_X1 U16773 ( .A1(n13673), .A2(n20703), .ZN(n13681) );
  AND2_X1 U16774 ( .A1(n20616), .A2(n20521), .ZN(n13678) );
  INV_X1 U16775 ( .A(n13676), .ZN(n13677) );
  NOR2_X1 U16776 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13677), .ZN(
        n13712) );
  INV_X1 U16777 ( .A(n13678), .ZN(n13680) );
  AOI21_X1 U16778 ( .B1(n13681), .B2(n13680), .A(n13679), .ZN(n13682) );
  OAI211_X1 U16779 ( .C1(n13712), .C2(n16512), .A(n20593), .B(n13682), .ZN(
        n13711) );
  AOI22_X1 U16780 ( .A1(n20701), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n13711), .ZN(n13683) );
  OAI21_X1 U16781 ( .B1(n13714), .B2(n20711), .A(n13683), .ZN(n13684) );
  AOI21_X1 U16782 ( .B1(n20645), .B2(n20708), .A(n13684), .ZN(n13685) );
  OAI21_X1 U16783 ( .B1(n13718), .B2(n13686), .A(n13685), .ZN(P1_U3081) );
  AOI22_X1 U16784 ( .A1(n20713), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n13711), .ZN(n13687) );
  OAI21_X1 U16785 ( .B1(n13714), .B2(n20717), .A(n13687), .ZN(n13688) );
  AOI21_X1 U16786 ( .B1(n20645), .B2(n20714), .A(n13688), .ZN(n13689) );
  OAI21_X1 U16787 ( .B1(n13718), .B2(n13690), .A(n13689), .ZN(P1_U3082) );
  AOI22_X1 U16788 ( .A1(n20725), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n13711), .ZN(n13691) );
  OAI21_X1 U16789 ( .B1(n13714), .B2(n20729), .A(n13691), .ZN(n13692) );
  AOI21_X1 U16790 ( .B1(n20645), .B2(n20726), .A(n13692), .ZN(n13693) );
  OAI21_X1 U16791 ( .B1(n13718), .B2(n13694), .A(n13693), .ZN(P1_U3084) );
  AOI22_X1 U16792 ( .A1(n20743), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n13711), .ZN(n13695) );
  OAI21_X1 U16793 ( .B1(n13714), .B2(n20747), .A(n13695), .ZN(n13696) );
  AOI21_X1 U16794 ( .B1(n20645), .B2(n20744), .A(n13696), .ZN(n13697) );
  OAI21_X1 U16795 ( .B1(n13718), .B2(n13698), .A(n13697), .ZN(P1_U3087) );
  AOI22_X1 U16796 ( .A1(n20751), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n13711), .ZN(n13699) );
  OAI21_X1 U16797 ( .B1(n13714), .B2(n20758), .A(n13699), .ZN(n13700) );
  AOI21_X1 U16798 ( .B1(n20645), .B2(n20752), .A(n13700), .ZN(n13701) );
  OAI21_X1 U16799 ( .B1(n13718), .B2(n13702), .A(n13701), .ZN(P1_U3088) );
  AOI22_X1 U16800 ( .A1(n20719), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n13711), .ZN(n13703) );
  OAI21_X1 U16801 ( .B1(n13714), .B2(n20723), .A(n13703), .ZN(n13704) );
  AOI21_X1 U16802 ( .B1(n20645), .B2(n20720), .A(n13704), .ZN(n13705) );
  OAI21_X1 U16803 ( .B1(n13718), .B2(n13706), .A(n13705), .ZN(P1_U3083) );
  AOI22_X1 U16804 ( .A1(n20737), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n13711), .ZN(n13707) );
  OAI21_X1 U16805 ( .B1(n13714), .B2(n20741), .A(n13707), .ZN(n13708) );
  AOI21_X1 U16806 ( .B1(n20645), .B2(n20738), .A(n13708), .ZN(n13709) );
  OAI21_X1 U16807 ( .B1(n13718), .B2(n13710), .A(n13709), .ZN(P1_U3086) );
  AOI22_X1 U16808 ( .A1(n20731), .A2(n13712), .B1(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n13711), .ZN(n13713) );
  OAI21_X1 U16809 ( .B1(n13714), .B2(n20735), .A(n13713), .ZN(n13715) );
  AOI21_X1 U16810 ( .B1(n20645), .B2(n20732), .A(n13715), .ZN(n13716) );
  OAI21_X1 U16811 ( .B1(n13718), .B2(n13717), .A(n13716), .ZN(P1_U3085) );
  INV_X1 U16812 ( .A(n13720), .ZN(n13721) );
  NAND2_X1 U16813 ( .A1(n13721), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13722) );
  XNOR2_X1 U16814 ( .A(n14877), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13724) );
  XNOR2_X1 U16815 ( .A(n14424), .B(n13724), .ZN(n13738) );
  NOR3_X1 U16816 ( .A1(n16468), .A2(n16469), .A3(n20999), .ZN(n14890) );
  NAND2_X1 U16817 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20462) );
  NOR2_X1 U16818 ( .A1(n13725), .A2(n20462), .ZN(n13726) );
  OAI21_X1 U16819 ( .B1(n9985), .B2(n20500), .A(n20870), .ZN(n20497) );
  NAND2_X1 U16820 ( .A1(n13726), .A2(n20497), .ZN(n14985) );
  INV_X1 U16821 ( .A(n13726), .ZN(n13730) );
  NAND2_X1 U16822 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20465) );
  NOR2_X1 U16823 ( .A1(n13730), .A2(n20465), .ZN(n14986) );
  INV_X1 U16824 ( .A(n14986), .ZN(n15000) );
  OAI21_X1 U16825 ( .B1(n20483), .B2(n14985), .A(n15000), .ZN(n13728) );
  OAI21_X1 U16826 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13727), .A(
        n20506), .ZN(n16443) );
  INV_X1 U16827 ( .A(n16443), .ZN(n20487) );
  OAI221_X1 U16828 ( .B1(n16476), .B2(n14890), .C1(n16476), .C2(n13728), .A(
        n20487), .ZN(n16463) );
  NAND2_X1 U16829 ( .A1(n16482), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n13734) );
  OAI21_X1 U16830 ( .B1(n20317), .B2(n20503), .A(n13734), .ZN(n13732) );
  NAND2_X1 U16831 ( .A1(n14890), .A2(n16491), .ZN(n16467) );
  NOR2_X1 U16832 ( .A1(n16467), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13731) );
  AOI211_X1 U16833 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16463), .A(
        n13732), .B(n13731), .ZN(n13733) );
  OAI21_X1 U16834 ( .B1(n13738), .B2(n16457), .A(n13733), .ZN(P1_U3022) );
  OAI21_X1 U16835 ( .B1(n16333), .B2(n20315), .A(n13734), .ZN(n13736) );
  NOR2_X1 U16836 ( .A1(n20320), .A2(n14888), .ZN(n13735) );
  AOI211_X1 U16837 ( .C1(n16365), .C2(n20321), .A(n13736), .B(n13735), .ZN(
        n13737) );
  OAI21_X1 U16838 ( .B1(n13738), .B2(n20299), .A(n13737), .ZN(P1_U2990) );
  AOI22_X1 U16839 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U16840 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U16841 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13740) );
  AOI22_X1 U16842 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13739) );
  NAND4_X1 U16843 ( .A1(n13742), .A2(n13741), .A3(n13740), .A4(n13739), .ZN(
        n13748) );
  AOI22_X1 U16844 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13746) );
  AOI22_X1 U16845 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13745) );
  AOI22_X1 U16846 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13744) );
  AOI22_X1 U16847 ( .A1(n14356), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13743) );
  NAND4_X1 U16848 ( .A1(n13746), .A2(n13745), .A3(n13744), .A4(n13743), .ZN(
        n13747) );
  OR2_X1 U16849 ( .A1(n13748), .A2(n13747), .ZN(n13749) );
  NAND2_X1 U16850 ( .A1(n13859), .A2(n13749), .ZN(n13832) );
  INV_X1 U16851 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13841) );
  OAI21_X1 U16852 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13751), .A(
        n13779), .ZN(n16372) );
  AOI22_X1 U16853 ( .A1(n14345), .A2(n16372), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13752) );
  OAI21_X1 U16854 ( .B1(n14285), .B2(n13841), .A(n13752), .ZN(n13753) );
  INV_X1 U16855 ( .A(n13753), .ZN(n13818) );
  XNOR2_X1 U16856 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n13754), .ZN(
        n14872) );
  INV_X1 U16857 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13845) );
  INV_X1 U16858 ( .A(n14444), .ZN(n14111) );
  OAI22_X1 U16859 ( .A1(n14285), .A2(n13845), .B1(n14111), .B2(n14590), .ZN(
        n13755) );
  INV_X1 U16860 ( .A(n13755), .ZN(n13767) );
  AOI22_X1 U16861 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14293), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13759) );
  AOI22_X1 U16862 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U16863 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13757) );
  AOI22_X1 U16864 ( .A1(n14357), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13756) );
  NAND4_X1 U16865 ( .A1(n13759), .A2(n13758), .A3(n13757), .A4(n13756), .ZN(
        n13765) );
  AOI22_X1 U16866 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U16867 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14219), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13762) );
  AOI22_X1 U16868 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U16869 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13760) );
  NAND4_X1 U16870 ( .A1(n13763), .A2(n13762), .A3(n13761), .A4(n13760), .ZN(
        n13764) );
  OAI21_X1 U16871 ( .B1(n13765), .B2(n13764), .A(n13859), .ZN(n13766) );
  OAI211_X1 U16872 ( .C1(n14872), .C2(n14351), .A(n13767), .B(n13766), .ZN(
        n13824) );
  INV_X1 U16873 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U16874 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12199), .B1(
        n9681), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U16875 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14358), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U16876 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11948), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U16877 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13768) );
  NAND4_X1 U16878 ( .A1(n13771), .A2(n13770), .A3(n13769), .A4(n13768), .ZN(
        n13777) );
  AOI22_X1 U16879 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13775) );
  AOI22_X1 U16880 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13774) );
  AOI22_X1 U16881 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U16882 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13772) );
  NAND4_X1 U16883 ( .A1(n13775), .A2(n13774), .A3(n13773), .A4(n13772), .ZN(
        n13776) );
  OR2_X1 U16884 ( .A1(n13777), .A2(n13776), .ZN(n13778) );
  NAND2_X1 U16885 ( .A1(n13859), .A2(n13778), .ZN(n13782) );
  XNOR2_X1 U16886 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13779), .ZN(
        n16364) );
  INV_X1 U16887 ( .A(n16364), .ZN(n13780) );
  AOI22_X1 U16888 ( .A1(n14444), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n14345), .B2(n13780), .ZN(n13781) );
  OAI211_X1 U16889 ( .C1(n14285), .C2(n14746), .A(n13782), .B(n13781), .ZN(
        n14739) );
  NAND2_X1 U16890 ( .A1(n13824), .A2(n14739), .ZN(n13783) );
  XNOR2_X1 U16891 ( .A(n13784), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14860) );
  NAND2_X1 U16892 ( .A1(n14860), .A2(n12477), .ZN(n13799) );
  INV_X1 U16893 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13805) );
  INV_X1 U16894 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14584) );
  OAI22_X1 U16895 ( .A1(n14285), .A2(n13805), .B1(n14111), .B2(n14584), .ZN(
        n13785) );
  INV_X1 U16896 ( .A(n13785), .ZN(n13797) );
  AOI22_X1 U16897 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U16898 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U16899 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U16900 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13786) );
  NAND4_X1 U16901 ( .A1(n13789), .A2(n13788), .A3(n13787), .A4(n13786), .ZN(
        n13795) );
  AOI22_X1 U16902 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13793) );
  AOI22_X1 U16903 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13792) );
  AOI22_X1 U16904 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13791) );
  AOI22_X1 U16905 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13790) );
  NAND4_X1 U16906 ( .A1(n13793), .A2(n13792), .A3(n13791), .A4(n13790), .ZN(
        n13794) );
  OAI21_X1 U16907 ( .B1(n13795), .B2(n13794), .A(n13859), .ZN(n13796) );
  AND2_X1 U16908 ( .A1(n13797), .A2(n13796), .ZN(n13798) );
  NAND2_X1 U16909 ( .A1(n13799), .A2(n13798), .ZN(n13800) );
  NOR2_X1 U16910 ( .A1(n13822), .A2(n13800), .ZN(n13801) );
  OR2_X1 U16911 ( .A1(n13862), .A2(n13801), .ZN(n14864) );
  INV_X1 U16912 ( .A(DATAI_14_), .ZN(n13803) );
  NAND2_X1 U16913 ( .A1(n14482), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13802) );
  OAI21_X1 U16914 ( .B1(n14482), .B2(n13803), .A(n13802), .ZN(n20431) );
  INV_X1 U16915 ( .A(n20431), .ZN(n13804) );
  OAI222_X1 U16916 ( .A1(n14864), .A2(n14717), .B1(n13805), .B2(n14745), .C1(
        n14744), .C2(n13804), .ZN(P1_U2890) );
  INV_X1 U16917 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16305) );
  NAND2_X1 U16918 ( .A1(n14412), .A2(n16305), .ZN(n13809) );
  INV_X1 U16919 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U16920 ( .A1(n12753), .A2(n13806), .ZN(n13807) );
  OAI211_X1 U16921 ( .C1(n14456), .C2(P1_EBX_REG_11__SCAN_IN), .A(n13807), .B(
        n14454), .ZN(n13808) );
  INV_X1 U16922 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16317) );
  NAND2_X1 U16923 ( .A1(n14399), .A2(n16317), .ZN(n13812) );
  INV_X1 U16924 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16453) );
  NAND2_X1 U16925 ( .A1(n9988), .A2(n16317), .ZN(n13810) );
  OAI211_X1 U16926 ( .C1(n14419), .C2(n16453), .A(n13810), .B(n12753), .ZN(
        n13811) );
  NAND2_X1 U16927 ( .A1(n13812), .A2(n13811), .ZN(n16297) );
  INV_X1 U16928 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16448) );
  NAND2_X1 U16929 ( .A1(n12753), .A2(n16448), .ZN(n13813) );
  OAI211_X1 U16930 ( .C1(n14456), .C2(P1_EBX_REG_13__SCAN_IN), .A(n13813), .B(
        n14454), .ZN(n13814) );
  OAI21_X1 U16931 ( .B1(n14410), .B2(P1_EBX_REG_13__SCAN_IN), .A(n13814), .ZN(
        n13825) );
  MUX2_X1 U16932 ( .A(n14417), .B(n14454), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13815) );
  OAI21_X1 U16933 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14457), .A(
        n13815), .ZN(n13816) );
  NAND2_X1 U16934 ( .A1(n13826), .A2(n13816), .ZN(n13817) );
  NAND2_X1 U16935 ( .A1(n13869), .A2(n13817), .ZN(n16430) );
  INV_X1 U16936 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14581) );
  OAI222_X1 U16937 ( .A1(n16430), .A2(n20385), .B1(n14581), .B2(n20390), .C1(
        n14864), .C2(n14666), .ZN(P1_U2858) );
  NAND2_X1 U16938 ( .A1(n13750), .A2(n13818), .ZN(n13819) );
  NAND2_X1 U16939 ( .A1(n13820), .A2(n13819), .ZN(n13831) );
  OR2_X1 U16940 ( .A1(n13831), .A2(n13832), .ZN(n13821) );
  NAND2_X1 U16941 ( .A1(n13821), .A2(n13820), .ZN(n14738) );
  INV_X1 U16942 ( .A(n13822), .ZN(n13823) );
  OR2_X1 U16943 ( .A1(n16295), .A2(n13825), .ZN(n13827) );
  AND2_X1 U16944 ( .A1(n13827), .A2(n13826), .ZN(n16445) );
  INV_X1 U16945 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13828) );
  NOR2_X1 U16946 ( .A1(n20390), .A2(n13828), .ZN(n13829) );
  AOI21_X1 U16947 ( .B1(n16445), .B2(n16315), .A(n13829), .ZN(n13830) );
  OAI21_X1 U16948 ( .B1(n14875), .B2(n14666), .A(n13830), .ZN(P1_U2859) );
  XOR2_X1 U16949 ( .A(n13832), .B(n13831), .Z(n16368) );
  NAND2_X1 U16950 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  NAND2_X1 U16951 ( .A1(n16296), .A2(n13835), .ZN(n16306) );
  OAI22_X1 U16952 ( .A1(n16306), .A2(n20385), .B1(n16305), .B2(n20390), .ZN(
        n13836) );
  AOI21_X1 U16953 ( .B1(n16368), .B2(n20387), .A(n13836), .ZN(n13837) );
  INV_X1 U16954 ( .A(n13837), .ZN(P1_U2861) );
  INV_X1 U16955 ( .A(n16368), .ZN(n13842) );
  INV_X1 U16956 ( .A(DATAI_11_), .ZN(n13839) );
  NAND2_X1 U16957 ( .A1(n14482), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13838) );
  OAI21_X1 U16958 ( .B1(n14482), .B2(n13839), .A(n13838), .ZN(n20425) );
  INV_X1 U16959 ( .A(n20425), .ZN(n13840) );
  OAI222_X1 U16960 ( .A1(n13842), .A2(n14717), .B1(n13841), .B2(n14745), .C1(
        n14744), .C2(n13840), .ZN(P1_U2893) );
  INV_X1 U16961 ( .A(DATAI_13_), .ZN(n13844) );
  NAND2_X1 U16962 ( .A1(n14482), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13843) );
  OAI21_X1 U16963 ( .B1(n14482), .B2(n13844), .A(n13843), .ZN(n20429) );
  INV_X1 U16964 ( .A(n20429), .ZN(n13846) );
  OAI222_X1 U16965 ( .A1(n14717), .A2(n14875), .B1(n14744), .B2(n13846), .C1(
        n13845), .C2(n14745), .ZN(P1_U2891) );
  XOR2_X1 U16966 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n13847), .Z(
        n16356) );
  AOI22_X1 U16967 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13851) );
  AOI22_X1 U16968 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U16969 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13849) );
  AOI22_X1 U16970 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13848) );
  NAND4_X1 U16971 ( .A1(n13851), .A2(n13850), .A3(n13849), .A4(n13848), .ZN(
        n13857) );
  AOI22_X1 U16972 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13337), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U16973 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U16974 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U16975 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13852) );
  NAND4_X1 U16976 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13856) );
  OR2_X1 U16977 ( .A1(n13857), .A2(n13856), .ZN(n13858) );
  AOI22_X1 U16978 ( .A1(n13859), .A2(n13858), .B1(n14444), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13861) );
  NAND2_X1 U16979 ( .A1(n14445), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13860) );
  OAI211_X1 U16980 ( .C1(n16356), .C2(n14351), .A(n13861), .B(n13860), .ZN(
        n13863) );
  OR2_X1 U16981 ( .A1(n13862), .A2(n13863), .ZN(n13864) );
  AND2_X1 U16982 ( .A1(n14099), .A2(n13864), .ZN(n16357) );
  INV_X1 U16983 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n13872) );
  NAND2_X1 U16984 ( .A1(n14412), .A2(n13872), .ZN(n13867) );
  INV_X1 U16985 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U16986 ( .A1(n12753), .A2(n14431), .ZN(n13865) );
  OAI211_X1 U16987 ( .C1(n14456), .C2(P1_EBX_REG_15__SCAN_IN), .A(n13865), .B(
        n14454), .ZN(n13866) );
  INV_X1 U16988 ( .A(n14567), .ZN(n13871) );
  NAND2_X1 U16989 ( .A1(n13869), .A2(n13868), .ZN(n13870) );
  NAND2_X1 U16990 ( .A1(n13871), .A2(n13870), .ZN(n16424) );
  OAI22_X1 U16991 ( .A1(n16424), .A2(n20385), .B1(n13872), .B2(n20390), .ZN(
        n13873) );
  AOI21_X1 U16992 ( .B1(n16357), .B2(n20387), .A(n13873), .ZN(n13874) );
  INV_X1 U16993 ( .A(n13874), .ZN(P1_U2857) );
  AOI22_X1 U16994 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U16995 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13877) );
  INV_X2 U16996 ( .A(n13957), .ZN(n17583) );
  AOI22_X1 U16997 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U16998 ( .A1(n16041), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13875) );
  NAND4_X1 U16999 ( .A1(n13878), .A2(n13877), .A3(n13876), .A4(n13875), .ZN(
        n13890) );
  NOR2_X2 U17000 ( .A1(n13879), .A2(n13881), .ZN(n17405) );
  AOI22_X1 U17001 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13888) );
  INV_X2 U17002 ( .A(n9714), .ZN(n17572) );
  AOI22_X1 U17003 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13887) );
  NOR2_X2 U17004 ( .A1(n13882), .A2(n19061), .ZN(n13986) );
  AOI22_X1 U17005 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17581), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13886) );
  NOR2_X2 U17006 ( .A1(n13882), .A2(n13881), .ZN(n13949) );
  AOI22_X1 U17007 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13885) );
  NAND4_X1 U17008 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13889) );
  AOI22_X1 U17009 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17010 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17011 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17012 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17554), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13892) );
  NAND4_X1 U17013 ( .A1(n13895), .A2(n13894), .A3(n13893), .A4(n13892), .ZN(
        n13902) );
  AOI22_X1 U17014 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17015 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13899) );
  INV_X1 U17016 ( .A(n13896), .ZN(n17538) );
  AOI22_X1 U17017 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13898) );
  INV_X2 U17018 ( .A(n17458), .ZN(n17574) );
  AOI22_X1 U17019 ( .A1(n17584), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13897) );
  NAND4_X1 U17020 ( .A1(n13900), .A2(n13899), .A3(n13898), .A4(n13897), .ZN(
        n13901) );
  AOI22_X1 U17021 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9667), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U17022 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17581), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13905) );
  AOI22_X1 U17023 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17024 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13903) );
  NAND4_X1 U17025 ( .A1(n13906), .A2(n13905), .A3(n13904), .A4(n13903), .ZN(
        n13912) );
  AOI22_X1 U17026 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n17573), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13910) );
  INV_X2 U17027 ( .A(n10251), .ZN(n17582) );
  AOI22_X1 U17028 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17029 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13908) );
  BUF_X2 U17030 ( .A(n13950), .Z(n16009) );
  AOI22_X1 U17031 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13907) );
  NAND4_X1 U17032 ( .A1(n13910), .A2(n13909), .A3(n13908), .A4(n13907), .ZN(
        n13911) );
  AOI22_X1 U17033 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13923) );
  AOI22_X1 U17034 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U17035 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13913) );
  OAI21_X1 U17036 ( .B1(n13962), .B2(n17618), .A(n13913), .ZN(n13920) );
  AOI22_X1 U17037 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17038 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U17039 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U17040 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13915) );
  NAND4_X1 U17041 ( .A1(n13918), .A2(n13917), .A3(n13916), .A4(n13915), .ZN(
        n13919) );
  AOI22_X1 U17042 ( .A1(n9676), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U17043 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13932) );
  INV_X1 U17044 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n20895) );
  AOI22_X1 U17045 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U17046 ( .B1(n20895), .B2(n14037), .A(n13924), .ZN(n13930) );
  AOI22_X1 U17047 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U17048 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U17049 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13926) );
  INV_X2 U17050 ( .A(n16040), .ZN(n17573) );
  AOI22_X1 U17051 ( .A1(n17405), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13925) );
  NAND4_X1 U17052 ( .A1(n13928), .A2(n13927), .A3(n13926), .A4(n13925), .ZN(
        n13929) );
  AOI22_X1 U17053 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U17054 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17055 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U17056 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n17572), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13934) );
  NAND4_X1 U17057 ( .A1(n13937), .A2(n13936), .A3(n13935), .A4(n13934), .ZN(
        n13943) );
  AOI22_X1 U17058 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13941) );
  AOI22_X1 U17059 ( .A1(n17584), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U17060 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17061 ( .A1(n17405), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13938) );
  NAND4_X1 U17062 ( .A1(n13941), .A2(n13940), .A3(n13939), .A4(n13938), .ZN(
        n13942) );
  NAND2_X1 U17063 ( .A1(n16102), .A2(n18629), .ZN(n15937) );
  INV_X1 U17064 ( .A(n15937), .ZN(n13944) );
  NAND2_X1 U17065 ( .A1(n19052), .A2(n13944), .ZN(n15954) );
  AOI22_X1 U17066 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U17067 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U17068 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13946) );
  AOI22_X1 U17069 ( .A1(n9676), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13945) );
  NAND4_X1 U17070 ( .A1(n13948), .A2(n13947), .A3(n13946), .A4(n13945), .ZN(
        n13956) );
  AOI22_X1 U17071 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n17580), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17072 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17556), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U17073 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17074 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13951) );
  NAND4_X1 U17075 ( .A1(n13954), .A2(n13953), .A3(n13952), .A4(n13951), .ZN(
        n13955) );
  INV_X2 U17076 ( .A(n13957), .ZN(n17555) );
  AOI22_X1 U17077 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U17078 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9667), .B1(n9679), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13960) );
  AOI22_X1 U17079 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13959) );
  AOI22_X1 U17080 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17581), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13958) );
  NAND4_X1 U17081 ( .A1(n13961), .A2(n13960), .A3(n13959), .A4(n13958), .ZN(
        n13970) );
  AOI22_X1 U17082 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13914), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13968) );
  INV_X2 U17083 ( .A(n13962), .ZN(n17562) );
  AOI22_X1 U17084 ( .A1(n17584), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U17085 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U17086 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13965) );
  NAND4_X1 U17087 ( .A1(n13968), .A2(n13967), .A3(n13966), .A4(n13965), .ZN(
        n13969) );
  AOI22_X1 U17088 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19074), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19227), .ZN(n15931) );
  AOI22_X1 U17089 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n19079), .B2(n19219), .ZN(
        n13976) );
  NOR2_X1 U17090 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19227), .ZN(
        n13971) );
  OAI22_X1 U17091 ( .A1(n15932), .A2(n13971), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19074), .ZN(n13975) );
  NOR2_X1 U17092 ( .A1(n13976), .A2(n13975), .ZN(n13972) );
  AOI21_X1 U17093 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19079), .A(
        n13972), .ZN(n13973) );
  AOI22_X1 U17094 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21004), .B1(
        n13973), .B2(n19207), .ZN(n13979) );
  NOR2_X1 U17095 ( .A1(n13973), .A2(n19207), .ZN(n13980) );
  NAND2_X1 U17096 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21004), .ZN(
        n13974) );
  OAI22_X1 U17097 ( .A1(n13979), .A2(n19082), .B1(n13980), .B2(n13974), .ZN(
        n13978) );
  AOI211_X1 U17098 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n19232), .A(
        n15932), .B(n13978), .ZN(n16105) );
  XOR2_X1 U17099 ( .A(n13976), .B(n13975), .Z(n16106) );
  INV_X1 U17100 ( .A(n16106), .ZN(n13977) );
  OAI21_X1 U17101 ( .B1(n13980), .B2(n19082), .A(n13979), .ZN(n13981) );
  INV_X1 U17102 ( .A(n19038), .ZN(n13982) );
  NOR2_X1 U17103 ( .A1(n18625), .A2(n16102), .ZN(n19053) );
  NAND3_X1 U17104 ( .A1(n15966), .A2(n16110), .A3(n19053), .ZN(n15965) );
  INV_X1 U17105 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n13985) );
  INV_X1 U17106 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17469) );
  INV_X1 U17107 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17148) );
  INV_X1 U17108 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17168) );
  INV_X1 U17109 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17194) );
  INV_X1 U17110 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17220) );
  INV_X1 U17111 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17602) );
  INV_X1 U17112 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n13984) );
  NAND4_X1 U17113 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(P3_EBX_REG_2__SCAN_IN), .ZN(n17594) );
  NAND2_X1 U17114 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17603), .ZN(n17599) );
  NOR2_X1 U17115 ( .A1(n17625), .A2(n17342), .ZN(n17454) );
  AOI22_X1 U17116 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13996) );
  AOI22_X1 U17117 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13995) );
  AOI22_X1 U17118 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13987) );
  OAI21_X1 U17119 ( .B1(n17458), .B2(n17618), .A(n13987), .ZN(n13993) );
  AOI22_X1 U17120 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13991) );
  AOI22_X1 U17121 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U17122 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U17123 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13988) );
  NAND4_X1 U17124 ( .A1(n13991), .A2(n13990), .A3(n13989), .A4(n13988), .ZN(
        n13992) );
  AOI211_X1 U17125 ( .C1(n17562), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n13993), .B(n13992), .ZN(n13994) );
  NAND3_X1 U17126 ( .A1(n13996), .A2(n13995), .A3(n13994), .ZN(n17695) );
  AOI22_X1 U17127 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17454), .B1(n17625), 
        .B2(n17695), .ZN(n13999) );
  NAND3_X1 U17128 ( .A1(n18639), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n9749), .ZN(
        n17470) );
  INV_X1 U17129 ( .A(n17470), .ZN(n13997) );
  NAND3_X1 U17130 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n13985), .A3(n13997), 
        .ZN(n13998) );
  NAND2_X1 U17131 ( .A1(n13999), .A2(n13998), .ZN(P3_U2685) );
  NOR2_X1 U17132 ( .A1(n19219), .A2(n19227), .ZN(n19060) );
  AOI21_X1 U17133 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19060), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15963) );
  NAND2_X1 U17134 ( .A1(n15963), .A2(n17458), .ZN(n18597) );
  NOR2_X1 U17135 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18597), .ZN(n14000) );
  INV_X1 U17136 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19249) );
  NOR2_X1 U17137 ( .A1(n19212), .A2(n19249), .ZN(n19106) );
  NAND2_X1 U17138 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19106), .ZN(n19200) );
  NAND2_X1 U17139 ( .A1(n19212), .A2(n19261), .ZN(n19248) );
  NAND2_X1 U17140 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18596) );
  OAI21_X1 U17141 ( .B1(n14000), .B2(n19200), .A(n18842), .ZN(n18604) );
  INV_X1 U17142 ( .A(n18604), .ZN(n14001) );
  AOI21_X1 U17143 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19255)
         );
  NOR2_X1 U17144 ( .A1(n19212), .A2(n16967), .ZN(n19107) );
  INV_X1 U17145 ( .A(n19107), .ZN(n18160) );
  AOI22_X1 U17146 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n19255), .B2(n18160), .ZN(n15929) );
  NOR2_X1 U17147 ( .A1(n14001), .A2(n15929), .ZN(n14003) );
  NOR3_X1 U17148 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16967), .ZN(n18662) );
  NOR2_X1 U17149 ( .A1(n19202), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18643) );
  OR2_X1 U17150 ( .A1(n18643), .A2(n14001), .ZN(n15927) );
  OR2_X1 U17151 ( .A1(n18662), .A2(n15927), .ZN(n14002) );
  MUX2_X1 U17152 ( .A(n14003), .B(n14002), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17153 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .ZN(n17341) );
  NAND2_X1 U17154 ( .A1(n18639), .A2(n17621), .ZN(n17627) );
  INV_X1 U17155 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17041) );
  INV_X1 U17156 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17343) );
  NAND3_X1 U17157 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17426), .ZN(n17395) );
  OAI21_X1 U17158 ( .B1(n17341), .B2(n17627), .A(n17383), .ZN(n17378) );
  AOI22_X1 U17159 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U17160 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17161 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14005) );
  AOI22_X1 U17162 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14004) );
  NAND4_X1 U17163 ( .A1(n14007), .A2(n14006), .A3(n14005), .A4(n14004), .ZN(
        n14013) );
  AOI22_X1 U17164 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n13986), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14011) );
  AOI22_X1 U17165 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U17166 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U17167 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14008) );
  NAND4_X1 U17168 ( .A1(n14011), .A2(n14010), .A3(n14009), .A4(n14008), .ZN(
        n14012) );
  NOR2_X1 U17169 ( .A1(n14013), .A2(n14012), .ZN(n17375) );
  AOI22_X1 U17170 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14017) );
  AOI22_X1 U17171 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14016) );
  AOI22_X1 U17172 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n17571), .B1(
        n9669), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14015) );
  AOI22_X1 U17173 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14014) );
  NAND4_X1 U17174 ( .A1(n14017), .A2(n14016), .A3(n14015), .A4(n14014), .ZN(
        n14023) );
  AOI22_X1 U17175 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14021) );
  AOI22_X1 U17176 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U17177 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U17178 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14018) );
  NAND4_X1 U17179 ( .A1(n14021), .A2(n14020), .A3(n14019), .A4(n14018), .ZN(
        n14022) );
  NOR2_X1 U17180 ( .A1(n14023), .A2(n14022), .ZN(n17386) );
  AOI22_X1 U17181 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17561), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14028) );
  AOI22_X1 U17182 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17555), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9667), .ZN(n14027) );
  AOI22_X1 U17183 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n16041), .ZN(n14026) );
  AOI22_X1 U17184 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17554), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14025) );
  NAND4_X1 U17185 ( .A1(n14028), .A2(n14027), .A3(n14026), .A4(n14025), .ZN(
        n14034) );
  AOI22_X1 U17186 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17575), .ZN(n14032) );
  AOI22_X1 U17187 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17571), .ZN(n14031) );
  AOI22_X1 U17188 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n13986), .ZN(n14030) );
  AOI22_X1 U17189 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14029) );
  NAND4_X1 U17190 ( .A1(n14032), .A2(n14031), .A3(n14030), .A4(n14029), .ZN(
        n14033) );
  NOR2_X1 U17191 ( .A1(n14034), .A2(n14033), .ZN(n17393) );
  AOI22_X1 U17192 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17573), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U17193 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14045) );
  INV_X1 U17194 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14036) );
  AOI22_X1 U17195 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14035) );
  OAI21_X1 U17196 ( .B1(n14037), .B2(n14036), .A(n14035), .ZN(n14043) );
  AOI22_X1 U17197 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U17198 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U17199 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U17200 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13986), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14038) );
  NAND4_X1 U17201 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14042) );
  AOI211_X1 U17202 ( .C1(n9669), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n14043), .B(n14042), .ZN(n14044) );
  NAND3_X1 U17203 ( .A1(n14046), .A2(n14045), .A3(n14044), .ZN(n17397) );
  AOI22_X1 U17204 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14056) );
  AOI22_X1 U17205 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14055) );
  INV_X1 U17206 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n21001) );
  AOI22_X1 U17207 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14047) );
  OAI21_X1 U17208 ( .B1(n21001), .B2(n17538), .A(n14047), .ZN(n14053) );
  AOI22_X1 U17209 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13986), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17210 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U17211 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U17212 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14048) );
  NAND4_X1 U17213 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14052) );
  AOI211_X1 U17214 ( .C1(n17556), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n14053), .B(n14052), .ZN(n14054) );
  NAND3_X1 U17215 ( .A1(n14056), .A2(n14055), .A3(n14054), .ZN(n17398) );
  NAND2_X1 U17216 ( .A1(n17397), .A2(n17398), .ZN(n17396) );
  NOR2_X1 U17217 ( .A1(n17393), .A2(n17396), .ZN(n17391) );
  AOI22_X1 U17218 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14066) );
  AOI22_X1 U17219 ( .A1(n9676), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13986), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14065) );
  AOI22_X1 U17220 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14057) );
  OAI21_X1 U17221 ( .B1(n13957), .B2(n17618), .A(n14057), .ZN(n14063) );
  AOI22_X1 U17222 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U17223 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U17224 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U17225 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14058) );
  NAND4_X1 U17226 ( .A1(n14061), .A2(n14060), .A3(n14059), .A4(n14058), .ZN(
        n14062) );
  AOI211_X1 U17227 ( .C1(n9669), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n14063), .B(n14062), .ZN(n14064) );
  NAND3_X1 U17228 ( .A1(n14066), .A2(n14065), .A3(n14064), .ZN(n17390) );
  NAND2_X1 U17229 ( .A1(n17391), .A2(n17390), .ZN(n17389) );
  NOR2_X1 U17230 ( .A1(n17386), .A2(n17389), .ZN(n17650) );
  AOI22_X1 U17231 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U17232 ( .A1(n13949), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14075) );
  INV_X1 U17233 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n21027) );
  AOI22_X1 U17234 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14067) );
  OAI21_X1 U17235 ( .B1(n21027), .B2(n10251), .A(n14067), .ZN(n14073) );
  AOI22_X1 U17236 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14071) );
  AOI22_X1 U17237 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U17238 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17562), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14069) );
  AOI22_X1 U17239 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14068) );
  NAND4_X1 U17240 ( .A1(n14071), .A2(n14070), .A3(n14069), .A4(n14068), .ZN(
        n14072) );
  AOI211_X1 U17241 ( .C1(n17539), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n14073), .B(n14072), .ZN(n14074) );
  NAND3_X1 U17242 ( .A1(n14076), .A2(n14075), .A3(n14074), .ZN(n17649) );
  NAND2_X1 U17243 ( .A1(n17650), .A2(n17649), .ZN(n17648) );
  XOR2_X1 U17244 ( .A(n17375), .B(n17648), .Z(n17643) );
  AOI22_X1 U17245 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17378), .B1(n17625), 
        .B2(n17643), .ZN(n14079) );
  INV_X1 U17246 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14077) );
  INV_X1 U17247 ( .A(n17385), .ZN(n17388) );
  NAND3_X1 U17248 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14077), .A3(n17388), 
        .ZN(n14078) );
  NAND2_X1 U17249 ( .A1(n14079), .A2(n14078), .ZN(P3_U2675) );
  XNOR2_X1 U17250 ( .A(n14080), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14846) );
  NAND2_X1 U17251 ( .A1(n14846), .A2(n12477), .ZN(n14098) );
  AOI22_X1 U17252 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U17253 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9672), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17254 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17255 ( .A1(n14338), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14081) );
  NAND4_X1 U17256 ( .A1(n14084), .A2(n14083), .A3(n14082), .A4(n14081), .ZN(
        n14093) );
  AOI22_X1 U17257 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14293), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U17258 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U17259 ( .A1(n14356), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14088) );
  NAND2_X1 U17260 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n14086) );
  AOI21_X1 U17261 ( .B1(n11984), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n14345), .ZN(n14085) );
  AND2_X1 U17262 ( .A1(n14086), .A2(n14085), .ZN(n14087) );
  NAND4_X1 U17263 ( .A1(n14090), .A2(n14089), .A3(n14088), .A4(n14087), .ZN(
        n14092) );
  NAND2_X1 U17264 ( .A1(n14348), .A2(n14351), .ZN(n14197) );
  OAI21_X1 U17265 ( .B1(n14093), .B2(n14092), .A(n14197), .ZN(n14096) );
  NAND2_X1 U17266 ( .A1(n14445), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n14095) );
  NAND2_X1 U17267 ( .A1(n20697), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14094) );
  NAND3_X1 U17268 ( .A1(n14096), .A2(n14095), .A3(n14094), .ZN(n14097) );
  NAND2_X1 U17269 ( .A1(n14098), .A2(n14097), .ZN(n14561) );
  XNOR2_X1 U17270 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n14100), .ZN(
        n16348) );
  AOI22_X1 U17271 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17272 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14103) );
  AOI22_X1 U17273 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U17274 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14101) );
  NAND4_X1 U17275 ( .A1(n14104), .A2(n14103), .A3(n14102), .A4(n14101), .ZN(
        n14110) );
  AOI22_X1 U17276 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17277 ( .A1(n14356), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U17278 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U17279 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14105) );
  NAND4_X1 U17280 ( .A1(n14108), .A2(n14107), .A3(n14106), .A4(n14105), .ZN(
        n14109) );
  OR2_X1 U17281 ( .A1(n14110), .A2(n14109), .ZN(n14113) );
  OAI22_X1 U17282 ( .A1(n14285), .A2(n12164), .B1(n14111), .B2(n16289), .ZN(
        n14112) );
  AOI21_X1 U17283 ( .B1(n14375), .B2(n14113), .A(n14112), .ZN(n14114) );
  OAI21_X1 U17284 ( .B1(n16348), .B2(n14351), .A(n14114), .ZN(n14115) );
  INV_X1 U17285 ( .A(n14115), .ZN(n14659) );
  XNOR2_X1 U17286 ( .A(n14116), .B(n16280), .ZN(n16277) );
  AOI22_X1 U17287 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14120) );
  AOI22_X1 U17288 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14119) );
  AOI22_X1 U17289 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U17290 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14117) );
  NAND4_X1 U17291 ( .A1(n14120), .A2(n14119), .A3(n14118), .A4(n14117), .ZN(
        n14128) );
  AOI22_X1 U17292 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17293 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U17294 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14122) );
  AOI21_X1 U17295 ( .B1(n11984), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n12477), .ZN(n14121) );
  AND2_X1 U17296 ( .A1(n14122), .A2(n14121), .ZN(n14124) );
  AOI22_X1 U17297 ( .A1(n14357), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14123) );
  NAND4_X1 U17298 ( .A1(n14126), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        n14127) );
  OAI21_X1 U17299 ( .B1(n14128), .B2(n14127), .A(n14197), .ZN(n14131) );
  NAND2_X1 U17300 ( .A1(n14445), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n14130) );
  NAND2_X1 U17301 ( .A1(n20697), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14129) );
  NAND3_X1 U17302 ( .A1(n14131), .A2(n14130), .A3(n14129), .ZN(n14132) );
  OAI21_X1 U17303 ( .B1(n16277), .B2(n14351), .A(n14132), .ZN(n14652) );
  OR2_X1 U17304 ( .A1(n14134), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14135) );
  NAND2_X1 U17305 ( .A1(n14135), .A2(n14164), .ZN(n16340) );
  INV_X1 U17306 ( .A(n16340), .ZN(n16267) );
  AOI22_X1 U17307 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14219), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14139) );
  AOI22_X1 U17308 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U17309 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17310 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14136) );
  NAND4_X1 U17311 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14145) );
  AOI22_X1 U17312 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17313 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14142) );
  AOI22_X1 U17314 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U17315 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14140) );
  NAND4_X1 U17316 ( .A1(n14143), .A2(n14142), .A3(n14141), .A4(n14140), .ZN(
        n14144) );
  OR2_X1 U17317 ( .A1(n14145), .A2(n14144), .ZN(n14149) );
  INV_X1 U17318 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14147) );
  NAND2_X1 U17319 ( .A1(n20697), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14146) );
  OAI211_X1 U17320 ( .C1(n14285), .C2(n14147), .A(n14351), .B(n14146), .ZN(
        n14148) );
  AOI21_X1 U17321 ( .B1(n14375), .B2(n14149), .A(n14148), .ZN(n14150) );
  AOI21_X1 U17322 ( .B1(n16267), .B2(n14345), .A(n14150), .ZN(n16268) );
  AOI22_X1 U17323 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9686), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U17324 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17325 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14152) );
  AOI22_X1 U17326 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11923), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14151) );
  NAND4_X1 U17327 ( .A1(n14154), .A2(n14153), .A3(n14152), .A4(n14151), .ZN(
        n14160) );
  AOI22_X1 U17328 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9681), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U17329 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14157) );
  AOI22_X1 U17330 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U17331 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14155) );
  NAND4_X1 U17332 ( .A1(n14158), .A2(n14157), .A3(n14156), .A4(n14155), .ZN(
        n14159) );
  NOR2_X1 U17333 ( .A1(n14160), .A2(n14159), .ZN(n14163) );
  AOI21_X1 U17334 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n16261), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14161) );
  AOI21_X1 U17335 ( .B1(n14445), .B2(P1_EAX_REG_20__SCAN_IN), .A(n14161), .ZN(
        n14162) );
  OAI21_X1 U17336 ( .B1(n14348), .B2(n14163), .A(n14162), .ZN(n14166) );
  XNOR2_X1 U17337 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n14164), .ZN(
        n16252) );
  NAND2_X1 U17338 ( .A1(n14345), .A2(n16252), .ZN(n14165) );
  NAND2_X1 U17339 ( .A1(n14166), .A2(n14165), .ZN(n14643) );
  OR2_X1 U17340 ( .A1(n14167), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14168) );
  NAND2_X1 U17341 ( .A1(n14168), .A2(n14199), .ZN(n16327) );
  AOI22_X1 U17342 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13337), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14172) );
  AOI22_X1 U17343 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U17344 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U17345 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14169) );
  NAND4_X1 U17346 ( .A1(n14172), .A2(n14171), .A3(n14170), .A4(n14169), .ZN(
        n14178) );
  AOI22_X1 U17347 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14176) );
  AOI22_X1 U17348 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U17349 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U17350 ( .A1(n14356), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14173) );
  NAND4_X1 U17351 ( .A1(n14176), .A2(n14175), .A3(n14174), .A4(n14173), .ZN(
        n14177) );
  NOR2_X1 U17352 ( .A1(n14178), .A2(n14177), .ZN(n14181) );
  OAI21_X1 U17353 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20702), .A(
        n20697), .ZN(n14180) );
  NAND2_X1 U17354 ( .A1(n14445), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n14179) );
  OAI211_X1 U17355 ( .C1(n14348), .C2(n14181), .A(n14180), .B(n14179), .ZN(
        n14182) );
  OAI21_X1 U17356 ( .B1(n16327), .B2(n14351), .A(n14182), .ZN(n14635) );
  AOI22_X1 U17357 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U17358 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14188) );
  AOI22_X1 U17359 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U17360 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14185) );
  AOI21_X1 U17361 ( .B1(n11984), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n14345), .ZN(n14184) );
  AND2_X1 U17362 ( .A1(n14185), .A2(n14184), .ZN(n14186) );
  NAND4_X1 U17363 ( .A1(n14189), .A2(n14188), .A3(n14187), .A4(n14186), .ZN(
        n14195) );
  AOI22_X1 U17364 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14193) );
  AOI22_X1 U17365 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U17366 ( .A1(n14338), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14191) );
  AOI22_X1 U17367 ( .A1(n11923), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14190) );
  NAND4_X1 U17368 ( .A1(n14193), .A2(n14192), .A3(n14191), .A4(n14190), .ZN(
        n14194) );
  OR2_X1 U17369 ( .A1(n14195), .A2(n14194), .ZN(n14196) );
  NAND2_X1 U17370 ( .A1(n14197), .A2(n14196), .ZN(n14202) );
  OAI22_X1 U17371 ( .A1(n14285), .A2(n12146), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13002), .ZN(n14198) );
  INV_X1 U17372 ( .A(n14198), .ZN(n14201) );
  XNOR2_X1 U17373 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n14199), .ZN(
        n16235) );
  AOI21_X1 U17374 ( .B1(n14202), .B2(n14201), .A(n14200), .ZN(n14629) );
  OR2_X1 U17375 ( .A1(n14203), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14204) );
  NAND2_X1 U17376 ( .A1(n14231), .A2(n14204), .ZN(n16326) );
  AOI22_X1 U17377 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14208) );
  AOI22_X1 U17378 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14338), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14207) );
  AOI22_X1 U17379 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14206) );
  AOI22_X1 U17380 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14205) );
  NAND4_X1 U17381 ( .A1(n14208), .A2(n14207), .A3(n14206), .A4(n14205), .ZN(
        n14214) );
  AOI22_X1 U17382 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14212) );
  AOI22_X1 U17383 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14219), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14211) );
  AOI22_X1 U17384 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14210) );
  AOI22_X1 U17385 ( .A1(n14337), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14209) );
  NAND4_X1 U17386 ( .A1(n14212), .A2(n14211), .A3(n14210), .A4(n14209), .ZN(
        n14213) );
  NOR2_X1 U17387 ( .A1(n14214), .A2(n14213), .ZN(n14232) );
  AOI22_X1 U17388 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14218) );
  AOI22_X1 U17389 ( .A1(n14356), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14217) );
  AOI22_X1 U17390 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14216) );
  AOI22_X1 U17391 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14215) );
  NAND4_X1 U17392 ( .A1(n14218), .A2(n14217), .A3(n14216), .A4(n14215), .ZN(
        n14225) );
  AOI22_X1 U17393 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14223) );
  AOI22_X1 U17394 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14222) );
  AOI22_X1 U17395 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14221) );
  AOI22_X1 U17396 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14220) );
  NAND4_X1 U17397 ( .A1(n14223), .A2(n14222), .A3(n14221), .A4(n14220), .ZN(
        n14224) );
  NOR2_X1 U17398 ( .A1(n14225), .A2(n14224), .ZN(n14233) );
  XNOR2_X1 U17399 ( .A(n14232), .B(n14233), .ZN(n14226) );
  NOR2_X1 U17400 ( .A1(n14226), .A2(n14348), .ZN(n14229) );
  NAND2_X1 U17401 ( .A1(n20697), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14227) );
  OAI211_X1 U17402 ( .C1(n14285), .C2(n12160), .A(n14351), .B(n14227), .ZN(
        n14228) );
  OAI22_X1 U17403 ( .A1(n16326), .A2(n14351), .B1(n14229), .B2(n14228), .ZN(
        n14621) );
  INV_X1 U17404 ( .A(n14621), .ZN(n14230) );
  XNOR2_X1 U17405 ( .A(n14231), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16215) );
  NAND2_X1 U17406 ( .A1(n16215), .A2(n12477), .ZN(n14249) );
  NOR2_X1 U17407 ( .A1(n14233), .A2(n14232), .ZN(n14264) );
  AOI22_X1 U17408 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U17409 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U17410 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14235) );
  AOI22_X1 U17411 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14234) );
  NAND4_X1 U17412 ( .A1(n14237), .A2(n14236), .A3(n14235), .A4(n14234), .ZN(
        n14243) );
  AOI22_X1 U17413 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U17414 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14240) );
  AOI22_X1 U17415 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U17416 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14238) );
  NAND4_X1 U17417 ( .A1(n14241), .A2(n14240), .A3(n14239), .A4(n14238), .ZN(
        n14242) );
  OR2_X1 U17418 ( .A1(n14243), .A2(n14242), .ZN(n14263) );
  XNOR2_X1 U17419 ( .A(n14264), .B(n14263), .ZN(n14247) );
  NAND2_X1 U17420 ( .A1(n20697), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14244) );
  OAI211_X1 U17421 ( .C1(n14285), .C2(n12144), .A(n14351), .B(n14244), .ZN(
        n14245) );
  INV_X1 U17422 ( .A(n14245), .ZN(n14246) );
  OAI21_X1 U17423 ( .B1(n14247), .B2(n14348), .A(n14246), .ZN(n14248) );
  NAND2_X1 U17424 ( .A1(n14249), .A2(n14248), .ZN(n14614) );
  NAND2_X1 U17425 ( .A1(n14251), .A2(n14250), .ZN(n14252) );
  NAND2_X1 U17426 ( .A1(n14270), .A2(n14252), .ZN(n14801) );
  AOI22_X1 U17427 ( .A1(n14356), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14256) );
  AOI22_X1 U17428 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14255) );
  AOI22_X1 U17429 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14254) );
  AOI22_X1 U17430 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14253) );
  NAND4_X1 U17431 ( .A1(n14256), .A2(n14255), .A3(n14254), .A4(n14253), .ZN(
        n14262) );
  AOI22_X1 U17432 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14260) );
  AOI22_X1 U17433 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14259) );
  AOI22_X1 U17434 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14258) );
  AOI22_X1 U17435 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14257) );
  NAND4_X1 U17436 ( .A1(n14260), .A2(n14259), .A3(n14258), .A4(n14257), .ZN(
        n14261) );
  NOR2_X1 U17437 ( .A1(n14262), .A2(n14261), .ZN(n14272) );
  NAND2_X1 U17438 ( .A1(n14264), .A2(n14263), .ZN(n14271) );
  XNOR2_X1 U17439 ( .A(n14272), .B(n14271), .ZN(n14265) );
  NOR2_X1 U17440 ( .A1(n14265), .A2(n14348), .ZN(n14269) );
  INV_X1 U17441 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14267) );
  NAND2_X1 U17442 ( .A1(n20697), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14266) );
  OAI211_X1 U17443 ( .C1(n14285), .C2(n14267), .A(n14351), .B(n14266), .ZN(
        n14268) );
  XNOR2_X1 U17444 ( .A(n14270), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14795) );
  NOR2_X1 U17445 ( .A1(n14272), .A2(n14271), .ZN(n14305) );
  AOI22_X1 U17446 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14276) );
  AOI22_X1 U17447 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14275) );
  AOI22_X1 U17448 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14274) );
  AOI22_X1 U17449 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14273) );
  NAND4_X1 U17450 ( .A1(n14276), .A2(n14275), .A3(n14274), .A4(n14273), .ZN(
        n14282) );
  AOI22_X1 U17451 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14280) );
  AOI22_X1 U17452 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14279) );
  AOI22_X1 U17453 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14278) );
  AOI22_X1 U17454 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14277) );
  NAND4_X1 U17455 ( .A1(n14280), .A2(n14279), .A3(n14278), .A4(n14277), .ZN(
        n14281) );
  OR2_X1 U17456 ( .A1(n14282), .A2(n14281), .ZN(n14304) );
  INV_X1 U17457 ( .A(n14304), .ZN(n14283) );
  XNOR2_X1 U17458 ( .A(n14305), .B(n14283), .ZN(n14287) );
  OAI21_X1 U17459 ( .B1(n20702), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n20697), .ZN(n14284) );
  OAI21_X1 U17460 ( .B1(n14285), .B2(n12156), .A(n14284), .ZN(n14286) );
  AOI21_X1 U17461 ( .B1(n14287), .B2(n14375), .A(n14286), .ZN(n14288) );
  INV_X1 U17462 ( .A(n14289), .ZN(n14291) );
  INV_X1 U17463 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14290) );
  NAND2_X1 U17464 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  NAND2_X1 U17465 ( .A1(n14310), .A2(n14292), .ZN(n14784) );
  AOI22_X1 U17466 ( .A1(n14293), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U17467 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n14356), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U17468 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14295) );
  AOI22_X1 U17469 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14294) );
  NAND4_X1 U17470 ( .A1(n14297), .A2(n14296), .A3(n14295), .A4(n14294), .ZN(
        n14303) );
  AOI22_X1 U17471 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12199), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14301) );
  AOI22_X1 U17472 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14300) );
  AOI22_X1 U17473 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17474 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14298) );
  NAND4_X1 U17475 ( .A1(n14301), .A2(n14300), .A3(n14299), .A4(n14298), .ZN(
        n14302) );
  NOR2_X1 U17476 ( .A1(n14303), .A2(n14302), .ZN(n14323) );
  NAND2_X1 U17477 ( .A1(n14305), .A2(n14304), .ZN(n14322) );
  XNOR2_X1 U17478 ( .A(n14323), .B(n14322), .ZN(n14308) );
  AOI21_X1 U17479 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20697), .A(
        n12477), .ZN(n14307) );
  NAND2_X1 U17480 ( .A1(n14445), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n14306) );
  OAI211_X1 U17481 ( .C1(n14308), .C2(n14348), .A(n14307), .B(n14306), .ZN(
        n14309) );
  OAI21_X1 U17482 ( .B1(n14784), .B2(n14351), .A(n14309), .ZN(n14522) );
  XNOR2_X1 U17483 ( .A(n14310), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14776) );
  INV_X1 U17484 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14773) );
  AOI21_X1 U17485 ( .B1(n14773), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14311) );
  AOI21_X1 U17486 ( .B1(n14445), .B2(P1_EAX_REG_28__SCAN_IN), .A(n14311), .ZN(
        n14326) );
  AOI22_X1 U17487 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14315) );
  INV_X1 U17488 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n21031) );
  AOI22_X1 U17489 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U17490 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U17491 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14312) );
  NAND4_X1 U17492 ( .A1(n14315), .A2(n14314), .A3(n14313), .A4(n14312), .ZN(
        n14321) );
  AOI22_X1 U17493 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U17494 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U17495 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U17496 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14316) );
  NAND4_X1 U17497 ( .A1(n14319), .A2(n14318), .A3(n14317), .A4(n14316), .ZN(
        n14320) );
  OR2_X1 U17498 ( .A1(n14321), .A2(n14320), .ZN(n14331) );
  NOR2_X1 U17499 ( .A1(n14323), .A2(n14322), .ZN(n14332) );
  XOR2_X1 U17500 ( .A(n14331), .B(n14332), .Z(n14324) );
  NAND2_X1 U17501 ( .A1(n14324), .A2(n14375), .ZN(n14325) );
  AOI22_X1 U17502 ( .A1(n14776), .A2(n12477), .B1(n14326), .B2(n14325), .ZN(
        n14473) );
  INV_X1 U17503 ( .A(n14327), .ZN(n14329) );
  INV_X1 U17504 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14328) );
  NAND2_X1 U17505 ( .A1(n14329), .A2(n14328), .ZN(n14330) );
  NAND2_X1 U17506 ( .A1(n14352), .A2(n14330), .ZN(n14761) );
  NAND2_X1 U17507 ( .A1(n14332), .A2(n14331), .ZN(n14354) );
  AOI22_X1 U17508 ( .A1(n13337), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14336) );
  AOI22_X1 U17509 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14335) );
  AOI22_X1 U17510 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U17511 ( .A1(n12219), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14333) );
  NAND4_X1 U17512 ( .A1(n14336), .A2(n14335), .A3(n14334), .A4(n14333), .ZN(
        n14344) );
  AOI22_X1 U17513 ( .A1(n14365), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14342) );
  AOI22_X1 U17514 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14337), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17515 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U17516 ( .A1(n14338), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14339) );
  NAND4_X1 U17517 ( .A1(n14342), .A2(n14341), .A3(n14340), .A4(n14339), .ZN(
        n14343) );
  NOR2_X1 U17518 ( .A1(n14344), .A2(n14343), .ZN(n14355) );
  XNOR2_X1 U17519 ( .A(n14354), .B(n14355), .ZN(n14349) );
  AOI21_X1 U17520 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20697), .A(
        n14345), .ZN(n14347) );
  NAND2_X1 U17521 ( .A1(n14445), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n14346) );
  OAI211_X1 U17522 ( .C1(n14349), .C2(n14348), .A(n14347), .B(n14346), .ZN(
        n14350) );
  OAI21_X1 U17523 ( .B1(n14761), .B2(n14351), .A(n14350), .ZN(n14512) );
  XNOR2_X1 U17524 ( .A(n14352), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14751) );
  NOR2_X1 U17525 ( .A1(n14753), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14353) );
  AOI211_X1 U17526 ( .C1(n14445), .C2(P1_EAX_REG_30__SCAN_IN), .A(n14353), .B(
        n12477), .ZN(n14378) );
  NOR2_X1 U17527 ( .A1(n14355), .A2(n14354), .ZN(n14374) );
  AOI22_X1 U17528 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14356), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U17529 ( .A1(n14358), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14357), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U17530 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U17531 ( .A1(n14337), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14359), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14360) );
  NAND4_X1 U17532 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14360), .ZN(
        n14372) );
  AOI22_X1 U17533 ( .A1(n14364), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11989), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U17534 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14369) );
  AOI22_X1 U17535 ( .A1(n12198), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14365), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U17536 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14367) );
  NAND4_X1 U17537 ( .A1(n14370), .A2(n14369), .A3(n14368), .A4(n14367), .ZN(
        n14371) );
  NOR2_X1 U17538 ( .A1(n14372), .A2(n14371), .ZN(n14373) );
  XNOR2_X1 U17539 ( .A(n14374), .B(n14373), .ZN(n14376) );
  NAND2_X1 U17540 ( .A1(n14376), .A2(n14375), .ZN(n14377) );
  AOI22_X1 U17541 ( .A1(n14751), .A2(n12477), .B1(n14378), .B2(n14377), .ZN(
        n14443) );
  XNOR2_X1 U17542 ( .A(n14510), .B(n14443), .ZN(n14502) );
  INV_X1 U17543 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14423) );
  NAND2_X1 U17544 ( .A1(n14457), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14380) );
  NAND2_X1 U17545 ( .A1(n14456), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14379) );
  NAND2_X1 U17546 ( .A1(n14380), .A2(n14379), .ZN(n14452) );
  MUX2_X1 U17547 ( .A(n14417), .B(n14454), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n14383) );
  INV_X1 U17548 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14381) );
  NAND2_X1 U17549 ( .A1(n14405), .A2(n14381), .ZN(n14382) );
  NAND2_X1 U17550 ( .A1(n12753), .A2(n16413), .ZN(n14384) );
  OAI211_X1 U17551 ( .C1(n14456), .C2(P1_EBX_REG_17__SCAN_IN), .A(n14384), .B(
        n14454), .ZN(n14385) );
  OAI21_X1 U17552 ( .B1(n14410), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14385), .ZN(
        n14660) );
  INV_X1 U17553 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14991) );
  NAND2_X1 U17554 ( .A1(n14991), .A2(n14405), .ZN(n14387) );
  MUX2_X1 U17555 ( .A(n14417), .B(n14454), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14386) );
  NAND2_X1 U17556 ( .A1(n14387), .A2(n14386), .ZN(n14653) );
  INV_X1 U17557 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14388) );
  NAND2_X1 U17558 ( .A1(n14399), .A2(n14388), .ZN(n14391) );
  INV_X1 U17559 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16178) );
  NAND2_X1 U17560 ( .A1(n9988), .A2(n14388), .ZN(n14389) );
  OAI211_X1 U17561 ( .C1(n14419), .C2(n16178), .A(n14389), .B(n12753), .ZN(
        n14390) );
  AND2_X1 U17562 ( .A1(n14391), .A2(n14390), .ZN(n14646) );
  INV_X1 U17563 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16314) );
  NAND2_X1 U17564 ( .A1(n14412), .A2(n16314), .ZN(n14395) );
  INV_X1 U17565 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U17566 ( .A1(n12753), .A2(n14392), .ZN(n14393) );
  OAI211_X1 U17567 ( .C1(n14456), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14393), .B(
        n14454), .ZN(n14394) );
  NAND2_X1 U17568 ( .A1(n14395), .A2(n14394), .ZN(n16271) );
  NAND2_X1 U17569 ( .A1(n14646), .A2(n16271), .ZN(n14396) );
  INV_X1 U17570 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16180) );
  NAND2_X1 U17571 ( .A1(n12753), .A2(n16180), .ZN(n14397) );
  OAI211_X1 U17572 ( .C1(n14456), .C2(P1_EBX_REG_21__SCAN_IN), .A(n14397), .B(
        n14454), .ZN(n14398) );
  OAI21_X1 U17573 ( .B1(n14410), .B2(P1_EBX_REG_21__SCAN_IN), .A(n14398), .ZN(
        n14636) );
  AND2_X2 U17574 ( .A1(n14647), .A2(n14636), .ZN(n14638) );
  MUX2_X1 U17575 ( .A(n14399), .B(n14419), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14401) );
  NOR2_X1 U17576 ( .A1(n14457), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14400) );
  NOR2_X1 U17577 ( .A1(n14401), .A2(n14400), .ZN(n14631) );
  INV_X1 U17578 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14625) );
  NAND2_X1 U17579 ( .A1(n14412), .A2(n14625), .ZN(n14404) );
  INV_X1 U17580 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14980) );
  NAND2_X1 U17581 ( .A1(n12753), .A2(n14980), .ZN(n14402) );
  OAI211_X1 U17582 ( .C1(n14456), .C2(P1_EBX_REG_23__SCAN_IN), .A(n14402), .B(
        n14454), .ZN(n14403) );
  INV_X1 U17583 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14809) );
  NAND2_X1 U17584 ( .A1(n14809), .A2(n14405), .ZN(n14407) );
  MUX2_X1 U17585 ( .A(n14417), .B(n14454), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14406) );
  NAND2_X1 U17586 ( .A1(n14407), .A2(n14406), .ZN(n14615) );
  INV_X1 U17587 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14953) );
  NAND2_X1 U17588 ( .A1(n12753), .A2(n14953), .ZN(n14408) );
  OAI211_X1 U17589 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14456), .A(n14408), .B(
        n14454), .ZN(n14409) );
  OAI21_X1 U17590 ( .B1(n14410), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14409), .ZN(
        n14549) );
  MUX2_X1 U17591 ( .A(n14417), .B(n14454), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14411) );
  OAI21_X1 U17592 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14457), .A(
        n14411), .ZN(n14535) );
  INV_X1 U17593 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21016) );
  NAND2_X1 U17594 ( .A1(n14412), .A2(n21016), .ZN(n14416) );
  INV_X1 U17595 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14413) );
  OAI21_X1 U17596 ( .B1(n14419), .B2(n14413), .A(n12753), .ZN(n14414) );
  OAI21_X1 U17597 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(n14456), .A(n14414), .ZN(
        n14415) );
  AND2_X1 U17598 ( .A1(n14416), .A2(n14415), .ZN(n14523) );
  MUX2_X1 U17599 ( .A(n14417), .B(n14454), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14418) );
  OAI21_X1 U17600 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14457), .A(
        n14418), .ZN(n14488) );
  MUX2_X1 U17601 ( .A(n14419), .B(n14452), .S(n14513), .Z(n14422) );
  AND2_X1 U17602 ( .A1(n14456), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14420) );
  AOI21_X1 U17603 ( .B1(n14457), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14420), .ZN(
        n14455) );
  INV_X1 U17604 ( .A(n14455), .ZN(n14421) );
  XNOR2_X1 U17605 ( .A(n14422), .B(n14421), .ZN(n14917) );
  OAI222_X1 U17606 ( .A1(n14666), .A2(n14502), .B1(n14423), .B2(n20390), .C1(
        n20385), .C2(n14917), .ZN(P1_U2842) );
  INV_X4 U17607 ( .A(n14806), .ZN(n14877) );
  NAND2_X1 U17608 ( .A1(n14877), .A2(n14425), .ZN(n14426) );
  NAND2_X1 U17609 ( .A1(n14806), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14856) );
  NAND2_X1 U17610 ( .A1(n13723), .A2(n16448), .ZN(n14427) );
  NAND2_X1 U17611 ( .A1(n14856), .A2(n14427), .ZN(n14869) );
  NOR2_X1 U17612 ( .A1(n14869), .A2(n14868), .ZN(n14855) );
  NAND3_X1 U17613 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U17614 ( .A1(n13723), .A2(n14428), .ZN(n14429) );
  NAND2_X1 U17615 ( .A1(n14806), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14430) );
  NAND2_X1 U17616 ( .A1(n14856), .A2(n14430), .ZN(n14432) );
  NOR2_X1 U17617 ( .A1(n13723), .A2(n14431), .ZN(n14842) );
  NOR2_X1 U17618 ( .A1(n14432), .A2(n14842), .ZN(n16341) );
  XNOR2_X1 U17619 ( .A(n14877), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14845) );
  NAND2_X1 U17620 ( .A1(n13723), .A2(n14431), .ZN(n14843) );
  INV_X1 U17621 ( .A(n14432), .ZN(n14434) );
  NOR2_X1 U17622 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14865) );
  NAND2_X1 U17623 ( .A1(n14865), .A2(n16453), .ZN(n14433) );
  NAND2_X1 U17624 ( .A1(n14806), .A2(n14433), .ZN(n14852) );
  NAND2_X1 U17625 ( .A1(n14434), .A2(n14852), .ZN(n14839) );
  INV_X1 U17626 ( .A(n14839), .ZN(n14435) );
  NAND2_X1 U17627 ( .A1(n9668), .A2(n14991), .ZN(n16335) );
  NAND2_X1 U17628 ( .A1(n13723), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14437) );
  NAND2_X1 U17629 ( .A1(n16335), .A2(n14437), .ZN(n14832) );
  NAND2_X1 U17630 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16197) );
  NAND2_X1 U17631 ( .A1(n14953), .A2(n14809), .ZN(n14765) );
  AND2_X1 U17632 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14954) );
  NAND2_X1 U17633 ( .A1(n14954), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14949) );
  INV_X1 U17634 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20885) );
  NAND2_X1 U17635 ( .A1(n14777), .A2(n14877), .ZN(n14797) );
  NOR2_X1 U17636 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14931) );
  AND2_X1 U17637 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14932) );
  AND2_X1 U17638 ( .A1(n14877), .A2(n14932), .ZN(n14440) );
  INV_X1 U17639 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14441) );
  MUX2_X2 U17640 ( .A(n14749), .B(n14748), .S(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n14442) );
  XNOR2_X1 U17641 ( .A(n14442), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14911) );
  AOI22_X1 U17642 ( .A1(n14445), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n14444), .ZN(n14446) );
  INV_X1 U17643 ( .A(n14446), .ZN(n14447) );
  INV_X1 U17644 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20833) );
  NOR2_X1 U17645 ( .A1(n16489), .A2(n20833), .ZN(n14893) );
  AOI21_X1 U17646 ( .B1(n20450), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14893), .ZN(n14448) );
  OAI21_X1 U17647 ( .B1(n14449), .B2(n20461), .A(n14448), .ZN(n14450) );
  OAI21_X1 U17648 ( .B1(n14911), .B2(n20299), .A(n14451), .ZN(P1_U2968) );
  XNOR2_X1 U17649 ( .A(n14452), .B(n14454), .ZN(n14514) );
  NAND2_X1 U17650 ( .A1(n14513), .A2(n14514), .ZN(n14453) );
  MUX2_X1 U17651 ( .A(n14455), .B(n14454), .S(n14453), .Z(n14459) );
  AOI22_X1 U17652 ( .A1(n14457), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14456), .ZN(n14458) );
  XNOR2_X1 U17653 ( .A(n14459), .B(n14458), .ZN(n14889) );
  NAND2_X1 U17654 ( .A1(n14499), .A2(n20348), .ZN(n14471) );
  NOR2_X1 U17655 ( .A1(n16239), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16223) );
  INV_X1 U17656 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20817) );
  INV_X1 U17657 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20814) );
  NAND4_X1 U17658 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .A4(P1_REIP_REG_12__SCAN_IN), .ZN(n14463) );
  NAND4_X1 U17659 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14462)
         );
  NAND4_X1 U17660 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_17__SCAN_IN), .A4(P1_REIP_REG_16__SCAN_IN), .ZN(n14461) );
  NAND4_X1 U17661 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_20__SCAN_IN), .ZN(n14460)
         );
  NOR4_X1 U17662 ( .A1(n14463), .A2(n14462), .A3(n14461), .A4(n14460), .ZN(
        n14464) );
  NAND2_X1 U17663 ( .A1(n14465), .A2(n14464), .ZN(n16237) );
  NOR2_X1 U17664 ( .A1(n20814), .A2(n16237), .ZN(n16234) );
  NAND2_X1 U17665 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n16234), .ZN(n16227) );
  NOR2_X1 U17666 ( .A1(n20817), .A2(n16227), .ZN(n16222) );
  OAI21_X1 U17667 ( .B1(n16239), .B2(n16222), .A(n16238), .ZN(n16229) );
  NOR2_X1 U17668 ( .A1(n16223), .A2(n16229), .ZN(n14553) );
  NAND3_X1 U17669 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .A3(n14553), .ZN(n14466) );
  NOR2_X1 U17670 ( .A1(n16239), .A2(n14466), .ZN(n14538) );
  NAND2_X1 U17671 ( .A1(n14538), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14526) );
  INV_X1 U17672 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14491) );
  INV_X1 U17673 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20829) );
  NOR2_X1 U17674 ( .A1(n14517), .A2(n20829), .ZN(n14504) );
  NAND2_X1 U17675 ( .A1(n14504), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14468) );
  AND2_X1 U17676 ( .A1(n14468), .A2(n16303), .ZN(n14503) );
  AOI22_X1 U17677 ( .A1(n20354), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20374), .ZN(n14467) );
  OAI21_X1 U17678 ( .B1(n14468), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14467), 
        .ZN(n14469) );
  AOI21_X1 U17679 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(n14503), .A(n14469), 
        .ZN(n14470) );
  OAI211_X1 U17680 ( .C1(n14889), .C2(n20376), .A(n14471), .B(n14470), .ZN(
        P1_U2809) );
  NOR2_X1 U17681 ( .A1(n21063), .A2(n14474), .ZN(n14476) );
  INV_X1 U17682 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n14485) );
  NAND2_X1 U17683 ( .A1(n21062), .A2(DATAI_28_), .ZN(n14484) );
  NAND2_X1 U17684 ( .A1(n14478), .A2(n14477), .ZN(n14479) );
  NOR2_X2 U17685 ( .A1(n21063), .A2(n14479), .ZN(n21065) );
  INV_X1 U17686 ( .A(DATAI_12_), .ZN(n14481) );
  NAND2_X1 U17687 ( .A1(n14482), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14480) );
  OAI21_X1 U17688 ( .B1(n14482), .B2(n14481), .A(n14480), .ZN(n20427) );
  AOI22_X1 U17689 ( .A1(n21065), .A2(n20427), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n21063), .ZN(n14483) );
  OAI211_X1 U17690 ( .C1(n21068), .C2(n14485), .A(n14484), .B(n14483), .ZN(
        n14486) );
  INV_X1 U17691 ( .A(n14486), .ZN(n14487) );
  OAI21_X1 U17692 ( .B1(n14774), .B2(n14717), .A(n14487), .ZN(P1_U2876) );
  AND2_X1 U17693 ( .A1(n14525), .A2(n14488), .ZN(n14489) );
  NOR2_X1 U17694 ( .A1(n14513), .A2(n14489), .ZN(n14935) );
  AOI22_X1 U17695 ( .A1(n14935), .A2(n16315), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14649), .ZN(n14490) );
  OAI21_X1 U17696 ( .B1(n14774), .B2(n14666), .A(n14490), .ZN(P1_U2844) );
  INV_X1 U17697 ( .A(n14776), .ZN(n14495) );
  AOI22_X1 U17698 ( .A1(n20354), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20374), .ZN(n14494) );
  OAI21_X1 U17699 ( .B1(n20329), .B2(n14491), .A(n14526), .ZN(n14492) );
  NAND2_X1 U17700 ( .A1(n14517), .A2(n14492), .ZN(n14493) );
  OAI211_X1 U17701 ( .C1(n20384), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        n14496) );
  AOI21_X1 U17702 ( .B1(n14935), .B2(n20356), .A(n14496), .ZN(n14497) );
  OAI21_X1 U17703 ( .B1(n14774), .B2(n16255), .A(n14497), .ZN(P1_U2812) );
  INV_X1 U17704 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19588) );
  NAND3_X1 U17705 ( .A1(n14499), .A2(n14498), .A3(n14745), .ZN(n14501) );
  AOI22_X1 U17706 ( .A1(n21062), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n21063), .ZN(n14500) );
  OAI211_X1 U17707 ( .C1(n21068), .C2(n19588), .A(n14501), .B(n14500), .ZN(
        P1_U2873) );
  INV_X1 U17708 ( .A(n14502), .ZN(n14755) );
  NAND2_X1 U17709 ( .A1(n14755), .A2(n20348), .ZN(n14509) );
  OAI21_X1 U17710 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14504), .A(n14503), 
        .ZN(n14506) );
  AOI22_X1 U17711 ( .A1(n20354), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20374), .ZN(n14505) );
  NAND2_X1 U17712 ( .A1(n14506), .A2(n14505), .ZN(n14507) );
  AOI21_X1 U17713 ( .B1(n20322), .B2(n14751), .A(n14507), .ZN(n14508) );
  OAI211_X1 U17714 ( .C1(n14917), .C2(n20376), .A(n14509), .B(n14508), .ZN(
        P1_U2810) );
  AOI21_X1 U17715 ( .B1(n14512), .B2(n14511), .A(n14510), .ZN(n14763) );
  INV_X1 U17716 ( .A(n14763), .ZN(n14677) );
  XOR2_X1 U17717 ( .A(n14514), .B(n14513), .Z(n14924) );
  NOR2_X1 U17718 ( .A1(n20384), .A2(n14761), .ZN(n14519) );
  NAND3_X1 U17719 ( .A1(n14517), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n16303), 
        .ZN(n14516) );
  AOI22_X1 U17720 ( .A1(n20354), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20374), .ZN(n14515) );
  OAI211_X1 U17721 ( .C1(n14517), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14516), 
        .B(n14515), .ZN(n14518) );
  AOI211_X1 U17722 ( .C1(n14924), .C2(n20356), .A(n14519), .B(n14518), .ZN(
        n14520) );
  OAI21_X1 U17723 ( .B1(n14677), .B2(n16255), .A(n14520), .ZN(P1_U2811) );
  AOI21_X1 U17724 ( .B1(n14522), .B2(n14521), .A(n14472), .ZN(n14786) );
  NAND2_X1 U17725 ( .A1(n14786), .A2(n20348), .ZN(n14532) );
  NAND2_X1 U17726 ( .A1(n14537), .A2(n14523), .ZN(n14524) );
  AND2_X1 U17727 ( .A1(n14525), .A2(n14524), .ZN(n14942) );
  AOI21_X1 U17728 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n16303), .A(n14538), 
        .ZN(n14529) );
  INV_X1 U17729 ( .A(n14526), .ZN(n14528) );
  AOI22_X1 U17730 ( .A1(n20354), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20374), .ZN(n14527) );
  OAI21_X1 U17731 ( .B1(n14529), .B2(n14528), .A(n14527), .ZN(n14530) );
  AOI21_X1 U17732 ( .B1(n14942), .B2(n20356), .A(n14530), .ZN(n14531) );
  OAI211_X1 U17733 ( .C1(n20384), .C2(n14784), .A(n14532), .B(n14531), .ZN(
        P1_U2813) );
  OAI21_X1 U17734 ( .B1(n14533), .B2(n14534), .A(n14521), .ZN(n14792) );
  NAND2_X1 U17735 ( .A1(n14551), .A2(n14535), .ZN(n14536) );
  NAND2_X1 U17736 ( .A1(n14537), .A2(n14536), .ZN(n14947) );
  AOI22_X1 U17737 ( .A1(n20354), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20374), .ZN(n14544) );
  INV_X1 U17738 ( .A(n14538), .ZN(n14542) );
  NAND3_X1 U17739 ( .A1(n20331), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14553), 
        .ZN(n14540) );
  NAND2_X1 U17740 ( .A1(n16303), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14539) );
  NAND2_X1 U17741 ( .A1(n14540), .A2(n14539), .ZN(n14541) );
  NAND2_X1 U17742 ( .A1(n14542), .A2(n14541), .ZN(n14543) );
  OAI211_X1 U17743 ( .C1(n14947), .C2(n20376), .A(n14544), .B(n14543), .ZN(
        n14545) );
  AOI21_X1 U17744 ( .B1(n14795), .B2(n20322), .A(n14545), .ZN(n14546) );
  OAI21_X1 U17745 ( .B1(n14792), .B2(n16255), .A(n14546), .ZN(P1_U2814) );
  AOI21_X1 U17746 ( .B1(n14548), .B2(n9854), .A(n14533), .ZN(n14803) );
  INV_X1 U17747 ( .A(n14803), .ZN(n14694) );
  INV_X1 U17748 ( .A(n14801), .ZN(n14558) );
  OR2_X1 U17749 ( .A1(n9758), .A2(n14549), .ZN(n14550) );
  AND2_X1 U17750 ( .A1(n14551), .A2(n14550), .ZN(n14961) );
  INV_X1 U17751 ( .A(n14961), .ZN(n14611) );
  INV_X1 U17752 ( .A(n14553), .ZN(n14552) );
  NOR3_X1 U17753 ( .A1(n16239), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14552), 
        .ZN(n14555) );
  INV_X1 U17754 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20820) );
  OAI22_X1 U17755 ( .A1(n20316), .A2(n14250), .B1(n14553), .B2(n20820), .ZN(
        n14554) );
  AOI211_X1 U17756 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n20354), .A(n14555), .B(
        n14554), .ZN(n14556) );
  OAI21_X1 U17757 ( .B1(n14611), .B2(n20376), .A(n14556), .ZN(n14557) );
  AOI21_X1 U17758 ( .B1(n14558), .B2(n20322), .A(n14557), .ZN(n14559) );
  OAI21_X1 U17759 ( .B1(n14694), .B2(n16255), .A(n14559), .ZN(P1_U2815) );
  INV_X1 U17760 ( .A(n14658), .ZN(n14560) );
  AOI21_X1 U17761 ( .B1(n14099), .B2(n14561), .A(n14560), .ZN(n14850) );
  INV_X1 U17762 ( .A(n14850), .ZN(n14667) );
  INV_X1 U17763 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20803) );
  INV_X1 U17764 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20798) );
  NAND2_X1 U17765 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n14562) );
  NAND2_X1 U17766 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n16312), .ZN(n16298) );
  INV_X1 U17767 ( .A(n16253), .ZN(n14565) );
  AND2_X1 U17768 ( .A1(n16303), .A2(n14563), .ZN(n14580) );
  NOR2_X1 U17769 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14563), .ZN(n14578) );
  NOR2_X1 U17770 ( .A1(n14580), .A2(n14578), .ZN(n14564) );
  MUX2_X1 U17771 ( .A(n14565), .B(n14564), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14574) );
  NOR2_X1 U17772 ( .A1(n14567), .A2(n14566), .ZN(n14568) );
  OR2_X1 U17773 ( .A1(n14661), .A2(n14568), .ZN(n16416) );
  INV_X1 U17774 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14665) );
  OAI22_X1 U17775 ( .A1(n16416), .A2(n20376), .B1(n20372), .B2(n14665), .ZN(
        n14569) );
  INV_X1 U17776 ( .A(n14569), .ZN(n14570) );
  OAI211_X1 U17777 ( .C1(n20316), .C2(n14571), .A(n14570), .B(n16489), .ZN(
        n14572) );
  AOI21_X1 U17778 ( .B1(n20322), .B2(n14846), .A(n14572), .ZN(n14573) );
  OAI211_X1 U17779 ( .C1(n14667), .C2(n16255), .A(n14574), .B(n14573), .ZN(
        P1_U2824) );
  INV_X1 U17780 ( .A(n16357), .ZN(n14737) );
  AOI21_X1 U17781 ( .B1(n20374), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16482), .ZN(n14576) );
  AOI22_X1 U17782 ( .A1(n20322), .A2(n16356), .B1(n20354), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14575) );
  OAI211_X1 U17783 ( .C1(n20376), .C2(n16424), .A(n14576), .B(n14575), .ZN(
        n14577) );
  AOI211_X1 U17784 ( .C1(n14580), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14578), 
        .B(n14577), .ZN(n14579) );
  OAI21_X1 U17785 ( .B1(n14737), .B2(n16255), .A(n14579), .ZN(P1_U2825) );
  OAI21_X1 U17786 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14589), .A(n14580), 
        .ZN(n14588) );
  INV_X1 U17787 ( .A(n14860), .ZN(n14586) );
  OAI22_X1 U17788 ( .A1(n16430), .A2(n20376), .B1(n20372), .B2(n14581), .ZN(
        n14582) );
  INV_X1 U17789 ( .A(n14582), .ZN(n14583) );
  OAI211_X1 U17790 ( .C1(n20316), .C2(n14584), .A(n14583), .B(n16489), .ZN(
        n14585) );
  AOI21_X1 U17791 ( .B1(n20322), .B2(n14586), .A(n14585), .ZN(n14587) );
  OAI211_X1 U17792 ( .C1(n14864), .C2(n16255), .A(n14588), .B(n14587), .ZN(
        P1_U2826) );
  INV_X1 U17793 ( .A(n14589), .ZN(n14597) );
  OAI21_X1 U17794 ( .B1(n20329), .B2(n20798), .A(n16298), .ZN(n14596) );
  INV_X1 U17795 ( .A(n16445), .ZN(n14594) );
  NAND2_X1 U17796 ( .A1(n20322), .A2(n14872), .ZN(n14593) );
  OAI21_X1 U17797 ( .B1(n20316), .B2(n14590), .A(n16489), .ZN(n14591) );
  AOI21_X1 U17798 ( .B1(n20354), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14591), .ZN(
        n14592) );
  OAI211_X1 U17799 ( .C1(n14594), .C2(n20376), .A(n14593), .B(n14592), .ZN(
        n14595) );
  AOI21_X1 U17800 ( .B1(n14597), .B2(n14596), .A(n14595), .ZN(n14598) );
  OAI21_X1 U17801 ( .B1(n14875), .B2(n16255), .A(n14598), .ZN(P1_U2827) );
  INV_X1 U17802 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20796) );
  INV_X1 U17803 ( .A(n14599), .ZN(n16304) );
  NOR2_X1 U17804 ( .A1(n20329), .A2(n16304), .ZN(n20324) );
  AOI21_X1 U17805 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n20324), .A(n16482), 
        .ZN(n14601) );
  NAND2_X1 U17806 ( .A1(n20374), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14600) );
  OAI211_X1 U17807 ( .C1(n14602), .C2(n20372), .A(n14601), .B(n14600), .ZN(
        n14603) );
  AOI21_X1 U17808 ( .B1(n16461), .B2(n20356), .A(n14603), .ZN(n14604) );
  OAI21_X1 U17809 ( .B1(n20384), .B2(n14883), .A(n14604), .ZN(n14605) );
  AOI21_X1 U17810 ( .B1(n20796), .B2(n16304), .A(n14605), .ZN(n14606) );
  OAI21_X1 U17811 ( .B1(n14887), .B2(n16255), .A(n14606), .ZN(P1_U2830) );
  INV_X1 U17812 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14607) );
  OAI22_X1 U17813 ( .A1(n14889), .A2(n20385), .B1(n20390), .B2(n14607), .ZN(
        P1_U2841) );
  AOI22_X1 U17814 ( .A1(n14924), .A2(n16315), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14649), .ZN(n14608) );
  OAI21_X1 U17815 ( .B1(n14677), .B2(n14666), .A(n14608), .ZN(P1_U2843) );
  INV_X1 U17816 ( .A(n14786), .ZN(n14683) );
  INV_X1 U17817 ( .A(n14942), .ZN(n14609) );
  OAI222_X1 U17818 ( .A1(n14666), .A2(n14683), .B1(n21016), .B2(n20390), .C1(
        n14609), .C2(n20385), .ZN(P1_U2845) );
  INV_X1 U17819 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14610) );
  OAI222_X1 U17820 ( .A1(n14666), .A2(n14792), .B1(n14610), .B2(n20390), .C1(
        n14947), .C2(n20385), .ZN(P1_U2846) );
  INV_X1 U17821 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14612) );
  OAI222_X1 U17822 ( .A1(n14666), .A2(n14694), .B1(n14612), .B2(n20390), .C1(
        n14611), .C2(n20385), .ZN(P1_U2847) );
  AOI21_X1 U17823 ( .B1(n14614), .B2(n14613), .A(n14547), .ZN(n14811) );
  INV_X1 U17824 ( .A(n14811), .ZN(n16219) );
  INV_X1 U17825 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14617) );
  AND2_X1 U17826 ( .A1(n14624), .A2(n14615), .ZN(n14616) );
  OR2_X1 U17827 ( .A1(n14616), .A2(n9758), .ZN(n16225) );
  OAI222_X1 U17828 ( .A1(n14666), .A2(n16219), .B1(n20390), .B2(n14617), .C1(
        n16225), .C2(n20385), .ZN(P1_U2848) );
  INV_X1 U17829 ( .A(n14618), .ZN(n14620) );
  INV_X1 U17830 ( .A(n14613), .ZN(n14619) );
  AOI21_X1 U17831 ( .B1(n14621), .B2(n14620), .A(n14619), .ZN(n16323) );
  NAND2_X1 U17832 ( .A1(n14633), .A2(n14622), .ZN(n14623) );
  NAND2_X1 U17833 ( .A1(n14624), .A2(n14623), .ZN(n16232) );
  OAI22_X1 U17834 ( .A1(n16232), .A2(n20385), .B1(n14625), .B2(n20390), .ZN(
        n14626) );
  AOI21_X1 U17835 ( .B1(n16323), .B2(n20387), .A(n14626), .ZN(n14627) );
  INV_X1 U17836 ( .A(n14627), .ZN(P1_U2849) );
  NOR2_X1 U17837 ( .A1(n14628), .A2(n14629), .ZN(n14630) );
  OR2_X1 U17838 ( .A1(n14618), .A2(n14630), .ZN(n21071) );
  INV_X1 U17839 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14634) );
  OR2_X1 U17840 ( .A1(n14638), .A2(n14631), .ZN(n14632) );
  NAND2_X1 U17841 ( .A1(n14633), .A2(n14632), .ZN(n16395) );
  OAI222_X1 U17842 ( .A1(n14666), .A2(n21071), .B1(n14634), .B2(n20390), .C1(
        n16395), .C2(n20385), .ZN(P1_U2850) );
  AOI21_X1 U17843 ( .B1(n14635), .B2(n9688), .A(n14628), .ZN(n16329) );
  NOR2_X1 U17844 ( .A1(n14647), .A2(n14636), .ZN(n14637) );
  OR2_X1 U17845 ( .A1(n14638), .A2(n14637), .ZN(n16246) );
  INV_X1 U17846 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14639) );
  OAI22_X1 U17847 ( .A1(n16246), .A2(n20385), .B1(n14639), .B2(n20390), .ZN(
        n14640) );
  AOI21_X1 U17848 ( .B1(n16329), .B2(n20387), .A(n14640), .ZN(n14641) );
  INV_X1 U17849 ( .A(n14641), .ZN(P1_U2851) );
  INV_X1 U17850 ( .A(n14642), .ZN(n14645) );
  INV_X1 U17851 ( .A(n14643), .ZN(n14644) );
  OAI21_X1 U17852 ( .B1(n14645), .B2(n14644), .A(n9688), .ZN(n16256) );
  AOI21_X1 U17853 ( .B1(n10007), .B2(n16271), .A(n14646), .ZN(n14648) );
  OR2_X1 U17854 ( .A1(n14648), .A2(n14647), .ZN(n16254) );
  INV_X1 U17855 ( .A(n16254), .ZN(n16198) );
  AOI22_X1 U17856 ( .A1(n16198), .A2(n16315), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n14649), .ZN(n14650) );
  OAI21_X1 U17857 ( .B1(n16256), .B2(n14666), .A(n14650), .ZN(P1_U2852) );
  INV_X1 U17858 ( .A(n14651), .ZN(n14657) );
  XOR2_X1 U17859 ( .A(n14652), .B(n14657), .Z(n16284) );
  INV_X1 U17860 ( .A(n16284), .ZN(n14656) );
  INV_X1 U17861 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14655) );
  NAND2_X1 U17862 ( .A1(n9760), .A2(n14653), .ZN(n14654) );
  AND2_X1 U17863 ( .A1(n16272), .A2(n14654), .ZN(n16282) );
  INV_X1 U17864 ( .A(n16282), .ZN(n14983) );
  OAI222_X1 U17865 ( .A1(n14656), .A2(n14666), .B1(n14655), .B2(n20390), .C1(
        n14983), .C2(n20385), .ZN(P1_U2854) );
  AOI21_X1 U17866 ( .B1(n14659), .B2(n14658), .A(n14651), .ZN(n16349) );
  OR2_X1 U17867 ( .A1(n14661), .A2(n14660), .ZN(n14662) );
  NAND2_X1 U17868 ( .A1(n9760), .A2(n14662), .ZN(n16408) );
  INV_X1 U17869 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16288) );
  OAI22_X1 U17870 ( .A1(n16408), .A2(n20385), .B1(n16288), .B2(n20390), .ZN(
        n14663) );
  AOI21_X1 U17871 ( .B1(n16349), .B2(n20387), .A(n14663), .ZN(n14664) );
  INV_X1 U17872 ( .A(n14664), .ZN(P1_U2855) );
  OAI222_X1 U17873 ( .A1(n14667), .A2(n14666), .B1(n14665), .B2(n20390), .C1(
        n16416), .C2(n20385), .ZN(P1_U2856) );
  INV_X1 U17874 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U17875 ( .A1(n21062), .A2(DATAI_30_), .ZN(n14669) );
  AOI22_X1 U17876 ( .A1(n21065), .A2(n20431), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n21063), .ZN(n14668) );
  OAI211_X1 U17877 ( .C1(n21068), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14671) );
  INV_X1 U17878 ( .A(n14671), .ZN(n14672) );
  OAI21_X1 U17879 ( .B1(n14502), .B2(n14717), .A(n14672), .ZN(P1_U2874) );
  INV_X1 U17880 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16852) );
  NAND2_X1 U17881 ( .A1(n21062), .A2(DATAI_29_), .ZN(n14674) );
  AOI22_X1 U17882 ( .A1(n21065), .A2(n20429), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n21063), .ZN(n14673) );
  OAI211_X1 U17883 ( .C1(n21068), .C2(n16852), .A(n14674), .B(n14673), .ZN(
        n14675) );
  INV_X1 U17884 ( .A(n14675), .ZN(n14676) );
  OAI21_X1 U17885 ( .B1(n14677), .B2(n14717), .A(n14676), .ZN(P1_U2875) );
  INV_X1 U17886 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14680) );
  NAND2_X1 U17887 ( .A1(n21062), .A2(DATAI_27_), .ZN(n14679) );
  AOI22_X1 U17888 ( .A1(n21065), .A2(n20425), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n21063), .ZN(n14678) );
  OAI211_X1 U17889 ( .C1(n21068), .C2(n14680), .A(n14679), .B(n14678), .ZN(
        n14681) );
  INV_X1 U17890 ( .A(n14681), .ZN(n14682) );
  OAI21_X1 U17891 ( .B1(n14683), .B2(n14717), .A(n14682), .ZN(P1_U2877) );
  INV_X1 U17892 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n14686) );
  NAND2_X1 U17893 ( .A1(n21062), .A2(DATAI_26_), .ZN(n14685) );
  AOI22_X1 U17894 ( .A1(n21065), .A2(n20423), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n21063), .ZN(n14684) );
  OAI211_X1 U17895 ( .C1(n21068), .C2(n14686), .A(n14685), .B(n14684), .ZN(
        n14687) );
  INV_X1 U17896 ( .A(n14687), .ZN(n14688) );
  OAI21_X1 U17897 ( .B1(n14792), .B2(n14717), .A(n14688), .ZN(P1_U2878) );
  INV_X1 U17898 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14691) );
  NAND2_X1 U17899 ( .A1(n21062), .A2(DATAI_25_), .ZN(n14690) );
  AOI22_X1 U17900 ( .A1(n21065), .A2(n20421), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n21063), .ZN(n14689) );
  OAI211_X1 U17901 ( .C1(n21068), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        n14692) );
  INV_X1 U17902 ( .A(n14692), .ZN(n14693) );
  OAI21_X1 U17903 ( .B1(n14694), .B2(n14717), .A(n14693), .ZN(P1_U2879) );
  INV_X1 U17904 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14697) );
  NAND2_X1 U17905 ( .A1(n21062), .A2(DATAI_24_), .ZN(n14696) );
  AOI22_X1 U17906 ( .A1(n21065), .A2(n20419), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n21063), .ZN(n14695) );
  OAI211_X1 U17907 ( .C1(n21068), .C2(n14697), .A(n14696), .B(n14695), .ZN(
        n14698) );
  INV_X1 U17908 ( .A(n14698), .ZN(n14699) );
  OAI21_X1 U17909 ( .B1(n16219), .B2(n14717), .A(n14699), .ZN(P1_U2880) );
  INV_X1 U17910 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14703) );
  NAND2_X1 U17911 ( .A1(n21062), .A2(DATAI_23_), .ZN(n14702) );
  AOI22_X1 U17912 ( .A1(n21065), .A2(n14700), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n21063), .ZN(n14701) );
  OAI211_X1 U17913 ( .C1(n14703), .C2(n21068), .A(n14702), .B(n14701), .ZN(
        n14704) );
  AOI21_X1 U17914 ( .B1(n16323), .B2(n16319), .A(n14704), .ZN(n14705) );
  INV_X1 U17915 ( .A(n14705), .ZN(P1_U2881) );
  NAND2_X1 U17916 ( .A1(n21062), .A2(DATAI_21_), .ZN(n14708) );
  AOI22_X1 U17917 ( .A1(n21065), .A2(n14706), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n21063), .ZN(n14707) );
  OAI211_X1 U17918 ( .C1(n16861), .C2(n21068), .A(n14708), .B(n14707), .ZN(
        n14709) );
  AOI21_X1 U17919 ( .B1(n16329), .B2(n16319), .A(n14709), .ZN(n14710) );
  INV_X1 U17920 ( .A(n14710), .ZN(P1_U2883) );
  INV_X1 U17921 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14714) );
  NAND2_X1 U17922 ( .A1(n21062), .A2(DATAI_20_), .ZN(n14713) );
  AOI22_X1 U17923 ( .A1(n21065), .A2(n14711), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n21063), .ZN(n14712) );
  OAI211_X1 U17924 ( .C1(n14714), .C2(n21068), .A(n14713), .B(n14712), .ZN(
        n14715) );
  INV_X1 U17925 ( .A(n14715), .ZN(n14716) );
  OAI21_X1 U17926 ( .B1(n16256), .B2(n14717), .A(n14716), .ZN(P1_U2884) );
  INV_X1 U17927 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14721) );
  NAND2_X1 U17928 ( .A1(n21062), .A2(DATAI_18_), .ZN(n14720) );
  AOI22_X1 U17929 ( .A1(n21065), .A2(n14718), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n21063), .ZN(n14719) );
  OAI211_X1 U17930 ( .C1(n14721), .C2(n21068), .A(n14720), .B(n14719), .ZN(
        n14722) );
  AOI21_X1 U17931 ( .B1(n16284), .B2(n16319), .A(n14722), .ZN(n14723) );
  INV_X1 U17932 ( .A(n14723), .ZN(P1_U2886) );
  INV_X1 U17933 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14727) );
  NAND2_X1 U17934 ( .A1(n21062), .A2(DATAI_17_), .ZN(n14726) );
  AOI22_X1 U17935 ( .A1(n21065), .A2(n14724), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n21063), .ZN(n14725) );
  OAI211_X1 U17936 ( .C1(n14727), .C2(n21068), .A(n14726), .B(n14725), .ZN(
        n14728) );
  AOI21_X1 U17937 ( .B1(n16349), .B2(n16319), .A(n14728), .ZN(n14729) );
  INV_X1 U17938 ( .A(n14729), .ZN(P1_U2887) );
  NAND2_X1 U17939 ( .A1(n21062), .A2(DATAI_16_), .ZN(n14732) );
  AOI22_X1 U17940 ( .A1(n21065), .A2(n14730), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n21063), .ZN(n14731) );
  OAI211_X1 U17941 ( .C1(n14733), .C2(n21068), .A(n14732), .B(n14731), .ZN(
        n14734) );
  AOI21_X1 U17942 ( .B1(n14850), .B2(n16319), .A(n14734), .ZN(n14735) );
  INV_X1 U17943 ( .A(n14735), .ZN(P1_U2888) );
  OAI222_X1 U17944 ( .A1(n14737), .A2(n14717), .B1(n14745), .B2(n12397), .C1(
        n14744), .C2(n14736), .ZN(P1_U2889) );
  INV_X1 U17945 ( .A(n14738), .ZN(n14742) );
  INV_X1 U17946 ( .A(n14739), .ZN(n14741) );
  INV_X1 U17947 ( .A(n16363), .ZN(n14747) );
  INV_X1 U17948 ( .A(n20427), .ZN(n14743) );
  OAI222_X1 U17949 ( .A1(n14747), .A2(n14717), .B1(n14746), .B2(n14745), .C1(
        n14744), .C2(n14743), .ZN(P1_U2892) );
  NOR2_X1 U17950 ( .A1(n14749), .A2(n14748), .ZN(n14750) );
  NAND2_X1 U17951 ( .A1(n14751), .A2(n16365), .ZN(n14752) );
  NAND2_X1 U17952 ( .A1(n16482), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14915) );
  OAI211_X1 U17953 ( .C1(n16333), .C2(n14753), .A(n14752), .B(n14915), .ZN(
        n14754) );
  OAI21_X1 U17954 ( .B1(n9721), .B2(n20299), .A(n14756), .ZN(P1_U2969) );
  NAND2_X1 U17955 ( .A1(n14758), .A2(n14757), .ZN(n14759) );
  XNOR2_X1 U17956 ( .A(n14759), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14929) );
  NOR2_X1 U17957 ( .A1(n16489), .A2(n20829), .ZN(n14923) );
  AOI21_X1 U17958 ( .B1(n20450), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14923), .ZN(n14760) );
  OAI21_X1 U17959 ( .B1(n14761), .B2(n20461), .A(n14760), .ZN(n14762) );
  AOI21_X1 U17960 ( .B1(n14763), .B2(n20456), .A(n14762), .ZN(n14764) );
  OAI21_X1 U17961 ( .B1(n14929), .B2(n20299), .A(n14764), .ZN(P1_U2970) );
  NAND3_X1 U17962 ( .A1(n14877), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14771) );
  NOR4_X1 U17963 ( .A1(n14765), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U17964 ( .A1(n10206), .A2(n14766), .ZN(n14770) );
  INV_X1 U17965 ( .A(n14949), .ZN(n14768) );
  OAI21_X1 U17966 ( .B1(n10206), .B2(n14768), .A(n14767), .ZN(n14769) );
  MUX2_X1 U17967 ( .A(n14771), .B(n14770), .S(n14769), .Z(n14772) );
  XOR2_X1 U17968 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14772), .Z(
        n14938) );
  NAND2_X1 U17969 ( .A1(n16482), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14930) );
  OAI21_X1 U17970 ( .B1(n16333), .B2(n14773), .A(n14930), .ZN(n14775) );
  INV_X1 U17971 ( .A(n14777), .ZN(n14778) );
  NAND2_X1 U17972 ( .A1(n14779), .A2(n14778), .ZN(n14780) );
  MUX2_X1 U17973 ( .A(n14781), .B(n14780), .S(n14877), .Z(n14782) );
  XOR2_X1 U17974 ( .A(n14782), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(
        n14946) );
  INV_X1 U17975 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20824) );
  NOR2_X1 U17976 ( .A1(n16489), .A2(n20824), .ZN(n14941) );
  AOI21_X1 U17977 ( .B1(n20450), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14941), .ZN(n14783) );
  OAI21_X1 U17978 ( .B1(n14784), .B2(n20461), .A(n14783), .ZN(n14785) );
  AOI21_X1 U17979 ( .B1(n14786), .B2(n20456), .A(n14785), .ZN(n14787) );
  OAI21_X1 U17980 ( .B1(n20299), .B2(n14946), .A(n14787), .ZN(P1_U2972) );
  INV_X1 U17981 ( .A(n14767), .ZN(n14805) );
  OAI21_X1 U17982 ( .B1(n14805), .B2(n14949), .A(n14877), .ZN(n14788) );
  NAND2_X1 U17983 ( .A1(n14789), .A2(n14788), .ZN(n14790) );
  XOR2_X1 U17984 ( .A(n14790), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(
        n14958) );
  NAND2_X1 U17985 ( .A1(n16482), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14948) );
  OAI21_X1 U17986 ( .B1(n16333), .B2(n14791), .A(n14948), .ZN(n14794) );
  NOR2_X1 U17987 ( .A1(n14792), .A2(n14888), .ZN(n14793) );
  AOI211_X1 U17988 ( .C1(n16365), .C2(n14795), .A(n14794), .B(n14793), .ZN(
        n14796) );
  OAI21_X1 U17989 ( .B1(n20299), .B2(n14958), .A(n14796), .ZN(P1_U2973) );
  NAND2_X1 U17990 ( .A1(n14797), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14808) );
  MUX2_X1 U17991 ( .A(n9748), .B(n14809), .S(n14877), .Z(n14798) );
  AOI21_X1 U17992 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14808), .A(
        n14798), .ZN(n14799) );
  XNOR2_X1 U17993 ( .A(n14799), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14965) );
  NOR2_X1 U17994 ( .A1(n16489), .A2(n20820), .ZN(n14960) );
  AOI21_X1 U17995 ( .B1(n20450), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14960), .ZN(n14800) );
  OAI21_X1 U17996 ( .B1(n14801), .B2(n20461), .A(n14800), .ZN(n14802) );
  AOI21_X1 U17997 ( .B1(n14803), .B2(n20456), .A(n14802), .ZN(n14804) );
  OAI21_X1 U17998 ( .B1(n20299), .B2(n14965), .A(n14804), .ZN(P1_U2974) );
  NAND2_X1 U17999 ( .A1(n14805), .A2(n14808), .ZN(n14807) );
  MUX2_X1 U18000 ( .A(n14808), .B(n14807), .S(n10206), .Z(n14810) );
  XNOR2_X1 U18001 ( .A(n14810), .B(n14809), .ZN(n14973) );
  NAND2_X1 U18002 ( .A1(n14811), .A2(n20456), .ZN(n14815) );
  INV_X1 U18003 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14812) );
  NOR2_X1 U18004 ( .A1(n16489), .A2(n14812), .ZN(n14967) );
  INV_X1 U18005 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16218) );
  NOR2_X1 U18006 ( .A1(n16333), .A2(n16218), .ZN(n14813) );
  AOI211_X1 U18007 ( .C1(n16215), .C2(n16365), .A(n14967), .B(n14813), .ZN(
        n14814) );
  OAI211_X1 U18008 ( .C1(n14973), .C2(n20299), .A(n14815), .B(n14814), .ZN(
        P1_U2975) );
  NAND2_X1 U18009 ( .A1(n14817), .A2(n14816), .ZN(n14818) );
  XOR2_X1 U18010 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14818), .Z(
        n16394) );
  INV_X1 U18011 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14819) );
  OAI22_X1 U18012 ( .A1(n16333), .A2(n13002), .B1(n16489), .B2(n14819), .ZN(
        n14821) );
  NOR2_X1 U18013 ( .A1(n21071), .A2(n14888), .ZN(n14820) );
  AOI211_X1 U18014 ( .C1(n16365), .C2(n16235), .A(n14821), .B(n14820), .ZN(
        n14822) );
  OAI21_X1 U18015 ( .B1(n20299), .B2(n16394), .A(n14822), .ZN(P1_U2977) );
  INV_X1 U18016 ( .A(n14823), .ZN(n14824) );
  NAND3_X1 U18017 ( .A1(n14824), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14877), .ZN(n16179) );
  INV_X1 U18018 ( .A(n14833), .ZN(n14826) );
  INV_X1 U18019 ( .A(n16335), .ZN(n14825) );
  NAND3_X1 U18020 ( .A1(n14826), .A2(n14825), .A3(n14392), .ZN(n16177) );
  NAND2_X1 U18021 ( .A1(n16179), .A2(n16177), .ZN(n14827) );
  XNOR2_X1 U18022 ( .A(n14827), .B(n16178), .ZN(n16199) );
  NAND2_X1 U18023 ( .A1(n16199), .A2(n20457), .ZN(n14831) );
  INV_X1 U18024 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14828) );
  OAI22_X1 U18025 ( .A1(n16333), .A2(n16261), .B1(n16489), .B2(n14828), .ZN(
        n14829) );
  AOI21_X1 U18026 ( .B1(n16365), .B2(n16252), .A(n14829), .ZN(n14830) );
  OAI211_X1 U18027 ( .C1(n14888), .C2(n16256), .A(n14831), .B(n14830), .ZN(
        P1_U2979) );
  OAI21_X1 U18028 ( .B1(n14833), .B2(n14832), .A(n14823), .ZN(n14994) );
  NAND2_X1 U18029 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14834) );
  NAND2_X1 U18030 ( .A1(n16482), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14982) );
  OAI211_X1 U18031 ( .C1(n16277), .C2(n20461), .A(n14834), .B(n14982), .ZN(
        n14835) );
  AOI21_X1 U18032 ( .B1(n16284), .B2(n20456), .A(n14835), .ZN(n14836) );
  OAI21_X1 U18033 ( .B1(n20299), .B2(n14994), .A(n14836), .ZN(P1_U2981) );
  INV_X1 U18034 ( .A(n14837), .ZN(n14876) );
  INV_X1 U18035 ( .A(n14838), .ZN(n14840) );
  AOI21_X1 U18036 ( .B1(n14876), .B2(n14840), .A(n14839), .ZN(n16354) );
  INV_X1 U18037 ( .A(n14843), .ZN(n14841) );
  NOR2_X1 U18038 ( .A1(n14842), .A2(n14841), .ZN(n16353) );
  NAND2_X1 U18039 ( .A1(n16354), .A2(n16353), .ZN(n16352) );
  NAND2_X1 U18040 ( .A1(n16352), .A2(n14843), .ZN(n14844) );
  XOR2_X1 U18041 ( .A(n14845), .B(n14844), .Z(n16415) );
  INV_X1 U18042 ( .A(n14846), .ZN(n14848) );
  AOI22_X1 U18043 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14847) );
  OAI21_X1 U18044 ( .B1(n14848), .B2(n20461), .A(n14847), .ZN(n14849) );
  AOI21_X1 U18045 ( .B1(n14850), .B2(n20456), .A(n14849), .ZN(n14851) );
  OAI21_X1 U18046 ( .B1(n16415), .B2(n20299), .A(n14851), .ZN(P1_U2983) );
  NAND2_X1 U18047 ( .A1(n14837), .A2(n14852), .ZN(n16344) );
  NAND2_X1 U18048 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14853) );
  AND2_X1 U18049 ( .A1(n14877), .A2(n14853), .ZN(n14866) );
  INV_X1 U18050 ( .A(n14866), .ZN(n14854) );
  NAND3_X1 U18051 ( .A1(n16344), .A2(n14855), .A3(n14854), .ZN(n14857) );
  NAND2_X1 U18052 ( .A1(n14857), .A2(n14856), .ZN(n14859) );
  XNOR2_X1 U18053 ( .A(n10206), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14858) );
  XNOR2_X1 U18054 ( .A(n14859), .B(n14858), .ZN(n16435) );
  NAND2_X1 U18055 ( .A1(n16435), .A2(n20457), .ZN(n14863) );
  AND2_X1 U18056 ( .A1(n16482), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16431) );
  NOR2_X1 U18057 ( .A1(n20461), .A2(n14860), .ZN(n14861) );
  AOI211_X1 U18058 ( .C1(n20450), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16431), .B(n14861), .ZN(n14862) );
  OAI211_X1 U18059 ( .C1(n14888), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        P1_U2985) );
  OAI22_X1 U18060 ( .A1(n14837), .A2(n14866), .B1(n14865), .B2(n14877), .ZN(
        n16361) );
  INV_X1 U18061 ( .A(n14868), .ZN(n14867) );
  OAI21_X1 U18062 ( .B1(n16453), .B2(n14877), .A(n14867), .ZN(n16362) );
  NOR2_X1 U18063 ( .A1(n16361), .A2(n16362), .ZN(n16360) );
  NOR2_X1 U18064 ( .A1(n16360), .A2(n14868), .ZN(n14870) );
  XNOR2_X1 U18065 ( .A(n14870), .B(n14869), .ZN(n16444) );
  NAND2_X1 U18066 ( .A1(n16444), .A2(n20457), .ZN(n14874) );
  OAI22_X1 U18067 ( .A1(n16333), .A2(n14590), .B1(n16489), .B2(n20798), .ZN(
        n14871) );
  AOI21_X1 U18068 ( .B1(n16365), .B2(n14872), .A(n14871), .ZN(n14873) );
  OAI211_X1 U18069 ( .C1(n14888), .C2(n14875), .A(n14874), .B(n14873), .ZN(
        P1_U2986) );
  NAND2_X1 U18070 ( .A1(n14880), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14879) );
  XNOR2_X1 U18071 ( .A(n14876), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14878) );
  MUX2_X1 U18072 ( .A(n14879), .B(n14878), .S(n14877), .Z(n14882) );
  INV_X1 U18073 ( .A(n14880), .ZN(n14881) );
  NAND3_X1 U18074 ( .A1(n14881), .A2(n10206), .A3(n14995), .ZN(n14997) );
  NAND2_X1 U18075 ( .A1(n14882), .A2(n14997), .ZN(n16462) );
  NAND2_X1 U18076 ( .A1(n16462), .A2(n20457), .ZN(n14886) );
  AND2_X1 U18077 ( .A1(n16482), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16460) );
  NOR2_X1 U18078 ( .A1(n20461), .A2(n14883), .ZN(n14884) );
  AOI211_X1 U18079 ( .C1(n20450), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16460), .B(n14884), .ZN(n14885) );
  OAI211_X1 U18080 ( .C1(n14888), .C2(n14887), .A(n14886), .B(n14885), .ZN(
        P1_U2989) );
  INV_X1 U18081 ( .A(n14889), .ZN(n14895) );
  INV_X1 U18082 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16413) );
  NAND3_X1 U18083 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n14890), .ZN(n15001) );
  NOR2_X1 U18084 ( .A1(n13806), .A2(n15001), .ZN(n16454) );
  NAND2_X1 U18085 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16454), .ZN(
        n14984) );
  NOR2_X1 U18086 ( .A1(n14985), .A2(n14984), .ZN(n16441) );
  INV_X1 U18087 ( .A(n20493), .ZN(n14891) );
  NOR2_X1 U18088 ( .A1(n14984), .A2(n15000), .ZN(n16440) );
  AOI22_X1 U18089 ( .A1(n20484), .A2(n16441), .B1(n14891), .B2(n16440), .ZN(
        n16449) );
  INV_X1 U18090 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16438) );
  NAND3_X1 U18091 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n16427), .ZN(n16412) );
  NOR2_X1 U18092 ( .A1(n16413), .A2(n16412), .ZN(n14992) );
  NAND2_X1 U18093 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14992), .ZN(
        n16407) );
  AND2_X1 U18094 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16401) );
  NAND2_X1 U18095 ( .A1(n16390), .A2(n16401), .ZN(n14975) );
  NOR3_X1 U18096 ( .A1(n14975), .A2(n20885), .A3(n14949), .ZN(n14920) );
  NAND3_X1 U18097 ( .A1(n14920), .A2(n14932), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14912) );
  INV_X1 U18098 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14892) );
  NOR3_X1 U18099 ( .A1(n14912), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14892), .ZN(n14894) );
  AOI211_X1 U18100 ( .C1(n14895), .C2(n20481), .A(n14894), .B(n14893), .ZN(
        n14910) );
  INV_X1 U18101 ( .A(n14932), .ZN(n14921) );
  NAND3_X1 U18102 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14988) );
  NOR4_X1 U18103 ( .A1(n14991), .A2(n16448), .A3(n16438), .A4(n14988), .ZN(
        n14898) );
  OAI221_X1 U18104 ( .B1(n16440), .B2(n16473), .C1(n14898), .C2(n16473), .A(
        n20487), .ZN(n14896) );
  INV_X1 U18105 ( .A(n14896), .ZN(n14897) );
  OAI221_X1 U18106 ( .B1(n20498), .B2(n16441), .C1(n20498), .C2(n14898), .A(
        n14897), .ZN(n16402) );
  NAND2_X1 U18107 ( .A1(n16476), .A2(n20487), .ZN(n14899) );
  OAI21_X1 U18108 ( .B1(n16197), .B2(n16402), .A(n14899), .ZN(n16391) );
  INV_X1 U18109 ( .A(n16401), .ZN(n14900) );
  NAND2_X1 U18110 ( .A1(n20499), .A2(n14900), .ZN(n14901) );
  INV_X1 U18111 ( .A(n14902), .ZN(n14903) );
  NAND2_X1 U18112 ( .A1(n14903), .A2(n14949), .ZN(n14904) );
  OAI211_X1 U18113 ( .C1(n14954), .C2(n20507), .A(n14981), .B(n14904), .ZN(
        n14962) );
  NOR2_X1 U18114 ( .A1(n14962), .A2(n20499), .ZN(n14905) );
  INV_X1 U18115 ( .A(n14905), .ZN(n14908) );
  INV_X1 U18116 ( .A(n14962), .ZN(n14907) );
  NOR2_X1 U18117 ( .A1(n20885), .A2(n14953), .ZN(n14906) );
  AOI21_X1 U18118 ( .B1(n14907), .B2(n14906), .A(n14905), .ZN(n14943) );
  AOI21_X1 U18119 ( .B1(n14921), .B2(n14908), .A(n14943), .ZN(n14925) );
  OAI211_X1 U18120 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16476), .A(
        n14925), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14913) );
  NAND3_X1 U18121 ( .A1(n14913), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14908), .ZN(n14909) );
  OAI211_X1 U18122 ( .C1(n14911), .C2(n16457), .A(n14910), .B(n14909), .ZN(
        P1_U3000) );
  INV_X1 U18123 ( .A(n14912), .ZN(n14914) );
  OAI21_X1 U18124 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14914), .A(
        n14913), .ZN(n14916) );
  OAI211_X1 U18125 ( .C1(n14917), .C2(n20503), .A(n14916), .B(n14915), .ZN(
        n14918) );
  INV_X1 U18126 ( .A(n14918), .ZN(n14919) );
  OAI21_X1 U18127 ( .B1(n9721), .B2(n16457), .A(n14919), .ZN(P1_U3001) );
  INV_X1 U18128 ( .A(n14920), .ZN(n14939) );
  NOR3_X1 U18129 ( .A1(n14939), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14921), .ZN(n14922) );
  AOI211_X1 U18130 ( .C1(n14924), .C2(n20481), .A(n14923), .B(n14922), .ZN(
        n14928) );
  INV_X1 U18131 ( .A(n14925), .ZN(n14926) );
  NAND2_X1 U18132 ( .A1(n14926), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14927) );
  OAI211_X1 U18133 ( .C1(n14929), .C2(n16457), .A(n14928), .B(n14927), .ZN(
        P1_U3002) );
  INV_X1 U18134 ( .A(n14930), .ZN(n14934) );
  NOR3_X1 U18135 ( .A1(n14939), .A2(n14932), .A3(n14931), .ZN(n14933) );
  AOI211_X1 U18136 ( .C1(n14935), .C2(n20481), .A(n14934), .B(n14933), .ZN(
        n14937) );
  NAND2_X1 U18137 ( .A1(n14943), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14936) );
  OAI211_X1 U18138 ( .C1(n14938), .C2(n16457), .A(n14937), .B(n14936), .ZN(
        P1_U3003) );
  NOR2_X1 U18139 ( .A1(n14939), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14940) );
  AOI211_X1 U18140 ( .C1(n14942), .C2(n20481), .A(n14941), .B(n14940), .ZN(
        n14945) );
  NAND2_X1 U18141 ( .A1(n14943), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14944) );
  OAI211_X1 U18142 ( .C1(n14946), .C2(n16457), .A(n14945), .B(n14944), .ZN(
        P1_U3004) );
  INV_X1 U18143 ( .A(n14947), .ZN(n14952) );
  INV_X1 U18144 ( .A(n14948), .ZN(n14951) );
  NOR3_X1 U18145 ( .A1(n14975), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14949), .ZN(n14950) );
  AOI211_X1 U18146 ( .C1(n14952), .C2(n20481), .A(n14951), .B(n14950), .ZN(
        n14957) );
  NAND2_X1 U18147 ( .A1(n14954), .A2(n14953), .ZN(n14955) );
  NOR2_X1 U18148 ( .A1(n14975), .A2(n14955), .ZN(n14959) );
  OAI21_X1 U18149 ( .B1(n14962), .B2(n14959), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14956) );
  OAI211_X1 U18150 ( .C1(n14958), .C2(n16457), .A(n14957), .B(n14956), .ZN(
        P1_U3005) );
  AOI211_X1 U18151 ( .C1(n14961), .C2(n20481), .A(n14960), .B(n14959), .ZN(
        n14964) );
  NAND2_X1 U18152 ( .A1(n14962), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14963) );
  OAI211_X1 U18153 ( .C1(n14965), .C2(n16457), .A(n14964), .B(n14963), .ZN(
        P1_U3006) );
  INV_X1 U18154 ( .A(n16225), .ZN(n14968) );
  NOR3_X1 U18155 ( .A1(n14975), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14980), .ZN(n14966) );
  AOI211_X1 U18156 ( .C1(n14968), .C2(n20481), .A(n14967), .B(n14966), .ZN(
        n14972) );
  INV_X1 U18157 ( .A(n14981), .ZN(n14970) );
  AOI21_X1 U18158 ( .B1(n20493), .B2(n20498), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14969) );
  OAI21_X1 U18159 ( .B1(n14970), .B2(n14969), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14971) );
  OAI211_X1 U18160 ( .C1(n14973), .C2(n16457), .A(n14972), .B(n14971), .ZN(
        P1_U3007) );
  XNOR2_X1 U18161 ( .A(n14877), .B(n14980), .ZN(n14974) );
  XNOR2_X1 U18162 ( .A(n14767), .B(n14974), .ZN(n16322) );
  NAND2_X1 U18163 ( .A1(n16322), .A2(n20509), .ZN(n14979) );
  INV_X1 U18164 ( .A(n16232), .ZN(n14977) );
  OAI22_X1 U18165 ( .A1(n16489), .A2(n20817), .B1(n14975), .B2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14976) );
  AOI21_X1 U18166 ( .B1(n14977), .B2(n20481), .A(n14976), .ZN(n14978) );
  OAI211_X1 U18167 ( .C1(n14981), .C2(n14980), .A(n14979), .B(n14978), .ZN(
        P1_U3008) );
  OAI21_X1 U18168 ( .B1(n14983), .B2(n20503), .A(n14982), .ZN(n14990) );
  OR2_X1 U18169 ( .A1(n16448), .A2(n14984), .ZN(n16433) );
  AOI21_X1 U18170 ( .B1(n20484), .B2(n14985), .A(n16443), .ZN(n16472) );
  OAI21_X1 U18171 ( .B1(n16473), .B2(n14986), .A(n16472), .ZN(n14987) );
  AOI21_X1 U18172 ( .B1(n20499), .B2(n16433), .A(n14987), .ZN(n16439) );
  OAI21_X1 U18173 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16476), .A(
        n16439), .ZN(n16426) );
  AOI21_X1 U18174 ( .B1(n20499), .B2(n14988), .A(n16426), .ZN(n16414) );
  NOR2_X1 U18175 ( .A1(n16414), .A2(n14991), .ZN(n14989) );
  AOI211_X1 U18176 ( .C1(n14992), .C2(n14991), .A(n14990), .B(n14989), .ZN(
        n14993) );
  OAI21_X1 U18177 ( .B1(n14994), .B2(n16457), .A(n14993), .ZN(P1_U3013) );
  OR3_X1 U18178 ( .A1(n14837), .A2(n10206), .A3(n14995), .ZN(n14996) );
  NAND2_X1 U18179 ( .A1(n14997), .A2(n14996), .ZN(n14998) );
  XNOR2_X1 U18180 ( .A(n14998), .B(n13806), .ZN(n16369) );
  NAND2_X1 U18181 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16459) );
  NOR2_X1 U18182 ( .A1(n16459), .A2(n16467), .ZN(n15003) );
  OAI21_X1 U18183 ( .B1(n16454), .B2(n20498), .A(n16472), .ZN(n14999) );
  AOI221_X1 U18184 ( .B1(n15001), .B2(n20483), .C1(n15000), .C2(n20483), .A(
        n14999), .ZN(n16450) );
  INV_X1 U18185 ( .A(n16450), .ZN(n15002) );
  MUX2_X1 U18186 ( .A(n15003), .B(n15002), .S(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(n15006) );
  INV_X1 U18187 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15004) );
  OAI22_X1 U18188 ( .A1(n16306), .A2(n20503), .B1(n16489), .B2(n15004), .ZN(
        n15005) );
  AOI211_X1 U18189 ( .C1(n16369), .C2(n20509), .A(n15006), .B(n15005), .ZN(
        n15007) );
  INV_X1 U18190 ( .A(n15007), .ZN(P1_U3020) );
  OAI211_X1 U18191 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n15009), .A(n15008), 
        .B(n20622), .ZN(n15010) );
  OAI21_X1 U18192 ( .B1(n20591), .B2(n15017), .A(n15010), .ZN(n15011) );
  MUX2_X1 U18193 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15011), .S(
        n20515), .Z(P1_U3477) );
  INV_X1 U18194 ( .A(n12677), .ZN(n15018) );
  INV_X1 U18195 ( .A(n15012), .ZN(n15015) );
  OAI21_X1 U18196 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15016) );
  OAI21_X1 U18197 ( .B1(n15018), .B2(n15017), .A(n15016), .ZN(n15019) );
  MUX2_X1 U18198 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15019), .S(
        n20515), .Z(P1_U3475) );
  INV_X1 U18199 ( .A(n15020), .ZN(n15024) );
  INV_X1 U18200 ( .A(n15021), .ZN(n15023) );
  AOI22_X1 U18201 ( .A1(n15024), .A2(n16172), .B1(n15023), .B2(n15022), .ZN(
        n15025) );
  OAI21_X1 U18202 ( .B1(n15026), .B2(n15030), .A(n15025), .ZN(n15027) );
  MUX2_X1 U18203 ( .A(n15027), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15032), .Z(P1_U3472) );
  OAI22_X1 U18204 ( .A1(n15031), .A2(n15030), .B1(n15029), .B2(n15028), .ZN(
        n15033) );
  MUX2_X1 U18205 ( .A(n15033), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15032), .Z(P1_U3469) );
  NAND2_X1 U18206 ( .A1(n20675), .A2(n20623), .ZN(n15047) );
  OR2_X1 U18207 ( .A1(n20585), .A2(n20651), .ZN(n15036) );
  INV_X1 U18208 ( .A(n15036), .ZN(n15073) );
  OR2_X1 U18209 ( .A1(n20650), .A2(n20521), .ZN(n15037) );
  OAI21_X1 U18210 ( .B1(n20675), .B2(n15075), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15038) );
  NAND2_X1 U18211 ( .A1(n15040), .A2(n15038), .ZN(n15039) );
  AOI22_X1 U18212 ( .A1(n20701), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__0__SCAN_IN), .B2(n15072), .ZN(n15046) );
  OR2_X1 U18213 ( .A1(n15040), .A2(n20703), .ZN(n15043) );
  NAND2_X1 U18214 ( .A1(n15041), .A2(n20529), .ZN(n15042) );
  NAND2_X1 U18215 ( .A1(n15043), .A2(n15042), .ZN(n15074) );
  NAND2_X1 U18216 ( .A1(n15074), .A2(n20700), .ZN(n15045) );
  NAND2_X1 U18217 ( .A1(n15075), .A2(n20708), .ZN(n15044) );
  NAND4_X1 U18218 ( .A1(n15047), .A2(n15046), .A3(n15045), .A4(n15044), .ZN(
        P1_U3097) );
  NAND2_X1 U18219 ( .A1(n20675), .A2(n20661), .ZN(n15051) );
  AOI22_X1 U18220 ( .A1(n20713), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n15072), .ZN(n15050) );
  NAND2_X1 U18221 ( .A1(n15074), .A2(n20712), .ZN(n15049) );
  NAND2_X1 U18222 ( .A1(n15075), .A2(n20714), .ZN(n15048) );
  NAND4_X1 U18223 ( .A1(n15051), .A2(n15050), .A3(n15049), .A4(n15048), .ZN(
        P1_U3098) );
  NAND2_X1 U18224 ( .A1(n20675), .A2(n20665), .ZN(n15055) );
  AOI22_X1 U18225 ( .A1(n20719), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n15072), .ZN(n15054) );
  NAND2_X1 U18226 ( .A1(n15074), .A2(n20718), .ZN(n15053) );
  NAND2_X1 U18227 ( .A1(n15075), .A2(n20720), .ZN(n15052) );
  NAND4_X1 U18228 ( .A1(n15055), .A2(n15054), .A3(n15053), .A4(n15052), .ZN(
        P1_U3099) );
  NAND2_X1 U18229 ( .A1(n20675), .A2(n20669), .ZN(n15059) );
  AOI22_X1 U18230 ( .A1(n20725), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n15072), .ZN(n15058) );
  NAND2_X1 U18231 ( .A1(n15074), .A2(n20724), .ZN(n15057) );
  NAND2_X1 U18232 ( .A1(n15075), .A2(n20726), .ZN(n15056) );
  NAND4_X1 U18233 ( .A1(n15059), .A2(n15058), .A3(n15057), .A4(n15056), .ZN(
        P1_U3100) );
  NAND2_X1 U18234 ( .A1(n20675), .A2(n20633), .ZN(n15063) );
  AOI22_X1 U18235 ( .A1(n20731), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n15072), .ZN(n15062) );
  NAND2_X1 U18236 ( .A1(n15074), .A2(n20730), .ZN(n15061) );
  NAND2_X1 U18237 ( .A1(n15075), .A2(n20732), .ZN(n15060) );
  NAND4_X1 U18238 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        P1_U3101) );
  NAND2_X1 U18239 ( .A1(n20675), .A2(n20637), .ZN(n15067) );
  AOI22_X1 U18240 ( .A1(n20737), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__5__SCAN_IN), .B2(n15072), .ZN(n15066) );
  NAND2_X1 U18241 ( .A1(n15074), .A2(n20736), .ZN(n15065) );
  NAND2_X1 U18242 ( .A1(n15075), .A2(n20738), .ZN(n15064) );
  NAND4_X1 U18243 ( .A1(n15067), .A2(n15066), .A3(n15065), .A4(n15064), .ZN(
        P1_U3102) );
  NAND2_X1 U18244 ( .A1(n20675), .A2(n20679), .ZN(n15071) );
  AOI22_X1 U18245 ( .A1(n21074), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n15072), .ZN(n15070) );
  NAND2_X1 U18246 ( .A1(n15074), .A2(n20742), .ZN(n15069) );
  NAND2_X1 U18247 ( .A1(n15075), .A2(n20744), .ZN(n15068) );
  NAND4_X1 U18248 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        P1_U3103) );
  NAND2_X1 U18249 ( .A1(n20675), .A2(n20685), .ZN(n15079) );
  AOI22_X1 U18250 ( .A1(n20751), .A2(n15073), .B1(
        P1_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n15072), .ZN(n15078) );
  NAND2_X1 U18251 ( .A1(n15074), .A2(n20749), .ZN(n15077) );
  NAND2_X1 U18252 ( .A1(n15075), .A2(n20752), .ZN(n15076) );
  NAND4_X1 U18253 ( .A1(n15079), .A2(n15078), .A3(n15077), .A4(n15076), .ZN(
        P1_U3104) );
  OR2_X1 U18254 ( .A1(n15117), .A2(n15080), .ZN(n15081) );
  NAND2_X1 U18255 ( .A1(n15264), .A2(n15081), .ZN(n15666) );
  INV_X1 U18256 ( .A(n15666), .ZN(n15082) );
  NAND2_X1 U18257 ( .A1(n15082), .A2(n19396), .ZN(n15113) );
  AND2_X1 U18258 ( .A1(n15085), .A2(n15084), .ZN(n15086) );
  NOR2_X1 U18259 ( .A1(n15083), .A2(n15086), .ZN(n16612) );
  NAND2_X1 U18260 ( .A1(n19411), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15110) );
  INV_X1 U18261 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20189) );
  OAI22_X1 U18262 ( .A1(n10043), .A2(n19389), .B1(n20189), .B2(n19405), .ZN(
        n15087) );
  INV_X1 U18263 ( .A(n15087), .ZN(n15109) );
  NOR2_X1 U18264 ( .A1(n9771), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15088) );
  OR2_X1 U18265 ( .A1(n9772), .A2(n15088), .ZN(n15436) );
  AND2_X1 U18266 ( .A1(n15089), .A2(n15091), .ZN(n15090) );
  OR2_X1 U18267 ( .A1(n15090), .A2(n9771), .ZN(n15447) );
  OAI21_X1 U18268 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n15092), .A(
        n15091), .ZN(n15471) );
  OAI21_X1 U18269 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15094), .A(
        n15093), .ZN(n19300) );
  AOI21_X1 U18270 ( .B1(n15494), .B2(n15105), .A(n15094), .ZN(n15496) );
  NAND2_X1 U18271 ( .A1(n15515), .A2(n15103), .ZN(n15096) );
  INV_X1 U18272 ( .A(n15106), .ZN(n15095) );
  AND2_X1 U18273 ( .A1(n15096), .A2(n15095), .ZN(n15517) );
  AND2_X1 U18274 ( .A1(n15102), .A2(n15538), .ZN(n15097) );
  OR2_X1 U18275 ( .A1(n15104), .A2(n15097), .ZN(n15174) );
  INV_X1 U18276 ( .A(n15174), .ZN(n15540) );
  INV_X1 U18277 ( .A(n15100), .ZN(n15098) );
  AOI21_X1 U18278 ( .B1(n15563), .B2(n15099), .A(n15098), .ZN(n15565) );
  NAND2_X1 U18279 ( .A1(n15194), .A2(n15577), .ZN(n15183) );
  NOR2_X1 U18280 ( .A1(n15565), .A2(n15183), .ZN(n19327) );
  NAND2_X1 U18281 ( .A1(n15100), .A2(n19328), .ZN(n15101) );
  NAND2_X1 U18282 ( .A1(n15102), .A2(n15101), .ZN(n19334) );
  NAND2_X1 U18283 ( .A1(n19327), .A2(n19334), .ZN(n15169) );
  NOR2_X1 U18284 ( .A1(n15540), .A2(n15169), .ZN(n15168) );
  OAI21_X1 U18285 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15104), .A(
        n15103), .ZN(n19320) );
  NAND2_X1 U18286 ( .A1(n15168), .A2(n19320), .ZN(n15160) );
  NOR2_X1 U18287 ( .A1(n15517), .A2(n15160), .ZN(n19308) );
  OAI21_X1 U18288 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n15106), .A(
        n15105), .ZN(n19309) );
  NAND2_X1 U18289 ( .A1(n9661), .A2(n15144), .ZN(n19299) );
  NAND2_X1 U18290 ( .A1(n19300), .A2(n19299), .ZN(n19298) );
  NAND2_X1 U18291 ( .A1(n9661), .A2(n19298), .ZN(n15129) );
  NAND2_X1 U18292 ( .A1(n15471), .A2(n15129), .ZN(n15128) );
  NAND2_X1 U18293 ( .A1(n9661), .A2(n15128), .ZN(n15120) );
  NAND2_X1 U18294 ( .A1(n15447), .A2(n15120), .ZN(n15119) );
  OAI211_X1 U18295 ( .C1(n15436), .C2(n15107), .A(n9671), .B(n16514), .ZN(
        n15108) );
  NAND3_X1 U18296 ( .A1(n15110), .A2(n15109), .A3(n15108), .ZN(n15111) );
  AOI21_X1 U18297 ( .B1(n16612), .B2(n19377), .A(n15111), .ZN(n15112) );
  OAI211_X1 U18298 ( .C1(n19404), .C2(n15114), .A(n15113), .B(n15112), .ZN(
        P2_U2832) );
  NOR2_X1 U18299 ( .A1(n15132), .A2(n15115), .ZN(n15116) );
  OR2_X1 U18300 ( .A1(n15117), .A2(n15116), .ZN(n15678) );
  XNOR2_X1 U18301 ( .A(n15135), .B(n15118), .ZN(n15680) );
  INV_X1 U18302 ( .A(n15680), .ZN(n16619) );
  INV_X1 U18303 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20187) );
  OAI22_X1 U18304 ( .A1(n15089), .A2(n19389), .B1(n20187), .B2(n19405), .ZN(
        n15124) );
  INV_X1 U18305 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15122) );
  OAI211_X1 U18306 ( .C1(n15447), .C2(n15120), .A(n9671), .B(n15119), .ZN(
        n15121) );
  OAI21_X1 U18307 ( .B1(n19352), .B2(n15122), .A(n15121), .ZN(n15123) );
  AOI211_X1 U18308 ( .C1(n16619), .C2(n19377), .A(n15124), .B(n15123), .ZN(
        n15127) );
  NAND2_X1 U18309 ( .A1(n15125), .A2(n19294), .ZN(n15126) );
  OAI211_X1 U18310 ( .C1(n15678), .C2(n19413), .A(n15127), .B(n15126), .ZN(
        P2_U2833) );
  OAI211_X1 U18311 ( .C1(n15129), .C2(n15471), .A(n9671), .B(n15128), .ZN(
        n15140) );
  AND2_X1 U18312 ( .A1(n15287), .A2(n15130), .ZN(n15131) );
  NOR2_X1 U18313 ( .A1(n15132), .A2(n15131), .ZN(n15690) );
  OR2_X1 U18314 ( .A1(n15362), .A2(n15133), .ZN(n15134) );
  NAND2_X1 U18315 ( .A1(n15135), .A2(n15134), .ZN(n15693) );
  OAI22_X1 U18316 ( .A1(n10042), .A2(n19389), .B1(n20185), .B2(n19405), .ZN(
        n15136) );
  AOI21_X1 U18317 ( .B1(n19411), .B2(P2_EBX_REG_21__SCAN_IN), .A(n15136), .ZN(
        n15137) );
  OAI21_X1 U18318 ( .B1(n15693), .B2(n19408), .A(n15137), .ZN(n15138) );
  AOI21_X1 U18319 ( .B1(n15690), .B2(n19396), .A(n15138), .ZN(n15139) );
  OAI211_X1 U18320 ( .C1(n15141), .C2(n19404), .A(n15140), .B(n15139), .ZN(
        P2_U2834) );
  AOI21_X1 U18321 ( .B1(n15496), .B2(n15142), .A(n20126), .ZN(n15143) );
  NAND2_X1 U18322 ( .A1(n15144), .A2(n15143), .ZN(n15156) );
  NAND2_X1 U18323 ( .A1(n15146), .A2(n15145), .ZN(n15147) );
  AND2_X1 U18324 ( .A1(n15363), .A2(n15147), .ZN(n15716) );
  INV_X1 U18325 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n15493) );
  NAND2_X1 U18326 ( .A1(n19411), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15149) );
  AOI21_X1 U18327 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19417), .A(
        n19529), .ZN(n15148) );
  OAI211_X1 U18328 ( .C1(n15493), .C2(n19405), .A(n15149), .B(n15148), .ZN(
        n15154) );
  OR2_X1 U18329 ( .A1(n15151), .A2(n15150), .ZN(n15152) );
  NAND2_X1 U18330 ( .A1(n15289), .A2(n15152), .ZN(n15718) );
  NOR2_X1 U18331 ( .A1(n15718), .A2(n19413), .ZN(n15153) );
  AOI211_X1 U18332 ( .C1(n19377), .C2(n15716), .A(n15154), .B(n15153), .ZN(
        n15155) );
  OAI211_X1 U18333 ( .C1(n19404), .C2(n15157), .A(n15156), .B(n15155), .ZN(
        P2_U2836) );
  INV_X1 U18334 ( .A(n15744), .ZN(n15165) );
  INV_X1 U18335 ( .A(n15517), .ZN(n15159) );
  INV_X1 U18336 ( .A(n19397), .ZN(n15173) );
  AOI22_X1 U18337 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19417), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19411), .ZN(n15158) );
  OAI211_X1 U18338 ( .C1(n15159), .C2(n15173), .A(n15727), .B(n15158), .ZN(
        n15162) );
  NAND2_X1 U18339 ( .A1(n9671), .A2(n13308), .ZN(n16528) );
  AOI211_X1 U18340 ( .C1(n15160), .C2(n15517), .A(n16528), .B(n19308), .ZN(
        n15161) );
  AOI211_X1 U18341 ( .C1(n19392), .C2(P2_REIP_REG_17__SCAN_IN), .A(n15162), 
        .B(n15161), .ZN(n15163) );
  OAI21_X1 U18342 ( .B1(n15746), .B2(n19408), .A(n15163), .ZN(n15164) );
  AOI21_X1 U18343 ( .B1(n15165), .B2(n19396), .A(n15164), .ZN(n15166) );
  OAI21_X1 U18344 ( .B1(n15167), .B2(n19404), .A(n15166), .ZN(P2_U2838) );
  OR2_X1 U18345 ( .A1(n19379), .A2(n15168), .ZN(n19321) );
  AOI211_X1 U18346 ( .C1(n15540), .C2(n15169), .A(n20126), .B(n19321), .ZN(
        n15182) );
  AND2_X1 U18347 ( .A1(n15782), .A2(n15170), .ZN(n15171) );
  NOR2_X1 U18348 ( .A1(n9759), .A2(n15171), .ZN(n19425) );
  INV_X1 U18349 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20174) );
  NOR2_X1 U18350 ( .A1(n19405), .A2(n20174), .ZN(n15176) );
  AOI22_X1 U18351 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n19411), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19417), .ZN(n15172) );
  OAI211_X1 U18352 ( .C1(n15174), .C2(n15173), .A(n15172), .B(n15727), .ZN(
        n15175) );
  AOI211_X1 U18353 ( .C1(n19425), .C2(n19377), .A(n15176), .B(n15175), .ZN(
        n15180) );
  OAI211_X1 U18354 ( .C1(n15178), .C2(n15177), .A(n10760), .B(n19294), .ZN(
        n15179) );
  OAI211_X1 U18355 ( .C1(n15769), .C2(n19413), .A(n15180), .B(n15179), .ZN(
        n15181) );
  OR2_X1 U18356 ( .A1(n15182), .A2(n15181), .ZN(P2_U2840) );
  NAND2_X1 U18357 ( .A1(n15565), .A2(n15183), .ZN(n15188) );
  NOR2_X1 U18358 ( .A1(n19327), .A2(n16528), .ZN(n19335) );
  OAI22_X1 U18359 ( .A1(n19352), .A2(n10928), .B1(n15563), .B2(n19389), .ZN(
        n15187) );
  AOI22_X1 U18360 ( .A1(n19397), .A2(n15565), .B1(n19294), .B2(n15184), .ZN(
        n15185) );
  OAI211_X1 U18361 ( .C1(n20170), .C2(n19405), .A(n15185), .B(n19363), .ZN(
        n15186) );
  AOI211_X1 U18362 ( .C1(n15188), .C2(n19335), .A(n15187), .B(n15186), .ZN(
        n15193) );
  OAI21_X1 U18363 ( .B1(n15190), .B2(n15189), .A(n15781), .ZN(n19435) );
  INV_X1 U18364 ( .A(n19435), .ZN(n15191) );
  NAND2_X1 U18365 ( .A1(n15191), .A2(n19377), .ZN(n15192) );
  OAI211_X1 U18366 ( .C1(n15795), .C2(n19413), .A(n15193), .B(n15192), .ZN(
        P2_U2842) );
  AOI211_X1 U18367 ( .C1(n16624), .C2(n15195), .A(n15194), .B(n16528), .ZN(
        n15196) );
  INV_X1 U18368 ( .A(n15196), .ZN(n15208) );
  INV_X1 U18369 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15205) );
  INV_X1 U18370 ( .A(n15197), .ZN(n15200) );
  INV_X1 U18371 ( .A(n15198), .ZN(n15199) );
  AOI21_X1 U18372 ( .B1(n15200), .B2(n9753), .A(n15199), .ZN(n19439) );
  NAND2_X1 U18373 ( .A1(n19377), .A2(n19439), .ZN(n15204) );
  OAI22_X1 U18374 ( .A1(n19352), .A2(n15201), .B1(n16635), .B2(n19389), .ZN(
        n15202) );
  AOI211_X1 U18375 ( .C1(n19397), .C2(n16624), .A(n15202), .B(n19529), .ZN(
        n15203) );
  OAI211_X1 U18376 ( .C1(n19405), .C2(n15205), .A(n15204), .B(n15203), .ZN(
        n15206) );
  AOI21_X1 U18377 ( .B1(n16672), .B2(n19396), .A(n15206), .ZN(n15207) );
  OAI211_X1 U18378 ( .C1(n19404), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        P2_U2844) );
  INV_X1 U18379 ( .A(n15212), .ZN(n15213) );
  NOR2_X1 U18380 ( .A1(n19379), .A2(n15210), .ZN(n15873) );
  INV_X1 U18381 ( .A(n15873), .ZN(n15211) );
  AOI221_X1 U18382 ( .B1(n15213), .B2(n15873), .C1(n15212), .C2(n15211), .A(
        n20126), .ZN(n15214) );
  INV_X1 U18383 ( .A(n15214), .ZN(n15221) );
  NAND2_X1 U18384 ( .A1(n19411), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U18385 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19417), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19392), .ZN(n15215) );
  OAI211_X1 U18386 ( .C1(n19404), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15219) );
  NOR2_X1 U18387 ( .A1(n12075), .A2(n19413), .ZN(n15218) );
  AOI211_X1 U18388 ( .C1(n19377), .C2(n20241), .A(n15219), .B(n15218), .ZN(
        n15220) );
  OAI211_X1 U18389 ( .C1(n20239), .C2(n19382), .A(n15221), .B(n15220), .ZN(
        P2_U2853) );
  MUX2_X1 U18390 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16525), .S(n15291), .Z(
        P2_U2856) );
  OR2_X1 U18391 ( .A1(n15223), .A2(n15222), .ZN(n15224) );
  NAND2_X1 U18392 ( .A1(n15225), .A2(n15224), .ZN(n16542) );
  OR2_X1 U18393 ( .A1(n9699), .A2(n15226), .ZN(n15303) );
  NAND3_X1 U18394 ( .A1(n15303), .A2(n15227), .A3(n15281), .ZN(n15229) );
  NAND2_X1 U18395 ( .A1(n15279), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15228) );
  OAI211_X1 U18396 ( .C1(n15279), .C2(n16542), .A(n15229), .B(n15228), .ZN(
        P2_U2858) );
  NOR2_X1 U18397 ( .A1(n15231), .A2(n15230), .ZN(n15233) );
  XNOR2_X1 U18398 ( .A(n15233), .B(n15232), .ZN(n15309) );
  NAND2_X1 U18399 ( .A1(n15309), .A2(n15281), .ZN(n15235) );
  NAND2_X1 U18400 ( .A1(n15279), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15234) );
  OAI211_X1 U18401 ( .C1(n15279), .C2(n16553), .A(n15235), .B(n15234), .ZN(
        P2_U2859) );
  OAI21_X1 U18402 ( .B1(n15238), .B2(n15237), .A(n15236), .ZN(n15323) );
  NAND2_X1 U18403 ( .A1(n15247), .A2(n15239), .ZN(n15240) );
  NAND2_X1 U18404 ( .A1(n15241), .A2(n15240), .ZN(n16567) );
  NOR2_X1 U18405 ( .A1(n16567), .A2(n15279), .ZN(n15242) );
  AOI21_X1 U18406 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15279), .A(n15242), .ZN(
        n15243) );
  OAI21_X1 U18407 ( .B1(n15323), .B2(n15298), .A(n15243), .ZN(P2_U2860) );
  OAI21_X1 U18408 ( .B1(n15246), .B2(n15245), .A(n15244), .ZN(n15333) );
  OAI21_X1 U18409 ( .B1(n9726), .B2(n15248), .A(n15247), .ZN(n16577) );
  NOR2_X1 U18410 ( .A1(n16577), .A2(n15279), .ZN(n15249) );
  AOI21_X1 U18411 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15279), .A(n15249), .ZN(
        n15250) );
  OAI21_X1 U18412 ( .B1(n15333), .B2(n15298), .A(n15250), .ZN(P2_U2861) );
  OAI21_X1 U18413 ( .B1(n15253), .B2(n15252), .A(n15251), .ZN(n15342) );
  AND2_X1 U18414 ( .A1(n15266), .A2(n15254), .ZN(n15255) );
  OR2_X1 U18415 ( .A1(n15255), .A2(n9726), .ZN(n16590) );
  NOR2_X1 U18416 ( .A1(n16590), .A2(n15279), .ZN(n15256) );
  AOI21_X1 U18417 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15279), .A(n15256), .ZN(
        n15257) );
  OAI21_X1 U18418 ( .B1(n15342), .B2(n15298), .A(n15257), .ZN(P2_U2862) );
  AOI21_X1 U18419 ( .B1(n15260), .B2(n15259), .A(n15258), .ZN(n15261) );
  XOR2_X1 U18420 ( .A(n15262), .B(n15261), .Z(n15354) );
  NAND2_X1 U18421 ( .A1(n15264), .A2(n15263), .ZN(n15265) );
  NAND2_X1 U18422 ( .A1(n15266), .A2(n15265), .ZN(n16602) );
  NOR2_X1 U18423 ( .A1(n16602), .A2(n15279), .ZN(n15267) );
  AOI21_X1 U18424 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15279), .A(n15267), .ZN(
        n15268) );
  OAI21_X1 U18425 ( .B1(n15354), .B2(n15298), .A(n15268), .ZN(P2_U2863) );
  NOR2_X1 U18426 ( .A1(n15270), .A2(n15269), .ZN(n15272) );
  NOR2_X1 U18427 ( .A1(n15272), .A2(n15271), .ZN(n16613) );
  NAND2_X1 U18428 ( .A1(n16613), .A2(n15281), .ZN(n15274) );
  NAND2_X1 U18429 ( .A1(n15279), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15273) );
  OAI211_X1 U18430 ( .C1(n15666), .C2(n15279), .A(n15274), .B(n15273), .ZN(
        P2_U2864) );
  AOI21_X1 U18431 ( .B1(n15276), .B2(n10232), .A(n9727), .ZN(n16620) );
  NAND2_X1 U18432 ( .A1(n16620), .A2(n15281), .ZN(n15278) );
  NAND2_X1 U18433 ( .A1(n15279), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15277) );
  OAI211_X1 U18434 ( .C1(n15678), .C2(n15279), .A(n15278), .B(n15277), .ZN(
        P2_U2865) );
  AOI21_X1 U18435 ( .B1(n15280), .B2(n15285), .A(n15275), .ZN(n15355) );
  NAND2_X1 U18436 ( .A1(n15355), .A2(n15281), .ZN(n15283) );
  NAND2_X1 U18437 ( .A1(n15690), .A2(n15291), .ZN(n15282) );
  OAI211_X1 U18438 ( .C1(n15291), .C2(n10955), .A(n15283), .B(n15282), .ZN(
        P2_U2866) );
  OAI21_X1 U18439 ( .B1(n15284), .B2(n15286), .A(n15285), .ZN(n15369) );
  INV_X1 U18440 ( .A(n15287), .ZN(n15288) );
  AOI21_X1 U18441 ( .B1(n15290), .B2(n15289), .A(n15288), .ZN(n19297) );
  INV_X1 U18442 ( .A(n19297), .ZN(n15705) );
  MUX2_X1 U18443 ( .A(n10951), .B(n15705), .S(n15291), .Z(n15292) );
  OAI21_X1 U18444 ( .B1(n15369), .B2(n15298), .A(n15292), .ZN(P2_U2867) );
  INV_X1 U18445 ( .A(n15284), .ZN(n15293) );
  OAI21_X1 U18446 ( .B1(n15295), .B2(n15294), .A(n15293), .ZN(n15374) );
  NOR2_X1 U18447 ( .A1(n15718), .A2(n15279), .ZN(n15296) );
  AOI21_X1 U18448 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15279), .A(n15296), .ZN(
        n15297) );
  OAI21_X1 U18449 ( .B1(n15374), .B2(n15298), .A(n15297), .ZN(P2_U2868) );
  OR2_X1 U18450 ( .A1(n15300), .A2(n15299), .ZN(n15301) );
  NAND3_X1 U18451 ( .A1(n15303), .A2(n15227), .A3(n19487), .ZN(n15308) );
  INV_X1 U18452 ( .A(n19427), .ZN(n16618) );
  INV_X1 U18453 ( .A(n19463), .ZN(n19485) );
  AOI22_X1 U18454 ( .A1(n16618), .A2(n19433), .B1(n19485), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15304) );
  OAI21_X1 U18455 ( .B1(n15305), .B2(n16852), .A(n15304), .ZN(n15306) );
  AOI21_X1 U18456 ( .B1(n19422), .B2(BUF2_REG_29__SCAN_IN), .A(n15306), .ZN(
        n15307) );
  OAI211_X1 U18457 ( .C1(n15314), .C2(n16541), .A(n15308), .B(n15307), .ZN(
        P2_U2890) );
  NAND2_X1 U18458 ( .A1(n15309), .A2(n19487), .ZN(n15313) );
  OAI22_X1 U18459 ( .A1(n19427), .A2(n19437), .B1(n19463), .B2(n21039), .ZN(
        n15311) );
  AND2_X1 U18460 ( .A1(n19420), .A2(BUF1_REG_28__SCAN_IN), .ZN(n15310) );
  AOI211_X1 U18461 ( .C1(BUF2_REG_28__SCAN_IN), .C2(n19422), .A(n15311), .B(
        n15310), .ZN(n15312) );
  OAI211_X1 U18462 ( .C1(n15314), .C2(n16552), .A(n15313), .B(n15312), .ZN(
        P2_U2891) );
  AND2_X1 U18463 ( .A1(n15324), .A2(n15315), .ZN(n15316) );
  NOR2_X1 U18464 ( .A1(n15317), .A2(n15316), .ZN(n16565) );
  INV_X1 U18465 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U18466 ( .A1(n16618), .A2(n19440), .B1(n19485), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15319) );
  NAND2_X1 U18467 ( .A1(n19420), .A2(BUF1_REG_27__SCAN_IN), .ZN(n15318) );
  OAI211_X1 U18468 ( .C1(n15350), .C2(n15320), .A(n15319), .B(n15318), .ZN(
        n15321) );
  AOI21_X1 U18469 ( .B1(n16565), .B2(n19486), .A(n15321), .ZN(n15322) );
  OAI21_X1 U18470 ( .B1(n15323), .B2(n19458), .A(n15322), .ZN(P2_U2892) );
  INV_X1 U18471 ( .A(n15324), .ZN(n15325) );
  AOI21_X1 U18472 ( .B1(n15326), .B2(n15336), .A(n15325), .ZN(n16578) );
  INV_X1 U18473 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n15330) );
  OAI22_X1 U18474 ( .A1(n19427), .A2(n19443), .B1(n19463), .B2(n15327), .ZN(
        n15328) );
  AOI21_X1 U18475 ( .B1(n19420), .B2(BUF1_REG_26__SCAN_IN), .A(n15328), .ZN(
        n15329) );
  OAI21_X1 U18476 ( .B1(n15350), .B2(n15330), .A(n15329), .ZN(n15331) );
  AOI21_X1 U18477 ( .B1(n16578), .B2(n19486), .A(n15331), .ZN(n15332) );
  OAI21_X1 U18478 ( .B1(n15333), .B2(n19458), .A(n15332), .ZN(P2_U2893) );
  OR2_X1 U18479 ( .A1(n15345), .A2(n15334), .ZN(n15335) );
  AND2_X1 U18480 ( .A1(n15336), .A2(n15335), .ZN(n16588) );
  INV_X1 U18481 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15339) );
  AOI22_X1 U18482 ( .A1(n16618), .A2(n19447), .B1(n19485), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15338) );
  NAND2_X1 U18483 ( .A1(n19420), .A2(BUF1_REG_25__SCAN_IN), .ZN(n15337) );
  OAI211_X1 U18484 ( .C1(n15350), .C2(n15339), .A(n15338), .B(n15337), .ZN(
        n15340) );
  AOI21_X1 U18485 ( .B1(n16588), .B2(n19486), .A(n15340), .ZN(n15341) );
  OAI21_X1 U18486 ( .B1(n15342), .B2(n19458), .A(n15341), .ZN(P2_U2894) );
  NOR2_X1 U18487 ( .A1(n15083), .A2(n15343), .ZN(n15344) );
  OR2_X1 U18488 ( .A1(n15345), .A2(n15344), .ZN(n16601) );
  INV_X1 U18489 ( .A(n16601), .ZN(n15352) );
  INV_X1 U18490 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n15349) );
  OAI22_X1 U18491 ( .A1(n19427), .A2(n19450), .B1(n19463), .B2(n15346), .ZN(
        n15347) );
  AOI21_X1 U18492 ( .B1(n19420), .B2(BUF1_REG_24__SCAN_IN), .A(n15347), .ZN(
        n15348) );
  OAI21_X1 U18493 ( .B1(n15350), .B2(n15349), .A(n15348), .ZN(n15351) );
  AOI21_X1 U18494 ( .B1(n15352), .B2(n19486), .A(n15351), .ZN(n15353) );
  OAI21_X1 U18495 ( .B1(n15354), .B2(n19458), .A(n15353), .ZN(P2_U2895) );
  INV_X1 U18496 ( .A(n15355), .ZN(n15361) );
  INV_X1 U18497 ( .A(n15693), .ZN(n15358) );
  OAI22_X1 U18498 ( .A1(n19427), .A2(n19577), .B1(n15356), .B2(n19463), .ZN(
        n15357) );
  AOI21_X1 U18499 ( .B1(n15358), .B2(n19486), .A(n15357), .ZN(n15360) );
  AOI22_X1 U18500 ( .A1(n19422), .A2(BUF2_REG_21__SCAN_IN), .B1(n19420), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15359) );
  OAI211_X1 U18501 ( .C1(n15361), .C2(n19458), .A(n15360), .B(n15359), .ZN(
        P2_U2898) );
  AOI21_X1 U18502 ( .B1(n15364), .B2(n15363), .A(n15362), .ZN(n19296) );
  OAI22_X1 U18503 ( .A1(n19427), .A2(n19574), .B1(n15365), .B2(n19463), .ZN(
        n15366) );
  AOI21_X1 U18504 ( .B1(n19296), .B2(n19486), .A(n15366), .ZN(n15368) );
  AOI22_X1 U18505 ( .A1(n19422), .A2(BUF2_REG_20__SCAN_IN), .B1(n19420), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15367) );
  OAI211_X1 U18506 ( .C1(n15369), .C2(n19458), .A(n15368), .B(n15367), .ZN(
        P2_U2899) );
  OAI22_X1 U18507 ( .A1(n19427), .A2(n19570), .B1(n15370), .B2(n19463), .ZN(
        n15371) );
  AOI21_X1 U18508 ( .B1(n15716), .B2(n19486), .A(n15371), .ZN(n15373) );
  AOI22_X1 U18509 ( .A1(n19422), .A2(BUF2_REG_19__SCAN_IN), .B1(n19420), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15372) );
  OAI211_X1 U18510 ( .C1(n15374), .C2(n19458), .A(n15373), .B(n15372), .ZN(
        P2_U2900) );
  NAND2_X1 U18511 ( .A1(n15376), .A2(n15375), .ZN(n15378) );
  XOR2_X1 U18512 ( .A(n15378), .B(n15377), .Z(n15616) );
  AOI21_X1 U18513 ( .B1(n15611), .B2(n15380), .A(n15379), .ZN(n15614) );
  AND2_X1 U18514 ( .A1(n15381), .A2(n15384), .ZN(n15382) );
  NOR2_X1 U18515 ( .A1(n9768), .A2(n15382), .ZN(n16517) );
  INV_X1 U18516 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n15383) );
  OR2_X1 U18517 ( .A1(n19363), .A2(n15383), .ZN(n15606) );
  OAI21_X1 U18518 ( .B1(n16666), .B2(n15384), .A(n15606), .ZN(n15385) );
  AOI21_X1 U18519 ( .B1(n16658), .B2(n16517), .A(n15385), .ZN(n15386) );
  OAI21_X1 U18520 ( .B1(n16542), .B2(n16648), .A(n15386), .ZN(n15387) );
  AOI21_X1 U18521 ( .B1(n15614), .B2(n16660), .A(n15387), .ZN(n15388) );
  OAI21_X1 U18522 ( .B1(n15616), .B2(n19534), .A(n15388), .ZN(P2_U2985) );
  NAND2_X1 U18523 ( .A1(n15389), .A2(n15626), .ZN(n15619) );
  NAND2_X1 U18524 ( .A1(n15619), .A2(n16662), .ZN(n15400) );
  AOI21_X1 U18525 ( .B1(n15626), .B2(n15390), .A(n10887), .ZN(n15617) );
  NOR2_X1 U18526 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n15391), .ZN(
        n15392) );
  NOR2_X1 U18527 ( .A1(n15393), .A2(n15392), .ZN(n16516) );
  INV_X1 U18528 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15395) );
  INV_X1 U18529 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n15394) );
  OR2_X1 U18530 ( .A1(n19363), .A2(n15394), .ZN(n15623) );
  OAI21_X1 U18531 ( .B1(n16666), .B2(n15395), .A(n15623), .ZN(n15396) );
  AOI21_X1 U18532 ( .B1(n16658), .B2(n16516), .A(n15396), .ZN(n15397) );
  OAI21_X1 U18533 ( .B1(n16567), .B2(n16648), .A(n15397), .ZN(n15398) );
  AOI21_X1 U18534 ( .B1(n15617), .B2(n16660), .A(n15398), .ZN(n15399) );
  OAI21_X1 U18535 ( .B1(n15618), .B2(n15400), .A(n15399), .ZN(P2_U2987) );
  OAI21_X1 U18536 ( .B1(n15401), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15390), .ZN(n15641) );
  NOR2_X1 U18537 ( .A1(n15402), .A2(n15410), .ZN(n15404) );
  XNOR2_X1 U18538 ( .A(n15404), .B(n15403), .ZN(n15639) );
  INV_X1 U18539 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20195) );
  NOR2_X1 U18540 ( .A1(n15727), .A2(n20195), .ZN(n15634) );
  OAI21_X1 U18541 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n15414), .A(
        n15405), .ZN(n16582) );
  NOR2_X1 U18542 ( .A1(n19542), .A2(n16582), .ZN(n15406) );
  AOI211_X1 U18543 ( .C1(n19530), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15634), .B(n15406), .ZN(n15407) );
  OAI21_X1 U18544 ( .B1(n16577), .B2(n16648), .A(n15407), .ZN(n15408) );
  AOI21_X1 U18545 ( .B1(n15639), .B2(n16662), .A(n15408), .ZN(n15409) );
  OAI21_X1 U18546 ( .B1(n19532), .B2(n15641), .A(n15409), .ZN(P2_U2988) );
  NOR2_X1 U18547 ( .A1(n15411), .A2(n15410), .ZN(n15413) );
  XOR2_X1 U18548 ( .A(n15413), .B(n15412), .Z(n15653) );
  AOI21_X1 U18549 ( .B1(n15415), .B2(n15425), .A(n15414), .ZN(n16515) );
  NAND2_X1 U18550 ( .A1(n19529), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15645) );
  OAI21_X1 U18551 ( .B1(n16666), .B2(n15415), .A(n15645), .ZN(n15417) );
  NOR2_X1 U18552 ( .A1(n16590), .A2(n16648), .ZN(n15416) );
  AOI211_X1 U18553 ( .C1(n16658), .C2(n16515), .A(n15417), .B(n15416), .ZN(
        n15420) );
  AOI21_X1 U18554 ( .B1(n15648), .B2(n15418), .A(n15401), .ZN(n15650) );
  NAND2_X1 U18555 ( .A1(n15650), .A2(n16660), .ZN(n15419) );
  OAI211_X1 U18556 ( .C1(n15653), .C2(n19534), .A(n15420), .B(n15419), .ZN(
        P2_U2989) );
  OAI21_X1 U18557 ( .B1(n15421), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15418), .ZN(n15664) );
  XOR2_X1 U18558 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15422), .Z(
        n15423) );
  XNOR2_X1 U18559 ( .A(n15424), .B(n15423), .ZN(n15662) );
  NOR2_X1 U18560 ( .A1(n15727), .A2(n20191), .ZN(n15656) );
  OAI21_X1 U18561 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n9772), .A(
        n15425), .ZN(n16606) );
  NOR2_X1 U18562 ( .A1(n19542), .A2(n16606), .ZN(n15426) );
  AOI211_X1 U18563 ( .C1(n19530), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15656), .B(n15426), .ZN(n15427) );
  OAI21_X1 U18564 ( .B1(n16602), .B2(n16648), .A(n15427), .ZN(n15428) );
  AOI21_X1 U18565 ( .B1(n15662), .B2(n16662), .A(n15428), .ZN(n15429) );
  OAI21_X1 U18566 ( .B1(n19532), .B2(n15664), .A(n15429), .ZN(P2_U2990) );
  NOR2_X1 U18567 ( .A1(n15430), .A2(n15431), .ZN(n15433) );
  INV_X1 U18568 ( .A(n15421), .ZN(n15432) );
  OAI21_X1 U18569 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15433), .A(
        n15432), .ZN(n15675) );
  XOR2_X1 U18570 ( .A(n15435), .B(n15434), .Z(n15673) );
  NOR2_X1 U18571 ( .A1(n15727), .A2(n20189), .ZN(n15668) );
  NOR2_X1 U18572 ( .A1(n19542), .A2(n15436), .ZN(n15437) );
  AOI211_X1 U18573 ( .C1(n19530), .C2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15668), .B(n15437), .ZN(n15438) );
  OAI21_X1 U18574 ( .B1(n15666), .B2(n16648), .A(n15438), .ZN(n15439) );
  AOI21_X1 U18575 ( .B1(n15673), .B2(n16662), .A(n15439), .ZN(n15440) );
  OAI21_X1 U18576 ( .B1(n19532), .B2(n15675), .A(n15440), .ZN(P2_U2991) );
  XOR2_X1 U18577 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15430), .Z(
        n15688) );
  INV_X1 U18578 ( .A(n15441), .ZN(n15442) );
  NOR2_X1 U18579 ( .A1(n15443), .A2(n15442), .ZN(n15444) );
  XNOR2_X1 U18580 ( .A(n15445), .B(n15444), .ZN(n15686) );
  NOR2_X1 U18581 ( .A1(n15678), .A2(n16648), .ZN(n15449) );
  NAND2_X1 U18582 ( .A1(n19529), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n15679) );
  NAND2_X1 U18583 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15446) );
  OAI211_X1 U18584 ( .C1(n19542), .C2(n15447), .A(n15679), .B(n15446), .ZN(
        n15448) );
  AOI211_X1 U18585 ( .C1(n15686), .C2(n16662), .A(n15449), .B(n15448), .ZN(
        n15450) );
  OAI21_X1 U18586 ( .B1(n15688), .B2(n19532), .A(n15450), .ZN(P2_U2992) );
  OAI21_X1 U18587 ( .B1(n15485), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15430), .ZN(n15700) );
  INV_X1 U18588 ( .A(n15533), .ZN(n15532) );
  NAND2_X1 U18589 ( .A1(n15532), .A2(n15452), .ZN(n15455) );
  OAI211_X1 U18590 ( .C1(n15451), .C2(n15455), .A(n15454), .B(n15453), .ZN(
        n15457) );
  INV_X1 U18591 ( .A(n15456), .ZN(n15535) );
  NAND2_X1 U18592 ( .A1(n15457), .A2(n15535), .ZN(n15524) );
  INV_X1 U18593 ( .A(n15523), .ZN(n15459) );
  OAI21_X1 U18594 ( .B1(n15524), .B2(n15459), .A(n15458), .ZN(n15514) );
  INV_X1 U18595 ( .A(n15460), .ZN(n15462) );
  NAND2_X1 U18596 ( .A1(n15462), .A2(n15461), .ZN(n15513) );
  OAI21_X1 U18597 ( .B1(n15514), .B2(n15513), .A(n15462), .ZN(n15503) );
  NAND2_X1 U18598 ( .A1(n15503), .A2(n15501), .ZN(n15490) );
  INV_X1 U18599 ( .A(n15488), .ZN(n15465) );
  INV_X1 U18600 ( .A(n15463), .ZN(n15464) );
  OAI21_X1 U18601 ( .B1(n15490), .B2(n15465), .A(n15464), .ZN(n15476) );
  NOR2_X1 U18602 ( .A1(n15476), .A2(n15477), .ZN(n15475) );
  NOR2_X1 U18603 ( .A1(n15475), .A2(n15479), .ZN(n15469) );
  NOR2_X1 U18604 ( .A1(n15467), .A2(n15466), .ZN(n15468) );
  XNOR2_X1 U18605 ( .A(n15469), .B(n15468), .ZN(n15689) );
  NAND2_X1 U18606 ( .A1(n15689), .A2(n16662), .ZN(n15474) );
  NAND2_X1 U18607 ( .A1(n19529), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15691) );
  NAND2_X1 U18608 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15470) );
  OAI211_X1 U18609 ( .C1(n19542), .C2(n15471), .A(n15691), .B(n15470), .ZN(
        n15472) );
  AOI21_X1 U18610 ( .B1(n15690), .B2(n19538), .A(n15472), .ZN(n15473) );
  OAI211_X1 U18611 ( .C1(n19532), .C2(n15700), .A(n15474), .B(n15473), .ZN(
        P2_U2993) );
  INV_X1 U18612 ( .A(n15475), .ZN(n15480) );
  OAI21_X1 U18613 ( .B1(n15477), .B2(n15479), .A(n15476), .ZN(n15478) );
  OAI21_X1 U18614 ( .B1(n15480), .B2(n15479), .A(n15478), .ZN(n15714) );
  INV_X1 U18615 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20183) );
  NOR2_X1 U18616 ( .A1(n15727), .A2(n20183), .ZN(n15703) );
  AOI21_X1 U18617 ( .B1(n19530), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15703), .ZN(n15481) );
  OAI21_X1 U18618 ( .B1(n19542), .B2(n19300), .A(n15481), .ZN(n15482) );
  AOI21_X1 U18619 ( .B1(n19297), .B2(n19538), .A(n15482), .ZN(n15487) );
  NAND2_X1 U18620 ( .A1(n15694), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15484) );
  OAI22_X1 U18621 ( .A1(n15485), .A2(n15708), .B1(n15483), .B2(n15484), .ZN(
        n15711) );
  NAND2_X1 U18622 ( .A1(n15711), .A2(n16660), .ZN(n15486) );
  OAI211_X1 U18623 ( .C1(n15714), .C2(n19534), .A(n15487), .B(n15486), .ZN(
        P2_U2994) );
  XNOR2_X1 U18624 ( .A(n15483), .B(n15707), .ZN(n15725) );
  NAND2_X1 U18625 ( .A1(n15489), .A2(n15488), .ZN(n15492) );
  NAND2_X1 U18626 ( .A1(n15490), .A2(n15500), .ZN(n15491) );
  XOR2_X1 U18627 ( .A(n15492), .B(n15491), .Z(n15723) );
  NOR2_X1 U18628 ( .A1(n15727), .A2(n15493), .ZN(n15715) );
  NOR2_X1 U18629 ( .A1(n16666), .A2(n15494), .ZN(n15495) );
  AOI211_X1 U18630 ( .C1(n15496), .C2(n16658), .A(n15715), .B(n15495), .ZN(
        n15497) );
  OAI21_X1 U18631 ( .B1(n15718), .B2(n16648), .A(n15497), .ZN(n15498) );
  AOI21_X1 U18632 ( .B1(n15723), .B2(n16662), .A(n15498), .ZN(n15499) );
  OAI21_X1 U18633 ( .B1(n19532), .B2(n15725), .A(n15499), .ZN(P2_U2995) );
  NAND2_X1 U18634 ( .A1(n15501), .A2(n15500), .ZN(n15502) );
  XNOR2_X1 U18635 ( .A(n15503), .B(n15502), .ZN(n15738) );
  INV_X1 U18636 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20180) );
  OAI22_X1 U18637 ( .A1(n20180), .A2(n19363), .B1(n19542), .B2(n19309), .ZN(
        n15505) );
  NOR2_X1 U18638 ( .A1(n15732), .A2(n16648), .ZN(n15504) );
  AOI211_X1 U18639 ( .C1(n19530), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15505), .B(n15504), .ZN(n15509) );
  INV_X1 U18640 ( .A(n15483), .ZN(n15507) );
  AOI21_X1 U18641 ( .B1(n11366), .B2(n15506), .A(n15507), .ZN(n15735) );
  NAND2_X1 U18642 ( .A1(n15735), .A2(n16660), .ZN(n15508) );
  OAI211_X1 U18643 ( .C1(n15738), .C2(n19534), .A(n15509), .B(n15508), .ZN(
        P2_U2996) );
  NOR2_X1 U18644 ( .A1(n15510), .A2(n15511), .ZN(n15522) );
  NAND2_X1 U18645 ( .A1(n15522), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15739) );
  INV_X1 U18646 ( .A(n15739), .ZN(n15512) );
  AOI22_X1 U18647 ( .A1(n15512), .A2(n15726), .B1(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15506), .ZN(n15521) );
  XNOR2_X1 U18648 ( .A(n15514), .B(n15513), .ZN(n15749) );
  OR2_X1 U18649 ( .A1(n19363), .A2(n20178), .ZN(n15745) );
  OAI21_X1 U18650 ( .B1(n16666), .B2(n15515), .A(n15745), .ZN(n15516) );
  AOI21_X1 U18651 ( .B1(n16658), .B2(n15517), .A(n15516), .ZN(n15518) );
  OAI21_X1 U18652 ( .B1(n15744), .B2(n16648), .A(n15518), .ZN(n15519) );
  AOI21_X1 U18653 ( .B1(n15749), .B2(n16662), .A(n15519), .ZN(n15520) );
  OAI21_X1 U18654 ( .B1(n15521), .B2(n19532), .A(n15520), .ZN(P2_U2997) );
  XNOR2_X1 U18655 ( .A(n15522), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15529) );
  XNOR2_X1 U18656 ( .A(n15524), .B(n15523), .ZN(n15760) );
  NOR2_X1 U18657 ( .A1(n19319), .A2(n16648), .ZN(n15527) );
  NAND2_X1 U18658 ( .A1(n19529), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15757) );
  NAND2_X1 U18659 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15525) );
  OAI211_X1 U18660 ( .C1(n19542), .C2(n19320), .A(n15757), .B(n15525), .ZN(
        n15526) );
  AOI211_X1 U18661 ( .C1(n15760), .C2(n16662), .A(n15527), .B(n15526), .ZN(
        n15528) );
  OAI21_X1 U18662 ( .B1(n15529), .B2(n19532), .A(n15528), .ZN(P2_U2998) );
  XOR2_X1 U18663 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n15510), .Z(
        n15777) );
  NAND2_X1 U18664 ( .A1(n15530), .A2(n15559), .ZN(n15546) );
  NAND2_X1 U18665 ( .A1(n15532), .A2(n15531), .ZN(n15545) );
  NOR2_X1 U18666 ( .A1(n15546), .A2(n15545), .ZN(n15544) );
  NOR2_X1 U18667 ( .A1(n15544), .A2(n15533), .ZN(n15537) );
  NAND2_X1 U18668 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  XNOR2_X1 U18669 ( .A(n15537), .B(n15536), .ZN(n15775) );
  NOR2_X1 U18670 ( .A1(n15727), .A2(n20174), .ZN(n15767) );
  NOR2_X1 U18671 ( .A1(n16666), .A2(n15538), .ZN(n15539) );
  AOI211_X1 U18672 ( .C1(n15540), .C2(n16658), .A(n15767), .B(n15539), .ZN(
        n15541) );
  OAI21_X1 U18673 ( .B1(n15769), .B2(n16648), .A(n15541), .ZN(n15542) );
  AOI21_X1 U18674 ( .B1(n15775), .B2(n16662), .A(n15542), .ZN(n15543) );
  OAI21_X1 U18675 ( .B1(n19532), .B2(n15777), .A(n15543), .ZN(P2_U2999) );
  AOI21_X1 U18676 ( .B1(n15546), .B2(n15545), .A(n15544), .ZN(n15791) );
  INV_X1 U18677 ( .A(n15547), .ZN(n19336) );
  NAND2_X1 U18678 ( .A1(n19529), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n15783) );
  NAND2_X1 U18679 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15548) );
  OAI211_X1 U18680 ( .C1(n19542), .C2(n19334), .A(n15783), .B(n15548), .ZN(
        n15549) );
  AOI21_X1 U18681 ( .B1(n19336), .B2(n19538), .A(n15549), .ZN(n15554) );
  INV_X1 U18682 ( .A(n15785), .ZN(n15780) );
  NAND2_X1 U18683 ( .A1(n16631), .A2(n15780), .ZN(n15556) );
  INV_X1 U18684 ( .A(n15510), .ZN(n15551) );
  AOI21_X1 U18685 ( .B1(n15556), .B2(n15552), .A(n15551), .ZN(n15788) );
  NAND2_X1 U18686 ( .A1(n15788), .A2(n16660), .ZN(n15553) );
  OAI211_X1 U18687 ( .C1(n15791), .C2(n19534), .A(n15554), .B(n15553), .ZN(
        P2_U3000) );
  INV_X1 U18688 ( .A(n16631), .ZN(n15555) );
  INV_X1 U18689 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15792) );
  NOR2_X1 U18690 ( .A1(n15555), .A2(n15792), .ZN(n15557) );
  OAI21_X1 U18691 ( .B1(n15557), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15556), .ZN(n15803) );
  NAND2_X1 U18692 ( .A1(n15559), .A2(n15558), .ZN(n15562) );
  NAND2_X1 U18693 ( .A1(n15560), .A2(n15571), .ZN(n15561) );
  XOR2_X1 U18694 ( .A(n15562), .B(n15561), .Z(n15801) );
  NOR2_X1 U18695 ( .A1(n15727), .A2(n20170), .ZN(n15796) );
  NOR2_X1 U18696 ( .A1(n16666), .A2(n15563), .ZN(n15564) );
  AOI211_X1 U18697 ( .C1(n15565), .C2(n16658), .A(n15796), .B(n15564), .ZN(
        n15566) );
  OAI21_X1 U18698 ( .B1(n15795), .B2(n16648), .A(n15566), .ZN(n15567) );
  AOI21_X1 U18699 ( .B1(n15801), .B2(n16662), .A(n15567), .ZN(n15568) );
  OAI21_X1 U18700 ( .B1(n15803), .B2(n19532), .A(n15568), .ZN(P2_U3001) );
  XNOR2_X1 U18701 ( .A(n16631), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15815) );
  INV_X1 U18702 ( .A(n15451), .ZN(n15570) );
  NOR2_X1 U18703 ( .A1(n15570), .A2(n15569), .ZN(n15575) );
  INV_X1 U18704 ( .A(n15571), .ZN(n15572) );
  NOR2_X1 U18705 ( .A1(n15573), .A2(n15572), .ZN(n15574) );
  XNOR2_X1 U18706 ( .A(n15575), .B(n15574), .ZN(n15813) );
  NOR2_X1 U18707 ( .A1(n15807), .A2(n16648), .ZN(n15579) );
  NAND2_X1 U18708 ( .A1(n19529), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n15805) );
  NAND2_X1 U18709 ( .A1(n19530), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15576) );
  OAI211_X1 U18710 ( .C1(n19542), .C2(n15577), .A(n15805), .B(n15576), .ZN(
        n15578) );
  AOI211_X1 U18711 ( .C1(n15813), .C2(n16662), .A(n15579), .B(n15578), .ZN(
        n15580) );
  OAI21_X1 U18712 ( .B1(n19532), .B2(n15815), .A(n15580), .ZN(P2_U3002) );
  INV_X1 U18713 ( .A(n15550), .ZN(n15581) );
  XNOR2_X1 U18714 ( .A(n16638), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15827) );
  NAND2_X1 U18715 ( .A1(n15582), .A2(n15828), .ZN(n15585) );
  NAND2_X1 U18716 ( .A1(n9776), .A2(n15583), .ZN(n15584) );
  XNOR2_X1 U18717 ( .A(n15585), .B(n15584), .ZN(n15825) );
  NAND2_X1 U18718 ( .A1(n19347), .A2(n19538), .ZN(n15587) );
  INV_X1 U18719 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20166) );
  NOR2_X1 U18720 ( .A1(n15727), .A2(n20166), .ZN(n15821) );
  AOI21_X1 U18721 ( .B1(n19530), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15821), .ZN(n15586) );
  OAI211_X1 U18722 ( .C1(n19542), .C2(n19345), .A(n15587), .B(n15586), .ZN(
        n15588) );
  AOI21_X1 U18723 ( .B1(n15825), .B2(n16662), .A(n15588), .ZN(n15589) );
  OAI21_X1 U18724 ( .B1(n15827), .B2(n19532), .A(n15589), .ZN(P2_U3004) );
  OAI21_X1 U18725 ( .B1(n15592), .B2(n15591), .A(n15590), .ZN(n15593) );
  INV_X1 U18726 ( .A(n15593), .ZN(n16691) );
  INV_X1 U18727 ( .A(n15842), .ZN(n15595) );
  OR2_X1 U18728 ( .A1(n15594), .A2(n15595), .ZN(n15596) );
  NAND2_X1 U18729 ( .A1(n15596), .A2(n15843), .ZN(n15600) );
  AND2_X1 U18730 ( .A1(n15598), .A2(n15597), .ZN(n15599) );
  XNOR2_X1 U18731 ( .A(n15600), .B(n15599), .ZN(n16694) );
  AOI22_X1 U18732 ( .A1(n19538), .A2(n19359), .B1(n19530), .B2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15603) );
  INV_X1 U18733 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20162) );
  OAI22_X1 U18734 ( .A1(n20162), .A2(n19363), .B1(n19542), .B2(n19357), .ZN(
        n15601) );
  INV_X1 U18735 ( .A(n15601), .ZN(n15602) );
  OAI211_X1 U18736 ( .C1(n16694), .C2(n19534), .A(n15603), .B(n15602), .ZN(
        n15604) );
  AOI21_X1 U18737 ( .B1(n16691), .B2(n16660), .A(n15604), .ZN(n15605) );
  INV_X1 U18738 ( .A(n15605), .ZN(P2_U3006) );
  INV_X1 U18739 ( .A(n16542), .ZN(n15610) );
  INV_X1 U18740 ( .A(n15627), .ZN(n15608) );
  NOR3_X1 U18741 ( .A1(n15608), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15607), .ZN(n15609) );
  AOI21_X1 U18742 ( .B1(n15614), .B2(n16690), .A(n15613), .ZN(n15615) );
  OAI21_X1 U18743 ( .B1(n15616), .B2(n16697), .A(n15615), .ZN(P2_U3017) );
  INV_X1 U18744 ( .A(n15617), .ZN(n15630) );
  INV_X1 U18745 ( .A(n15618), .ZN(n15620) );
  NAND3_X1 U18746 ( .A1(n15620), .A2(n16673), .A3(n15619), .ZN(n15629) );
  NOR2_X1 U18747 ( .A1(n15621), .A2(n15626), .ZN(n15625) );
  NAND2_X1 U18748 ( .A1(n16565), .A2(n16669), .ZN(n15622) );
  OAI211_X1 U18749 ( .C1(n16567), .C2(n16702), .A(n15623), .B(n15622), .ZN(
        n15624) );
  AOI211_X1 U18750 ( .C1(n15627), .C2(n15626), .A(n15625), .B(n15624), .ZN(
        n15628) );
  OAI211_X1 U18751 ( .C1(n15630), .C2(n16710), .A(n15629), .B(n15628), .ZN(
        P2_U3019) );
  INV_X1 U18752 ( .A(n15631), .ZN(n15632) );
  AOI211_X1 U18753 ( .C1(n15633), .C2(n15648), .A(n15632), .B(n15642), .ZN(
        n15638) );
  AOI21_X1 U18754 ( .B1(n16578), .B2(n16669), .A(n15634), .ZN(n15636) );
  NAND3_X1 U18755 ( .A1(n15643), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15816), .ZN(n15635) );
  OAI211_X1 U18756 ( .C1(n16577), .C2(n16702), .A(n15636), .B(n15635), .ZN(
        n15637) );
  AOI211_X1 U18757 ( .C1(n15639), .C2(n16673), .A(n15638), .B(n15637), .ZN(
        n15640) );
  OAI21_X1 U18758 ( .B1(n16710), .B2(n15641), .A(n15640), .ZN(P2_U3020) );
  INV_X1 U18759 ( .A(n15642), .ZN(n15649) );
  INV_X1 U18760 ( .A(n15643), .ZN(n15659) );
  NOR3_X1 U18761 ( .A1(n15659), .A2(n15701), .A3(n15648), .ZN(n15647) );
  NAND2_X1 U18762 ( .A1(n16588), .A2(n16669), .ZN(n15644) );
  OAI211_X1 U18763 ( .C1(n16590), .C2(n16702), .A(n15645), .B(n15644), .ZN(
        n15646) );
  AOI211_X1 U18764 ( .C1(n15649), .C2(n15648), .A(n15647), .B(n15646), .ZN(
        n15652) );
  NAND2_X1 U18765 ( .A1(n15650), .A2(n16690), .ZN(n15651) );
  OAI211_X1 U18766 ( .C1(n15653), .C2(n16697), .A(n15652), .B(n15651), .ZN(
        P2_U3021) );
  AOI21_X1 U18767 ( .B1(n15676), .B2(n15654), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15660) );
  INV_X1 U18768 ( .A(n16602), .ZN(n15657) );
  NOR2_X1 U18769 ( .A1(n16601), .A2(n16701), .ZN(n15655) );
  AOI211_X1 U18770 ( .C1(n15657), .C2(n16689), .A(n15656), .B(n15655), .ZN(
        n15658) );
  OAI21_X1 U18771 ( .B1(n15660), .B2(n15659), .A(n15658), .ZN(n15661) );
  AOI21_X1 U18772 ( .B1(n15662), .B2(n16673), .A(n15661), .ZN(n15663) );
  OAI21_X1 U18773 ( .B1(n16710), .B2(n15664), .A(n15663), .ZN(P2_U3022) );
  OAI211_X1 U18774 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15676), .B(n15665), .ZN(
        n15670) );
  NOR2_X1 U18775 ( .A1(n15666), .A2(n16702), .ZN(n15667) );
  AOI211_X1 U18776 ( .C1(n16669), .C2(n16612), .A(n15668), .B(n15667), .ZN(
        n15669) );
  OAI211_X1 U18777 ( .C1(n15677), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        n15672) );
  AOI21_X1 U18778 ( .B1(n15673), .B2(n16673), .A(n15672), .ZN(n15674) );
  OAI21_X1 U18779 ( .B1(n16710), .B2(n15675), .A(n15674), .ZN(P2_U3023) );
  INV_X1 U18780 ( .A(n15676), .ZN(n15684) );
  INV_X1 U18781 ( .A(n15677), .ZN(n15697) );
  NOR2_X1 U18782 ( .A1(n15678), .A2(n16702), .ZN(n15682) );
  OAI21_X1 U18783 ( .B1(n15680), .B2(n16701), .A(n15679), .ZN(n15681) );
  AOI211_X1 U18784 ( .C1(n15697), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15682), .B(n15681), .ZN(n15683) );
  OAI21_X1 U18785 ( .B1(n15684), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15683), .ZN(n15685) );
  AOI21_X1 U18786 ( .B1(n15686), .B2(n16673), .A(n15685), .ZN(n15687) );
  OAI21_X1 U18787 ( .B1(n15688), .B2(n16710), .A(n15687), .ZN(P2_U3024) );
  NAND2_X1 U18788 ( .A1(n15689), .A2(n16673), .ZN(n15699) );
  NAND2_X1 U18789 ( .A1(n15690), .A2(n16689), .ZN(n15692) );
  OAI211_X1 U18790 ( .C1(n16701), .C2(n15693), .A(n15692), .B(n15691), .ZN(
        n15696) );
  NOR3_X1 U18791 ( .A1(n15721), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15694), .ZN(n15695) );
  AOI211_X1 U18792 ( .C1(n15697), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15696), .B(n15695), .ZN(n15698) );
  OAI211_X1 U18793 ( .C1(n15700), .C2(n16710), .A(n15699), .B(n15698), .ZN(
        P2_U3025) );
  AOI21_X1 U18794 ( .B1(n15831), .B2(n15702), .A(n15701), .ZN(n15734) );
  AOI21_X1 U18795 ( .B1(n19296), .B2(n16669), .A(n15703), .ZN(n15704) );
  OAI21_X1 U18796 ( .B1(n15705), .B2(n16702), .A(n15704), .ZN(n15710) );
  AOI211_X1 U18797 ( .C1(n15708), .C2(n15707), .A(n15706), .B(n15721), .ZN(
        n15709) );
  AOI211_X1 U18798 ( .C1(n15734), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15710), .B(n15709), .ZN(n15713) );
  NAND2_X1 U18799 ( .A1(n15711), .A2(n16690), .ZN(n15712) );
  OAI211_X1 U18800 ( .C1(n15714), .C2(n16697), .A(n15713), .B(n15712), .ZN(
        P2_U3026) );
  AOI21_X1 U18801 ( .B1(n15716), .B2(n16669), .A(n15715), .ZN(n15717) );
  OAI21_X1 U18802 ( .B1(n15718), .B2(n16702), .A(n15717), .ZN(n15719) );
  AOI21_X1 U18803 ( .B1(n15734), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15719), .ZN(n15720) );
  OAI21_X1 U18804 ( .B1(n15721), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15720), .ZN(n15722) );
  AOI21_X1 U18805 ( .B1(n15723), .B2(n16673), .A(n15722), .ZN(n15724) );
  OAI21_X1 U18806 ( .B1(n16710), .B2(n15725), .A(n15724), .ZN(P2_U3027) );
  NOR3_X1 U18807 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15750), .A3(
        n15818), .ZN(n15730) );
  NOR2_X1 U18808 ( .A1(n20180), .A2(n15727), .ZN(n15729) );
  NOR2_X1 U18809 ( .A1(n19315), .A2(n16701), .ZN(n15728) );
  AOI211_X1 U18810 ( .C1(n10885), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        n15731) );
  OAI21_X1 U18811 ( .B1(n15732), .B2(n16702), .A(n15731), .ZN(n15733) );
  AOI21_X1 U18812 ( .B1(n15734), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15733), .ZN(n15737) );
  NAND2_X1 U18813 ( .A1(n15735), .A2(n16690), .ZN(n15736) );
  OAI211_X1 U18814 ( .C1(n15738), .C2(n16697), .A(n15737), .B(n15736), .ZN(
        P2_U3028) );
  OAI21_X1 U18815 ( .B1(n16690), .B2(n15740), .A(n15739), .ZN(n15742) );
  NAND2_X1 U18816 ( .A1(n16705), .A2(n15750), .ZN(n15741) );
  AND2_X1 U18817 ( .A1(n15831), .A2(n15741), .ZN(n15766) );
  OAI211_X1 U18818 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15743), .A(
        n15742), .B(n15766), .ZN(n15756) );
  AOI21_X1 U18819 ( .B1(n15764), .B2(n16705), .A(n15756), .ZN(n15755) );
  NOR2_X1 U18820 ( .A1(n15744), .A2(n16702), .ZN(n15748) );
  OAI21_X1 U18821 ( .B1(n15746), .B2(n16701), .A(n15745), .ZN(n15747) );
  AOI211_X1 U18822 ( .C1(n15749), .C2(n16673), .A(n15748), .B(n15747), .ZN(
        n15753) );
  OR2_X1 U18823 ( .A1(n15818), .A2(n15750), .ZN(n15773) );
  OAI21_X1 U18824 ( .B1(n15510), .B2(n16710), .A(n15773), .ZN(n15761) );
  NAND3_X1 U18825 ( .A1(n15761), .A2(n15751), .A3(n15754), .ZN(n15752) );
  OAI211_X1 U18826 ( .C1(n15755), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        P2_U3029) );
  INV_X1 U18827 ( .A(n15756), .ZN(n15765) );
  NOR2_X1 U18828 ( .A1(n19319), .A2(n16702), .ZN(n15759) );
  OAI21_X1 U18829 ( .B1(n16701), .B2(n19326), .A(n15757), .ZN(n15758) );
  AOI211_X1 U18830 ( .C1(n15760), .C2(n16673), .A(n15759), .B(n15758), .ZN(
        n15763) );
  NAND3_X1 U18831 ( .A1(n15761), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n15764), .ZN(n15762) );
  OAI211_X1 U18832 ( .C1(n15765), .C2(n15764), .A(n15763), .B(n15762), .ZN(
        P2_U3030) );
  INV_X1 U18833 ( .A(n15766), .ZN(n15771) );
  AOI21_X1 U18834 ( .B1(n16669), .B2(n19425), .A(n15767), .ZN(n15768) );
  OAI21_X1 U18835 ( .B1(n15769), .B2(n16702), .A(n15768), .ZN(n15770) );
  AOI21_X1 U18836 ( .B1(n15771), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15770), .ZN(n15772) );
  OAI21_X1 U18837 ( .B1(n15773), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15772), .ZN(n15774) );
  AOI21_X1 U18838 ( .B1(n15775), .B2(n16673), .A(n15774), .ZN(n15776) );
  OAI21_X1 U18839 ( .B1(n16710), .B2(n15777), .A(n15776), .ZN(P2_U3031) );
  INV_X1 U18840 ( .A(n15818), .ZN(n15837) );
  NAND2_X1 U18841 ( .A1(n15837), .A2(n15778), .ZN(n15811) );
  NAND2_X1 U18842 ( .A1(n15831), .A2(n15778), .ZN(n15779) );
  NAND2_X1 U18843 ( .A1(n15779), .A2(n15816), .ZN(n15804) );
  OAI21_X1 U18844 ( .B1(n15811), .B2(n15780), .A(n15804), .ZN(n15793) );
  OAI21_X1 U18845 ( .B1(n11284), .B2(n10254), .A(n15782), .ZN(n19432) );
  NAND2_X1 U18846 ( .A1(n19336), .A2(n16689), .ZN(n15784) );
  OAI211_X1 U18847 ( .C1(n16701), .C2(n19432), .A(n15784), .B(n15783), .ZN(
        n15787) );
  NOR3_X1 U18848 ( .A1(n15811), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15785), .ZN(n15786) );
  AOI211_X1 U18849 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15793), .A(
        n15787), .B(n15786), .ZN(n15790) );
  NAND2_X1 U18850 ( .A1(n15788), .A2(n16690), .ZN(n15789) );
  OAI211_X1 U18851 ( .C1(n15791), .C2(n16697), .A(n15790), .B(n15789), .ZN(
        P2_U3032) );
  NOR2_X1 U18852 ( .A1(n15811), .A2(n15792), .ZN(n15794) );
  OAI21_X1 U18853 ( .B1(n15794), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15793), .ZN(n15799) );
  INV_X1 U18854 ( .A(n15795), .ZN(n15797) );
  AOI21_X1 U18855 ( .B1(n15797), .B2(n16689), .A(n15796), .ZN(n15798) );
  OAI211_X1 U18856 ( .C1(n16701), .C2(n19435), .A(n15799), .B(n15798), .ZN(
        n15800) );
  AOI21_X1 U18857 ( .B1(n15801), .B2(n16673), .A(n15800), .ZN(n15802) );
  OAI21_X1 U18858 ( .B1(n15803), .B2(n16710), .A(n15802), .ZN(P2_U3033) );
  INV_X1 U18859 ( .A(n15804), .ZN(n15809) );
  NAND2_X1 U18860 ( .A1(n16669), .A2(n19436), .ZN(n15806) );
  OAI211_X1 U18861 ( .C1(n15807), .C2(n16702), .A(n15806), .B(n15805), .ZN(
        n15808) );
  AOI21_X1 U18862 ( .B1(n15809), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15808), .ZN(n15810) );
  OAI21_X1 U18863 ( .B1(n15811), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15810), .ZN(n15812) );
  AOI21_X1 U18864 ( .B1(n15813), .B2(n16673), .A(n15812), .ZN(n15814) );
  OAI21_X1 U18865 ( .B1(n15815), .B2(n16710), .A(n15814), .ZN(P2_U3034) );
  INV_X1 U18866 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16676) );
  INV_X1 U18867 ( .A(n15831), .ZN(n15817) );
  OAI21_X1 U18868 ( .B1(n15817), .B2(n15836), .A(n15816), .ZN(n16668) );
  NOR2_X1 U18869 ( .A1(n15818), .A2(n15836), .ZN(n16675) );
  NAND2_X1 U18870 ( .A1(n16675), .A2(n16676), .ZN(n15823) );
  OAI21_X1 U18871 ( .B1(n13325), .B2(n15819), .A(n9753), .ZN(n19444) );
  NOR2_X1 U18872 ( .A1(n16701), .A2(n19444), .ZN(n15820) );
  AOI211_X1 U18873 ( .C1(n19347), .C2(n16689), .A(n15821), .B(n15820), .ZN(
        n15822) );
  OAI211_X1 U18874 ( .C1(n16676), .C2(n16668), .A(n15823), .B(n15822), .ZN(
        n15824) );
  AOI21_X1 U18875 ( .B1(n15825), .B2(n16673), .A(n15824), .ZN(n15826) );
  OAI21_X1 U18876 ( .B1(n15827), .B2(n16710), .A(n15826), .ZN(P2_U3036) );
  NAND2_X1 U18877 ( .A1(n15829), .A2(n15828), .ZN(n15830) );
  XOR2_X1 U18878 ( .A(n15830), .B(n9747), .Z(n16640) );
  NOR2_X1 U18879 ( .A1(n15550), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16637) );
  OR3_X1 U18880 ( .A1(n16638), .A2(n16637), .A3(n16710), .ZN(n15839) );
  NOR2_X1 U18881 ( .A1(n15831), .A2(n15836), .ZN(n15835) );
  NAND2_X1 U18882 ( .A1(n16669), .A2(n19445), .ZN(n15833) );
  NAND2_X1 U18883 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19529), .ZN(n15832) );
  OAI211_X1 U18884 ( .C1(n16639), .C2(n16702), .A(n15833), .B(n15832), .ZN(
        n15834) );
  AOI211_X1 U18885 ( .C1(n15837), .C2(n15836), .A(n15835), .B(n15834), .ZN(
        n15838) );
  OAI211_X1 U18886 ( .C1(n16640), .C2(n16697), .A(n15839), .B(n15838), .ZN(
        P2_U3037) );
  OR2_X1 U18887 ( .A1(n15840), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16647) );
  NAND3_X1 U18888 ( .A1(n16647), .A2(n16690), .A3(n15841), .ZN(n15852) );
  AND2_X1 U18889 ( .A1(n15843), .A2(n15842), .ZN(n15844) );
  XNOR2_X1 U18890 ( .A(n15594), .B(n15844), .ZN(n16651) );
  NAND2_X1 U18891 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15847), .ZN(
        n16681) );
  AOI21_X1 U18892 ( .B1(n15847), .B2(n15846), .A(n15845), .ZN(n16686) );
  NAND2_X1 U18893 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19529), .ZN(n15848) );
  OAI221_X1 U18894 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16681), .C1(
        n16682), .C2(n16686), .A(n15848), .ZN(n15850) );
  OAI22_X1 U18895 ( .A1(n19452), .A2(n16701), .B1(n16702), .B2(n16649), .ZN(
        n15849) );
  AOI211_X1 U18896 ( .C1(n16651), .C2(n16673), .A(n15850), .B(n15849), .ZN(
        n15851) );
  NAND2_X1 U18897 ( .A1(n15852), .A2(n15851), .ZN(P2_U3039) );
  INV_X1 U18898 ( .A(n20219), .ZN(n20225) );
  AND2_X1 U18899 ( .A1(n15854), .A2(n15853), .ZN(n15877) );
  INV_X1 U18900 ( .A(n15877), .ZN(n15855) );
  MUX2_X1 U18901 ( .A(n15855), .B(n10390), .S(n15871), .Z(n15856) );
  AOI21_X1 U18902 ( .B1(n15857), .B2(n15912), .A(n15856), .ZN(n16734) );
  INV_X1 U18903 ( .A(n15875), .ZN(n19401) );
  AOI22_X1 U18904 ( .A1(n19379), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19401), .B2(n9661), .ZN(n15872) );
  INV_X1 U18905 ( .A(n15872), .ZN(n15858) );
  OAI222_X1 U18906 ( .A1(n20256), .A2(n16761), .B1(n20225), .B2(n16734), .C1(
        n15859), .C2(n15858), .ZN(n15870) );
  OR2_X1 U18907 ( .A1(n15860), .A2(n16729), .ZN(n15867) );
  NAND2_X1 U18908 ( .A1(n16728), .A2(n16726), .ZN(n15861) );
  OR2_X1 U18909 ( .A1(n16725), .A2(n15861), .ZN(n15862) );
  AND4_X1 U18910 ( .A1(n15865), .A2(n15864), .A3(n15863), .A4(n15862), .ZN(
        n15866) );
  NAND2_X1 U18911 ( .A1(n15867), .A2(n15866), .ZN(n16752) );
  NAND2_X1 U18912 ( .A1(n16752), .A2(n20122), .ZN(n15869) );
  NOR2_X1 U18913 ( .A1(n20278), .A2(n20253), .ZN(n16769) );
  AOI22_X1 U18914 ( .A1(n16769), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n20278), .ZN(n15868) );
  NAND2_X1 U18915 ( .A1(n15869), .A2(n15868), .ZN(n20222) );
  MUX2_X1 U18916 ( .A(n15871), .B(n15870), .S(n20222), .Z(P2_U3601) );
  NOR2_X1 U18917 ( .A1(n15872), .A2(n15859), .ZN(n15896) );
  INV_X1 U18918 ( .A(n15896), .ZN(n15880) );
  OAI21_X1 U18919 ( .B1(n15875), .B2(n15874), .A(n15873), .ZN(n19400) );
  OAI21_X1 U18920 ( .B1(n9661), .B2(n10594), .A(n19400), .ZN(n15897) );
  INV_X1 U18921 ( .A(n10390), .ZN(n15908) );
  NOR2_X1 U18922 ( .A1(n15908), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15879) );
  NOR3_X1 U18923 ( .A1(n15877), .A2(n15876), .A3(n15883), .ZN(n15878) );
  AOI211_X1 U18924 ( .C1(n10437), .C2(n15912), .A(n15879), .B(n15878), .ZN(
        n16733) );
  OAI222_X1 U18925 ( .A1(n16761), .A2(n20227), .B1(n15880), .B2(n15897), .C1(
        n20225), .C2(n16733), .ZN(n15881) );
  MUX2_X1 U18926 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15881), .S(
        n20222), .Z(P2_U3600) );
  OR2_X1 U18927 ( .A1(n15882), .A2(n16718), .ZN(n15900) );
  INV_X1 U18928 ( .A(n15883), .ZN(n15884) );
  NAND2_X1 U18929 ( .A1(n15884), .A2(n10572), .ZN(n15905) );
  NAND2_X1 U18930 ( .A1(n15903), .A2(n15905), .ZN(n15887) );
  NAND2_X1 U18931 ( .A1(n15900), .A2(n15887), .ZN(n15892) );
  NAND2_X1 U18932 ( .A1(n15886), .A2(n15885), .ZN(n15904) );
  INV_X1 U18933 ( .A(n15887), .ZN(n15890) );
  NOR2_X1 U18934 ( .A1(n15888), .A2(n15907), .ZN(n15889) );
  AOI22_X1 U18935 ( .A1(n15904), .A2(n15890), .B1(n10390), .B2(n15889), .ZN(
        n15891) );
  NAND2_X1 U18936 ( .A1(n15892), .A2(n15891), .ZN(n15893) );
  AOI21_X1 U18937 ( .B1(n15894), .B2(n15912), .A(n15893), .ZN(n16737) );
  OAI22_X1 U18938 ( .A1(n20239), .A2(n16761), .B1(n16737), .B2(n20225), .ZN(
        n15895) );
  AOI21_X1 U18939 ( .B1(n15897), .B2(n15896), .A(n15895), .ZN(n15898) );
  MUX2_X1 U18940 ( .A(n10572), .B(n15898), .S(n20222), .Z(n15899) );
  INV_X1 U18941 ( .A(n15899), .ZN(P2_U3599) );
  INV_X1 U18942 ( .A(n15907), .ZN(n15902) );
  NAND2_X1 U18943 ( .A1(n15900), .A2(n15905), .ZN(n15901) );
  OAI211_X1 U18944 ( .C1(n15908), .C2(n15902), .A(n15901), .B(n15903), .ZN(
        n15910) );
  NAND2_X1 U18945 ( .A1(n15904), .A2(n15903), .ZN(n15906) );
  OAI211_X1 U18946 ( .C1(n15908), .C2(n15907), .A(n15906), .B(n15905), .ZN(
        n15909) );
  MUX2_X1 U18947 ( .A(n15910), .B(n15909), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15911) );
  OAI22_X1 U18948 ( .A1(n19860), .A2(n16761), .B1(n16740), .B2(n20225), .ZN(
        n15913) );
  MUX2_X1 U18949 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15913), .S(
        n20222), .Z(P2_U3596) );
  AOI22_X1 U18950 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15917) );
  AOI22_X1 U18951 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n17574), .B1(
        n17562), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15916) );
  AOI22_X1 U18952 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15915) );
  AOI22_X1 U18953 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15914) );
  NAND4_X1 U18954 ( .A1(n15917), .A2(n15916), .A3(n15915), .A4(n15914), .ZN(
        n15923) );
  AOI22_X1 U18955 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15921) );
  AOI22_X1 U18956 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15920) );
  AOI22_X1 U18957 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15919) );
  AOI22_X1 U18958 ( .A1(n13949), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15918) );
  NAND4_X1 U18959 ( .A1(n15921), .A2(n15920), .A3(n15919), .A4(n15918), .ZN(
        n15922) );
  NOR2_X1 U18960 ( .A1(n15923), .A2(n15922), .ZN(n17727) );
  INV_X1 U18961 ( .A(n17521), .ZN(n15924) );
  OAI33_X1 U18962 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17717), .A3(n17521), 
        .B1(n17168), .B2(n17625), .B3(n15924), .ZN(n15925) );
  INV_X1 U18963 ( .A(n15925), .ZN(n15926) );
  OAI21_X1 U18964 ( .B1(n17727), .B2(n17619), .A(n15926), .ZN(P3_U2690) );
  NAND2_X1 U18965 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18749) );
  INV_X1 U18966 ( .A(n19255), .ZN(n18600) );
  NOR2_X1 U18967 ( .A1(n19107), .A2(n18600), .ZN(n15928) );
  AOI221_X1 U18968 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18749), .C1(n15928), 
        .C2(n18749), .A(n15927), .ZN(n18603) );
  NOR2_X1 U18969 ( .A1(n15929), .A2(n19074), .ZN(n15930) );
  OAI21_X1 U18970 ( .B1(n15930), .B2(n18662), .A(n18604), .ZN(n18601) );
  AOI22_X1 U18971 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18603), .B1(
        n18601), .B2(n19079), .ZN(P3_U2865) );
  NAND2_X1 U18972 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19093) );
  INV_X1 U18973 ( .A(n19093), .ZN(n19252) );
  XOR2_X1 U18974 ( .A(n15932), .B(n15931), .Z(n15935) );
  INV_X1 U18975 ( .A(n19041), .ZN(n16109) );
  NOR2_X1 U18976 ( .A1(n19252), .A2(n16109), .ZN(n15948) );
  NAND4_X1 U18977 ( .A1(n15966), .A2(n18629), .A3(n15950), .A4(n17786), .ZN(
        n15956) );
  OR2_X2 U18978 ( .A1(n18629), .A2(n18633), .ZN(n15941) );
  NOR4_X2 U18979 ( .A1(n15953), .A2(n16114), .A3(n15955), .A4(n15941), .ZN(
        n19050) );
  NAND2_X1 U18980 ( .A1(n19050), .A2(n16101), .ZN(n15945) );
  NAND2_X1 U18981 ( .A1(n15956), .A2(n15945), .ZN(n16945) );
  INV_X1 U18982 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19122) );
  INV_X2 U18983 ( .A(n19258), .ZN(n19260) );
  NAND2_X2 U18984 ( .A1(n19260), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19187) );
  OAI211_X1 U18985 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19122), .B(n19187), .ZN(n19116) );
  INV_X1 U18986 ( .A(n19069), .ZN(n15936) );
  INV_X1 U18987 ( .A(n16101), .ZN(n18617) );
  OAI21_X1 U18988 ( .B1(n18613), .B2(n17786), .A(n18617), .ZN(n15940) );
  AOI21_X1 U18989 ( .B1(n16114), .B2(n15936), .A(n15940), .ZN(n15938) );
  NAND3_X1 U18990 ( .A1(n15966), .A2(n15938), .A3(n15937), .ZN(n16103) );
  AOI22_X1 U18991 ( .A1(n18621), .A2(n15955), .B1(n18625), .B2(n19069), .ZN(
        n15944) );
  AOI21_X1 U18992 ( .B1(n17717), .B2(n15941), .A(n18625), .ZN(n15939) );
  AOI21_X1 U18993 ( .B1(n15941), .B2(n15940), .A(n15939), .ZN(n15943) );
  NOR2_X1 U18994 ( .A1(n16101), .A2(n15941), .ZN(n16115) );
  OAI21_X1 U18995 ( .B1(n15950), .B2(n16115), .A(n18609), .ZN(n15942) );
  NAND3_X1 U18996 ( .A1(n15944), .A2(n15943), .A3(n15942), .ZN(n15951) );
  OAI21_X1 U18997 ( .B1(n16103), .B2(n15951), .A(n15945), .ZN(n15946) );
  NOR2_X1 U18998 ( .A1(n18639), .A2(n19069), .ZN(n16213) );
  OR3_X1 U18999 ( .A1(n19246), .A2(n18609), .A3(n16213), .ZN(n15949) );
  NAND2_X1 U19000 ( .A1(n15946), .A2(n15949), .ZN(n16111) );
  AOI211_X1 U19001 ( .C1(n15948), .C2(n17784), .A(n15947), .B(n16111), .ZN(
        n15960) );
  OAI21_X1 U19002 ( .B1(n16110), .B2(n15950), .A(n15949), .ZN(n15952) );
  NAND2_X1 U19003 ( .A1(n19050), .A2(n15969), .ZN(n15970) );
  NOR2_X1 U19004 ( .A1(n15955), .A2(n15954), .ZN(n15958) );
  NAND2_X1 U19005 ( .A1(n17827), .A2(n19246), .ZN(n15959) );
  NAND2_X1 U19006 ( .A1(n16960), .A2(n15959), .ZN(n15957) );
  INV_X1 U19007 ( .A(n19055), .ZN(n15962) );
  NAND3_X1 U19008 ( .A1(n19041), .A2(n19093), .A3(n16961), .ZN(n16212) );
  NAND2_X1 U19009 ( .A1(n15960), .A2(n16212), .ZN(n19067) );
  NOR2_X1 U19010 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19202), .ZN(n18608) );
  INV_X1 U19011 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18598) );
  NOR2_X1 U19012 ( .A1(n18598), .A2(n19200), .ZN(n15961) );
  AOI211_X1 U19013 ( .C1(n19090), .C2(n19067), .A(n18608), .B(n15961), .ZN(
        n19233) );
  INV_X1 U19014 ( .A(n19233), .ZN(n19230) );
  NOR2_X1 U19015 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19262) );
  NOR3_X1 U19016 ( .A1(n15963), .A2(n15962), .A3(n15970), .ZN(n19089) );
  NAND3_X1 U19017 ( .A1(n19230), .A2(n19262), .A3(n19089), .ZN(n15964) );
  OAI21_X1 U19018 ( .B1(n19230), .B2(n21004), .A(n15964), .ZN(P3_U3284) );
  INV_X1 U19019 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18286) );
  INV_X1 U19020 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17935) );
  NOR2_X1 U19021 ( .A1(n18286), .A2(n17935), .ZN(n18260) );
  NOR2_X2 U19022 ( .A1(n19265), .A2(n15965), .ZN(n19066) );
  INV_X1 U19023 ( .A(n19066), .ZN(n18537) );
  INV_X1 U19024 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18380) );
  INV_X1 U19025 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18378) );
  NOR2_X1 U19026 ( .A1(n18380), .A2(n18378), .ZN(n18370) );
  INV_X1 U19027 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18030) );
  INV_X1 U19028 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18364) );
  INV_X1 U19029 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18351) );
  NOR2_X1 U19030 ( .A1(n18364), .A2(n18351), .ZN(n18336) );
  NAND2_X1 U19031 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18336), .ZN(
        n18318) );
  INV_X1 U19032 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18327) );
  NOR3_X1 U19033 ( .A1(n18030), .A2(n18318), .A3(n18327), .ZN(n16135) );
  NAND2_X1 U19034 ( .A1(n18370), .A2(n16135), .ZN(n18310) );
  INV_X1 U19035 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18142) );
  NOR2_X1 U19036 ( .A1(n18484), .A2(n18142), .ZN(n18456) );
  NAND2_X1 U19037 ( .A1(n18456), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18444) );
  NAND2_X1 U19038 ( .A1(n18411), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18417) );
  INV_X1 U19039 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18420) );
  NOR2_X1 U19040 ( .A1(n18417), .A2(n18420), .ZN(n16100) );
  INV_X1 U19041 ( .A(n16100), .ZN(n18399) );
  INV_X1 U19042 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18410) );
  INV_X1 U19043 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18526) );
  INV_X1 U19044 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18524) );
  NOR3_X1 U19045 ( .A1(n18526), .A2(n18524), .A3(n18549), .ZN(n18493) );
  INV_X1 U19046 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20997) );
  INV_X1 U19047 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19211) );
  INV_X1 U19048 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18562) );
  OAI21_X1 U19049 ( .B1(n20997), .B2(n19211), .A(n18562), .ZN(n18536) );
  NAND2_X1 U19050 ( .A1(n18493), .A2(n18536), .ZN(n18486) );
  NOR4_X1 U19051 ( .A1(n21015), .A2(n18514), .A3(n18518), .A4(n18486), .ZN(
        n18386) );
  NAND2_X1 U19052 ( .A1(n18366), .A2(n18386), .ZN(n18367) );
  NOR2_X1 U19053 ( .A1(n18310), .A2(n18367), .ZN(n18299) );
  INV_X1 U19054 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18316) );
  INV_X1 U19055 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18302) );
  NOR2_X1 U19056 ( .A1(n18316), .A2(n18302), .ZN(n17934) );
  NAND2_X1 U19057 ( .A1(n18299), .A2(n17934), .ZN(n18279) );
  INV_X1 U19058 ( .A(n15966), .ZN(n15967) );
  NAND3_X1 U19059 ( .A1(n15967), .A2(n19246), .A3(n16960), .ZN(n15968) );
  NAND2_X1 U19060 ( .A1(n15969), .A2(n15968), .ZN(n19051) );
  AOI21_X1 U19061 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19068), .A(
        n18585), .ZN(n18492) );
  INV_X1 U19062 ( .A(n18493), .ZN(n18516) );
  NAND2_X1 U19063 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18534) );
  NOR2_X1 U19064 ( .A1(n18516), .A2(n18534), .ZN(n18489) );
  NAND3_X1 U19065 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n18489), .ZN(n18387) );
  NOR2_X1 U19066 ( .A1(n21015), .A2(n18387), .ZN(n18319) );
  NAND2_X1 U19067 ( .A1(n18366), .A2(n18319), .ZN(n18372) );
  NOR2_X1 U19068 ( .A1(n18310), .A2(n18372), .ZN(n18295) );
  NAND2_X1 U19069 ( .A1(n17934), .A2(n18295), .ZN(n18264) );
  OAI22_X1 U19070 ( .A1(n18537), .A2(n18279), .B1(n18492), .B2(n18264), .ZN(
        n18283) );
  NAND2_X1 U19071 ( .A1(n18260), .A2(n18283), .ZN(n16821) );
  INV_X1 U19072 ( .A(n16821), .ZN(n16119) );
  NOR2_X4 U19073 ( .A1(n18434), .A2(n19068), .ZN(n18491) );
  AOI22_X1 U19074 ( .A1(n17405), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15974) );
  AOI22_X1 U19075 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15973) );
  AOI22_X1 U19076 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15972) );
  AOI22_X1 U19077 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17562), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15971) );
  NAND4_X1 U19078 ( .A1(n15974), .A2(n15973), .A3(n15972), .A4(n15971), .ZN(
        n15980) );
  AOI22_X1 U19079 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15978) );
  AOI22_X1 U19080 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15977) );
  AOI22_X1 U19081 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15976) );
  AOI22_X1 U19082 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15975) );
  NAND4_X1 U19083 ( .A1(n15978), .A2(n15977), .A3(n15976), .A4(n15975), .ZN(
        n15979) );
  AOI22_X1 U19084 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15984) );
  AOI22_X1 U19085 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15983) );
  AOI22_X1 U19086 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n17571), .B1(
        n17562), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15982) );
  AOI22_X1 U19087 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15981) );
  NAND4_X1 U19088 ( .A1(n15984), .A2(n15983), .A3(n15982), .A4(n15981), .ZN(
        n15990) );
  AOI22_X1 U19089 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15988) );
  AOI22_X1 U19090 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17573), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15987) );
  AOI22_X1 U19091 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15986) );
  AOI22_X1 U19092 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15985) );
  NAND4_X1 U19093 ( .A1(n15988), .A2(n15987), .A3(n15986), .A4(n15985), .ZN(
        n15989) );
  AOI22_X1 U19094 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15994) );
  AOI22_X1 U19095 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16010), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15993) );
  AOI22_X1 U19096 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15992) );
  AOI22_X1 U19097 ( .A1(n13949), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13914), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15991) );
  NAND4_X1 U19098 ( .A1(n15994), .A2(n15993), .A3(n15992), .A4(n15991), .ZN(
        n15998) );
  AOI22_X1 U19099 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15997) );
  AOI22_X1 U19100 ( .A1(n17584), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17581), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15996) );
  AOI22_X1 U19101 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14024), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15995) );
  AOI22_X1 U19102 ( .A1(n13949), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n16010), .ZN(n16002) );
  AOI22_X1 U19103 ( .A1(n9676), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16001) );
  AOI22_X1 U19104 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16000) );
  AOI22_X1 U19105 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n13914), .ZN(n15999) );
  NAND4_X1 U19106 ( .A1(n16002), .A2(n16001), .A3(n16000), .A4(n15999), .ZN(
        n16008) );
  AOI22_X1 U19107 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U19108 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17580), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U19109 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n13896), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14024), .ZN(n16004) );
  AOI22_X1 U19110 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17554), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17555), .ZN(n16003) );
  NAND4_X1 U19111 ( .A1(n16006), .A2(n16005), .A3(n16004), .A4(n16003), .ZN(
        n16007) );
  NOR2_X2 U19112 ( .A1(n16008), .A2(n16007), .ZN(n16081) );
  NOR2_X1 U19113 ( .A1(n16056), .A2(n16081), .ZN(n16060) );
  AOI22_X1 U19114 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16017) );
  AOI22_X1 U19115 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17581), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16016) );
  AOI22_X1 U19116 ( .A1(n16010), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16011) );
  AOI22_X1 U19117 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13896), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16015) );
  AOI22_X1 U19118 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16014) );
  AOI22_X1 U19119 ( .A1(n16022), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13914), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16013) );
  AOI22_X1 U19120 ( .A1(n17584), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13891), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16012) );
  NOR2_X1 U19121 ( .A1(n16060), .A2(n16078), .ZN(n16054) );
  AOI22_X1 U19122 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16021) );
  AOI22_X1 U19123 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n9667), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16020) );
  AOI22_X1 U19124 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U19125 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16018) );
  NAND4_X1 U19126 ( .A1(n16021), .A2(n16020), .A3(n16019), .A4(n16018), .ZN(
        n16028) );
  AOI22_X1 U19127 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16026) );
  AOI22_X1 U19128 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16025) );
  AOI22_X1 U19129 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16024) );
  AOI22_X1 U19130 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16022), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16023) );
  NAND4_X1 U19131 ( .A1(n16026), .A2(n16025), .A3(n16024), .A4(n16023), .ZN(
        n16027) );
  NOR2_X1 U19132 ( .A1(n16054), .A2(n17765), .ZN(n16063) );
  AOI22_X1 U19133 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16038) );
  AOI22_X1 U19134 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U19135 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16029) );
  OAI21_X1 U19136 ( .B1(n21027), .B2(n9720), .A(n16029), .ZN(n16035) );
  AOI22_X1 U19137 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16033) );
  AOI22_X1 U19138 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17581), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16032) );
  AOI22_X1 U19139 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16031) );
  AOI22_X1 U19140 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16030) );
  NAND4_X1 U19141 ( .A1(n16033), .A2(n16032), .A3(n16031), .A4(n16030), .ZN(
        n16034) );
  AOI211_X1 U19142 ( .C1(n17574), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n16035), .B(n16034), .ZN(n16036) );
  NAND3_X1 U19143 ( .A1(n16038), .A2(n16037), .A3(n16036), .ZN(n16079) );
  NAND2_X1 U19144 ( .A1(n16063), .A2(n16079), .ZN(n16053) );
  NOR2_X1 U19145 ( .A1(n17758), .A2(n16053), .ZN(n16052) );
  AOI22_X1 U19146 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16050) );
  AOI22_X1 U19147 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16049) );
  AOI22_X1 U19148 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16039) );
  OAI21_X1 U19149 ( .B1(n20895), .B2(n16040), .A(n16039), .ZN(n16047) );
  AOI22_X1 U19150 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16045) );
  AOI22_X1 U19151 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16044) );
  AOI22_X1 U19152 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16043) );
  AOI22_X1 U19153 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16042) );
  NAND4_X1 U19154 ( .A1(n16045), .A2(n16044), .A3(n16043), .A4(n16042), .ZN(
        n16046) );
  AOI211_X1 U19155 ( .C1(n17575), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n16047), .B(n16046), .ZN(n16048) );
  NAND3_X1 U19156 ( .A1(n16050), .A2(n16049), .A3(n16048), .ZN(n16096) );
  NAND2_X1 U19157 ( .A1(n16052), .A2(n16096), .ZN(n16051) );
  NOR2_X1 U19158 ( .A1(n17751), .A2(n16051), .ZN(n16075) );
  XNOR2_X1 U19159 ( .A(n16051), .B(n16786), .ZN(n18176) );
  XNOR2_X1 U19160 ( .A(n16052), .B(n17755), .ZN(n16068) );
  XNOR2_X1 U19161 ( .A(n17758), .B(n16053), .ZN(n16066) );
  OR2_X1 U19162 ( .A1(n18526), .A2(n16066), .ZN(n16067) );
  XOR2_X1 U19163 ( .A(n17765), .B(n16054), .Z(n16055) );
  NAND2_X1 U19164 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16055), .ZN(
        n16062) );
  XNOR2_X1 U19165 ( .A(n18549), .B(n16055), .ZN(n18224) );
  AOI21_X1 U19166 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17775), .A(
        n18253), .ZN(n16058) );
  NOR2_X1 U19167 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17775), .ZN(
        n16057) );
  AOI221_X1 U19168 ( .B1(n18253), .B2(n17775), .C1(n16058), .C2(n20997), .A(
        n16057), .ZN(n16059) );
  NAND2_X1 U19169 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n16059), .ZN(
        n16061) );
  XNOR2_X1 U19170 ( .A(n18562), .B(n16059), .ZN(n18237) );
  XOR2_X1 U19171 ( .A(n17770), .B(n16060), .Z(n18236) );
  NAND2_X1 U19172 ( .A1(n18237), .A2(n18236), .ZN(n18235) );
  NAND2_X1 U19173 ( .A1(n16061), .A2(n18235), .ZN(n18223) );
  NAND2_X1 U19174 ( .A1(n18224), .A2(n18223), .ZN(n18222) );
  NOR2_X1 U19175 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n16064), .ZN(
        n16065) );
  INV_X1 U19176 ( .A(n16079), .ZN(n17762) );
  XNOR2_X1 U19177 ( .A(n16063), .B(n17762), .ZN(n18212) );
  XNOR2_X1 U19178 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n16064), .ZN(
        n18211) );
  NOR2_X1 U19179 ( .A1(n18212), .A2(n18211), .ZN(n18210) );
  NOR2_X1 U19180 ( .A1(n16065), .A2(n18210), .ZN(n18200) );
  XNOR2_X1 U19181 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n16066), .ZN(
        n18199) );
  NAND2_X1 U19182 ( .A1(n18200), .A2(n18199), .ZN(n18198) );
  NAND2_X1 U19183 ( .A1(n16067), .A2(n18198), .ZN(n16069) );
  NAND2_X1 U19184 ( .A1(n16068), .A2(n16069), .ZN(n16070) );
  XOR2_X1 U19185 ( .A(n16069), .B(n16068), .Z(n18191) );
  NAND2_X1 U19186 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18191), .ZN(
        n18190) );
  NAND2_X1 U19187 ( .A1(n16070), .A2(n18190), .ZN(n18177) );
  NOR2_X1 U19188 ( .A1(n18176), .A2(n18177), .ZN(n16071) );
  NOR2_X1 U19189 ( .A1(n16071), .A2(n18514), .ZN(n16072) );
  NAND2_X1 U19190 ( .A1(n16075), .A2(n16072), .ZN(n16077) );
  INV_X1 U19191 ( .A(n16072), .ZN(n16074) );
  NAND2_X1 U19192 ( .A1(n18176), .A2(n18177), .ZN(n18175) );
  NAND2_X1 U19193 ( .A1(n16075), .A2(n16074), .ZN(n16073) );
  OAI211_X1 U19194 ( .C1(n16075), .C2(n16074), .A(n18175), .B(n16073), .ZN(
        n18166) );
  NAND2_X1 U19195 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18166), .ZN(
        n16076) );
  NAND2_X2 U19196 ( .A1(n16077), .A2(n16076), .ZN(n18450) );
  NOR2_X1 U19197 ( .A1(n18316), .A2(n18310), .ZN(n16130) );
  NAND2_X1 U19198 ( .A1(n18396), .A2(n16130), .ZN(n18294) );
  NAND2_X1 U19199 ( .A1(n17944), .A2(n18260), .ZN(n17896) );
  NAND2_X1 U19200 ( .A1(n16078), .A2(n17775), .ZN(n16085) );
  NAND2_X1 U19201 ( .A1(n16080), .A2(n16079), .ZN(n16090) );
  XOR2_X1 U19202 ( .A(n16095), .B(n17755), .Z(n16094) );
  XNOR2_X1 U19203 ( .A(n16080), .B(n16079), .ZN(n16089) );
  NOR2_X1 U19204 ( .A1(n18562), .A2(n16083), .ZN(n16084) );
  NOR2_X1 U19205 ( .A1(n17775), .A2(n19211), .ZN(n16082) );
  XNOR2_X1 U19206 ( .A(n16081), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18246) );
  NAND2_X1 U19207 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18253), .ZN(
        n18252) );
  NOR2_X1 U19208 ( .A1(n18246), .A2(n18252), .ZN(n18245) );
  NOR2_X1 U19209 ( .A1(n16082), .A2(n18245), .ZN(n18234) );
  XNOR2_X1 U19210 ( .A(n17765), .B(n16085), .ZN(n16087) );
  NOR2_X1 U19211 ( .A1(n16086), .A2(n16087), .ZN(n16088) );
  XNOR2_X1 U19212 ( .A(n18524), .B(n16089), .ZN(n18216) );
  XNOR2_X1 U19213 ( .A(n17758), .B(n16090), .ZN(n16092) );
  XNOR2_X1 U19214 ( .A(n16092), .B(n16091), .ZN(n18202) );
  XNOR2_X1 U19215 ( .A(n18518), .B(n16094), .ZN(n18189) );
  NOR2_X1 U19216 ( .A1(n16097), .A2(n16098), .ZN(n16099) );
  NAND2_X1 U19217 ( .A1(n16100), .A2(n18453), .ZN(n18082) );
  NAND2_X1 U19218 ( .A1(n16130), .A2(n18397), .ZN(n18293) );
  NOR2_X1 U19219 ( .A1(n18613), .A2(n16101), .ZN(n16108) );
  NAND2_X1 U19220 ( .A1(n16108), .A2(n16102), .ZN(n16104) );
  NAND2_X1 U19221 ( .A1(n18507), .A2(n17751), .ZN(n18452) );
  OAI22_X1 U19222 ( .A1(n18451), .A2(n17896), .B1(n18263), .B2(n18452), .ZN(
        n16118) );
  INV_X1 U19223 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18267) );
  INV_X1 U19224 ( .A(n16104), .ZN(n16113) );
  AOI21_X1 U19225 ( .B1(n16106), .B2(n16105), .A(n16109), .ZN(n19042) );
  OAI21_X1 U19226 ( .B1(n18617), .B2(n19246), .A(n19116), .ZN(n16107) );
  OAI21_X1 U19227 ( .B1(n16108), .B2(n16107), .A(n19093), .ZN(n16944) );
  NOR3_X1 U19228 ( .A1(n16110), .A2(n16109), .A3(n16944), .ZN(n16112) );
  OAI21_X1 U19229 ( .B1(n16115), .B2(n16114), .A(n19038), .ZN(n16116) );
  NOR2_X1 U19230 ( .A1(n18267), .A2(n18498), .ZN(n18269) );
  OAI211_X1 U19231 ( .C1(n16119), .C2(n16118), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18269), .ZN(n16190) );
  NAND2_X1 U19232 ( .A1(n18260), .A2(n17934), .ZN(n16838) );
  INV_X1 U19233 ( .A(n16838), .ZN(n16793) );
  AOI21_X1 U19234 ( .B1(n18299), .B2(n16793), .A(n18537), .ZN(n18261) );
  NOR2_X1 U19235 ( .A1(n20997), .A2(n18267), .ZN(n16122) );
  NAND2_X1 U19236 ( .A1(n16793), .A2(n18295), .ZN(n16120) );
  OAI21_X1 U19237 ( .B1(n18585), .B2(n19068), .A(n16120), .ZN(n16121) );
  OAI21_X1 U19238 ( .B1(n9660), .B2(n16122), .A(n16121), .ZN(n16123) );
  NOR2_X1 U19239 ( .A1(n18261), .A2(n16123), .ZN(n16185) );
  OAI211_X1 U19240 ( .C1(n18465), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16185), .B(n18575), .ZN(n16836) );
  NOR2_X1 U19241 ( .A1(n18491), .A2(n18498), .ZN(n18538) );
  INV_X1 U19242 ( .A(n18538), .ZN(n18576) );
  NOR2_X1 U19243 ( .A1(n18498), .A2(n18452), .ZN(n18425) );
  NAND3_X1 U19244 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16822) );
  NOR2_X1 U19245 ( .A1(n16822), .A2(n18263), .ZN(n16787) );
  INV_X1 U19246 ( .A(n16787), .ZN(n16791) );
  NAND2_X1 U19247 ( .A1(n19037), .A2(n18586), .ZN(n18572) );
  INV_X1 U19248 ( .A(n18572), .ZN(n18590) );
  NOR2_X1 U19249 ( .A1(n17896), .A2(n16822), .ZN(n16771) );
  INV_X1 U19250 ( .A(n16771), .ZN(n16792) );
  AOI22_X1 U19251 ( .A1(n18425), .A2(n16791), .B1(n18590), .B2(n16792), .ZN(
        n16193) );
  OAI21_X1 U19252 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18576), .A(
        n16193), .ZN(n16124) );
  AOI21_X1 U19253 ( .B1(n18476), .B2(n16836), .A(n16124), .ZN(n16141) );
  INV_X1 U19254 ( .A(n18507), .ZN(n19043) );
  NOR3_X4 U19255 ( .A1(n17751), .A2(n19043), .A3(n18498), .ZN(n18480) );
  NOR2_X1 U19256 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18148) );
  NOR2_X2 U19257 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18120), .ZN(
        n18094) );
  INV_X1 U19258 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18098) );
  NAND2_X1 U19259 ( .A1(n18094), .A2(n18098), .ZN(n18085) );
  NOR2_X2 U19260 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18085), .ZN(
        n18066) );
  NAND3_X1 U19261 ( .A1(n18066), .A2(n21047), .A3(n18410), .ZN(n16125) );
  INV_X1 U19262 ( .A(n16126), .ZN(n18138) );
  NAND2_X1 U19263 ( .A1(n18095), .A2(n18366), .ZN(n16128) );
  NAND2_X2 U19264 ( .A1(n18041), .A2(n18168), .ZN(n17962) );
  NAND2_X1 U19265 ( .A1(n16129), .A2(n16128), .ZN(n18051) );
  INV_X1 U19266 ( .A(n18051), .ZN(n16133) );
  INV_X1 U19267 ( .A(n16130), .ZN(n16132) );
  NAND2_X1 U19268 ( .A1(n18036), .A2(n18364), .ZN(n16131) );
  NOR2_X1 U19269 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16131), .ZN(
        n18001) );
  INV_X1 U19270 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18341) );
  NAND2_X1 U19271 ( .A1(n18001), .A2(n18341), .ZN(n17979) );
  NAND2_X1 U19272 ( .A1(n18370), .A2(n18051), .ZN(n18000) );
  NAND2_X1 U19273 ( .A1(n16135), .A2(n18037), .ZN(n17963) );
  NOR2_X1 U19274 ( .A1(n18052), .A2(n16136), .ZN(n17941) );
  AOI21_X1 U19275 ( .B1(n18286), .B2(n17935), .A(n18052), .ZN(n16137) );
  INV_X1 U19276 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17898) );
  NOR2_X1 U19277 ( .A1(n16187), .A2(n16188), .ZN(n16139) );
  XNOR2_X1 U19278 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n16139), .ZN(
        n16817) );
  AOI22_X1 U19279 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18481), .B1(n18480), 
        .B2(n16817), .ZN(n16140) );
  OAI221_X1 U19280 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16190), 
        .C1(n9957), .C2(n16141), .A(n16140), .ZN(P3_U2833) );
  INV_X1 U19281 ( .A(n16142), .ZN(n16144) );
  NOR3_X1 U19282 ( .A1(n16144), .A2(n16143), .A3(n20693), .ZN(n16149) );
  INV_X1 U19283 ( .A(n16149), .ZN(n16147) );
  OAI211_X1 U19284 ( .C1(n16147), .C2(n20554), .A(n16146), .B(n16145), .ZN(
        n16148) );
  OAI21_X1 U19285 ( .B1(n16149), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16148), .ZN(n16150) );
  AOI222_X1 U19286 ( .A1(n16152), .A2(n16151), .B1(n16152), .B2(n16150), .C1(
        n16151), .C2(n16150), .ZN(n16153) );
  AOI222_X1 U19287 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16154), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16153), .C1(n16154), 
        .C2(n16153), .ZN(n16164) );
  NAND2_X1 U19288 ( .A1(n16156), .A2(n16155), .ZN(n16160) );
  OAI21_X1 U19289 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16157), .ZN(n16158) );
  NAND4_X1 U19290 ( .A1(n16161), .A2(n16160), .A3(n16159), .A4(n16158), .ZN(
        n16162) );
  AOI211_X1 U19291 ( .C1(n16164), .C2(n20516), .A(n16163), .B(n16162), .ZN(
        n16176) );
  INV_X1 U19292 ( .A(n16176), .ZN(n16169) );
  NAND2_X1 U19293 ( .A1(n20702), .A2(n20857), .ZN(n16168) );
  NAND3_X1 U19294 ( .A1(n16166), .A2(n12059), .A3(n16165), .ZN(n16167) );
  NAND2_X1 U19295 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20857), .ZN(n16502) );
  AOI21_X1 U19296 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .A(n20697), .ZN(n20759) );
  OAI211_X1 U19297 ( .C1(n16168), .C2(n16167), .A(n16502), .B(n20759), .ZN(
        n16508) );
  AOI221_X1 U19298 ( .B1(n16503), .B2(n16510), .C1(n16169), .C2(n16510), .A(
        n16508), .ZN(n16171) );
  NOR2_X1 U19299 ( .A1(n16171), .A2(n16503), .ZN(n16513) );
  NAND2_X1 U19300 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20861), .ZN(n16170) );
  OAI211_X1 U19301 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20857), .A(n16513), 
        .B(n16170), .ZN(n16509) );
  AOI21_X1 U19302 ( .B1(n16172), .B2(n20861), .A(n16171), .ZN(n16173) );
  OAI22_X1 U19303 ( .A1(n16174), .A2(n16509), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16173), .ZN(n16175) );
  OAI21_X1 U19304 ( .B1(n16176), .B2(n20293), .A(n16175), .ZN(P1_U3161) );
  AOI22_X1 U19305 ( .A1(n16179), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16178), .B2(n16177), .ZN(n16181) );
  XNOR2_X1 U19306 ( .A(n16181), .B(n16180), .ZN(n16330) );
  INV_X1 U19307 ( .A(n16330), .ZN(n16182) );
  OAI22_X1 U19308 ( .A1(n16182), .A2(n16457), .B1(n20503), .B2(n16246), .ZN(
        n16183) );
  AOI21_X1 U19309 ( .B1(n16390), .B2(n16180), .A(n16183), .ZN(n16184) );
  NAND2_X1 U19310 ( .A1(n16482), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16331) );
  OAI211_X1 U19311 ( .C1(n16391), .C2(n16180), .A(n16184), .B(n16331), .ZN(
        P1_U3010) );
  INV_X1 U19312 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16803) );
  OAI21_X1 U19313 ( .B1(n16185), .B2(n18498), .A(n18575), .ZN(n16186) );
  AOI21_X1 U19314 ( .B1(n18538), .B2(n16822), .A(n16186), .ZN(n16823) );
  NAND2_X1 U19315 ( .A1(n16189), .A2(n16803), .ZN(n16780) );
  OAI21_X1 U19316 ( .B1(n16189), .B2(n16803), .A(n16780), .ZN(n16801) );
  INV_X1 U19317 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19186) );
  NOR2_X1 U19318 ( .A1(n18476), .A2(n19186), .ZN(n16795) );
  NOR3_X1 U19319 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n9957), .A3(
        n16190), .ZN(n16191) );
  AOI211_X1 U19320 ( .C1(n18480), .C2(n16801), .A(n16795), .B(n16191), .ZN(
        n16192) );
  OAI221_X1 U19321 ( .B1(n16803), .B2(n16823), .C1(n16803), .C2(n16193), .A(
        n16192), .ZN(P3_U2832) );
  INV_X1 U19322 ( .A(HOLD), .ZN(n20769) );
  INV_X1 U19323 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20780) );
  NAND2_X1 U19324 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20764) );
  OAI21_X1 U19325 ( .B1(n20769), .B2(n20763), .A(n20764), .ZN(n16194) );
  OAI21_X1 U19326 ( .B1(n20769), .B2(n20780), .A(n16194), .ZN(n16196) );
  NOR2_X1 U19327 ( .A1(n20763), .A2(n20857), .ZN(n20772) );
  INV_X1 U19328 ( .A(n20772), .ZN(n20762) );
  NAND3_X1 U19329 ( .A1(n16196), .A2(n16195), .A3(n20762), .ZN(P1_U3195) );
  INV_X1 U19330 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16933) );
  NOR2_X1 U19331 ( .A1(n20395), .A2(n16933), .ZN(P1_U2905) );
  OAI21_X1 U19332 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16197), .ZN(n16202) );
  AOI22_X1 U19333 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16402), .B1(
        n16482), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n16201) );
  AOI22_X1 U19334 ( .A1(n16199), .A2(n20509), .B1(n20481), .B2(n16198), .ZN(
        n16200) );
  OAI211_X1 U19335 ( .C1(n16407), .C2(n16202), .A(n16201), .B(n16200), .ZN(
        P1_U3011) );
  NOR2_X1 U19336 ( .A1(n20274), .A2(n20278), .ZN(n20123) );
  INV_X1 U19337 ( .A(n16203), .ZN(n20245) );
  INV_X1 U19338 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20269) );
  OAI21_X1 U19339 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n20245), .A(n20269), 
        .ZN(n16204) );
  AOI21_X1 U19340 ( .B1(n20123), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n16204), 
        .ZN(n16205) );
  NOR2_X1 U19341 ( .A1(n16769), .A2(n16205), .ZN(P2_U3178) );
  AOI21_X1 U19342 ( .B1(n20269), .B2(n15859), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20275) );
  NAND2_X1 U19343 ( .A1(n20275), .A2(n20253), .ZN(n16206) );
  AOI221_X1 U19344 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16769), .C1(n16208), .C2(
        n16769), .A(n20067), .ZN(n20264) );
  INV_X1 U19345 ( .A(n20264), .ZN(n20261) );
  NOR2_X1 U19346 ( .A1(n16209), .A2(n20261), .ZN(P2_U3047) );
  NAND2_X1 U19347 ( .A1(n18639), .A2(n17631), .ZN(n17778) );
  INV_X1 U19348 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17858) );
  NAND2_X1 U19349 ( .A1(n16213), .A2(n17631), .ZN(n17774) );
  INV_X1 U19350 ( .A(n17774), .ZN(n17777) );
  AOI22_X1 U19351 ( .A1(n17777), .A2(BUF2_REG_0__SCAN_IN), .B1(n17776), .B2(
        n18253), .ZN(n16214) );
  OAI221_X1 U19352 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17778), .C1(n17858), 
        .C2(n17631), .A(n16214), .ZN(P3_U2735) );
  NAND2_X1 U19353 ( .A1(n20354), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n16217) );
  AOI22_X1 U19354 ( .A1(n16215), .A2(n20322), .B1(P1_REIP_REG_24__SCAN_IN), 
        .B2(n16229), .ZN(n16216) );
  OAI211_X1 U19355 ( .C1(n20316), .C2(n16218), .A(n16217), .B(n16216), .ZN(
        n16221) );
  NOR2_X1 U19356 ( .A1(n16219), .A2(n16255), .ZN(n16220) );
  AOI211_X1 U19357 ( .C1(n16223), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        n16224) );
  OAI21_X1 U19358 ( .B1(n20376), .B2(n16225), .A(n16224), .ZN(P1_U2816) );
  INV_X1 U19359 ( .A(n16326), .ZN(n16226) );
  AOI222_X1 U19360 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20374), .B1(
        n20354), .B2(P1_EBX_REG_23__SCAN_IN), .C1(n16226), .C2(n20322), .ZN(
        n16231) );
  OAI21_X1 U19361 ( .B1(n16239), .B2(n16227), .A(n20817), .ZN(n16228) );
  AOI22_X1 U19362 ( .A1(n16323), .A2(n20348), .B1(n16229), .B2(n16228), .ZN(
        n16230) );
  OAI211_X1 U19363 ( .C1(n20376), .C2(n16232), .A(n16231), .B(n16230), .ZN(
        P1_U2817) );
  NOR2_X1 U19364 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n16239), .ZN(n16233) );
  AOI22_X1 U19365 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20374), .B1(
        n16234), .B2(n16233), .ZN(n16243) );
  AOI22_X1 U19366 ( .A1(n20322), .A2(n16235), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n20354), .ZN(n16242) );
  OAI22_X1 U19367 ( .A1(n21071), .A2(n16255), .B1(n20376), .B2(n16395), .ZN(
        n16236) );
  INV_X1 U19368 ( .A(n16236), .ZN(n16241) );
  INV_X1 U19369 ( .A(n16237), .ZN(n16244) );
  OAI21_X1 U19370 ( .B1(n16244), .B2(n16239), .A(n16238), .ZN(n16258) );
  NOR2_X1 U19371 ( .A1(n16239), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16245) );
  OAI21_X1 U19372 ( .B1(n16258), .B2(n16245), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n16240) );
  NAND4_X1 U19373 ( .A1(n16243), .A2(n16242), .A3(n16241), .A4(n16240), .ZN(
        P1_U2818) );
  INV_X1 U19374 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16334) );
  AOI22_X1 U19375 ( .A1(n16245), .A2(n16244), .B1(n20354), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n16251) );
  NOR2_X1 U19376 ( .A1(n16327), .A2(n20384), .ZN(n16249) );
  INV_X1 U19377 ( .A(n16329), .ZN(n16247) );
  OAI22_X1 U19378 ( .A1(n16247), .A2(n16255), .B1(n20376), .B2(n16246), .ZN(
        n16248) );
  AOI211_X1 U19379 ( .C1(n16258), .C2(P1_REIP_REG_21__SCAN_IN), .A(n16249), 
        .B(n16248), .ZN(n16250) );
  OAI211_X1 U19380 ( .C1(n16334), .C2(n20316), .A(n16251), .B(n16250), .ZN(
        P1_U2819) );
  AOI22_X1 U19381 ( .A1(n20322), .A2(n16252), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n20354), .ZN(n16260) );
  INV_X1 U19382 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20811) );
  INV_X1 U19383 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20808) );
  NAND2_X1 U19384 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n16283), .ZN(n16262) );
  NOR2_X1 U19385 ( .A1(n20811), .A2(n16262), .ZN(n16276) );
  OAI22_X1 U19386 ( .A1(n16256), .A2(n16255), .B1(n20376), .B2(n16254), .ZN(
        n16257) );
  AOI221_X1 U19387 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n16258), .C1(n16276), 
        .C2(n16258), .A(n16257), .ZN(n16259) );
  OAI211_X1 U19388 ( .C1(n16261), .C2(n20316), .A(n16260), .B(n16259), .ZN(
        P1_U2820) );
  INV_X1 U19389 ( .A(n16262), .ZN(n16263) );
  AOI21_X1 U19390 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n16303), .A(n16263), 
        .ZN(n16275) );
  INV_X1 U19391 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16265) );
  NAND2_X1 U19392 ( .A1(n20354), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n16264) );
  OAI211_X1 U19393 ( .C1(n20316), .C2(n16265), .A(n16264), .B(n16489), .ZN(
        n16266) );
  AOI21_X1 U19394 ( .B1(n20322), .B2(n16267), .A(n16266), .ZN(n16274) );
  OR2_X1 U19395 ( .A1(n16269), .A2(n16268), .ZN(n16270) );
  AND2_X1 U19396 ( .A1(n14642), .A2(n16270), .ZN(n16337) );
  XNOR2_X1 U19397 ( .A(n16272), .B(n16271), .ZN(n16403) );
  AOI22_X1 U19398 ( .A1(n16337), .A2(n20348), .B1(n20356), .B2(n16403), .ZN(
        n16273) );
  OAI211_X1 U19399 ( .C1(n16276), .C2(n16275), .A(n16274), .B(n16273), .ZN(
        P1_U2821) );
  INV_X1 U19400 ( .A(n16283), .ZN(n16287) );
  INV_X1 U19401 ( .A(n16277), .ZN(n16278) );
  AOI22_X1 U19402 ( .A1(n20322), .A2(n16278), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n20354), .ZN(n16279) );
  OAI211_X1 U19403 ( .C1(n20316), .C2(n16280), .A(n16279), .B(n16489), .ZN(
        n16281) );
  AOI21_X1 U19404 ( .B1(n20356), .B2(n16282), .A(n16281), .ZN(n16286) );
  AOI22_X1 U19405 ( .A1(n16284), .A2(n20348), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n10239), .ZN(n16285) );
  OAI211_X1 U19406 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n16287), .A(n16286), 
        .B(n16285), .ZN(P1_U2822) );
  OAI22_X1 U19407 ( .A1(n20316), .A2(n16289), .B1(n20372), .B2(n16288), .ZN(
        n16290) );
  AOI211_X1 U19408 ( .C1(n20322), .C2(n16348), .A(n16482), .B(n16290), .ZN(
        n16294) );
  NAND2_X1 U19409 ( .A1(n20808), .A2(n16291), .ZN(n16292) );
  AOI22_X1 U19410 ( .A1(n16349), .A2(n20348), .B1(n10239), .B2(n16292), .ZN(
        n16293) );
  OAI211_X1 U19411 ( .C1(n20376), .C2(n16408), .A(n16294), .B(n16293), .ZN(
        P1_U2823) );
  AOI22_X1 U19412 ( .A1(n20354), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20374), .ZN(n16302) );
  AOI21_X1 U19413 ( .B1(n16297), .B2(n16296), .A(n16295), .ZN(n16451) );
  AOI21_X1 U19414 ( .B1(n16451), .B2(n20356), .A(n16482), .ZN(n16301) );
  AOI22_X1 U19415 ( .A1(n16364), .A2(n20322), .B1(n20348), .B2(n16363), .ZN(
        n16300) );
  OAI211_X1 U19416 ( .C1(P1_REIP_REG_12__SCAN_IN), .C2(n16312), .A(n16303), 
        .B(n16298), .ZN(n16299) );
  NAND4_X1 U19417 ( .A1(n16302), .A2(n16301), .A3(n16300), .A4(n16299), .ZN(
        P1_U2828) );
  AOI22_X1 U19418 ( .A1(n16304), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n16303), .ZN(n16311) );
  OAI22_X1 U19419 ( .A1(n16306), .A2(n20376), .B1(n16305), .B2(n20372), .ZN(
        n16307) );
  AOI211_X1 U19420 ( .C1(n20374), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16482), .B(n16307), .ZN(n16310) );
  INV_X1 U19421 ( .A(n16372), .ZN(n16308) );
  AOI22_X1 U19422 ( .A1(n16308), .A2(n20322), .B1(n20348), .B2(n16368), .ZN(
        n16309) );
  OAI211_X1 U19423 ( .C1(n16312), .C2(n16311), .A(n16310), .B(n16309), .ZN(
        P1_U2829) );
  AOI22_X1 U19424 ( .A1(n16337), .A2(n20387), .B1(n16315), .B2(n16403), .ZN(
        n16313) );
  OAI21_X1 U19425 ( .B1(n20390), .B2(n16314), .A(n16313), .ZN(P1_U2853) );
  AOI22_X1 U19426 ( .A1(n16363), .A2(n20387), .B1(n16315), .B2(n16451), .ZN(
        n16316) );
  OAI21_X1 U19427 ( .B1(n20390), .B2(n16317), .A(n16316), .ZN(P1_U2860) );
  INV_X1 U19428 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U19429 ( .A1(n21065), .A2(n16318), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n21063), .ZN(n16321) );
  AOI22_X1 U19430 ( .A1(n16337), .A2(n16319), .B1(n21062), .B2(DATAI_19_), 
        .ZN(n16320) );
  OAI211_X1 U19431 ( .C1(n21068), .C2(n16863), .A(n16321), .B(n16320), .ZN(
        P1_U2885) );
  AOI22_X1 U19432 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16325) );
  AOI22_X1 U19433 ( .A1(n16323), .A2(n20456), .B1(n20457), .B2(n16322), .ZN(
        n16324) );
  OAI211_X1 U19434 ( .C1(n20461), .C2(n16326), .A(n16325), .B(n16324), .ZN(
        P1_U2976) );
  INV_X1 U19435 ( .A(n16327), .ZN(n16328) );
  AOI222_X1 U19436 ( .A1(n20457), .A2(n16330), .B1(n16329), .B2(n20456), .C1(
        n16328), .C2(n16365), .ZN(n16332) );
  OAI211_X1 U19437 ( .C1(n16334), .C2(n16333), .A(n16332), .B(n16331), .ZN(
        P1_U2978) );
  AOI22_X1 U19438 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16339) );
  MUX2_X1 U19439 ( .A(n10206), .B(n16335), .S(n14823), .Z(n16336) );
  XNOR2_X1 U19440 ( .A(n16336), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16404) );
  AOI22_X1 U19441 ( .A1(n16404), .A2(n20457), .B1(n20456), .B2(n16337), .ZN(
        n16338) );
  OAI211_X1 U19442 ( .C1(n20461), .C2(n16340), .A(n16339), .B(n16338), .ZN(
        P1_U2980) );
  INV_X1 U19443 ( .A(n16341), .ZN(n16343) );
  OAI21_X1 U19444 ( .B1(n16344), .B2(n16343), .A(n16342), .ZN(n16346) );
  NAND2_X1 U19445 ( .A1(n16346), .A2(n14381), .ZN(n16345) );
  MUX2_X1 U19446 ( .A(n16346), .B(n16345), .S(n10206), .Z(n16347) );
  XNOR2_X1 U19447 ( .A(n16347), .B(n16413), .ZN(n16409) );
  AOI22_X1 U19448 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16351) );
  AOI22_X1 U19449 ( .A1(n16349), .A2(n20456), .B1(n16348), .B2(n16365), .ZN(
        n16350) );
  OAI211_X1 U19450 ( .C1(n20299), .C2(n16409), .A(n16351), .B(n16350), .ZN(
        P1_U2982) );
  OAI21_X1 U19451 ( .B1(n16354), .B2(n16353), .A(n16352), .ZN(n16355) );
  INV_X1 U19452 ( .A(n16355), .ZN(n16429) );
  AOI22_X1 U19453 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16359) );
  AOI22_X1 U19454 ( .A1(n16357), .A2(n20456), .B1(n16365), .B2(n16356), .ZN(
        n16358) );
  OAI211_X1 U19455 ( .C1(n16429), .C2(n20299), .A(n16359), .B(n16358), .ZN(
        P1_U2984) );
  AOI21_X1 U19456 ( .B1(n16362), .B2(n16361), .A(n16360), .ZN(n16458) );
  AOI22_X1 U19457 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19458 ( .A1(n16365), .A2(n16364), .B1(n20456), .B2(n16363), .ZN(
        n16366) );
  OAI211_X1 U19459 ( .C1(n16458), .C2(n20299), .A(n16367), .B(n16366), .ZN(
        P1_U2987) );
  AOI22_X1 U19460 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U19461 ( .A1(n20457), .A2(n16369), .B1(n20456), .B2(n16368), .ZN(
        n16370) );
  OAI211_X1 U19462 ( .C1(n20461), .C2(n16372), .A(n16371), .B(n16370), .ZN(
        P1_U2988) );
  AOI22_X1 U19463 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16378) );
  NAND2_X1 U19464 ( .A1(n16374), .A2(n16373), .ZN(n16375) );
  XNOR2_X1 U19465 ( .A(n16376), .B(n16375), .ZN(n16484) );
  AOI22_X1 U19466 ( .A1(n16484), .A2(n20457), .B1(n20456), .B2(n20338), .ZN(
        n16377) );
  OAI211_X1 U19467 ( .C1(n20461), .C2(n20334), .A(n16378), .B(n16377), .ZN(
        P1_U2992) );
  AOI22_X1 U19468 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16383) );
  XNOR2_X1 U19469 ( .A(n16379), .B(n20999), .ZN(n16380) );
  XNOR2_X1 U19470 ( .A(n16381), .B(n16380), .ZN(n16492) );
  AOI22_X1 U19471 ( .A1(n16492), .A2(n20457), .B1(n20456), .B2(n20347), .ZN(
        n16382) );
  OAI211_X1 U19472 ( .C1(n20461), .C2(n20353), .A(n16383), .B(n16382), .ZN(
        P1_U2993) );
  AOI22_X1 U19473 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16389) );
  OAI21_X1 U19474 ( .B1(n16386), .B2(n16385), .A(n16384), .ZN(n16387) );
  INV_X1 U19475 ( .A(n16387), .ZN(n16498) );
  AOI22_X1 U19476 ( .A1(n16498), .A2(n20457), .B1(n20456), .B2(n20360), .ZN(
        n16388) );
  OAI211_X1 U19477 ( .C1(n20461), .C2(n20358), .A(n16389), .B(n16388), .ZN(
        P1_U2994) );
  OAI21_X1 U19478 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16390), .ZN(n16400) );
  INV_X1 U19479 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16392) );
  OAI22_X1 U19480 ( .A1(n16392), .A2(n16391), .B1(n16489), .B2(n14819), .ZN(
        n16393) );
  INV_X1 U19481 ( .A(n16393), .ZN(n16399) );
  INV_X1 U19482 ( .A(n16394), .ZN(n16397) );
  INV_X1 U19483 ( .A(n16395), .ZN(n16396) );
  AOI22_X1 U19484 ( .A1(n16397), .A2(n20509), .B1(n20481), .B2(n16396), .ZN(
        n16398) );
  OAI211_X1 U19485 ( .C1(n16401), .C2(n16400), .A(n16399), .B(n16398), .ZN(
        P1_U3009) );
  AOI22_X1 U19486 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16402), .B1(
        n16482), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16406) );
  AOI22_X1 U19487 ( .A1(n16404), .A2(n20509), .B1(n20481), .B2(n16403), .ZN(
        n16405) );
  OAI211_X1 U19488 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16407), .A(
        n16406), .B(n16405), .ZN(P1_U3012) );
  OAI22_X1 U19489 ( .A1(n16409), .A2(n16457), .B1(n20503), .B2(n16408), .ZN(
        n16410) );
  AOI21_X1 U19490 ( .B1(n16482), .B2(P1_REIP_REG_17__SCAN_IN), .A(n16410), 
        .ZN(n16411) );
  OAI221_X1 U19491 ( .B1(n16414), .B2(n16413), .C1(n16414), .C2(n16412), .A(
        n16411), .ZN(P1_U3014) );
  INV_X1 U19492 ( .A(n16415), .ZN(n16418) );
  INV_X1 U19493 ( .A(n16416), .ZN(n16417) );
  AOI22_X1 U19494 ( .A1(n16418), .A2(n20509), .B1(n20481), .B2(n16417), .ZN(
        n16423) );
  NAND2_X1 U19495 ( .A1(n16482), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16422) );
  NAND2_X1 U19496 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16426), .ZN(
        n16421) );
  NAND2_X1 U19497 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16419) );
  OAI211_X1 U19498 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16427), .B(n16419), .ZN(
        n16420) );
  NAND4_X1 U19499 ( .A1(n16423), .A2(n16422), .A3(n16421), .A4(n16420), .ZN(
        P1_U3015) );
  OAI22_X1 U19500 ( .A1(n16424), .A2(n20503), .B1(n20803), .B2(n16489), .ZN(
        n16425) );
  AOI221_X1 U19501 ( .B1(n16427), .B2(n14431), .C1(n16426), .C2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16425), .ZN(n16428) );
  OAI21_X1 U19502 ( .B1(n16429), .B2(n16457), .A(n16428), .ZN(P1_U3016) );
  INV_X1 U19503 ( .A(n16430), .ZN(n16432) );
  AOI21_X1 U19504 ( .B1(n16432), .B2(n20481), .A(n16431), .ZN(n16437) );
  NOR2_X1 U19505 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16433), .ZN(
        n16434) );
  AOI22_X1 U19506 ( .A1(n20509), .A2(n16435), .B1(n16491), .B2(n16434), .ZN(
        n16436) );
  OAI211_X1 U19507 ( .C1(n16439), .C2(n16438), .A(n16437), .B(n16436), .ZN(
        P1_U3017) );
  OAI22_X1 U19508 ( .A1(n16441), .A2(n20498), .B1(n16473), .B2(n16440), .ZN(
        n16442) );
  NOR2_X1 U19509 ( .A1(n16443), .A2(n16442), .ZN(n16447) );
  AOI222_X1 U19510 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16482), .B1(n20481), 
        .B2(n16445), .C1(n20509), .C2(n16444), .ZN(n16446) );
  OAI221_X1 U19511 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16449), 
        .C1(n16448), .C2(n16447), .A(n16446), .ZN(P1_U3018) );
  OAI21_X1 U19512 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n20493), .A(
        n16450), .ZN(n16452) );
  AOI222_X1 U19513 ( .A1(n16452), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .B1(n20481), .B2(n16451), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n16482), 
        .ZN(n16456) );
  NAND3_X1 U19514 ( .A1(n16454), .A2(n16491), .A3(n16453), .ZN(n16455) );
  OAI211_X1 U19515 ( .C1(n16458), .C2(n16457), .A(n16456), .B(n16455), .ZN(
        P1_U3019) );
  OAI21_X1 U19516 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16459), .ZN(n16466) );
  AOI21_X1 U19517 ( .B1(n16461), .B2(n20481), .A(n16460), .ZN(n16465) );
  AOI22_X1 U19518 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16463), .B1(
        n20509), .B2(n16462), .ZN(n16464) );
  OAI211_X1 U19519 ( .C1(n16467), .C2(n16466), .A(n16465), .B(n16464), .ZN(
        P1_U3021) );
  NAND2_X1 U19520 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16491), .ZN(
        n16487) );
  AOI22_X1 U19521 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16469), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16468), .ZN(n16480) );
  AOI21_X1 U19522 ( .B1(n16471), .B2(n20481), .A(n16470), .ZN(n16479) );
  NOR2_X1 U19523 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20462), .ZN(
        n16496) );
  NOR2_X1 U19524 ( .A1(n20462), .A2(n20465), .ZN(n16474) );
  OAI21_X1 U19525 ( .B1(n16474), .B2(n16473), .A(n16472), .ZN(n16497) );
  AOI21_X1 U19526 ( .B1(n16475), .B2(n16496), .A(n16497), .ZN(n16495) );
  OAI21_X1 U19527 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16476), .A(
        n16495), .ZN(n16483) );
  AOI22_X1 U19528 ( .A1(n16477), .A2(n20509), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16483), .ZN(n16478) );
  OAI211_X1 U19529 ( .C1(n16487), .C2(n16480), .A(n16479), .B(n16478), .ZN(
        P1_U3023) );
  INV_X1 U19530 ( .A(n16481), .ZN(n20332) );
  AOI22_X1 U19531 ( .A1(n20332), .A2(n20481), .B1(n16482), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U19532 ( .A1(n16484), .A2(n20509), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16483), .ZN(n16485) );
  OAI211_X1 U19533 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16487), .A(
        n16486), .B(n16485), .ZN(P1_U3024) );
  INV_X1 U19534 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n16488) );
  OAI22_X1 U19535 ( .A1(n20342), .A2(n20503), .B1(n16489), .B2(n16488), .ZN(
        n16490) );
  INV_X1 U19536 ( .A(n16490), .ZN(n16494) );
  AOI22_X1 U19537 ( .A1(n16492), .A2(n20509), .B1(n20999), .B2(n16491), .ZN(
        n16493) );
  OAI211_X1 U19538 ( .C1(n16495), .C2(n20999), .A(n16494), .B(n16493), .ZN(
        P1_U3025) );
  INV_X1 U19539 ( .A(n16496), .ZN(n16501) );
  AOI22_X1 U19540 ( .A1(n20355), .A2(n20481), .B1(n16482), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16500) );
  AOI22_X1 U19541 ( .A1(n16498), .A2(n20509), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16497), .ZN(n16499) );
  OAI211_X1 U19542 ( .C1(n20478), .C2(n16501), .A(n16500), .B(n16499), .ZN(
        P1_U3026) );
  NOR3_X1 U19543 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n16503), .A3(n16502), 
        .ZN(n16505) );
  NOR2_X1 U19544 ( .A1(n16505), .A2(n16504), .ZN(n20760) );
  NAND2_X1 U19545 ( .A1(n20760), .A2(n16506), .ZN(n16507) );
  AOI22_X1 U19546 ( .A1(n16510), .A2(n16509), .B1(n16508), .B2(n16507), .ZN(
        P1_U3162) );
  OAI21_X1 U19547 ( .B1(n16513), .B2(n16512), .A(n16511), .ZN(P1_U3466) );
  INV_X1 U19548 ( .A(n16515), .ZN(n16594) );
  NAND2_X1 U19549 ( .A1(n9661), .A2(n16592), .ZN(n16581) );
  NAND2_X1 U19550 ( .A1(n16582), .A2(n16581), .ZN(n16580) );
  INV_X1 U19551 ( .A(n16516), .ZN(n16571) );
  NAND2_X1 U19552 ( .A1(n13308), .A2(n16569), .ZN(n16556) );
  NAND2_X1 U19553 ( .A1(n16557), .A2(n16556), .ZN(n16555) );
  INV_X1 U19554 ( .A(n16517), .ZN(n16546) );
  NAND2_X1 U19555 ( .A1(n9661), .A2(n16544), .ZN(n16534) );
  NAND2_X1 U19556 ( .A1(n16535), .A2(n16534), .ZN(n16533) );
  INV_X1 U19557 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16522) );
  INV_X1 U19558 ( .A(n16518), .ZN(n16519) );
  AOI22_X1 U19559 ( .A1(n16519), .A2(n19294), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n19392), .ZN(n16520) );
  OAI21_X1 U19560 ( .B1(n16522), .B2(n16521), .A(n16520), .ZN(n16523) );
  AOI21_X1 U19561 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19417), .A(
        n16523), .ZN(n16527) );
  INV_X1 U19562 ( .A(n16524), .ZN(n19421) );
  AOI22_X1 U19563 ( .A1(n16525), .A2(n19396), .B1(n19377), .B2(n19421), .ZN(
        n16526) );
  OAI211_X1 U19564 ( .C1(n16528), .C2(n16533), .A(n16527), .B(n16526), .ZN(
        P2_U2824) );
  AOI22_X1 U19565 ( .A1(n16529), .A2(n19294), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19417), .ZN(n16539) );
  AOI22_X1 U19566 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19411), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19392), .ZN(n16538) );
  INV_X1 U19567 ( .A(n16530), .ZN(n16531) );
  AOI22_X1 U19568 ( .A1(n16532), .A2(n19396), .B1(n19377), .B2(n16531), .ZN(
        n16537) );
  OAI211_X1 U19569 ( .C1(n16535), .C2(n16534), .A(n9671), .B(n16533), .ZN(
        n16536) );
  NAND4_X1 U19570 ( .A1(n16539), .A2(n16538), .A3(n16537), .A4(n16536), .ZN(
        P2_U2825) );
  AOI22_X1 U19571 ( .A1(n16540), .A2(n19294), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19417), .ZN(n16550) );
  AOI22_X1 U19572 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19411), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19392), .ZN(n16549) );
  OAI22_X1 U19573 ( .A1(n16542), .A2(n19413), .B1(n16541), .B2(n19408), .ZN(
        n16543) );
  INV_X1 U19574 ( .A(n16543), .ZN(n16548) );
  OAI211_X1 U19575 ( .C1(n16546), .C2(n16545), .A(n9671), .B(n16544), .ZN(
        n16547) );
  NAND4_X1 U19576 ( .A1(n16550), .A2(n16549), .A3(n16548), .A4(n16547), .ZN(
        P2_U2826) );
  AOI22_X1 U19577 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19417), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19392), .ZN(n16561) );
  AOI22_X1 U19578 ( .A1(n16551), .A2(n19294), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n19411), .ZN(n16560) );
  OAI22_X1 U19579 ( .A1(n16553), .A2(n19413), .B1(n16552), .B2(n19408), .ZN(
        n16554) );
  INV_X1 U19580 ( .A(n16554), .ZN(n16559) );
  OAI211_X1 U19581 ( .C1(n16557), .C2(n16556), .A(n9671), .B(n16555), .ZN(
        n16558) );
  NAND4_X1 U19582 ( .A1(n16561), .A2(n16560), .A3(n16559), .A4(n16558), .ZN(
        P2_U2827) );
  AOI22_X1 U19583 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19417), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19392), .ZN(n16575) );
  OAI22_X1 U19584 ( .A1(n16563), .A2(n19404), .B1(n19352), .B2(n16562), .ZN(
        n16564) );
  INV_X1 U19585 ( .A(n16564), .ZN(n16574) );
  INV_X1 U19586 ( .A(n16565), .ZN(n16566) );
  OAI22_X1 U19587 ( .A1(n16567), .A2(n19413), .B1(n16566), .B2(n19408), .ZN(
        n16568) );
  INV_X1 U19588 ( .A(n16568), .ZN(n16573) );
  OAI211_X1 U19589 ( .C1(n16571), .C2(n16570), .A(n9671), .B(n16569), .ZN(
        n16572) );
  NAND4_X1 U19590 ( .A1(n16575), .A2(n16574), .A3(n16573), .A4(n16572), .ZN(
        P2_U2828) );
  AOI22_X1 U19591 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19417), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19392), .ZN(n16586) );
  AOI22_X1 U19592 ( .A1(n16576), .A2(n19294), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19411), .ZN(n16585) );
  INV_X1 U19593 ( .A(n16577), .ZN(n16579) );
  AOI22_X1 U19594 ( .A1(n16579), .A2(n19396), .B1(n16578), .B2(n19377), .ZN(
        n16584) );
  OAI211_X1 U19595 ( .C1(n16582), .C2(n16581), .A(n9671), .B(n16580), .ZN(
        n16583) );
  NAND4_X1 U19596 ( .A1(n16586), .A2(n16585), .A3(n16584), .A4(n16583), .ZN(
        P2_U2829) );
  AOI22_X1 U19597 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19417), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19392), .ZN(n16598) );
  AOI22_X1 U19598 ( .A1(n16587), .A2(n19294), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n19411), .ZN(n16597) );
  INV_X1 U19599 ( .A(n16588), .ZN(n16589) );
  OAI22_X1 U19600 ( .A1(n16590), .A2(n19413), .B1(n16589), .B2(n19408), .ZN(
        n16591) );
  INV_X1 U19601 ( .A(n16591), .ZN(n16596) );
  OAI211_X1 U19602 ( .C1(n16594), .C2(n16593), .A(n9671), .B(n16592), .ZN(
        n16595) );
  NAND4_X1 U19603 ( .A1(n16598), .A2(n16597), .A3(n16596), .A4(n16595), .ZN(
        P2_U2830) );
  AOI22_X1 U19604 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19417), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19392), .ZN(n16610) );
  INV_X1 U19605 ( .A(n16599), .ZN(n16600) );
  AOI22_X1 U19606 ( .A1(n16600), .A2(n19294), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19411), .ZN(n16609) );
  OAI22_X1 U19607 ( .A1(n16602), .A2(n19413), .B1(n16601), .B2(n19408), .ZN(
        n16603) );
  INV_X1 U19608 ( .A(n16603), .ZN(n16608) );
  OAI211_X1 U19609 ( .C1(n16606), .C2(n16605), .A(n9671), .B(n16604), .ZN(
        n16607) );
  NAND4_X1 U19610 ( .A1(n16610), .A2(n16609), .A3(n16608), .A4(n16607), .ZN(
        P2_U2831) );
  AOI22_X1 U19611 ( .A1(n16618), .A2(n16611), .B1(n19485), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16616) );
  AOI22_X1 U19612 ( .A1(n19420), .A2(BUF1_REG_23__SCAN_IN), .B1(n19422), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16615) );
  AOI22_X1 U19613 ( .A1(n16613), .A2(n19487), .B1(n19486), .B2(n16612), .ZN(
        n16614) );
  NAND3_X1 U19614 ( .A1(n16616), .A2(n16615), .A3(n16614), .ZN(P2_U2896) );
  AOI22_X1 U19615 ( .A1(n16618), .A2(n16617), .B1(n19485), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16623) );
  AOI22_X1 U19616 ( .A1(n19420), .A2(BUF1_REG_22__SCAN_IN), .B1(n19422), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16622) );
  AOI22_X1 U19617 ( .A1(n16620), .A2(n19487), .B1(n19486), .B2(n16619), .ZN(
        n16621) );
  NAND3_X1 U19618 ( .A1(n16623), .A2(n16622), .A3(n16621), .ZN(P2_U2897) );
  AOI22_X1 U19619 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19529), .B1(n16658), 
        .B2(n16624), .ZN(n16634) );
  NAND2_X1 U19620 ( .A1(n16626), .A2(n16625), .ZN(n16630) );
  NOR2_X1 U19621 ( .A1(n16628), .A2(n16627), .ZN(n16629) );
  XOR2_X1 U19622 ( .A(n16630), .B(n16629), .Z(n16674) );
  AOI21_X1 U19623 ( .B1(n16638), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16632) );
  NOR2_X1 U19624 ( .A1(n16632), .A2(n16631), .ZN(n16671) );
  AOI222_X1 U19625 ( .A1(n16674), .A2(n16662), .B1(n19538), .B2(n16672), .C1(
        n16660), .C2(n16671), .ZN(n16633) );
  OAI211_X1 U19626 ( .C1(n16635), .C2(n16666), .A(n16634), .B(n16633), .ZN(
        P2_U3003) );
  AOI22_X1 U19627 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19529), .B1(n16658), 
        .B2(n16636), .ZN(n16644) );
  NOR3_X1 U19628 ( .A1(n16638), .A2(n16637), .A3(n19532), .ZN(n16642) );
  OAI22_X1 U19629 ( .A1(n16640), .A2(n19534), .B1(n16648), .B2(n16639), .ZN(
        n16641) );
  NOR2_X1 U19630 ( .A1(n16642), .A2(n16641), .ZN(n16643) );
  OAI211_X1 U19631 ( .C1(n16645), .C2(n16666), .A(n16644), .B(n16643), .ZN(
        P2_U3005) );
  AOI22_X1 U19632 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19529), .B1(n16658), 
        .B2(n16646), .ZN(n16655) );
  NAND3_X1 U19633 ( .A1(n16647), .A2(n16660), .A3(n15841), .ZN(n16653) );
  NOR2_X1 U19634 ( .A1(n16649), .A2(n16648), .ZN(n16650) );
  AOI21_X1 U19635 ( .B1(n16651), .B2(n16662), .A(n16650), .ZN(n16652) );
  AND2_X1 U19636 ( .A1(n16653), .A2(n16652), .ZN(n16654) );
  OAI211_X1 U19637 ( .C1(n16656), .C2(n16666), .A(n16655), .B(n16654), .ZN(
        P2_U3007) );
  AOI22_X1 U19638 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19529), .B1(n16658), 
        .B2(n16657), .ZN(n16665) );
  AOI222_X1 U19639 ( .A1(n16663), .A2(n16662), .B1(n16661), .B2(n16660), .C1(
        n19538), .C2(n16659), .ZN(n16664) );
  OAI211_X1 U19640 ( .C1(n16667), .C2(n16666), .A(n16665), .B(n16664), .ZN(
        P2_U3009) );
  INV_X1 U19641 ( .A(n16668), .ZN(n16670) );
  AOI22_X1 U19642 ( .A1(n16670), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16669), .B2(n19439), .ZN(n16680) );
  AOI222_X1 U19643 ( .A1(n16674), .A2(n16673), .B1(n16689), .B2(n16672), .C1(
        n16690), .C2(n16671), .ZN(n16679) );
  NAND2_X1 U19644 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19529), .ZN(n16678) );
  OAI221_X1 U19645 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n16676), .C2(n10921), .A(
        n16675), .ZN(n16677) );
  NAND4_X1 U19646 ( .A1(n16680), .A2(n16679), .A3(n16678), .A4(n16677), .ZN(
        P2_U3035) );
  AOI221_X1 U19647 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n16682), .C2(n16685), .A(
        n16681), .ZN(n16688) );
  OAI21_X1 U19648 ( .B1(n13304), .B2(n16684), .A(n16683), .ZN(n19451) );
  OAI22_X1 U19649 ( .A1(n16701), .A2(n19451), .B1(n16686), .B2(n16685), .ZN(
        n16687) );
  AOI211_X1 U19650 ( .C1(n19529), .C2(P2_REIP_REG_8__SCAN_IN), .A(n16688), .B(
        n16687), .ZN(n16693) );
  AOI22_X1 U19651 ( .A1(n16691), .A2(n16690), .B1(n16689), .B2(n19359), .ZN(
        n16692) );
  OAI211_X1 U19652 ( .C1(n16694), .C2(n16697), .A(n16693), .B(n16692), .ZN(
        P2_U3038) );
  OAI22_X1 U19653 ( .A1(n16697), .A2(n16696), .B1(n16695), .B2(n16706), .ZN(
        n16704) );
  INV_X1 U19654 ( .A(n16698), .ZN(n16700) );
  XNOR2_X1 U19655 ( .A(n16700), .B(n16699), .ZN(n19489) );
  INV_X1 U19656 ( .A(n19489), .ZN(n19407) );
  OAI22_X1 U19657 ( .A1(n19414), .A2(n16702), .B1(n16701), .B2(n19407), .ZN(
        n16703) );
  AOI211_X1 U19658 ( .C1(n16706), .C2(n16705), .A(n16704), .B(n16703), .ZN(
        n16708) );
  OAI211_X1 U19659 ( .C1(n16710), .C2(n16709), .A(n16708), .B(n16707), .ZN(
        P2_U3046) );
  NAND2_X1 U19660 ( .A1(n16725), .A2(n16728), .ZN(n16715) );
  INV_X1 U19661 ( .A(n16711), .ZN(n16712) );
  NAND2_X1 U19662 ( .A1(n16713), .A2(n16712), .ZN(n16714) );
  OAI211_X1 U19663 ( .C1(n16753), .C2(n16716), .A(n16715), .B(n16714), .ZN(
        n16717) );
  AOI21_X1 U19664 ( .B1(n16721), .B2(n16718), .A(n16717), .ZN(n16719) );
  OAI21_X1 U19665 ( .B1(n16721), .B2(n16720), .A(n16719), .ZN(n20267) );
  NAND2_X1 U19666 ( .A1(n9659), .A2(n16722), .ZN(n16724) );
  NOR2_X1 U19667 ( .A1(n11066), .A2(n16724), .ZN(n20218) );
  INV_X1 U19668 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n21041) );
  INV_X1 U19669 ( .A(n16725), .ZN(n16730) );
  INV_X1 U19670 ( .A(n16726), .ZN(n16727) );
  NAND4_X1 U19671 ( .A1(n16730), .A2(n16729), .A3(n16728), .A4(n16727), .ZN(
        n19274) );
  AOI21_X1 U19672 ( .B1(n19276), .B2(n21041), .A(n19274), .ZN(n16732) );
  NOR4_X1 U19673 ( .A1(n20267), .A2(n20218), .A3(n16732), .A4(n16731), .ZN(
        n16751) );
  INV_X1 U19674 ( .A(n16734), .ZN(n16736) );
  OAI211_X1 U19675 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16734), .A(
        n16733), .B(n19829), .ZN(n16735) );
  OAI211_X1 U19676 ( .C1(n19920), .C2(n16736), .A(n16735), .B(n16752), .ZN(
        n16743) );
  INV_X1 U19677 ( .A(n16743), .ZN(n16739) );
  MUX2_X1 U19678 ( .A(n10572), .B(n16737), .S(n16752), .Z(n16746) );
  OAI21_X1 U19679 ( .B1(n16743), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16746), .ZN(n16738) );
  NOR2_X1 U19680 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16744) );
  OAI211_X1 U19681 ( .C1(n16739), .C2(n20243), .A(n16738), .B(n16744), .ZN(
        n16742) );
  MUX2_X1 U19682 ( .A(n9802), .B(n16740), .S(n16752), .Z(n16741) );
  NAND2_X1 U19683 ( .A1(n16742), .A2(n16741), .ZN(n16749) );
  OR2_X1 U19684 ( .A1(n16743), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16747) );
  INV_X1 U19685 ( .A(n16744), .ZN(n16745) );
  OAI211_X1 U19686 ( .C1(n16747), .C2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16746), .B(n16745), .ZN(n16748) );
  NAND2_X1 U19687 ( .A1(n16749), .A2(n16748), .ZN(n16750) );
  OAI211_X1 U19688 ( .C1(n20221), .C2(n16752), .A(n16751), .B(n16750), .ZN(
        n16754) );
  AOI22_X1 U19689 ( .A1(n20122), .A2(n16754), .B1(n16753), .B2(n16769), .ZN(
        n16768) );
  NOR2_X1 U19690 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20278), .ZN(n20124) );
  OAI21_X1 U19691 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n16754), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16760) );
  NAND2_X1 U19692 ( .A1(n16723), .A2(n16755), .ZN(n16757) );
  OAI211_X1 U19693 ( .C1(n11866), .C2(n16757), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n16756), .ZN(n16758) );
  INV_X1 U19694 ( .A(n16758), .ZN(n16759) );
  AND2_X1 U19695 ( .A1(n16760), .A2(n16759), .ZN(n20128) );
  INV_X1 U19696 ( .A(n20128), .ZN(n16764) );
  NOR3_X1 U19697 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n16761), .ZN(n16763) );
  OAI21_X1 U19698 ( .B1(n20276), .B2(n16764), .A(n20278), .ZN(n16762) );
  OAI22_X1 U19699 ( .A1(n20278), .A2(n16764), .B1(n16763), .B2(n16762), .ZN(
        n16766) );
  AOI211_X1 U19700 ( .C1(n20274), .C2(n20124), .A(n16766), .B(n16765), .ZN(
        n16767) );
  NAND2_X1 U19701 ( .A1(n16768), .A2(n16767), .ZN(P2_U3176) );
  AOI221_X1 U19702 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20278), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n20128), .A(n16769), .ZN(n16770) );
  INV_X1 U19703 ( .A(n16770), .ZN(P2_U3593) );
  NAND2_X1 U19704 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16771), .ZN(
        n16772) );
  XOR2_X1 U19705 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16772), .Z(
        n16832) );
  NOR3_X4 U19706 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18251), .A3(n19212), 
        .ZN(n18093) );
  INV_X1 U19707 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21010) );
  NAND2_X1 U19708 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18209) );
  NAND2_X1 U19709 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17203) );
  NAND3_X1 U19710 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17161) );
  NOR2_X1 U19711 ( .A1(n17203), .A2(n17161), .ZN(n18078) );
  NAND2_X1 U19712 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18102) );
  NAND2_X1 U19713 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18056) );
  NAND2_X1 U19714 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18019) );
  NAND2_X1 U19715 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16977) );
  NAND2_X1 U19716 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17948) );
  INV_X1 U19717 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16971) );
  INV_X1 U19718 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19184) );
  NOR2_X1 U19719 ( .A1(n19184), .A2(n18476), .ZN(n16824) );
  INV_X1 U19720 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16773) );
  NOR2_X1 U19721 ( .A1(n16813), .A2(n16773), .ZN(n16774) );
  NOR2_X1 U19722 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19261), .ZN(n17985) );
  OAI21_X1 U19723 ( .B1(n17329), .B2(n18012), .A(n18843), .ZN(n17899) );
  NAND2_X1 U19724 ( .A1(n16774), .A2(n17899), .ZN(n16798) );
  XNOR2_X1 U19725 ( .A(n9963), .B(n21010), .ZN(n16775) );
  NOR2_X1 U19726 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18012), .ZN(
        n16810) );
  INV_X1 U19727 ( .A(n17985), .ZN(n18090) );
  OR2_X1 U19728 ( .A1(n18843), .A2(n16774), .ZN(n16814) );
  OAI211_X1 U19729 ( .C1(n16968), .C2(n18090), .A(n18242), .B(n16814), .ZN(
        n16807) );
  NOR2_X1 U19730 ( .A1(n16810), .A2(n16807), .ZN(n16797) );
  OAI22_X1 U19731 ( .A1(n16798), .A2(n16775), .B1(n9963), .B2(n16797), .ZN(
        n16776) );
  AOI211_X1 U19732 ( .C1(n18093), .C2(n17292), .A(n16824), .B(n16776), .ZN(
        n16790) );
  INV_X1 U19733 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19210) );
  AOI22_X1 U19734 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18168), .B1(
        n18052), .B2(n19210), .ZN(n16785) );
  NAND2_X1 U19735 ( .A1(n18168), .A2(n16777), .ZN(n17909) );
  OAI21_X1 U19736 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n18168), .ZN(n16778) );
  NAND3_X1 U19737 ( .A1(n17909), .A2(n16779), .A3(n16778), .ZN(n16781) );
  AOI22_X1 U19738 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18168), .B1(
        n16781), .B2(n16780), .ZN(n16784) );
  NOR2_X1 U19739 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16803), .ZN(
        n16827) );
  OAI22_X1 U19740 ( .A1(n16827), .A2(n16781), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18168), .ZN(n16782) );
  NAND2_X1 U19741 ( .A1(n16785), .A2(n16782), .ZN(n16783) );
  OAI21_X1 U19742 ( .B1(n16785), .B2(n16784), .A(n16783), .ZN(n16828) );
  NOR2_X2 U19743 ( .A1(n16946), .A2(n18613), .ZN(n18255) );
  NAND2_X1 U19744 ( .A1(n16787), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16788) );
  XNOR2_X1 U19745 ( .A(n16788), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16829) );
  NAND2_X1 U19746 ( .A1(n17751), .A2(n18255), .ZN(n18169) );
  INV_X2 U19747 ( .A(n18169), .ZN(n18123) );
  OAI211_X1 U19748 ( .C1(n18238), .C2(n16832), .A(n16790), .B(n16789), .ZN(
        P3_U2799) );
  NAND2_X1 U19749 ( .A1(n18123), .A2(n16791), .ZN(n16820) );
  NAND2_X1 U19750 ( .A1(n18254), .A2(n16792), .ZN(n16805) );
  AOI22_X1 U19751 ( .A1(n18450), .A2(n18254), .B1(n18123), .B2(n18453), .ZN(
        n18159) );
  INV_X1 U19752 ( .A(n18159), .ZN(n18125) );
  NOR2_X2 U19753 ( .A1(n18310), .A2(n18063), .ZN(n17961) );
  NAND2_X1 U19754 ( .A1(n16793), .A2(n17961), .ZN(n17921) );
  NOR3_X1 U19755 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16822), .A3(
        n17921), .ZN(n16800) );
  AOI21_X1 U19756 ( .B1(n21010), .B2(n16808), .A(n16794), .ZN(n16991) );
  AOI21_X1 U19757 ( .B1(n18093), .B2(n16991), .A(n16795), .ZN(n16796) );
  OAI221_X1 U19758 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16798), .C1(
        n21010), .C2(n16797), .A(n16796), .ZN(n16799) );
  AOI211_X1 U19759 ( .C1(n18156), .C2(n16801), .A(n16800), .B(n16799), .ZN(
        n16802) );
  OAI221_X1 U19760 ( .B1(n16803), .B2(n16820), .C1(n16803), .C2(n16805), .A(
        n16802), .ZN(P3_U2800) );
  NAND2_X1 U19761 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16804) );
  NOR2_X1 U19762 ( .A1(n16804), .A2(n18263), .ZN(n16834) );
  NOR2_X1 U19763 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16834), .ZN(
        n16819) );
  NOR2_X1 U19764 ( .A1(n17896), .A2(n16804), .ZN(n16833) );
  INV_X1 U19765 ( .A(n16833), .ZN(n16806) );
  AOI21_X1 U19766 ( .B1(n9957), .B2(n16806), .A(n16805), .ZN(n16816) );
  AOI22_X1 U19767 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18481), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16807), .ZN(n16812) );
  OAI21_X1 U19768 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16968), .A(
        n16808), .ZN(n16809) );
  INV_X1 U19769 ( .A(n16809), .ZN(n16998) );
  OAI21_X1 U19770 ( .B1(n16810), .B2(n18093), .A(n16998), .ZN(n16811) );
  OAI211_X1 U19771 ( .C1(n16814), .C2(n16813), .A(n16812), .B(n16811), .ZN(
        n16815) );
  AOI211_X1 U19772 ( .C1(n18156), .C2(n16817), .A(n16816), .B(n16815), .ZN(
        n16818) );
  OAI21_X1 U19773 ( .B1(n16820), .B2(n16819), .A(n16818), .ZN(P3_U2801) );
  NOR3_X1 U19774 ( .A1(n16822), .A2(n18498), .A3(n16821), .ZN(n16826) );
  AOI221_X1 U19775 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16823), 
        .C1(n18576), .C2(n16823), .A(n19210), .ZN(n16825) );
  AOI211_X1 U19776 ( .C1(n16827), .C2(n16826), .A(n16825), .B(n16824), .ZN(
        n16831) );
  AOI22_X1 U19777 ( .A1(n16829), .A2(n18425), .B1(n16828), .B2(n18480), .ZN(
        n16830) );
  OAI211_X1 U19778 ( .C1(n16832), .C2(n18572), .A(n16831), .B(n16830), .ZN(
        P3_U2831) );
  AOI211_X1 U19779 ( .C1(n16840), .C2(n16839), .A(n17751), .B(n19043), .ZN(
        n16837) );
  AOI22_X1 U19780 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18052), .B1(
        n18168), .B2(n17898), .ZN(n17912) );
  NAND3_X1 U19781 ( .A1(n17912), .A2(n17909), .A3(n17916), .ZN(n17910) );
  OAI22_X1 U19782 ( .A1(n16834), .A2(n18452), .B1(n16833), .B2(n18451), .ZN(
        n16835) );
  AOI211_X1 U19783 ( .C1(n16837), .C2(n17910), .A(n16836), .B(n16835), .ZN(
        n16846) );
  NAND2_X1 U19784 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18476), .ZN(
        n16845) );
  INV_X1 U19785 ( .A(n18370), .ZN(n18368) );
  NOR2_X1 U19786 ( .A1(n18368), .A2(n18030), .ZN(n18323) );
  AOI22_X1 U19787 ( .A1(n19037), .A2(n18450), .B1(n18453), .B2(n18432), .ZN(
        n18365) );
  INV_X1 U19788 ( .A(n18492), .ZN(n18563) );
  AOI22_X1 U19789 ( .A1(n19066), .A2(n18386), .B1(n18319), .B2(n18563), .ZN(
        n18416) );
  INV_X1 U19790 ( .A(n18366), .ZN(n18320) );
  AOI21_X1 U19791 ( .B1(n18365), .B2(n18416), .A(n18320), .ZN(n18311) );
  NAND3_X1 U19792 ( .A1(n18586), .A2(n18323), .A3(n18311), .ZN(n18358) );
  NOR2_X1 U19793 ( .A1(n18318), .A2(n18358), .ZN(n18332) );
  NAND2_X1 U19794 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18332), .ZN(
        n18273) );
  NOR2_X1 U19795 ( .A1(n16838), .A2(n18273), .ZN(n18268) );
  NOR2_X1 U19796 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18267), .ZN(
        n17895) );
  AOI22_X1 U19797 ( .A1(n18481), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18268), 
        .B2(n17895), .ZN(n16844) );
  NAND3_X1 U19798 ( .A1(n17898), .A2(n16840), .A3(n16839), .ZN(n16841) );
  AOI221_X1 U19799 ( .B1(n16841), .B2(n16777), .C1(n16841), .C2(n17912), .A(
        n18504), .ZN(n16842) );
  INV_X1 U19800 ( .A(n16842), .ZN(n16843) );
  OAI211_X1 U19801 ( .C1(n16846), .C2(n16845), .A(n16844), .B(n16843), .ZN(
        P3_U2834) );
  NOR3_X1 U19802 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16848) );
  NOR4_X1 U19803 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16847) );
  INV_X2 U19804 ( .A(n16932), .ZN(U215) );
  NAND4_X1 U19805 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16848), .A3(n16847), .A4(
        U215), .ZN(U213) );
  INV_X1 U19806 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19493) );
  INV_X2 U19807 ( .A(U214), .ZN(n16895) );
  OAI222_X1 U19808 ( .A1(U212), .A2(n19493), .B1(n16897), .B2(n19588), .C1(
        U214), .C2(n16933), .ZN(U216) );
  INV_X2 U19809 ( .A(U212), .ZN(n16894) );
  AOI22_X1 U19810 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16894), .ZN(n16850) );
  OAI21_X1 U19811 ( .B1(n14670), .B2(n16897), .A(n16850), .ZN(U217) );
  AOI22_X1 U19812 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16894), .ZN(n16851) );
  OAI21_X1 U19813 ( .B1(n16852), .B2(n16897), .A(n16851), .ZN(U218) );
  AOI22_X1 U19814 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16894), .ZN(n16853) );
  OAI21_X1 U19815 ( .B1(n14485), .B2(n16897), .A(n16853), .ZN(U219) );
  AOI22_X1 U19816 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16894), .ZN(n16854) );
  OAI21_X1 U19817 ( .B1(n14680), .B2(n16897), .A(n16854), .ZN(U220) );
  AOI22_X1 U19818 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16894), .ZN(n16855) );
  OAI21_X1 U19819 ( .B1(n14686), .B2(n16897), .A(n16855), .ZN(U221) );
  INV_X1 U19820 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16924) );
  INV_X1 U19821 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n21046) );
  OAI222_X1 U19822 ( .A1(U212), .A2(n16924), .B1(n16897), .B2(n14691), .C1(
        U214), .C2(n21046), .ZN(U222) );
  AOI22_X1 U19823 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16894), .ZN(n16856) );
  OAI21_X1 U19824 ( .B1(n14697), .B2(n16897), .A(n16856), .ZN(U223) );
  AOI22_X1 U19825 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16894), .ZN(n16857) );
  OAI21_X1 U19826 ( .B1(n14703), .B2(n16897), .A(n16857), .ZN(U224) );
  INV_X1 U19827 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U19828 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16894), .ZN(n16858) );
  OAI21_X1 U19829 ( .B1(n16859), .B2(n16897), .A(n16858), .ZN(U225) );
  INV_X1 U19830 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U19831 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16894), .ZN(n16860) );
  OAI21_X1 U19832 ( .B1(n16861), .B2(n16897), .A(n16860), .ZN(U226) );
  AOI22_X1 U19833 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16894), .ZN(n16862) );
  OAI21_X1 U19834 ( .B1(n14714), .B2(n16897), .A(n16862), .ZN(U227) );
  INV_X1 U19835 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16864) );
  INV_X1 U19836 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n21011) );
  OAI222_X1 U19837 ( .A1(U212), .A2(n16864), .B1(U214), .B2(n21011), .C1(
        n16863), .C2(n16897), .ZN(U228) );
  AOI22_X1 U19838 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16894), .ZN(n16865) );
  OAI21_X1 U19839 ( .B1(n14721), .B2(n16897), .A(n16865), .ZN(U229) );
  AOI22_X1 U19840 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16894), .ZN(n16866) );
  OAI21_X1 U19841 ( .B1(n14727), .B2(n16897), .A(n16866), .ZN(U230) );
  AOI22_X1 U19842 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16894), .ZN(n16867) );
  OAI21_X1 U19843 ( .B1(n14733), .B2(n16897), .A(n16867), .ZN(U231) );
  AOI22_X1 U19844 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16894), .ZN(n16868) );
  OAI21_X1 U19845 ( .B1(n12393), .B2(n16897), .A(n16868), .ZN(U232) );
  INV_X1 U19846 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16870) );
  AOI22_X1 U19847 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16894), .ZN(n16869) );
  OAI21_X1 U19848 ( .B1(n16870), .B2(n16897), .A(n16869), .ZN(U233) );
  AOI22_X1 U19849 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16894), .ZN(n16871) );
  OAI21_X1 U19850 ( .B1(n16872), .B2(n16897), .A(n16871), .ZN(U234) );
  INV_X1 U19851 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U19852 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16894), .ZN(n16873) );
  OAI21_X1 U19853 ( .B1(n16874), .B2(n16897), .A(n16873), .ZN(U235) );
  AOI22_X1 U19854 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16894), .ZN(n16875) );
  OAI21_X1 U19855 ( .B1(n16876), .B2(n16897), .A(n16875), .ZN(U236) );
  AOI22_X1 U19856 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16894), .ZN(n16877) );
  OAI21_X1 U19857 ( .B1(n12422), .B2(n16897), .A(n16877), .ZN(U237) );
  AOI22_X1 U19858 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16894), .ZN(n16878) );
  OAI21_X1 U19859 ( .B1(n16879), .B2(n16897), .A(n16878), .ZN(U238) );
  INV_X1 U19860 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n19508) );
  INV_X1 U19861 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n16880) );
  OAI222_X1 U19862 ( .A1(U212), .A2(n19508), .B1(n16897), .B2(n12427), .C1(
        U214), .C2(n16880), .ZN(U239) );
  INV_X1 U19863 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U19864 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16894), .ZN(n16881) );
  OAI21_X1 U19865 ( .B1(n21018), .B2(n16897), .A(n16881), .ZN(U240) );
  INV_X1 U19866 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16883) );
  AOI22_X1 U19867 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16894), .ZN(n16882) );
  OAI21_X1 U19868 ( .B1(n16883), .B2(n16897), .A(n16882), .ZN(U241) );
  INV_X1 U19869 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U19870 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16894), .ZN(n16884) );
  OAI21_X1 U19871 ( .B1(n16885), .B2(n16897), .A(n16884), .ZN(U242) );
  INV_X1 U19872 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U19873 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16894), .ZN(n16886) );
  OAI21_X1 U19874 ( .B1(n16887), .B2(n16897), .A(n16886), .ZN(U243) );
  INV_X1 U19875 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U19876 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16894), .ZN(n16888) );
  OAI21_X1 U19877 ( .B1(n16889), .B2(n16897), .A(n16888), .ZN(U244) );
  INV_X1 U19878 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U19879 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16894), .ZN(n16890) );
  OAI21_X1 U19880 ( .B1(n16891), .B2(n16897), .A(n16890), .ZN(U245) );
  INV_X1 U19881 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U19882 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16894), .ZN(n16892) );
  OAI21_X1 U19883 ( .B1(n16893), .B2(n16897), .A(n16892), .ZN(U246) );
  INV_X1 U19884 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U19885 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16895), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16894), .ZN(n16896) );
  OAI21_X1 U19886 ( .B1(n16898), .B2(n16897), .A(n16896), .ZN(U247) );
  OAI22_X1 U19887 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16932), .ZN(n16899) );
  INV_X1 U19888 ( .A(n16899), .ZN(U251) );
  INV_X1 U19889 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16900) );
  INV_X1 U19890 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18612) );
  AOI22_X1 U19891 ( .A1(n16932), .A2(n16900), .B1(n18612), .B2(U215), .ZN(U252) );
  INV_X1 U19892 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16901) );
  INV_X1 U19893 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18616) );
  AOI22_X1 U19894 ( .A1(n16932), .A2(n16901), .B1(n18616), .B2(U215), .ZN(U253) );
  INV_X1 U19895 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16902) );
  INV_X1 U19896 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18620) );
  AOI22_X1 U19897 ( .A1(n16932), .A2(n16902), .B1(n18620), .B2(U215), .ZN(U254) );
  INV_X1 U19898 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16903) );
  INV_X1 U19899 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18624) );
  AOI22_X1 U19900 ( .A1(n16932), .A2(n16903), .B1(n18624), .B2(U215), .ZN(U255) );
  INV_X1 U19901 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16904) );
  INV_X1 U19902 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18628) );
  AOI22_X1 U19903 ( .A1(n16932), .A2(n16904), .B1(n18628), .B2(U215), .ZN(U256) );
  INV_X1 U19904 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16905) );
  INV_X1 U19905 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18632) );
  AOI22_X1 U19906 ( .A1(n16928), .A2(n16905), .B1(n18632), .B2(U215), .ZN(U257) );
  INV_X1 U19907 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16906) );
  INV_X1 U19908 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18636) );
  AOI22_X1 U19909 ( .A1(n16928), .A2(n16906), .B1(n18636), .B2(U215), .ZN(U258) );
  INV_X1 U19910 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U19911 ( .A1(n16932), .A2(n19508), .B1(n16907), .B2(U215), .ZN(U259) );
  INV_X1 U19912 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16908) );
  INV_X1 U19913 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U19914 ( .A1(n16928), .A2(n16908), .B1(n17746), .B2(U215), .ZN(U260) );
  OAI22_X1 U19915 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16932), .ZN(n16909) );
  INV_X1 U19916 ( .A(n16909), .ZN(U261) );
  INV_X1 U19917 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16910) );
  INV_X1 U19918 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17738) );
  AOI22_X1 U19919 ( .A1(n16932), .A2(n16910), .B1(n17738), .B2(U215), .ZN(U262) );
  INV_X1 U19920 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16911) );
  INV_X1 U19921 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17734) );
  AOI22_X1 U19922 ( .A1(n16928), .A2(n16911), .B1(n17734), .B2(U215), .ZN(U263) );
  INV_X1 U19923 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16912) );
  INV_X1 U19924 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17730) );
  AOI22_X1 U19925 ( .A1(n16932), .A2(n16912), .B1(n17730), .B2(U215), .ZN(U264) );
  OAI22_X1 U19926 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16932), .ZN(n16913) );
  INV_X1 U19927 ( .A(n16913), .ZN(U265) );
  OAI22_X1 U19928 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16932), .ZN(n16914) );
  INV_X1 U19929 ( .A(n16914), .ZN(U266) );
  OAI22_X1 U19930 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16932), .ZN(n16915) );
  INV_X1 U19931 ( .A(n16915), .ZN(U267) );
  OAI22_X1 U19932 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16928), .ZN(n16916) );
  INV_X1 U19933 ( .A(n16916), .ZN(U268) );
  INV_X1 U19934 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16917) );
  INV_X1 U19935 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19563) );
  AOI22_X1 U19936 ( .A1(n16928), .A2(n16917), .B1(n19563), .B2(U215), .ZN(U269) );
  OAI22_X1 U19937 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16928), .ZN(n16918) );
  INV_X1 U19938 ( .A(n16918), .ZN(U270) );
  INV_X1 U19939 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16919) );
  INV_X1 U19940 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U19941 ( .A1(n16928), .A2(n16919), .B1(n17686), .B2(U215), .ZN(U271) );
  OAI22_X1 U19942 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16928), .ZN(n16920) );
  INV_X1 U19943 ( .A(n16920), .ZN(U272) );
  INV_X1 U19944 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16921) );
  INV_X1 U19945 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17675) );
  AOI22_X1 U19946 ( .A1(n16932), .A2(n16921), .B1(n17675), .B2(U215), .ZN(U273) );
  OAI22_X1 U19947 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16932), .ZN(n16922) );
  INV_X1 U19948 ( .A(n16922), .ZN(U274) );
  INV_X1 U19949 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U19950 ( .A1(n16932), .A2(n16923), .B1(n15349), .B2(U215), .ZN(U275) );
  AOI22_X1 U19951 ( .A1(n16932), .A2(n16924), .B1(n15339), .B2(U215), .ZN(U276) );
  OAI22_X1 U19952 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16932), .ZN(n16925) );
  INV_X1 U19953 ( .A(n16925), .ZN(U277) );
  OAI22_X1 U19954 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16932), .ZN(n16926) );
  INV_X1 U19955 ( .A(n16926), .ZN(U278) );
  INV_X1 U19956 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16927) );
  INV_X1 U19957 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19573) );
  AOI22_X1 U19958 ( .A1(n16928), .A2(n16927), .B1(n19573), .B2(U215), .ZN(U279) );
  OAI22_X1 U19959 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16932), .ZN(n16929) );
  INV_X1 U19960 ( .A(n16929), .ZN(U280) );
  OAI22_X1 U19961 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16932), .ZN(n16930) );
  INV_X1 U19962 ( .A(n16930), .ZN(U281) );
  INV_X1 U19963 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19586) );
  AOI22_X1 U19964 ( .A1(n16932), .A2(n19493), .B1(n19586), .B2(U215), .ZN(U282) );
  INV_X1 U19965 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17785) );
  AOI222_X1 U19966 ( .A1(n16933), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19493), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17785), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16934) );
  INV_X2 U19967 ( .A(n16936), .ZN(n16935) );
  INV_X1 U19968 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19144) );
  INV_X1 U19969 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20167) );
  AOI22_X1 U19970 ( .A1(n16935), .A2(n19144), .B1(n20167), .B2(n16936), .ZN(
        U347) );
  INV_X1 U19971 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19142) );
  INV_X1 U19972 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20165) );
  AOI22_X1 U19973 ( .A1(n16935), .A2(n19142), .B1(n20165), .B2(n16936), .ZN(
        U348) );
  INV_X1 U19974 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19140) );
  INV_X1 U19975 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20163) );
  AOI22_X1 U19976 ( .A1(n16935), .A2(n19140), .B1(n20163), .B2(n16936), .ZN(
        U349) );
  INV_X1 U19977 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19138) );
  INV_X1 U19978 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U19979 ( .A1(n16935), .A2(n19138), .B1(n20161), .B2(n16936), .ZN(
        U350) );
  INV_X1 U19980 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19136) );
  INV_X1 U19981 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20160) );
  AOI22_X1 U19982 ( .A1(n16935), .A2(n19136), .B1(n20160), .B2(n16936), .ZN(
        U351) );
  INV_X1 U19983 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19133) );
  INV_X1 U19984 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20158) );
  AOI22_X1 U19985 ( .A1(n16935), .A2(n19133), .B1(n20158), .B2(n16936), .ZN(
        U352) );
  INV_X1 U19986 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19132) );
  INV_X1 U19987 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20156) );
  AOI22_X1 U19988 ( .A1(n16935), .A2(n19132), .B1(n20156), .B2(n16936), .ZN(
        U353) );
  INV_X1 U19989 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19130) );
  AOI22_X1 U19990 ( .A1(n16935), .A2(n19130), .B1(n20153), .B2(n16936), .ZN(
        U354) );
  INV_X1 U19991 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19185) );
  INV_X1 U19992 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20205) );
  AOI22_X1 U19993 ( .A1(n16935), .A2(n19185), .B1(n20205), .B2(n16936), .ZN(
        U355) );
  INV_X1 U19994 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19182) );
  INV_X1 U19995 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20201) );
  AOI22_X1 U19996 ( .A1(n16935), .A2(n19182), .B1(n20201), .B2(n16936), .ZN(
        U356) );
  INV_X1 U19997 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19179) );
  INV_X1 U19998 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20200) );
  AOI22_X1 U19999 ( .A1(n16935), .A2(n19179), .B1(n20200), .B2(n16936), .ZN(
        U357) );
  INV_X1 U20000 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19178) );
  INV_X1 U20001 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20198) );
  AOI22_X1 U20002 ( .A1(n16935), .A2(n19178), .B1(n20198), .B2(n16936), .ZN(
        U358) );
  INV_X1 U20003 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19176) );
  INV_X1 U20004 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20196) );
  AOI22_X1 U20005 ( .A1(n16935), .A2(n19176), .B1(n20196), .B2(n16936), .ZN(
        U359) );
  INV_X1 U20006 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19174) );
  INV_X1 U20007 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20194) );
  AOI22_X1 U20008 ( .A1(n16935), .A2(n19174), .B1(n20194), .B2(n16936), .ZN(
        U360) );
  INV_X1 U20009 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19172) );
  INV_X1 U20010 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20192) );
  AOI22_X1 U20011 ( .A1(n16935), .A2(n19172), .B1(n20192), .B2(n16936), .ZN(
        U361) );
  INV_X1 U20012 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19169) );
  INV_X1 U20013 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20190) );
  AOI22_X1 U20014 ( .A1(n16935), .A2(n19169), .B1(n20190), .B2(n16936), .ZN(
        U362) );
  INV_X1 U20015 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19168) );
  INV_X1 U20016 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20188) );
  AOI22_X1 U20017 ( .A1(n16935), .A2(n19168), .B1(n20188), .B2(n16936), .ZN(
        U363) );
  INV_X1 U20018 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19166) );
  INV_X1 U20019 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20186) );
  AOI22_X1 U20020 ( .A1(n16935), .A2(n19166), .B1(n20186), .B2(n16936), .ZN(
        U364) );
  INV_X1 U20021 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19128) );
  INV_X1 U20022 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20151) );
  AOI22_X1 U20023 ( .A1(n16935), .A2(n19128), .B1(n20151), .B2(n16936), .ZN(
        U365) );
  INV_X1 U20024 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19163) );
  INV_X1 U20025 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20184) );
  AOI22_X1 U20026 ( .A1(n16935), .A2(n19163), .B1(n20184), .B2(n16936), .ZN(
        U366) );
  INV_X1 U20027 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19162) );
  INV_X1 U20028 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20182) );
  AOI22_X1 U20029 ( .A1(n16935), .A2(n19162), .B1(n20182), .B2(n16936), .ZN(
        U367) );
  INV_X1 U20030 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19160) );
  INV_X1 U20031 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20181) );
  AOI22_X1 U20032 ( .A1(n16935), .A2(n19160), .B1(n20181), .B2(n16936), .ZN(
        U368) );
  INV_X1 U20033 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19158) );
  INV_X1 U20034 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20179) );
  AOI22_X1 U20035 ( .A1(n16935), .A2(n19158), .B1(n20179), .B2(n16936), .ZN(
        U369) );
  INV_X1 U20036 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19156) );
  INV_X1 U20037 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20177) );
  AOI22_X1 U20038 ( .A1(n16935), .A2(n19156), .B1(n20177), .B2(n16936), .ZN(
        U370) );
  INV_X1 U20039 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19154) );
  INV_X1 U20040 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20175) );
  AOI22_X1 U20041 ( .A1(n16935), .A2(n19154), .B1(n20175), .B2(n16936), .ZN(
        U371) );
  INV_X1 U20042 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19151) );
  INV_X1 U20043 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20173) );
  AOI22_X1 U20044 ( .A1(n16935), .A2(n19151), .B1(n20173), .B2(n16936), .ZN(
        U372) );
  INV_X1 U20045 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19150) );
  INV_X1 U20046 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20171) );
  AOI22_X1 U20047 ( .A1(n16935), .A2(n19150), .B1(n20171), .B2(n16936), .ZN(
        U373) );
  INV_X1 U20048 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19148) );
  INV_X1 U20049 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20169) );
  AOI22_X1 U20050 ( .A1(n16935), .A2(n19148), .B1(n20169), .B2(n16936), .ZN(
        U374) );
  INV_X1 U20051 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19146) );
  INV_X1 U20052 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20168) );
  AOI22_X1 U20053 ( .A1(n16935), .A2(n19146), .B1(n20168), .B2(n16936), .ZN(
        U375) );
  INV_X1 U20054 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19126) );
  INV_X1 U20055 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U20056 ( .A1(n16935), .A2(n19126), .B1(n20150), .B2(n16936), .ZN(
        U376) );
  INV_X1 U20057 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16938) );
  INV_X1 U20058 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19125) );
  NAND2_X1 U20059 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19125), .ZN(n16937) );
  AOI22_X1 U20060 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n16937), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19110), .ZN(n19199) );
  OAI21_X1 U20061 ( .B1(n19122), .B2(n16938), .A(n19196), .ZN(P3_U2633) );
  NAND2_X1 U20062 ( .A1(n19262), .A2(n19261), .ZN(n16941) );
  INV_X1 U20063 ( .A(n16945), .ZN(n16939) );
  OAI21_X1 U20064 ( .B1(n16939), .B2(n17825), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16940) );
  OAI21_X1 U20065 ( .B1(n16941), .B2(n19249), .A(n16940), .ZN(P3_U2634) );
  NOR2_X1 U20066 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16943) );
  AOI22_X1 U20067 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n19258), .B1(n16943), .B2(
        n19122), .ZN(n16942) );
  OAI21_X1 U20068 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n19258), .A(n16942), 
        .ZN(P3_U2635) );
  OAI21_X1 U20069 ( .B1(n16943), .B2(BS16), .A(n19199), .ZN(n19197) );
  OAI21_X1 U20070 ( .B1(n19199), .B2(n16967), .A(n19197), .ZN(P3_U2636) );
  AND3_X1 U20071 ( .A1(n19041), .A2(n16945), .A3(n16944), .ZN(n19044) );
  NOR2_X1 U20072 ( .A1(n19044), .A2(n19254), .ZN(n19243) );
  OAI21_X1 U20073 ( .B1(n19243), .B2(n18598), .A(n16946), .ZN(P3_U2637) );
  NOR4_X1 U20074 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16950) );
  NOR4_X1 U20075 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16949) );
  NOR4_X1 U20076 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16948) );
  NOR4_X1 U20077 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16947) );
  NAND4_X1 U20078 ( .A1(n16950), .A2(n16949), .A3(n16948), .A4(n16947), .ZN(
        n16956) );
  NOR4_X1 U20079 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16954) );
  AOI211_X1 U20080 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16953) );
  NOR4_X1 U20081 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16952) );
  NOR4_X1 U20082 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16951) );
  NAND4_X1 U20083 ( .A1(n16954), .A2(n16953), .A3(n16952), .A4(n16951), .ZN(
        n16955) );
  NOR2_X1 U20084 ( .A1(n16956), .A2(n16955), .ZN(n19241) );
  INV_X1 U20085 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19192) );
  NOR3_X1 U20086 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16958) );
  OAI21_X1 U20087 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16958), .A(n19241), .ZN(
        n16957) );
  OAI21_X1 U20088 ( .B1(n19241), .B2(n19192), .A(n16957), .ZN(P3_U2638) );
  INV_X1 U20089 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19234) );
  INV_X1 U20090 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19198) );
  AOI21_X1 U20091 ( .B1(n19234), .B2(n19198), .A(n16958), .ZN(n16959) );
  INV_X1 U20092 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19189) );
  INV_X1 U20093 ( .A(n19241), .ZN(n19236) );
  AOI22_X1 U20094 ( .A1(n19241), .A2(n16959), .B1(n19189), .B2(n19236), .ZN(
        P3_U2639) );
  INV_X1 U20095 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19171) );
  INV_X1 U20096 ( .A(n16960), .ZN(n16962) );
  NOR4_X4 U20097 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n19212), .ZN(n17239) );
  NAND2_X1 U20098 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19261), .ZN(n18976) );
  NOR2_X1 U20099 ( .A1(n19102), .A2(n18976), .ZN(n19094) );
  INV_X1 U20100 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19161) );
  INV_X1 U20101 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19159) );
  INV_X1 U20102 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19147) );
  INV_X1 U20103 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19139) );
  INV_X1 U20104 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19131) );
  NAND3_X1 U20105 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17281) );
  NOR2_X1 U20106 ( .A1(n19131), .A2(n17281), .ZN(n17266) );
  NAND2_X1 U20107 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17266), .ZN(n17237) );
  NAND2_X1 U20108 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17242) );
  NOR3_X1 U20109 ( .A1(n19139), .A2(n17237), .A3(n17242), .ZN(n17200) );
  NAND4_X1 U20110 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_9__SCAN_IN), .A4(n17200), .ZN(n17186) );
  NOR2_X1 U20111 ( .A1(n19147), .A2(n17186), .ZN(n17166) );
  NAND3_X1 U20112 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17166), .ZN(n17091) );
  NAND3_X1 U20113 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n17107) );
  NOR4_X1 U20114 ( .A1(n19161), .A2(n19159), .A3(n17091), .A4(n17107), .ZN(
        n17088) );
  NAND2_X1 U20115 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17088), .ZN(n16982) );
  NOR2_X1 U20116 ( .A1(n17333), .A2(n16982), .ZN(n17073) );
  NAND4_X1 U20117 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17073), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n17048) );
  NOR2_X1 U20118 ( .A1(n19171), .A2(n17048), .ZN(n17037) );
  NAND3_X1 U20119 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n17037), .ZN(n17006) );
  NAND3_X1 U20120 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16963) );
  INV_X1 U20121 ( .A(n17333), .ZN(n17282) );
  INV_X1 U20122 ( .A(n19116), .ZN(n19245) );
  OAI211_X1 U20123 ( .C1(n19246), .C2(n19245), .A(n19093), .B(n16967), .ZN(
        n19092) );
  NAND2_X1 U20124 ( .A1(n17282), .A2(n17326), .ZN(n17335) );
  OAI21_X1 U20125 ( .B1(n17006), .B2(n16963), .A(n17335), .ZN(n16999) );
  INV_X1 U20126 ( .A(n19092), .ZN(n16964) );
  AOI211_X4 U20127 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19246), .A(n16964), .B(
        n16966), .ZN(n17337) );
  AOI22_X1 U20128 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n17305), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17337), .ZN(n16987) );
  NAND2_X1 U20129 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19246), .ZN(n16965) );
  AOI211_X4 U20130 ( .C1(n16967), .C2(n19093), .A(n16966), .B(n16965), .ZN(
        n17336) );
  NOR3_X1 U20131 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17311) );
  INV_X1 U20132 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17300) );
  NAND2_X1 U20133 ( .A1(n17311), .A2(n17300), .ZN(n17299) );
  INV_X1 U20134 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17595) );
  NAND2_X1 U20135 ( .A1(n17283), .A2(n17595), .ZN(n17272) );
  NAND2_X1 U20136 ( .A1(n17252), .A2(n20911), .ZN(n17246) );
  NAND2_X1 U20137 ( .A1(n17226), .A2(n17220), .ZN(n17219) );
  NAND2_X1 U20138 ( .A1(n17198), .A2(n17194), .ZN(n17193) );
  NAND2_X1 U20139 ( .A1(n17177), .A2(n17168), .ZN(n17167) );
  NAND2_X1 U20140 ( .A1(n17155), .A2(n17148), .ZN(n17147) );
  NAND2_X1 U20141 ( .A1(n17128), .A2(n17469), .ZN(n17117) );
  INV_X1 U20142 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17452) );
  NAND2_X1 U20143 ( .A1(n17104), .A2(n17452), .ZN(n17097) );
  INV_X1 U20144 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17428) );
  NAND2_X1 U20145 ( .A1(n17084), .A2(n17428), .ZN(n17078) );
  NAND2_X1 U20146 ( .A1(n17065), .A2(n17343), .ZN(n17060) );
  NAND2_X1 U20147 ( .A1(n17045), .A2(n17041), .ZN(n17040) );
  INV_X1 U20148 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17384) );
  NAND2_X1 U20149 ( .A1(n17024), .A2(n17384), .ZN(n17020) );
  NOR2_X1 U20150 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17020), .ZN(n17007) );
  INV_X1 U20151 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17374) );
  NAND2_X1 U20152 ( .A1(n17007), .A2(n17374), .ZN(n16988) );
  NOR2_X1 U20153 ( .A1(n17325), .A2(n16988), .ZN(n16994) );
  INV_X1 U20154 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17348) );
  NAND2_X1 U20155 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9769), .ZN(
        n16969) );
  AOI21_X1 U20156 ( .B1(n9975), .B2(n16969), .A(n16968), .ZN(n17908) );
  OR2_X1 U20157 ( .A1(n17329), .A2(n17902), .ZN(n16972) );
  INV_X1 U20158 ( .A(n16969), .ZN(n16970) );
  AOI21_X1 U20159 ( .B1(n16971), .B2(n16972), .A(n16970), .ZN(n17919) );
  NOR2_X1 U20160 ( .A1(n17329), .A2(n17947), .ZN(n16978) );
  INV_X1 U20161 ( .A(n16978), .ZN(n16976) );
  NOR2_X1 U20162 ( .A1(n17948), .A2(n16976), .ZN(n17900) );
  OAI21_X1 U20163 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17900), .A(
        n16972), .ZN(n16973) );
  INV_X1 U20164 ( .A(n16973), .ZN(n17933) );
  INV_X1 U20165 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16975) );
  NAND2_X1 U20166 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16978), .ZN(
        n16974) );
  AOI21_X1 U20167 ( .B1(n16975), .B2(n16974), .A(n17900), .ZN(n17940) );
  INV_X1 U20168 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U20169 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16978), .B1(
        n16976), .B2(n17954), .ZN(n17952) );
  INV_X1 U20170 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17973) );
  INV_X1 U20171 ( .A(n16977), .ZN(n17982) );
  INV_X1 U20172 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17987) );
  INV_X1 U20173 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18034) );
  NOR2_X1 U20174 ( .A1(n17329), .A2(n18055), .ZN(n18054) );
  INV_X1 U20175 ( .A(n18054), .ZN(n17140) );
  NOR2_X1 U20176 ( .A1(n18056), .A2(n17140), .ZN(n17114) );
  NAND2_X1 U20177 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17114), .ZN(
        n17113) );
  NOR2_X1 U20178 ( .A1(n18034), .A2(n17113), .ZN(n17093) );
  NAND2_X1 U20179 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17093), .ZN(
        n17984) );
  NOR2_X1 U20180 ( .A1(n17987), .A2(n17984), .ZN(n16981) );
  NAND2_X1 U20181 ( .A1(n17982), .A2(n16981), .ZN(n17939) );
  AOI21_X1 U20182 ( .B1(n17973), .B2(n17939), .A(n16978), .ZN(n17970) );
  INV_X1 U20183 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17990) );
  NAND2_X1 U20184 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16981), .ZN(
        n16979) );
  INV_X1 U20185 ( .A(n17939), .ZN(n17968) );
  AOI21_X1 U20186 ( .B1(n17990), .B2(n16979), .A(n17968), .ZN(n17988) );
  INV_X1 U20187 ( .A(n16981), .ZN(n16980) );
  INV_X1 U20188 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U20189 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16981), .B1(
        n16980), .B2(n17996), .ZN(n17999) );
  AOI21_X1 U20190 ( .B1(n17987), .B2(n17984), .A(n16981), .ZN(n18013) );
  INV_X1 U20191 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18257) );
  INV_X1 U20192 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18071) );
  NOR2_X1 U20193 ( .A1(n18071), .A2(n17140), .ZN(n17139) );
  NAND2_X1 U20194 ( .A1(n18257), .A2(n17139), .ZN(n17133) );
  NOR2_X1 U20195 ( .A1(n17999), .A2(n17075), .ZN(n17074) );
  NOR2_X1 U20196 ( .A1(n17074), .A2(n17261), .ZN(n17067) );
  NOR2_X1 U20197 ( .A1(n17988), .A2(n17067), .ZN(n17066) );
  NOR2_X1 U20198 ( .A1(n17066), .A2(n17261), .ZN(n17056) );
  NOR2_X1 U20199 ( .A1(n17970), .A2(n17056), .ZN(n17055) );
  NOR2_X1 U20200 ( .A1(n17055), .A2(n17261), .ZN(n17047) );
  NOR2_X1 U20201 ( .A1(n17952), .A2(n17047), .ZN(n17046) );
  NOR2_X1 U20202 ( .A1(n17046), .A2(n17261), .ZN(n17035) );
  NOR2_X1 U20203 ( .A1(n17940), .A2(n17035), .ZN(n17034) );
  NOR2_X1 U20204 ( .A1(n17034), .A2(n17261), .ZN(n17026) );
  NOR2_X1 U20205 ( .A1(n17933), .A2(n17026), .ZN(n17025) );
  NOR2_X1 U20206 ( .A1(n17008), .A2(n17261), .ZN(n16997) );
  NOR2_X1 U20207 ( .A1(n16998), .A2(n16997), .ZN(n16996) );
  NAND2_X1 U20208 ( .A1(n17292), .A2(n17239), .ZN(n17323) );
  NOR3_X1 U20209 ( .A1(n16991), .A2(n16990), .A3(n17323), .ZN(n16985) );
  INV_X1 U20210 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19175) );
  NAND2_X1 U20211 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16983) );
  NAND2_X1 U20212 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17054), .ZN(n17050) );
  NOR2_X1 U20213 ( .A1(n19171), .A2(n17050), .ZN(n17033) );
  NAND2_X1 U20214 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17033), .ZN(n17029) );
  NAND4_X1 U20215 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17015), .ZN(n16992) );
  AOI221_X1 U20216 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n19184), .C2(n19186), .A(n16992), .ZN(n16984) );
  AOI211_X1 U20217 ( .C1(n16994), .C2(n17348), .A(n16985), .B(n16984), .ZN(
        n16986) );
  OAI211_X1 U20218 ( .C1(n19184), .C2(n16999), .A(n16987), .B(n16986), .ZN(
        P3_U2640) );
  NAND2_X1 U20219 ( .A1(n17336), .A2(n16988), .ZN(n17004) );
  OAI21_X1 U20220 ( .B1(n16991), .B2(n16990), .A(n17239), .ZN(n16989) );
  AOI22_X1 U20221 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16999), .B1(n16992), 
        .B2(n19186), .ZN(n16993) );
  OAI21_X1 U20222 ( .B1(n17337), .B2(n16994), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16995) );
  NOR2_X1 U20223 ( .A1(n17007), .A2(n17374), .ZN(n17005) );
  AOI211_X1 U20224 ( .C1(n16998), .C2(n16997), .A(n16996), .B(n19105), .ZN(
        n17001) );
  INV_X1 U20225 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19181) );
  OAI22_X1 U20226 ( .A1(n19181), .A2(n16999), .B1(n17275), .B2(n17374), .ZN(
        n17000) );
  AOI211_X1 U20227 ( .C1(n17267), .C2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17001), .B(n17000), .ZN(n17003) );
  NAND4_X1 U20228 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17015), .A4(n19181), .ZN(n17002) );
  OAI211_X1 U20229 ( .C1(n17005), .C2(n17004), .A(n17003), .B(n17002), .ZN(
        P3_U2642) );
  INV_X1 U20230 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19180) );
  NAND2_X1 U20231 ( .A1(n17335), .A2(n17006), .ZN(n17028) );
  AOI22_X1 U20232 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17267), .B1(
        n17337), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17014) );
  INV_X1 U20233 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19177) );
  AOI22_X1 U20234 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .B1(n19177), .B2(n19180), .ZN(n17012) );
  AOI211_X1 U20235 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17020), .A(n17007), .B(
        n17325), .ZN(n17011) );
  AOI211_X1 U20236 ( .C1(n17908), .C2(n17009), .A(n17008), .B(n19105), .ZN(
        n17010) );
  AOI211_X1 U20237 ( .C1(n17015), .C2(n17012), .A(n17011), .B(n17010), .ZN(
        n17013) );
  OAI211_X1 U20238 ( .C1(n19180), .C2(n17028), .A(n17014), .B(n17013), .ZN(
        P3_U2643) );
  INV_X1 U20239 ( .A(n17015), .ZN(n17023) );
  AOI211_X1 U20240 ( .C1(n17919), .C2(n17017), .A(n17016), .B(n19105), .ZN(
        n17019) );
  OAI22_X1 U20241 ( .A1(n17384), .A2(n17275), .B1(n19177), .B2(n17028), .ZN(
        n17018) );
  AOI211_X1 U20242 ( .C1(n17267), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17019), .B(n17018), .ZN(n17022) );
  OAI211_X1 U20243 ( .C1(n17024), .C2(n17384), .A(n17336), .B(n17020), .ZN(
        n17021) );
  OAI211_X1 U20244 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17023), .A(n17022), 
        .B(n17021), .ZN(P3_U2644) );
  AOI211_X1 U20245 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17040), .A(n17024), .B(
        n17325), .ZN(n17032) );
  AOI211_X1 U20246 ( .C1(n17933), .C2(n17026), .A(n17025), .B(n19105), .ZN(
        n17031) );
  AOI22_X1 U20247 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17267), .B1(
        n17337), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17027) );
  OAI221_X1 U20248 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n17029), .C1(n19175), 
        .C2(n17028), .A(n17027), .ZN(n17030) );
  OR3_X1 U20249 ( .A1(n17032), .A2(n17031), .A3(n17030), .ZN(P3_U2645) );
  INV_X1 U20250 ( .A(n17033), .ZN(n17044) );
  AOI211_X1 U20251 ( .C1(n17940), .C2(n17035), .A(n17034), .B(n19105), .ZN(
        n17039) );
  NAND2_X1 U20252 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17335), .ZN(n17036) );
  OAI22_X1 U20253 ( .A1(n17037), .A2(n17036), .B1(n17275), .B2(n17041), .ZN(
        n17038) );
  AOI211_X1 U20254 ( .C1(n17267), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17039), .B(n17038), .ZN(n17043) );
  OAI211_X1 U20255 ( .C1(n17045), .C2(n17041), .A(n17336), .B(n17040), .ZN(
        n17042) );
  OAI211_X1 U20256 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n17044), .A(n17043), 
        .B(n17042), .ZN(P3_U2646) );
  AOI211_X1 U20257 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17060), .A(n17045), .B(
        n17325), .ZN(n17053) );
  AOI211_X1 U20258 ( .C1(n17952), .C2(n17047), .A(n17046), .B(n19105), .ZN(
        n17052) );
  NAND2_X1 U20259 ( .A1(n17335), .A2(n17048), .ZN(n17057) );
  AOI22_X1 U20260 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17267), .B1(
        n17337), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n17049) );
  OAI221_X1 U20261 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17050), .C1(n19171), 
        .C2(n17057), .A(n17049), .ZN(n17051) );
  OR3_X1 U20262 ( .A1(n17053), .A2(n17052), .A3(n17051), .ZN(P3_U2647) );
  INV_X1 U20263 ( .A(n17054), .ZN(n17063) );
  AOI211_X1 U20264 ( .C1(n17970), .C2(n17056), .A(n17055), .B(n19105), .ZN(
        n17059) );
  INV_X1 U20265 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19170) );
  OAI22_X1 U20266 ( .A1(n19170), .A2(n17057), .B1(n17275), .B2(n17343), .ZN(
        n17058) );
  AOI211_X1 U20267 ( .C1(n17267), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17059), .B(n17058), .ZN(n17062) );
  OAI211_X1 U20268 ( .C1(n17065), .C2(n17343), .A(n17336), .B(n17060), .ZN(
        n17061) );
  OAI211_X1 U20269 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n17063), .A(n17062), 
        .B(n17061), .ZN(P3_U2648) );
  NOR2_X1 U20270 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17081), .ZN(n17064) );
  AOI22_X1 U20271 ( .A1(n17337), .A2(P3_EBX_REG_22__SCAN_IN), .B1(
        P3_REIP_REG_21__SCAN_IN), .B2(n17064), .ZN(n17072) );
  INV_X1 U20272 ( .A(n17335), .ZN(n17092) );
  OAI22_X1 U20273 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n17081), .B1(n17092), 
        .B2(n17073), .ZN(n17070) );
  AOI211_X1 U20274 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17078), .A(n17065), .B(
        n17325), .ZN(n17069) );
  AOI211_X1 U20275 ( .C1(n17988), .C2(n17067), .A(n17066), .B(n19105), .ZN(
        n17068) );
  AOI211_X1 U20276 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17070), .A(n17069), 
        .B(n17068), .ZN(n17071) );
  OAI211_X1 U20277 ( .C1(n17990), .C2(n17322), .A(n17072), .B(n17071), .ZN(
        P3_U2649) );
  NOR2_X1 U20278 ( .A1(n17092), .A2(n17073), .ZN(n17087) );
  AOI211_X1 U20279 ( .C1(n17999), .C2(n17075), .A(n17074), .B(n19105), .ZN(
        n17077) );
  OAI22_X1 U20280 ( .A1(n17996), .A2(n17322), .B1(n17275), .B2(n17428), .ZN(
        n17076) );
  AOI211_X1 U20281 ( .C1(n17087), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17077), 
        .B(n17076), .ZN(n17080) );
  OAI211_X1 U20282 ( .C1(n17084), .C2(n17428), .A(n17336), .B(n17078), .ZN(
        n17079) );
  OAI211_X1 U20283 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n17081), .A(n17080), 
        .B(n17079), .ZN(P3_U2650) );
  AOI211_X1 U20284 ( .C1(n18013), .C2(n17083), .A(n17082), .B(n19105), .ZN(
        n17086) );
  AOI211_X1 U20285 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17097), .A(n17084), .B(
        n17325), .ZN(n17085) );
  AOI211_X1 U20286 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17337), .A(n17086), .B(
        n17085), .ZN(n17090) );
  OAI221_X1 U20287 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n17310), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n17088), .A(n17087), .ZN(n17089) );
  OAI211_X1 U20288 ( .C1(n17322), .C2(n17987), .A(n17090), .B(n17089), .ZN(
        P3_U2651) );
  AOI22_X1 U20289 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17305), .B1(
        n17337), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n17100) );
  NAND4_X1 U20290 ( .A1(n17310), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .A4(n17166), .ZN(n17143) );
  NOR3_X1 U20291 ( .A1(n19159), .A2(n17107), .A3(n17143), .ZN(n17096) );
  AOI21_X1 U20292 ( .B1(n17091), .B2(n17310), .A(n17333), .ZN(n17153) );
  INV_X1 U20293 ( .A(n17153), .ZN(n17127) );
  AOI21_X1 U20294 ( .B1(n17310), .B2(n17107), .A(n17127), .ZN(n17120) );
  OAI21_X1 U20295 ( .B1(n17092), .B2(P3_REIP_REG_18__SCAN_IN), .A(n17120), 
        .ZN(n17108) );
  OAI21_X1 U20296 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17093), .A(
        n17984), .ZN(n18021) );
  INV_X1 U20297 ( .A(n17093), .ZN(n17101) );
  OAI21_X1 U20298 ( .B1(n17101), .B2(n17133), .A(n17292), .ZN(n17103) );
  OAI21_X1 U20299 ( .B1(n18021), .B2(n17103), .A(n17239), .ZN(n17094) );
  AOI21_X1 U20300 ( .B1(n18021), .B2(n17103), .A(n17094), .ZN(n17095) );
  AOI221_X1 U20301 ( .B1(n17096), .B2(n19161), .C1(n17108), .C2(
        P3_REIP_REG_19__SCAN_IN), .A(n17095), .ZN(n17099) );
  OAI211_X1 U20302 ( .C1(n17104), .C2(n17452), .A(n17336), .B(n17097), .ZN(
        n17098) );
  NAND4_X1 U20303 ( .A1(n17100), .A2(n17099), .A3(n18476), .A4(n17098), .ZN(
        P3_U2652) );
  AOI21_X1 U20304 ( .B1(n17337), .B2(P3_EBX_REG_18__SCAN_IN), .A(n18481), .ZN(
        n17112) );
  INV_X1 U20305 ( .A(n17113), .ZN(n18017) );
  OAI21_X1 U20306 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18017), .A(
        n17101), .ZN(n18031) );
  NAND2_X1 U20307 ( .A1(n17239), .A2(n17261), .ZN(n17320) );
  INV_X1 U20308 ( .A(n17133), .ZN(n17138) );
  OAI221_X1 U20309 ( .B1(n18031), .B2(n17138), .C1(n18031), .C2(n18034), .A(
        n17239), .ZN(n17102) );
  AOI22_X1 U20310 ( .A1(n18031), .A2(n17103), .B1(n17320), .B2(n17102), .ZN(
        n17106) );
  AOI211_X1 U20311 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17117), .A(n17104), .B(
        n17325), .ZN(n17105) );
  AOI211_X1 U20312 ( .C1(n17305), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17106), .B(n17105), .ZN(n17111) );
  NOR2_X1 U20313 ( .A1(n17107), .A2(n17143), .ZN(n17109) );
  OAI21_X1 U20314 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17109), .A(n17108), 
        .ZN(n17110) );
  NAND3_X1 U20315 ( .A1(n17112), .A2(n17111), .A3(n17110), .ZN(P3_U2653) );
  OAI21_X1 U20316 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17114), .A(
        n17113), .ZN(n18050) );
  INV_X1 U20317 ( .A(n17114), .ZN(n17115) );
  OAI21_X1 U20318 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17139), .A(
        n17115), .ZN(n18059) );
  AOI21_X1 U20319 ( .B1(n17138), .B2(n18059), .A(n17261), .ZN(n17116) );
  XOR2_X1 U20320 ( .A(n18050), .B(n17116), .Z(n17126) );
  OAI211_X1 U20321 ( .C1(n17128), .C2(n17469), .A(n17336), .B(n17117), .ZN(
        n17118) );
  OAI211_X1 U20322 ( .C1(n17275), .C2(n17469), .A(n18476), .B(n17118), .ZN(
        n17124) );
  NAND2_X1 U20323 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17119) );
  NOR2_X1 U20324 ( .A1(n17119), .A2(n17143), .ZN(n17122) );
  INV_X1 U20325 ( .A(n17120), .ZN(n17121) );
  MUX2_X1 U20326 ( .A(n17122), .B(n17121), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n17123) );
  AOI211_X1 U20327 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n17267), .A(
        n17124), .B(n17123), .ZN(n17125) );
  OAI21_X1 U20328 ( .B1(n19105), .B2(n17126), .A(n17125), .ZN(P3_U2654) );
  INV_X1 U20329 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19153) );
  AOI21_X1 U20330 ( .B1(n17310), .B2(n19153), .A(n17127), .ZN(n17142) );
  INV_X1 U20331 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19155) );
  NOR3_X1 U20332 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n19153), .A3(n17143), 
        .ZN(n17132) );
  AOI211_X1 U20333 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17147), .A(n17128), .B(
        n17325), .ZN(n17131) );
  AOI22_X1 U20334 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17267), .B1(
        n17337), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n17129) );
  INV_X1 U20335 ( .A(n17129), .ZN(n17130) );
  NOR4_X1 U20336 ( .A1(n18481), .A2(n17132), .A3(n17131), .A4(n17130), .ZN(
        n17137) );
  NAND2_X1 U20337 ( .A1(n17292), .A2(n17133), .ZN(n17135) );
  OAI21_X1 U20338 ( .B1(n17138), .B2(n17261), .A(n18059), .ZN(n17134) );
  OAI211_X1 U20339 ( .C1(n18059), .C2(n17135), .A(n17239), .B(n17134), .ZN(
        n17136) );
  OAI211_X1 U20340 ( .C1(n17142), .C2(n19155), .A(n17137), .B(n17136), .ZN(
        P3_U2655) );
  AOI22_X1 U20341 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17267), .B1(
        n17337), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n17151) );
  NOR2_X1 U20342 ( .A1(n17138), .A2(n17323), .ZN(n17146) );
  AOI21_X1 U20343 ( .B1(n18071), .B2(n17140), .A(n17139), .ZN(n17141) );
  INV_X1 U20344 ( .A(n17141), .ZN(n18068) );
  OAI21_X1 U20345 ( .B1(n17261), .B2(n18257), .A(n17239), .ZN(n17324) );
  AOI211_X1 U20346 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17320), .A(
        n17324), .B(n18068), .ZN(n17145) );
  AOI21_X1 U20347 ( .B1(n19153), .B2(n17143), .A(n17142), .ZN(n17144) );
  AOI211_X1 U20348 ( .C1(n17146), .C2(n18068), .A(n17145), .B(n17144), .ZN(
        n17150) );
  OAI211_X1 U20349 ( .C1(n17155), .C2(n17148), .A(n17336), .B(n17147), .ZN(
        n17149) );
  NAND4_X1 U20350 ( .A1(n17151), .A2(n17150), .A3(n18476), .A4(n17149), .ZN(
        P3_U2656) );
  NAND2_X1 U20351 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17162), .ZN(
        n17152) );
  AOI21_X1 U20352 ( .B1(n9967), .B2(n17152), .A(n18054), .ZN(n18081) );
  NOR2_X1 U20353 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17329), .ZN(
        n17278) );
  AOI21_X1 U20354 ( .B1(n17162), .B2(n17278), .A(n17261), .ZN(n17164) );
  XNOR2_X1 U20355 ( .A(n18081), .B(n17164), .ZN(n17160) );
  AOI21_X1 U20356 ( .B1(n17337), .B2(P3_EBX_REG_14__SCAN_IN), .A(n18481), .ZN(
        n17159) );
  INV_X1 U20357 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19152) );
  NAND3_X1 U20358 ( .A1(n17310), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n17166), 
        .ZN(n17154) );
  AOI21_X1 U20359 ( .B1(n19152), .B2(n17154), .A(n17153), .ZN(n17157) );
  AOI211_X1 U20360 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17167), .A(n17155), .B(
        n17325), .ZN(n17156) );
  AOI211_X1 U20361 ( .C1(n17267), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17157), .B(n17156), .ZN(n17158) );
  OAI211_X1 U20362 ( .C1(n19105), .C2(n17160), .A(n17159), .B(n17158), .ZN(
        P3_U2657) );
  INV_X1 U20363 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17176) );
  NAND2_X1 U20364 ( .A1(n18161), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18163) );
  NOR2_X1 U20365 ( .A1(n17329), .A2(n18163), .ZN(n17238) );
  NAND2_X1 U20366 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17238), .ZN(
        n17228) );
  NOR2_X1 U20367 ( .A1(n17161), .A2(n17228), .ZN(n18091) );
  NAND2_X1 U20368 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18091), .ZN(
        n17178) );
  AOI22_X1 U20369 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17162), .B1(
        n17176), .B2(n17178), .ZN(n18092) );
  NOR2_X1 U20370 ( .A1(n18092), .A2(n19105), .ZN(n17163) );
  AOI22_X1 U20371 ( .A1(n17337), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n17164), 
        .B2(n17163), .ZN(n17175) );
  AOI21_X1 U20372 ( .B1(n17310), .B2(n17186), .A(n17333), .ZN(n17190) );
  OAI21_X1 U20373 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17326), .A(n17190), 
        .ZN(n17173) );
  INV_X1 U20374 ( .A(n18092), .ZN(n17165) );
  AOI211_X1 U20375 ( .C1(n17292), .C2(n17178), .A(n17324), .B(n17165), .ZN(
        n17172) );
  NAND2_X1 U20376 ( .A1(n17310), .A2(n17166), .ZN(n17170) );
  OAI211_X1 U20377 ( .C1(n17177), .C2(n17168), .A(n17336), .B(n17167), .ZN(
        n17169) );
  OAI211_X1 U20378 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17170), .A(n18476), 
        .B(n17169), .ZN(n17171) );
  AOI211_X1 U20379 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17173), .A(n17172), 
        .B(n17171), .ZN(n17174) );
  OAI211_X1 U20380 ( .C1(n17176), .C2(n17322), .A(n17175), .B(n17174), .ZN(
        P3_U2658) );
  NAND2_X1 U20381 ( .A1(n17310), .A2(n19147), .ZN(n17185) );
  AOI21_X1 U20382 ( .B1(n17337), .B2(P3_EBX_REG_12__SCAN_IN), .A(n18481), .ZN(
        n17184) );
  AOI211_X1 U20383 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17193), .A(n17177), .B(
        n17325), .ZN(n17182) );
  OAI21_X1 U20384 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18091), .A(
        n17178), .ZN(n18114) );
  INV_X1 U20385 ( .A(n17278), .ZN(n17307) );
  OAI21_X1 U20386 ( .B1(n18100), .B2(n17307), .A(n17292), .ZN(n17179) );
  XNOR2_X1 U20387 ( .A(n18114), .B(n17179), .ZN(n17180) );
  OAI22_X1 U20388 ( .A1(n17190), .A2(n19147), .B1(n19105), .B2(n17180), .ZN(
        n17181) );
  AOI211_X1 U20389 ( .C1(n17267), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17182), .B(n17181), .ZN(n17183) );
  OAI211_X1 U20390 ( .C1(n17186), .C2(n17185), .A(n17184), .B(n17183), .ZN(
        P3_U2659) );
  INV_X1 U20391 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17197) );
  INV_X1 U20392 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19141) );
  NAND2_X1 U20393 ( .A1(n17310), .A2(n17200), .ZN(n17212) );
  NOR2_X1 U20394 ( .A1(n19141), .A2(n17212), .ZN(n17209) );
  AOI21_X1 U20395 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17209), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n17191) );
  INV_X1 U20396 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18127) );
  INV_X1 U20397 ( .A(n17228), .ZN(n17215) );
  NAND2_X1 U20398 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17215), .ZN(
        n17214) );
  NOR2_X1 U20399 ( .A1(n18127), .A2(n17214), .ZN(n17202) );
  AOI21_X1 U20400 ( .B1(n17202), .B2(n18257), .A(n17261), .ZN(n17188) );
  INV_X1 U20401 ( .A(n18091), .ZN(n17187) );
  OAI21_X1 U20402 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17202), .A(
        n17187), .ZN(n18131) );
  XOR2_X1 U20403 ( .A(n17188), .B(n18131), .Z(n17189) );
  OAI22_X1 U20404 ( .A1(n17191), .A2(n17190), .B1(n19105), .B2(n17189), .ZN(
        n17192) );
  AOI211_X1 U20405 ( .C1(n17337), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18481), .B(
        n17192), .ZN(n17196) );
  OAI211_X1 U20406 ( .C1(n17198), .C2(n17194), .A(n17336), .B(n17193), .ZN(
        n17195) );
  OAI211_X1 U20407 ( .C1(n17322), .C2(n17197), .A(n17196), .B(n17195), .ZN(
        P3_U2660) );
  AOI211_X1 U20408 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17219), .A(n17198), .B(
        n17325), .ZN(n17199) );
  AOI211_X1 U20409 ( .C1(n17337), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18481), .B(
        n17199), .ZN(n17211) );
  INV_X1 U20410 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19143) );
  INV_X1 U20411 ( .A(n17200), .ZN(n17201) );
  AOI21_X1 U20412 ( .B1(n17310), .B2(n17201), .A(n17333), .ZN(n17232) );
  OAI21_X1 U20413 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n17212), .A(n17232), .ZN(
        n17208) );
  AOI21_X1 U20414 ( .B1(n18127), .B2(n17214), .A(n17202), .ZN(n18145) );
  INV_X1 U20415 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17204) );
  INV_X1 U20416 ( .A(n17203), .ZN(n18162) );
  NAND3_X1 U20417 ( .A1(n18161), .A2(n18162), .A3(n17278), .ZN(n17218) );
  NOR2_X1 U20418 ( .A1(n17204), .A2(n17218), .ZN(n17216) );
  NOR2_X1 U20419 ( .A1(n17216), .A2(n17261), .ZN(n17206) );
  OAI21_X1 U20420 ( .B1(n18145), .B2(n17206), .A(n17239), .ZN(n17205) );
  AOI21_X1 U20421 ( .B1(n18145), .B2(n17206), .A(n17205), .ZN(n17207) );
  AOI221_X1 U20422 ( .B1(n17209), .B2(n19143), .C1(n17208), .C2(
        P3_REIP_REG_10__SCAN_IN), .A(n17207), .ZN(n17210) );
  OAI211_X1 U20423 ( .C1(n18127), .C2(n17322), .A(n17211), .B(n17210), .ZN(
        P3_U2661) );
  NOR2_X1 U20424 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17212), .ZN(n17213) );
  AOI211_X1 U20425 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17267), .A(
        n18481), .B(n17213), .ZN(n17225) );
  OAI21_X1 U20426 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17215), .A(
        n17214), .ZN(n18151) );
  NAND2_X1 U20427 ( .A1(n17292), .A2(n18151), .ZN(n17217) );
  AOI211_X1 U20428 ( .C1(n17218), .C2(n17217), .A(n17216), .B(n19105), .ZN(
        n17223) );
  OAI211_X1 U20429 ( .C1(n17226), .C2(n17220), .A(n17336), .B(n17219), .ZN(
        n17221) );
  OAI21_X1 U20430 ( .B1(n17320), .B2(n18151), .A(n17221), .ZN(n17222) );
  AOI211_X1 U20431 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17337), .A(n17223), .B(
        n17222), .ZN(n17224) );
  OAI211_X1 U20432 ( .C1(n17232), .C2(n19141), .A(n17225), .B(n17224), .ZN(
        P3_U2662) );
  INV_X1 U20433 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17236) );
  AOI211_X1 U20434 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17246), .A(n17226), .B(
        n17325), .ZN(n17234) );
  INV_X1 U20435 ( .A(n17242), .ZN(n17227) );
  NOR2_X1 U20436 ( .A1(n17326), .A2(n17237), .ZN(n17257) );
  AOI21_X1 U20437 ( .B1(n17227), .B2(n17257), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n17231) );
  AOI21_X1 U20438 ( .B1(n17238), .B2(n18257), .A(n17261), .ZN(n17229) );
  OAI21_X1 U20439 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17238), .A(
        n17228), .ZN(n18174) );
  XOR2_X1 U20440 ( .A(n17229), .B(n18174), .Z(n17230) );
  OAI22_X1 U20441 ( .A1(n17232), .A2(n17231), .B1(n19105), .B2(n17230), .ZN(
        n17233) );
  AOI211_X1 U20442 ( .C1(n17305), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17234), .B(n17233), .ZN(n17235) );
  OAI211_X1 U20443 ( .C1(n17275), .C2(n17236), .A(n17235), .B(n18476), .ZN(
        P3_U2663) );
  INV_X1 U20444 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18180) );
  NAND2_X1 U20445 ( .A1(n17310), .A2(n17237), .ZN(n17264) );
  NAND2_X1 U20446 ( .A1(n17282), .A2(n17264), .ZN(n17271) );
  NAND2_X1 U20447 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18161), .ZN(
        n17251) );
  AOI21_X1 U20448 ( .B1(n18180), .B2(n17251), .A(n17238), .ZN(n18184) );
  AOI21_X1 U20449 ( .B1(n18161), .B2(n17278), .A(n17261), .ZN(n17241) );
  OAI21_X1 U20450 ( .B1(n18184), .B2(n17241), .A(n17239), .ZN(n17240) );
  AOI21_X1 U20451 ( .B1(n18184), .B2(n17241), .A(n17240), .ZN(n17245) );
  OAI211_X1 U20452 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n17257), .B(n17242), .ZN(n17243) );
  OAI211_X1 U20453 ( .C1(n20911), .C2(n17275), .A(n18476), .B(n17243), .ZN(
        n17244) );
  AOI211_X1 U20454 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n17271), .A(n17245), .B(
        n17244), .ZN(n17248) );
  OAI211_X1 U20455 ( .C1(n17252), .C2(n20911), .A(n17336), .B(n17246), .ZN(
        n17247) );
  OAI211_X1 U20456 ( .C1(n17322), .C2(n18180), .A(n17248), .B(n17247), .ZN(
        P3_U2664) );
  NOR2_X1 U20457 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19105), .ZN(
        n17250) );
  INV_X1 U20458 ( .A(n17320), .ZN(n17249) );
  AOI21_X1 U20459 ( .B1(n17250), .B2(n18193), .A(n17249), .ZN(n17260) );
  NOR2_X1 U20460 ( .A1(n17329), .A2(n18192), .ZN(n17262) );
  OAI21_X1 U20461 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17262), .A(
        n17251), .ZN(n18197) );
  AOI211_X1 U20462 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17272), .A(n17252), .B(
        n17325), .ZN(n17255) );
  INV_X1 U20463 ( .A(n18197), .ZN(n17253) );
  AOI211_X1 U20464 ( .C1(n18161), .C2(n17278), .A(n17253), .B(n17323), .ZN(
        n17254) );
  AOI211_X1 U20465 ( .C1(n17305), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17255), .B(n17254), .ZN(n17259) );
  INV_X1 U20466 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19135) );
  OAI21_X1 U20467 ( .B1(n17275), .B2(n17602), .A(n18476), .ZN(n17256) );
  AOI221_X1 U20468 ( .B1(n17257), .B2(n19135), .C1(n17271), .C2(
        P3_REIP_REG_6__SCAN_IN), .A(n17256), .ZN(n17258) );
  OAI211_X1 U20469 ( .C1(n17260), .C2(n18197), .A(n17259), .B(n17258), .ZN(
        P3_U2665) );
  AND2_X1 U20470 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18203), .ZN(
        n17276) );
  AOI21_X1 U20471 ( .B1(n17276), .B2(n18257), .A(n17261), .ZN(n17277) );
  INV_X1 U20472 ( .A(n17262), .ZN(n17263) );
  OAI21_X1 U20473 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17276), .A(
        n17263), .ZN(n18206) );
  XOR2_X1 U20474 ( .A(n17277), .B(n18206), .Z(n17269) );
  INV_X1 U20475 ( .A(n17264), .ZN(n17265) );
  AOI22_X1 U20476 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17267), .B1(
        n17266), .B2(n17265), .ZN(n17268) );
  OAI211_X1 U20477 ( .C1(n19105), .C2(n17269), .A(n17268), .B(n18476), .ZN(
        n17270) );
  AOI21_X1 U20478 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n17271), .A(n17270), .ZN(
        n17274) );
  OAI211_X1 U20479 ( .C1(n17283), .C2(n17595), .A(n17336), .B(n17272), .ZN(
        n17273) );
  OAI211_X1 U20480 ( .C1(n17595), .C2(n17275), .A(n17274), .B(n17273), .ZN(
        P3_U2666) );
  NOR2_X1 U20481 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18209), .ZN(
        n18214) );
  OR2_X1 U20482 ( .A1(n17329), .A2(n18209), .ZN(n17290) );
  AOI21_X1 U20483 ( .B1(n18221), .B2(n17290), .A(n17276), .ZN(n18218) );
  INV_X1 U20484 ( .A(n18218), .ZN(n17284) );
  AOI22_X1 U20485 ( .A1(n17278), .A2(n18214), .B1(n17277), .B2(n17284), .ZN(
        n17289) );
  NOR3_X1 U20486 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17326), .A3(n17281), .ZN(
        n17280) );
  NAND2_X1 U20487 ( .A1(n18609), .A2(n19264), .ZN(n17340) );
  OAI221_X1 U20488 ( .B1(n17340), .B2(n21004), .C1(n17340), .C2(n9714), .A(
        n18476), .ZN(n17279) );
  AOI211_X1 U20489 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17337), .A(n17280), .B(
        n17279), .ZN(n17288) );
  NAND2_X1 U20490 ( .A1(n17310), .A2(n17281), .ZN(n17296) );
  NAND2_X1 U20491 ( .A1(n17282), .A2(n17296), .ZN(n17298) );
  AOI211_X1 U20492 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17299), .A(n17283), .B(
        n17325), .ZN(n17286) );
  OAI22_X1 U20493 ( .A1(n18221), .A2(n17322), .B1(n17320), .B2(n17284), .ZN(
        n17285) );
  AOI211_X1 U20494 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n17298), .A(n17286), .B(
        n17285), .ZN(n17287) );
  OAI211_X1 U20495 ( .C1(n17289), .C2(n19105), .A(n17288), .B(n17287), .ZN(
        P3_U2667) );
  INV_X1 U20496 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17303) );
  NAND2_X1 U20497 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17309) );
  INV_X1 U20498 ( .A(n17340), .ZN(n19266) );
  NAND2_X1 U20499 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19060), .ZN(
        n19057) );
  AOI21_X1 U20500 ( .B1(n19207), .B2(n19057), .A(n17572), .ZN(n19203) );
  AOI22_X1 U20501 ( .A1(n17337), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n19266), .B2(
        n19203), .ZN(n17295) );
  INV_X1 U20502 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18243) );
  NOR2_X1 U20503 ( .A1(n17329), .A2(n18243), .ZN(n17291) );
  OAI21_X1 U20504 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17291), .A(
        n17290), .ZN(n18227) );
  INV_X1 U20505 ( .A(n17291), .ZN(n17304) );
  OAI21_X1 U20506 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17304), .A(
        n17292), .ZN(n17306) );
  AOI21_X1 U20507 ( .B1(n18227), .B2(n17306), .A(n19105), .ZN(n17293) );
  OAI21_X1 U20508 ( .B1(n18227), .B2(n17306), .A(n17293), .ZN(n17294) );
  OAI211_X1 U20509 ( .C1(n17296), .C2(n17309), .A(n17295), .B(n17294), .ZN(
        n17297) );
  AOI21_X1 U20510 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n17298), .A(n17297), .ZN(
        n17302) );
  OAI211_X1 U20511 ( .C1(n17311), .C2(n17300), .A(n17336), .B(n17299), .ZN(
        n17301) );
  OAI211_X1 U20512 ( .C1(n17322), .C2(n17303), .A(n17302), .B(n17301), .ZN(
        P3_U2668) );
  OAI21_X1 U20513 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17304), .ZN(n18239) );
  AOI22_X1 U20514 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17305), .B1(
        n17337), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n17319) );
  INV_X1 U20515 ( .A(n18239), .ZN(n17308) );
  AOI211_X1 U20516 ( .C1(n17308), .C2(n17307), .A(n19105), .B(n17306), .ZN(
        n17317) );
  NAND2_X1 U20517 ( .A1(n19219), .A2(n19061), .ZN(n19048) );
  NAND2_X1 U20518 ( .A1(n19048), .A2(n19057), .ZN(n19213) );
  OAI211_X1 U20519 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17310), .B(n17309), .ZN(n17315) );
  NOR2_X1 U20520 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17313) );
  INV_X1 U20521 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17610) );
  INV_X1 U20522 ( .A(n17311), .ZN(n17312) );
  OAI211_X1 U20523 ( .C1(n17313), .C2(n17610), .A(n17336), .B(n17312), .ZN(
        n17314) );
  OAI211_X1 U20524 ( .C1(n17340), .C2(n19213), .A(n17315), .B(n17314), .ZN(
        n17316) );
  AOI211_X1 U20525 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n17333), .A(n17317), .B(
        n17316), .ZN(n17318) );
  OAI211_X1 U20526 ( .C1(n17320), .C2(n18239), .A(n17319), .B(n17318), .ZN(
        P3_U2669) );
  NAND2_X1 U20527 ( .A1(n19061), .A2(n17321), .ZN(n19220) );
  AOI22_X1 U20528 ( .A1(n17337), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n17333), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17332) );
  OAI21_X1 U20529 ( .B1(n18257), .B2(n17323), .A(n17322), .ZN(n17330) );
  INV_X1 U20530 ( .A(n17324), .ZN(n17328) );
  NAND2_X1 U20531 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17614) );
  OAI21_X1 U20532 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17614), .ZN(n17623) );
  OAI22_X1 U20533 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17326), .B1(n17325), 
        .B2(n17623), .ZN(n17327) );
  AOI221_X1 U20534 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17330), .C1(
        n17329), .C2(n17328), .A(n17327), .ZN(n17331) );
  OAI211_X1 U20535 ( .C1(n19220), .C2(n17340), .A(n17332), .B(n17331), .ZN(
        P3_U2670) );
  NOR3_X1 U20536 ( .A1(n19262), .A2(n17333), .A3(n18257), .ZN(n17334) );
  AOI21_X1 U20537 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n17335), .A(n17334), .ZN(
        n17339) );
  OAI21_X1 U20538 ( .B1(n17337), .B2(n17336), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17338) );
  OAI211_X1 U20539 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17340), .A(
        n17339), .B(n17338), .ZN(P3_U2671) );
  NAND4_X1 U20540 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(n17341), .ZN(n17381) );
  NAND3_X1 U20541 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17342), .ZN(n17414) );
  NOR4_X1 U20542 ( .A1(n17374), .A2(n17343), .A3(n17381), .A4(n17414), .ZN(
        n17344) );
  NAND3_X1 U20543 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17344), .ZN(n17347) );
  NAND2_X1 U20544 ( .A1(n17619), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17346) );
  NAND2_X1 U20545 ( .A1(n17373), .A2(n18639), .ZN(n17345) );
  OAI22_X1 U20546 ( .A1(n17373), .A2(n17346), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17345), .ZN(P3_U2672) );
  NAND2_X1 U20547 ( .A1(n17348), .A2(n17347), .ZN(n17349) );
  NAND2_X1 U20548 ( .A1(n17349), .A2(n17619), .ZN(n17372) );
  AOI22_X1 U20549 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20550 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17574), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20551 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U20552 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17350) );
  NAND4_X1 U20553 ( .A1(n17353), .A2(n17352), .A3(n17351), .A4(n17350), .ZN(
        n17359) );
  AOI22_X1 U20554 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20555 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U20556 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U20557 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17354) );
  NAND4_X1 U20558 ( .A1(n17357), .A2(n17356), .A3(n17355), .A4(n17354), .ZN(
        n17358) );
  NOR2_X1 U20559 ( .A1(n17359), .A2(n17358), .ZN(n17371) );
  AOI22_X1 U20560 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U20561 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n17572), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U20562 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U20563 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17360) );
  NAND4_X1 U20564 ( .A1(n17363), .A2(n17362), .A3(n17361), .A4(n17360), .ZN(
        n17369) );
  AOI22_X1 U20565 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20566 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U20567 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20568 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17364) );
  NAND4_X1 U20569 ( .A1(n17367), .A2(n17366), .A3(n17365), .A4(n17364), .ZN(
        n17368) );
  NOR2_X1 U20570 ( .A1(n17369), .A2(n17368), .ZN(n17376) );
  NOR3_X1 U20571 ( .A1(n17376), .A2(n17648), .A3(n17375), .ZN(n17370) );
  XOR2_X1 U20572 ( .A(n17371), .B(n17370), .Z(n17638) );
  OAI22_X1 U20573 ( .A1(n17373), .A2(n17372), .B1(n17638), .B2(n17619), .ZN(
        P3_U2673) );
  NAND2_X1 U20574 ( .A1(n17400), .A2(n17374), .ZN(n17380) );
  NOR2_X1 U20575 ( .A1(n17648), .A2(n17375), .ZN(n17377) );
  XNOR2_X1 U20576 ( .A(n17377), .B(n17376), .ZN(n17639) );
  AOI22_X1 U20577 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17378), .B1(n17625), 
        .B2(n17639), .ZN(n17379) );
  OAI21_X1 U20578 ( .B1(n17381), .B2(n17380), .A(n17379), .ZN(P3_U2674) );
  OAI211_X1 U20579 ( .C1(n17650), .C2(n17649), .A(n17625), .B(n17648), .ZN(
        n17382) );
  OAI221_X1 U20580 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17385), .C1(n17384), 
        .C2(n17383), .A(n17382), .ZN(P3_U2676) );
  AOI21_X1 U20581 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17619), .A(n9751), .ZN(
        n17387) );
  XNOR2_X1 U20582 ( .A(n17386), .B(n17389), .ZN(n17659) );
  OAI22_X1 U20583 ( .A1(n17388), .A2(n17387), .B1(n17619), .B2(n17659), .ZN(
        P3_U2677) );
  AOI21_X1 U20584 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17619), .A(n9752), .ZN(
        n17392) );
  OAI21_X1 U20585 ( .B1(n17391), .B2(n17390), .A(n17389), .ZN(n17664) );
  OAI22_X1 U20586 ( .A1(n9751), .A2(n17392), .B1(n17619), .B2(n17664), .ZN(
        P3_U2678) );
  AOI21_X1 U20587 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17619), .A(n17400), .ZN(
        n17394) );
  XNOR2_X1 U20588 ( .A(n17393), .B(n17396), .ZN(n17669) );
  OAI22_X1 U20589 ( .A1(n9752), .A2(n17394), .B1(n17619), .B2(n17669), .ZN(
        P3_U2679) );
  INV_X1 U20590 ( .A(n17395), .ZN(n17413) );
  AOI21_X1 U20591 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17619), .A(n17413), .ZN(
        n17399) );
  OAI21_X1 U20592 ( .B1(n17398), .B2(n17397), .A(n17396), .ZN(n17674) );
  OAI22_X1 U20593 ( .A1(n17400), .A2(n17399), .B1(n17619), .B2(n17674), .ZN(
        P3_U2680) );
  AOI22_X1 U20594 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17619), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n17426), .ZN(n17412) );
  AOI22_X1 U20595 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20596 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17403) );
  AOI22_X1 U20597 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20598 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n17562), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17401) );
  NAND4_X1 U20599 ( .A1(n17404), .A2(n17403), .A3(n17402), .A4(n17401), .ZN(
        n17411) );
  AOI22_X1 U20600 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17409) );
  AOI22_X1 U20601 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20602 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17405), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U20603 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17406) );
  NAND4_X1 U20604 ( .A1(n17409), .A2(n17408), .A3(n17407), .A4(n17406), .ZN(
        n17410) );
  NOR2_X1 U20605 ( .A1(n17411), .A2(n17410), .ZN(n17676) );
  OAI22_X1 U20606 ( .A1(n17413), .A2(n17412), .B1(n17676), .B2(n17619), .ZN(
        P3_U2681) );
  NAND2_X1 U20607 ( .A1(n17619), .A2(n17414), .ZN(n17439) );
  AOI22_X1 U20608 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17425) );
  AOI22_X1 U20609 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17424) );
  INV_X1 U20610 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17416) );
  AOI22_X1 U20611 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17415) );
  OAI21_X1 U20612 ( .B1(n17416), .B2(n13957), .A(n17415), .ZN(n17422) );
  AOI22_X1 U20613 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20614 ( .A1(n9676), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17419) );
  AOI22_X1 U20615 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20616 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17417) );
  NAND4_X1 U20617 ( .A1(n17420), .A2(n17419), .A3(n17418), .A4(n17417), .ZN(
        n17421) );
  AOI211_X1 U20618 ( .C1(n17539), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n17422), .B(n17421), .ZN(n17423) );
  NAND3_X1 U20619 ( .A1(n17425), .A2(n17424), .A3(n17423), .ZN(n17681) );
  AOI22_X1 U20620 ( .A1(n17625), .A2(n17681), .B1(n17426), .B2(n17428), .ZN(
        n17427) );
  OAI21_X1 U20621 ( .B1(n17428), .B2(n17439), .A(n17427), .ZN(P3_U2682) );
  AOI21_X1 U20622 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17453), .A(
        P3_EBX_REG_20__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20623 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20624 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20625 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20626 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17429) );
  NAND4_X1 U20627 ( .A1(n17432), .A2(n17431), .A3(n17430), .A4(n17429), .ZN(
        n17438) );
  AOI22_X1 U20628 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20629 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n17561), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20630 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U20631 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17433) );
  NAND4_X1 U20632 ( .A1(n17436), .A2(n17435), .A3(n17434), .A4(n17433), .ZN(
        n17437) );
  NOR2_X1 U20633 ( .A1(n17438), .A2(n17437), .ZN(n17687) );
  OAI22_X1 U20634 ( .A1(n17440), .A2(n17439), .B1(n17687), .B2(n17619), .ZN(
        P3_U2683) );
  AOI22_X1 U20635 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U20636 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13914), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20637 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20638 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n17572), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17442) );
  NAND4_X1 U20639 ( .A1(n17445), .A2(n17444), .A3(n17443), .A4(n17442), .ZN(
        n17451) );
  AOI22_X1 U20640 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U20641 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13964), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20642 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U20643 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17446) );
  NAND4_X1 U20644 ( .A1(n17449), .A2(n17448), .A3(n17447), .A4(n17446), .ZN(
        n17450) );
  NOR2_X1 U20645 ( .A1(n17451), .A2(n17450), .ZN(n17694) );
  AOI22_X1 U20646 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17454), .B1(n17453), 
        .B2(n17452), .ZN(n17455) );
  OAI21_X1 U20647 ( .B1(n17694), .B2(n17619), .A(n17455), .ZN(P3_U2684) );
  NAND2_X1 U20648 ( .A1(n17619), .A2(n17456), .ZN(n17482) );
  AOI22_X1 U20649 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17555), .ZN(n17467) );
  AOI22_X1 U20650 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17466) );
  INV_X1 U20651 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U20652 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17554), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U20653 ( .B1(n17620), .B2(n17458), .A(n17457), .ZN(n17464) );
  AOI22_X1 U20654 ( .A1(n9676), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17580), .ZN(n17462) );
  AOI22_X1 U20655 ( .A1(n17405), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U20656 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9667), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20657 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17575), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17459) );
  NAND4_X1 U20658 ( .A1(n17462), .A2(n17461), .A3(n17460), .A4(n17459), .ZN(
        n17463) );
  AOI211_X1 U20659 ( .C1(n9679), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n17464), .B(n17463), .ZN(n17465) );
  NAND3_X1 U20660 ( .A1(n17467), .A2(n17466), .A3(n17465), .ZN(n17702) );
  NAND2_X1 U20661 ( .A1(n17625), .A2(n17702), .ZN(n17468) );
  OAI221_X1 U20662 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17470), .C1(n17469), 
        .C2(n17482), .A(n17468), .ZN(P3_U2686) );
  AOI22_X1 U20663 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17475) );
  AOI22_X1 U20664 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17474) );
  AOI22_X1 U20665 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13964), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U20666 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17472) );
  NAND4_X1 U20667 ( .A1(n17475), .A2(n17474), .A3(n17473), .A4(n17472), .ZN(
        n17481) );
  AOI22_X1 U20668 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U20669 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20670 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U20671 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17476) );
  NAND4_X1 U20672 ( .A1(n17479), .A2(n17478), .A3(n17477), .A4(n17476), .ZN(
        n17480) );
  NOR2_X1 U20673 ( .A1(n17481), .A2(n17480), .ZN(n17714) );
  NOR2_X1 U20674 ( .A1(n9749), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17483) );
  OAI22_X1 U20675 ( .A1(n17714), .A2(n17619), .B1(n17483), .B2(n17482), .ZN(
        P3_U2687) );
  INV_X1 U20676 ( .A(n17508), .ZN(n17484) );
  OAI21_X1 U20677 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17484), .A(n17619), .ZN(
        n17496) );
  AOI22_X1 U20678 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U20679 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17572), .B1(
        n9679), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U20680 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U20681 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17485) );
  NAND4_X1 U20682 ( .A1(n17488), .A2(n17487), .A3(n17486), .A4(n17485), .ZN(
        n17495) );
  AOI22_X1 U20683 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U20684 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20685 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17573), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17491) );
  AOI22_X1 U20686 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17490) );
  NAND4_X1 U20687 ( .A1(n17493), .A2(n17492), .A3(n17491), .A4(n17490), .ZN(
        n17494) );
  NOR2_X1 U20688 ( .A1(n17495), .A2(n17494), .ZN(n17721) );
  OAI22_X1 U20689 ( .A1(n9749), .A2(n17496), .B1(n17721), .B2(n17619), .ZN(
        P3_U2688) );
  AOI22_X1 U20690 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U20691 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U20692 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U20693 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17497) );
  NAND4_X1 U20694 ( .A1(n17500), .A2(n17499), .A3(n17498), .A4(n17497), .ZN(
        n17507) );
  AOI22_X1 U20695 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17505) );
  AOI22_X1 U20696 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n9667), .B1(n9666), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17504) );
  AOI22_X1 U20697 ( .A1(n9676), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20698 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17554), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17502) );
  NAND4_X1 U20699 ( .A1(n17505), .A2(n17504), .A3(n17503), .A4(n17502), .ZN(
        n17506) );
  NOR2_X1 U20700 ( .A1(n17507), .A2(n17506), .ZN(n17726) );
  OAI21_X1 U20701 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17509), .A(n17508), .ZN(
        n17510) );
  AOI22_X1 U20702 ( .A1(n17625), .A2(n17726), .B1(n17510), .B2(n17619), .ZN(
        P3_U2689) );
  AOI22_X1 U20703 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U20704 ( .A1(n17584), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20705 ( .A1(n17405), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U20706 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17511) );
  NAND4_X1 U20707 ( .A1(n17514), .A2(n17513), .A3(n17512), .A4(n17511), .ZN(
        n17520) );
  AOI22_X1 U20708 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U20709 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17517) );
  AOI22_X1 U20710 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n17554), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17516) );
  AOI22_X1 U20711 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17515) );
  NAND4_X1 U20712 ( .A1(n17518), .A2(n17517), .A3(n17516), .A4(n17515), .ZN(
        n17519) );
  NOR2_X1 U20713 ( .A1(n17520), .A2(n17519), .ZN(n17731) );
  OAI211_X1 U20714 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17536), .A(n17521), .B(
        n17619), .ZN(n17522) );
  OAI21_X1 U20715 ( .B1(n17731), .B2(n17619), .A(n17522), .ZN(P3_U2691) );
  INV_X1 U20716 ( .A(n17550), .ZN(n17523) );
  OAI21_X1 U20717 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17523), .A(n17619), .ZN(
        n17535) );
  AOI22_X1 U20718 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17528) );
  AOI22_X1 U20719 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n17562), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17527) );
  AOI22_X1 U20720 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U20721 ( .A1(n17524), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17525) );
  NAND4_X1 U20722 ( .A1(n17528), .A2(n17527), .A3(n17526), .A4(n17525), .ZN(
        n17534) );
  AOI22_X1 U20723 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17532) );
  AOI22_X1 U20724 ( .A1(n17556), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20725 ( .A1(n9669), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17530) );
  AOI22_X1 U20726 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17529) );
  NAND4_X1 U20727 ( .A1(n17532), .A2(n17531), .A3(n17530), .A4(n17529), .ZN(
        n17533) );
  NOR2_X1 U20728 ( .A1(n17534), .A2(n17533), .ZN(n17735) );
  OAI22_X1 U20729 ( .A1(n17536), .A2(n17535), .B1(n17735), .B2(n17619), .ZN(
        P3_U2692) );
  AOI22_X1 U20730 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17549) );
  AOI22_X1 U20731 ( .A1(n17582), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16041), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17548) );
  AOI22_X1 U20732 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17554), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17537) );
  OAI21_X1 U20733 ( .B1(n17538), .B2(n17618), .A(n17537), .ZN(n17546) );
  AOI22_X1 U20734 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17544) );
  AOI22_X1 U20735 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U20736 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U20737 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17555), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17541) );
  NAND4_X1 U20738 ( .A1(n17544), .A2(n17543), .A3(n17542), .A4(n17541), .ZN(
        n17545) );
  AOI211_X1 U20739 ( .C1(n17562), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17546), .B(n17545), .ZN(n17547) );
  NAND3_X1 U20740 ( .A1(n17549), .A2(n17548), .A3(n17547), .ZN(n17739) );
  INV_X1 U20741 ( .A(n17739), .ZN(n17552) );
  OAI21_X1 U20742 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17570), .A(n17550), .ZN(
        n17551) );
  AOI22_X1 U20743 ( .A1(n17625), .A2(n17552), .B1(n17551), .B2(n17619), .ZN(
        P3_U2693) );
  INV_X1 U20744 ( .A(n17591), .ZN(n17553) );
  OAI21_X1 U20745 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17553), .A(n17619), .ZN(
        n17569) );
  AOI22_X1 U20746 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17571), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17554), .ZN(n17560) );
  AOI22_X1 U20747 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17575), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17555), .ZN(n17559) );
  AOI22_X1 U20748 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17556), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17558) );
  AOI22_X1 U20749 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9667), .ZN(n17557) );
  NAND4_X1 U20750 ( .A1(n17560), .A2(n17559), .A3(n17558), .A4(n17557), .ZN(
        n17568) );
  AOI22_X1 U20751 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17574), .B1(
        n17581), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17566) );
  AOI22_X1 U20752 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9666), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17565) );
  AOI22_X1 U20753 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17564) );
  AOI22_X1 U20754 ( .A1(n17562), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17580), .ZN(n17563) );
  NAND4_X1 U20755 ( .A1(n17566), .A2(n17565), .A3(n17564), .A4(n17563), .ZN(
        n17567) );
  NOR2_X1 U20756 ( .A1(n17568), .A2(n17567), .ZN(n17743) );
  OAI22_X1 U20757 ( .A1(n17570), .A2(n17569), .B1(n17743), .B2(n17619), .ZN(
        P3_U2694) );
  AOI22_X1 U20758 ( .A1(n17572), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17571), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17579) );
  AOI22_X1 U20759 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16009), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17578) );
  AOI22_X1 U20760 ( .A1(n9679), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17577) );
  AOI22_X1 U20761 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17576) );
  NAND4_X1 U20762 ( .A1(n17579), .A2(n17578), .A3(n17577), .A4(n17576), .ZN(
        n17590) );
  AOI22_X1 U20763 ( .A1(n17581), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U20764 ( .A1(n13949), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17582), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17587) );
  AOI22_X1 U20765 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17583), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17586) );
  AOI22_X1 U20766 ( .A1(n17584), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13964), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17585) );
  NAND4_X1 U20767 ( .A1(n17588), .A2(n17587), .A3(n17586), .A4(n17585), .ZN(
        n17589) );
  NOR2_X1 U20768 ( .A1(n17590), .A2(n17589), .ZN(n17750) );
  OAI21_X1 U20769 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17593), .A(n17591), .ZN(
        n17592) );
  AOI22_X1 U20770 ( .A1(n17625), .A2(n17750), .B1(n17592), .B2(n17619), .ZN(
        P3_U2695) );
  OR2_X1 U20771 ( .A1(n20911), .A2(n17593), .ZN(n17598) );
  INV_X1 U20772 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17597) );
  NOR2_X1 U20773 ( .A1(n17594), .A2(n17627), .ZN(n17613) );
  NAND2_X1 U20774 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17613), .ZN(n17607) );
  NOR2_X1 U20775 ( .A1(n17595), .A2(n17607), .ZN(n17600) );
  NAND3_X1 U20776 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17600), .A3(n20911), .ZN(
        n17596) );
  OAI221_X1 U20777 ( .B1(n17625), .B2(n17598), .C1(n17619), .C2(n17597), .A(
        n17596), .ZN(P3_U2696) );
  NAND2_X1 U20778 ( .A1(n17619), .A2(n17599), .ZN(n17605) );
  AOI22_X1 U20779 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17625), .B1(
        n17600), .B2(n17602), .ZN(n17601) );
  OAI21_X1 U20780 ( .B1(n17602), .B2(n17605), .A(n17601), .ZN(P3_U2697) );
  NOR2_X1 U20781 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17603), .ZN(n17606) );
  INV_X1 U20782 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17604) );
  OAI22_X1 U20783 ( .A1(n17606), .A2(n17605), .B1(n17604), .B2(n17619), .ZN(
        P3_U2698) );
  INV_X1 U20784 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17609) );
  OAI211_X1 U20785 ( .C1(n17613), .C2(P3_EBX_REG_4__SCAN_IN), .A(n17619), .B(
        n17607), .ZN(n17608) );
  OAI21_X1 U20786 ( .B1(n17619), .B2(n17609), .A(n17608), .ZN(P3_U2699) );
  NOR3_X1 U20787 ( .A1(n17610), .A2(n17614), .A3(n17627), .ZN(n17616) );
  AOI21_X1 U20788 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17619), .A(n17616), .ZN(
        n17612) );
  INV_X1 U20789 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17611) );
  OAI22_X1 U20790 ( .A1(n17613), .A2(n17612), .B1(n17611), .B2(n17619), .ZN(
        P3_U2700) );
  INV_X1 U20791 ( .A(n17614), .ZN(n17615) );
  AOI221_X1 U20792 ( .B1(n17615), .B2(n17621), .C1(n17717), .C2(n17621), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17617) );
  AOI211_X1 U20793 ( .C1(n17625), .C2(n17618), .A(n17617), .B(n17616), .ZN(
        P3_U2701) );
  INV_X1 U20794 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17622) );
  OAI222_X1 U20795 ( .A1(n17623), .A2(n17627), .B1(n17622), .B2(n17621), .C1(
        n17620), .C2(n17619), .ZN(P3_U2702) );
  AOI22_X1 U20796 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17625), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17624), .ZN(n17626) );
  OAI21_X1 U20797 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17627), .A(n17626), .ZN(
        P3_U2703) );
  INV_X1 U20798 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17852) );
  INV_X1 U20799 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17848) );
  INV_X1 U20800 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20871) );
  INV_X1 U20801 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17894) );
  NAND2_X1 U20802 ( .A1(n17631), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17779) );
  NAND3_X1 U20803 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17629) );
  NAND4_X1 U20804 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17628) );
  INV_X1 U20805 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17889) );
  INV_X1 U20806 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17877) );
  INV_X1 U20807 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17875) );
  NAND4_X1 U20808 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17722)
         );
  NOR4_X1 U20809 ( .A1(n17889), .A2(n17877), .A3(n17875), .A4(n17722), .ZN(
        n17718) );
  NAND2_X1 U20810 ( .A1(n17716), .A2(n17718), .ZN(n17723) );
  INV_X1 U20811 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17840) );
  NAND4_X1 U20812 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17630)
         );
  NAND2_X1 U20813 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17671), .ZN(n17670) );
  NAND2_X1 U20814 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17666), .ZN(n17665) );
  NAND2_X1 U20815 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17655), .ZN(n17651) );
  NAND2_X1 U20816 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17644), .ZN(n17640) );
  NAND2_X1 U20817 ( .A1(n17635), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17634) );
  NAND2_X2 U20818 ( .A1(n17631), .A2(n17717), .ZN(n17769) );
  NOR2_X2 U20819 ( .A1(n18633), .A2(n17769), .ZN(n17708) );
  OAI22_X1 U20820 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17778), .B1(n17696), 
        .B2(n17635), .ZN(n17632) );
  AOI22_X1 U20821 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17708), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17632), .ZN(n17633) );
  OAI21_X1 U20822 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17634), .A(n17633), .ZN(
        P3_U2704) );
  NAND2_X1 U20823 ( .A1(n18629), .A2(n17696), .ZN(n17707) );
  AOI22_X1 U20824 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17708), .ZN(n17637) );
  OAI211_X1 U20825 ( .C1(n17635), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17769), .B(
        n17634), .ZN(n17636) );
  OAI211_X1 U20826 ( .C1(n17638), .C2(n17771), .A(n17637), .B(n17636), .ZN(
        P3_U2705) );
  AOI22_X1 U20827 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17708), .B1(n17639), .B2(
        n17776), .ZN(n17642) );
  OAI211_X1 U20828 ( .C1(n17644), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17769), .B(
        n17640), .ZN(n17641) );
  OAI211_X1 U20829 ( .C1(n17707), .C2(n17730), .A(n17642), .B(n17641), .ZN(
        P3_U2706) );
  INV_X1 U20830 ( .A(n17708), .ZN(n17701) );
  AOI22_X1 U20831 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17709), .B1(n17643), .B2(
        n17776), .ZN(n17647) );
  AOI211_X1 U20832 ( .C1(n17852), .C2(n17651), .A(n17644), .B(n17696), .ZN(
        n17645) );
  INV_X1 U20833 ( .A(n17645), .ZN(n17646) );
  OAI211_X1 U20834 ( .C1(n17701), .C2(n19573), .A(n17647), .B(n17646), .ZN(
        P3_U2707) );
  OAI21_X1 U20835 ( .B1(n17650), .B2(n17649), .A(n17648), .ZN(n17654) );
  AOI22_X1 U20836 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17708), .ZN(n17653) );
  OAI211_X1 U20837 ( .C1(n17655), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17769), .B(
        n17651), .ZN(n17652) );
  OAI211_X1 U20838 ( .C1(n17771), .C2(n17654), .A(n17653), .B(n17652), .ZN(
        P3_U2708) );
  AOI22_X1 U20839 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17708), .ZN(n17658) );
  AOI211_X1 U20840 ( .C1(n17848), .C2(n17660), .A(n17655), .B(n17696), .ZN(
        n17656) );
  INV_X1 U20841 ( .A(n17656), .ZN(n17657) );
  OAI211_X1 U20842 ( .C1(n17771), .C2(n17659), .A(n17658), .B(n17657), .ZN(
        P3_U2709) );
  AOI22_X1 U20843 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17708), .ZN(n17663) );
  OAI211_X1 U20844 ( .C1(n17661), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17769), .B(
        n17660), .ZN(n17662) );
  OAI211_X1 U20845 ( .C1(n17664), .C2(n17771), .A(n17663), .B(n17662), .ZN(
        P3_U2710) );
  AOI22_X1 U20846 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17708), .ZN(n17668) );
  OAI211_X1 U20847 ( .C1(n17666), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17769), .B(
        n17665), .ZN(n17667) );
  OAI211_X1 U20848 ( .C1(n17669), .C2(n17771), .A(n17668), .B(n17667), .ZN(
        P3_U2711) );
  AOI22_X1 U20849 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17708), .ZN(n17673) );
  OAI211_X1 U20850 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17671), .A(n17769), .B(
        n17670), .ZN(n17672) );
  OAI211_X1 U20851 ( .C1(n17674), .C2(n17771), .A(n17673), .B(n17672), .ZN(
        P3_U2712) );
  INV_X1 U20852 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17833) );
  NOR2_X1 U20853 ( .A1(n17717), .A2(n17710), .ZN(n17704) );
  NAND2_X1 U20854 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17704), .ZN(n17703) );
  NAND3_X1 U20855 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n17697), .ZN(n17682) );
  NOR2_X1 U20856 ( .A1(n20871), .A2(n17682), .ZN(n17679) );
  NAND2_X1 U20857 ( .A1(n17769), .A2(n17682), .ZN(n17690) );
  OAI21_X1 U20858 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17778), .A(n17690), .ZN(
        n17678) );
  OAI22_X1 U20859 ( .A1(n17676), .A2(n17771), .B1(n17675), .B2(n17701), .ZN(
        n17677) );
  AOI221_X1 U20860 ( .B1(n17679), .B2(n17840), .C1(n17678), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17677), .ZN(n17680) );
  OAI21_X1 U20861 ( .B1(n18632), .B2(n17707), .A(n17680), .ZN(P3_U2713) );
  AOI22_X1 U20862 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17708), .B1(n17776), .B2(
        n17681), .ZN(n17685) );
  OAI22_X1 U20863 ( .A1(n17707), .A2(n18628), .B1(n17682), .B2(
        P3_EAX_REG_21__SCAN_IN), .ZN(n17683) );
  INV_X1 U20864 ( .A(n17683), .ZN(n17684) );
  OAI211_X1 U20865 ( .C1(n20871), .C2(n17690), .A(n17685), .B(n17684), .ZN(
        P3_U2714) );
  NAND2_X1 U20866 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17697), .ZN(n17691) );
  INV_X1 U20867 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17837) );
  OAI22_X1 U20868 ( .A1(n17687), .A2(n17771), .B1(n17686), .B2(n17701), .ZN(
        n17688) );
  AOI21_X1 U20869 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n17709), .A(n17688), .ZN(
        n17689) );
  OAI221_X1 U20870 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n17691), .C1(n17837), 
        .C2(n17690), .A(n17689), .ZN(P3_U2715) );
  AOI22_X1 U20871 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17708), .ZN(n17693) );
  OAI211_X1 U20872 ( .C1(n17697), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17769), .B(
        n17691), .ZN(n17692) );
  OAI211_X1 U20873 ( .C1(n17694), .C2(n17771), .A(n17693), .B(n17692), .ZN(
        P3_U2716) );
  AOI22_X1 U20874 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17709), .B1(n17776), .B2(
        n17695), .ZN(n17700) );
  AOI211_X1 U20875 ( .C1(n17833), .C2(n17703), .A(n17697), .B(n17696), .ZN(
        n17698) );
  INV_X1 U20876 ( .A(n17698), .ZN(n17699) );
  OAI211_X1 U20877 ( .C1(n17701), .C2(n19563), .A(n17700), .B(n17699), .ZN(
        P3_U2717) );
  AOI22_X1 U20878 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n17708), .B1(n17776), .B2(
        n17702), .ZN(n17706) );
  OAI211_X1 U20879 ( .C1(n17704), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17769), .B(
        n17703), .ZN(n17705) );
  OAI211_X1 U20880 ( .C1(n17707), .C2(n18612), .A(n17706), .B(n17705), .ZN(
        P3_U2718) );
  AOI22_X1 U20881 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17709), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17708), .ZN(n17713) );
  OAI211_X1 U20882 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17711), .A(n17769), .B(
        n17710), .ZN(n17712) );
  OAI211_X1 U20883 ( .C1(n17714), .C2(n17771), .A(n17713), .B(n17712), .ZN(
        P3_U2719) );
  AND2_X1 U20884 ( .A1(n17769), .A2(n17723), .ZN(n17715) );
  AOI22_X1 U20885 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17777), .B1(
        P3_EAX_REG_15__SCAN_IN), .B2(n17715), .ZN(n17720) );
  INV_X1 U20886 ( .A(n17716), .ZN(n17747) );
  NAND3_X1 U20887 ( .A1(n17718), .A2(n17753), .A3(n17894), .ZN(n17719) );
  OAI211_X1 U20888 ( .C1(n17721), .C2(n17771), .A(n17720), .B(n17719), .ZN(
        P3_U2720) );
  NAND3_X1 U20889 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17753), .ZN(n17740) );
  NOR2_X1 U20890 ( .A1(n17722), .A2(n17740), .ZN(n17729) );
  AOI22_X1 U20891 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17777), .B1(n17729), .B2(
        n17889), .ZN(n17725) );
  NAND3_X1 U20892 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17769), .A3(n17723), 
        .ZN(n17724) );
  OAI211_X1 U20893 ( .C1(n17726), .C2(n17771), .A(n17725), .B(n17724), .ZN(
        P3_U2721) );
  INV_X1 U20894 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17881) );
  INV_X1 U20895 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17879) );
  NOR3_X1 U20896 ( .A1(n17881), .A2(n17879), .A3(n17740), .ZN(n17737) );
  AND2_X1 U20897 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17737), .ZN(n17733) );
  AOI21_X1 U20898 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17769), .A(n17733), .ZN(
        n17728) );
  OAI222_X1 U20899 ( .A1(n17774), .A2(n17730), .B1(n17729), .B2(n17728), .C1(
        n17771), .C2(n17727), .ZN(P3_U2722) );
  AOI21_X1 U20900 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17769), .A(n17737), .ZN(
        n17732) );
  OAI222_X1 U20901 ( .A1(n17774), .A2(n17734), .B1(n17733), .B2(n17732), .C1(
        n17771), .C2(n17731), .ZN(P3_U2723) );
  INV_X1 U20902 ( .A(n17740), .ZN(n17745) );
  AOI22_X1 U20903 ( .A1(n17745), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n17769), .ZN(n17736) );
  OAI222_X1 U20904 ( .A1(n17774), .A2(n17738), .B1(n17737), .B2(n17736), .C1(
        n17771), .C2(n17735), .ZN(P3_U2724) );
  AOI22_X1 U20905 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17777), .B1(n17776), .B2(
        n17739), .ZN(n17742) );
  OAI221_X1 U20906 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17745), .C1(n17879), 
        .C2(n17740), .A(n17769), .ZN(n17741) );
  NAND2_X1 U20907 ( .A1(n17742), .A2(n17741), .ZN(P3_U2725) );
  AOI22_X1 U20908 ( .A1(n17753), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17769), .ZN(n17744) );
  OAI222_X1 U20909 ( .A1(n17774), .A2(n17746), .B1(n17745), .B2(n17744), .C1(
        n17771), .C2(n17743), .ZN(P3_U2726) );
  AOI22_X1 U20910 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17777), .B1(n17753), .B2(
        n17875), .ZN(n17749) );
  NAND3_X1 U20911 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17769), .A3(n17747), .ZN(
        n17748) );
  OAI211_X1 U20912 ( .C1(n17750), .C2(n17771), .A(n17749), .B(n17748), .ZN(
        P3_U2727) );
  INV_X1 U20913 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17871) );
  INV_X1 U20914 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17867) );
  INV_X1 U20915 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17860) );
  NOR3_X1 U20916 ( .A1(n17860), .A2(n17858), .A3(n17778), .ZN(n17768) );
  AND2_X1 U20917 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17768), .ZN(n17773) );
  NAND2_X1 U20918 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17773), .ZN(n17761) );
  NOR2_X1 U20919 ( .A1(n17867), .A2(n17761), .ZN(n17764) );
  NAND2_X1 U20920 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17764), .ZN(n17754) );
  NOR2_X1 U20921 ( .A1(n17871), .A2(n17754), .ZN(n17757) );
  AOI21_X1 U20922 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17769), .A(n17757), .ZN(
        n17752) );
  OAI222_X1 U20923 ( .A1(n17774), .A2(n18636), .B1(n17753), .B2(n17752), .C1(
        n17771), .C2(n17751), .ZN(P3_U2728) );
  INV_X1 U20924 ( .A(n17754), .ZN(n17760) );
  AOI21_X1 U20925 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17769), .A(n17760), .ZN(
        n17756) );
  OAI222_X1 U20926 ( .A1(n17774), .A2(n18632), .B1(n17757), .B2(n17756), .C1(
        n17771), .C2(n17755), .ZN(P3_U2729) );
  AOI21_X1 U20927 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17769), .A(n17764), .ZN(
        n17759) );
  OAI222_X1 U20928 ( .A1(n18628), .A2(n17774), .B1(n17760), .B2(n17759), .C1(
        n17771), .C2(n17758), .ZN(P3_U2730) );
  INV_X1 U20929 ( .A(n17761), .ZN(n17767) );
  AOI21_X1 U20930 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17769), .A(n17767), .ZN(
        n17763) );
  OAI222_X1 U20931 ( .A1(n18624), .A2(n17774), .B1(n17764), .B2(n17763), .C1(
        n17771), .C2(n17762), .ZN(P3_U2731) );
  AOI21_X1 U20932 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17769), .A(n17773), .ZN(
        n17766) );
  OAI222_X1 U20933 ( .A1(n18620), .A2(n17774), .B1(n17767), .B2(n17766), .C1(
        n17771), .C2(n17765), .ZN(P3_U2732) );
  AOI21_X1 U20934 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17769), .A(n17768), .ZN(
        n17772) );
  OAI222_X1 U20935 ( .A1(n18616), .A2(n17774), .B1(n17773), .B2(n17772), .C1(
        n17771), .C2(n17770), .ZN(P3_U2733) );
  AOI22_X1 U20936 ( .A1(n17777), .A2(BUF2_REG_1__SCAN_IN), .B1(n17776), .B2(
        n17775), .ZN(n17783) );
  NOR2_X1 U20937 ( .A1(n17858), .A2(n17778), .ZN(n17781) );
  NOR2_X1 U20938 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17778), .ZN(n17780) );
  OAI22_X1 U20939 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17781), .B1(n17780), .B2(
        n17779), .ZN(n17782) );
  NAND2_X1 U20940 ( .A1(n17783), .A2(n17782), .ZN(P3_U2734) );
  NOR2_X1 U20941 ( .A1(n19212), .A2(n18090), .ZN(n17822) );
  INV_X1 U20942 ( .A(n17822), .ZN(n19251) );
  INV_X1 U20943 ( .A(n19251), .ZN(n19096) );
  INV_X1 U20944 ( .A(n17825), .ZN(n17826) );
  NOR2_X1 U20945 ( .A1(n17811), .A2(n17785), .ZN(P3_U2736) );
  INV_X1 U20946 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17856) );
  INV_X2 U20947 ( .A(n17811), .ZN(n17820) );
  AOI22_X1 U20948 ( .A1(n19096), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17787) );
  OAI21_X1 U20949 ( .B1(n17856), .B2(n17803), .A(n17787), .ZN(P3_U2737) );
  INV_X1 U20950 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17854) );
  AOI22_X1 U20951 ( .A1(n19096), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17788) );
  OAI21_X1 U20952 ( .B1(n17854), .B2(n17803), .A(n17788), .ZN(P3_U2738) );
  AOI22_X1 U20953 ( .A1(n19096), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17789) );
  OAI21_X1 U20954 ( .B1(n17852), .B2(n17803), .A(n17789), .ZN(P3_U2739) );
  INV_X1 U20955 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17850) );
  AOI22_X1 U20956 ( .A1(n19096), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17790) );
  OAI21_X1 U20957 ( .B1(n17850), .B2(n17803), .A(n17790), .ZN(P3_U2740) );
  INV_X1 U20958 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n20905) );
  INV_X1 U20959 ( .A(n17803), .ZN(n17791) );
  AOI22_X1 U20960 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17791), .B1(n19096), 
        .B2(P3_UWORD_REG_10__SCAN_IN), .ZN(n17792) );
  OAI21_X1 U20961 ( .B1(n20905), .B2(n17811), .A(n17792), .ZN(P3_U2741) );
  INV_X1 U20962 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17846) );
  AOI22_X1 U20963 ( .A1(n19096), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17793) );
  OAI21_X1 U20964 ( .B1(n17846), .B2(n17803), .A(n17793), .ZN(P3_U2742) );
  INV_X1 U20965 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17844) );
  AOI22_X1 U20966 ( .A1(n19096), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17794) );
  OAI21_X1 U20967 ( .B1(n17844), .B2(n17803), .A(n17794), .ZN(P3_U2743) );
  INV_X1 U20968 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17842) );
  AOI22_X1 U20969 ( .A1(n19096), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17795) );
  OAI21_X1 U20970 ( .B1(n17842), .B2(n17803), .A(n17795), .ZN(P3_U2744) );
  AOI22_X1 U20971 ( .A1(n19096), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17796) );
  OAI21_X1 U20972 ( .B1(n17840), .B2(n17803), .A(n17796), .ZN(P3_U2745) );
  AOI22_X1 U20973 ( .A1(n19096), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17797) );
  OAI21_X1 U20974 ( .B1(n20871), .B2(n17803), .A(n17797), .ZN(P3_U2746) );
  AOI22_X1 U20975 ( .A1(n19096), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17798) );
  OAI21_X1 U20976 ( .B1(n17837), .B2(n17803), .A(n17798), .ZN(P3_U2747) );
  INV_X1 U20977 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U20978 ( .A1(n19096), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17799) );
  OAI21_X1 U20979 ( .B1(n17835), .B2(n17803), .A(n17799), .ZN(P3_U2748) );
  AOI22_X1 U20980 ( .A1(n19096), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17800) );
  OAI21_X1 U20981 ( .B1(n17833), .B2(n17803), .A(n17800), .ZN(P3_U2749) );
  INV_X1 U20982 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17831) );
  AOI22_X1 U20983 ( .A1(n19096), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17801) );
  OAI21_X1 U20984 ( .B1(n17831), .B2(n17803), .A(n17801), .ZN(P3_U2750) );
  INV_X1 U20985 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17829) );
  AOI22_X1 U20986 ( .A1(n19096), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17802) );
  OAI21_X1 U20987 ( .B1(n17829), .B2(n17803), .A(n17802), .ZN(P3_U2751) );
  AOI22_X1 U20988 ( .A1(n19096), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17804) );
  OAI21_X1 U20989 ( .B1(n17894), .B2(n17824), .A(n17804), .ZN(P3_U2752) );
  AOI22_X1 U20990 ( .A1(n17822), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17805) );
  OAI21_X1 U20991 ( .B1(n17889), .B2(n17824), .A(n17805), .ZN(P3_U2753) );
  INV_X1 U20992 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17887) );
  AOI22_X1 U20993 ( .A1(n17822), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17806) );
  OAI21_X1 U20994 ( .B1(n17887), .B2(n17824), .A(n17806), .ZN(P3_U2754) );
  INV_X1 U20995 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17885) );
  AOI22_X1 U20996 ( .A1(n17822), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17807) );
  OAI21_X1 U20997 ( .B1(n17885), .B2(n17824), .A(n17807), .ZN(P3_U2755) );
  AOI22_X1 U20998 ( .A1(n17822), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17808) );
  OAI21_X1 U20999 ( .B1(n17881), .B2(n17824), .A(n17808), .ZN(P3_U2756) );
  INV_X1 U21000 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n21040) );
  AOI22_X1 U21001 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17817), .B1(n17820), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17809) );
  OAI21_X1 U21002 ( .B1(n21040), .B2(n19251), .A(n17809), .ZN(P3_U2757) );
  AOI22_X1 U21003 ( .A1(n17822), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17810) );
  OAI21_X1 U21004 ( .B1(n17877), .B2(n17824), .A(n17810), .ZN(P3_U2758) );
  INV_X1 U21005 ( .A(P3_LWORD_REG_8__SCAN_IN), .ZN(n17812) );
  INV_X1 U21006 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n20914) );
  OAI222_X1 U21007 ( .A1(n17812), .A2(n19251), .B1(n17811), .B2(n20914), .C1(
        n17875), .C2(n17824), .ZN(P3_U2759) );
  INV_X1 U21008 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17873) );
  AOI22_X1 U21009 ( .A1(n17822), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17813) );
  OAI21_X1 U21010 ( .B1(n17873), .B2(n17824), .A(n17813), .ZN(P3_U2760) );
  AOI22_X1 U21011 ( .A1(n19096), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17814) );
  OAI21_X1 U21012 ( .B1(n17871), .B2(n17824), .A(n17814), .ZN(P3_U2761) );
  INV_X1 U21013 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17869) );
  AOI22_X1 U21014 ( .A1(n17822), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17815) );
  OAI21_X1 U21015 ( .B1(n17869), .B2(n17824), .A(n17815), .ZN(P3_U2762) );
  AOI22_X1 U21016 ( .A1(n17822), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17816) );
  OAI21_X1 U21017 ( .B1(n17867), .B2(n17824), .A(n17816), .ZN(P3_U2763) );
  INV_X1 U21018 ( .A(P3_LWORD_REG_3__SCAN_IN), .ZN(n20906) );
  AOI22_X1 U21019 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17817), .B1(n17820), .B2(
        P3_DATAO_REG_3__SCAN_IN), .ZN(n17818) );
  OAI21_X1 U21020 ( .B1(n20906), .B2(n19251), .A(n17818), .ZN(P3_U2764) );
  INV_X1 U21021 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17862) );
  AOI22_X1 U21022 ( .A1(n17822), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17819) );
  OAI21_X1 U21023 ( .B1(n17862), .B2(n17824), .A(n17819), .ZN(P3_U2765) );
  AOI22_X1 U21024 ( .A1(n17822), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17821) );
  OAI21_X1 U21025 ( .B1(n17860), .B2(n17824), .A(n17821), .ZN(P3_U2766) );
  AOI22_X1 U21026 ( .A1(n17822), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17820), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17823) );
  OAI21_X1 U21027 ( .B1(n17858), .B2(n17824), .A(n17823), .ZN(P3_U2767) );
  NAND2_X1 U21028 ( .A1(n18613), .A2(n17827), .ZN(n19091) );
  NOR2_X1 U21029 ( .A1(n17825), .A2(n19091), .ZN(n17863) );
  AOI22_X1 U21030 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17891), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17890), .ZN(n17828) );
  OAI21_X1 U21031 ( .B1(n17829), .B2(n17893), .A(n17828), .ZN(P3_U2768) );
  AOI22_X1 U21032 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17891), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17890), .ZN(n17830) );
  OAI21_X1 U21033 ( .B1(n17831), .B2(n17893), .A(n17830), .ZN(P3_U2769) );
  AOI22_X1 U21034 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17890), .ZN(n17832) );
  OAI21_X1 U21035 ( .B1(n17833), .B2(n17893), .A(n17832), .ZN(P3_U2770) );
  AOI22_X1 U21036 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17890), .ZN(n17834) );
  OAI21_X1 U21037 ( .B1(n17835), .B2(n17893), .A(n17834), .ZN(P3_U2771) );
  AOI22_X1 U21038 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17890), .ZN(n17836) );
  OAI21_X1 U21039 ( .B1(n17837), .B2(n17893), .A(n17836), .ZN(P3_U2772) );
  AOI22_X1 U21040 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17890), .ZN(n17838) );
  OAI21_X1 U21041 ( .B1(n20871), .B2(n17893), .A(n17838), .ZN(P3_U2773) );
  AOI22_X1 U21042 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17890), .ZN(n17839) );
  OAI21_X1 U21043 ( .B1(n17840), .B2(n17893), .A(n17839), .ZN(P3_U2774) );
  AOI22_X1 U21044 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17890), .ZN(n17841) );
  OAI21_X1 U21045 ( .B1(n17842), .B2(n17893), .A(n17841), .ZN(P3_U2775) );
  AOI22_X1 U21046 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17890), .ZN(n17843) );
  OAI21_X1 U21047 ( .B1(n17844), .B2(n17893), .A(n17843), .ZN(P3_U2776) );
  AOI22_X1 U21048 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17890), .ZN(n17845) );
  OAI21_X1 U21049 ( .B1(n17846), .B2(n17893), .A(n17845), .ZN(P3_U2777) );
  AOI22_X1 U21050 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17883), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17890), .ZN(n17847) );
  OAI21_X1 U21051 ( .B1(n17848), .B2(n17893), .A(n17847), .ZN(P3_U2778) );
  AOI22_X1 U21052 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17891), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17882), .ZN(n17849) );
  OAI21_X1 U21053 ( .B1(n17850), .B2(n17893), .A(n17849), .ZN(P3_U2779) );
  AOI22_X1 U21054 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17891), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17882), .ZN(n17851) );
  OAI21_X1 U21055 ( .B1(n17852), .B2(n17893), .A(n17851), .ZN(P3_U2780) );
  AOI22_X1 U21056 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17891), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17882), .ZN(n17853) );
  OAI21_X1 U21057 ( .B1(n17854), .B2(n17893), .A(n17853), .ZN(P3_U2781) );
  AOI22_X1 U21058 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17891), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17882), .ZN(n17855) );
  OAI21_X1 U21059 ( .B1(n17856), .B2(n17893), .A(n17855), .ZN(P3_U2782) );
  AOI22_X1 U21060 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17882), .ZN(n17857) );
  OAI21_X1 U21061 ( .B1(n17858), .B2(n17893), .A(n17857), .ZN(P3_U2783) );
  AOI22_X1 U21062 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17882), .ZN(n17859) );
  OAI21_X1 U21063 ( .B1(n17860), .B2(n17893), .A(n17859), .ZN(P3_U2784) );
  AOI22_X1 U21064 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17882), .ZN(n17861) );
  OAI21_X1 U21065 ( .B1(n17862), .B2(n17893), .A(n17861), .ZN(P3_U2785) );
  AOI22_X1 U21066 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17891), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n17863), .ZN(n17864) );
  OAI21_X1 U21067 ( .B1(n17865), .B2(n20906), .A(n17864), .ZN(P3_U2786) );
  AOI22_X1 U21068 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17882), .ZN(n17866) );
  OAI21_X1 U21069 ( .B1(n17867), .B2(n17893), .A(n17866), .ZN(P3_U2787) );
  AOI22_X1 U21070 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17882), .ZN(n17868) );
  OAI21_X1 U21071 ( .B1(n17869), .B2(n17893), .A(n17868), .ZN(P3_U2788) );
  AOI22_X1 U21072 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17890), .ZN(n17870) );
  OAI21_X1 U21073 ( .B1(n17871), .B2(n17893), .A(n17870), .ZN(P3_U2789) );
  AOI22_X1 U21074 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17890), .ZN(n17872) );
  OAI21_X1 U21075 ( .B1(n17873), .B2(n17893), .A(n17872), .ZN(P3_U2790) );
  AOI22_X1 U21076 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17890), .ZN(n17874) );
  OAI21_X1 U21077 ( .B1(n17875), .B2(n17893), .A(n17874), .ZN(P3_U2791) );
  AOI22_X1 U21078 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17890), .ZN(n17876) );
  OAI21_X1 U21079 ( .B1(n17877), .B2(n17893), .A(n17876), .ZN(P3_U2792) );
  AOI22_X1 U21080 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17883), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17890), .ZN(n17878) );
  OAI21_X1 U21081 ( .B1(n17879), .B2(n17893), .A(n17878), .ZN(P3_U2793) );
  AOI22_X1 U21082 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17890), .ZN(n17880) );
  OAI21_X1 U21083 ( .B1(n17881), .B2(n17893), .A(n17880), .ZN(P3_U2794) );
  AOI22_X1 U21084 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17883), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17882), .ZN(n17884) );
  OAI21_X1 U21085 ( .B1(n17885), .B2(n17893), .A(n17884), .ZN(P3_U2795) );
  AOI22_X1 U21086 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17890), .ZN(n17886) );
  OAI21_X1 U21087 ( .B1(n17887), .B2(n17893), .A(n17886), .ZN(P3_U2796) );
  AOI22_X1 U21088 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17890), .ZN(n17888) );
  OAI21_X1 U21089 ( .B1(n17889), .B2(n17893), .A(n17888), .ZN(P3_U2797) );
  AOI22_X1 U21090 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17891), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17890), .ZN(n17892) );
  OAI21_X1 U21091 ( .B1(n17894), .B2(n17893), .A(n17892), .ZN(P3_U2798) );
  INV_X1 U21092 ( .A(n17895), .ZN(n17915) );
  NOR2_X1 U21093 ( .A1(n18254), .A2(n18123), .ZN(n18006) );
  INV_X1 U21094 ( .A(n17896), .ZN(n18266) );
  INV_X1 U21095 ( .A(n18263), .ZN(n17897) );
  OAI22_X1 U21096 ( .A1(n18266), .A2(n18238), .B1(n17897), .B2(n18169), .ZN(
        n17936) );
  NOR2_X1 U21097 ( .A1(n18267), .A2(n17936), .ZN(n17920) );
  NOR3_X1 U21098 ( .A1(n18006), .A2(n17920), .A3(n17898), .ZN(n17907) );
  NAND2_X1 U21099 ( .A1(n9769), .A2(n17899), .ZN(n17905) );
  NOR3_X1 U21100 ( .A1(n18101), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17902), .ZN(n17918) );
  OAI21_X1 U21101 ( .B1(n17900), .B2(n18090), .A(n18242), .ZN(n17901) );
  AOI21_X1 U21102 ( .B1(n19107), .B2(n17902), .A(n17901), .ZN(n17930) );
  OAI21_X1 U21103 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18012), .A(
        n17930), .ZN(n17923) );
  OAI21_X1 U21104 ( .B1(n17918), .B2(n17923), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17904) );
  NAND2_X1 U21105 ( .A1(n18481), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17903) );
  OAI211_X1 U21106 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17905), .A(
        n17904), .B(n17903), .ZN(n17906) );
  AOI211_X1 U21107 ( .C1(n18093), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        n17914) );
  AND2_X1 U21108 ( .A1(n17909), .A2(n17916), .ZN(n17911) );
  OAI211_X1 U21109 ( .C1(n17912), .C2(n17911), .A(n18156), .B(n17910), .ZN(
        n17913) );
  OAI211_X1 U21110 ( .C1(n17915), .C2(n17921), .A(n17914), .B(n17913), .ZN(
        P3_U2802) );
  NAND2_X1 U21111 ( .A1(n17916), .A2(n16777), .ZN(n17917) );
  XNOR2_X1 U21112 ( .A(n17917), .B(n18052), .ZN(n18272) );
  NOR2_X1 U21113 ( .A1(n18476), .A2(n19177), .ZN(n18259) );
  AOI211_X1 U21114 ( .C1(n18093), .C2(n17919), .A(n18259), .B(n17918), .ZN(
        n17925) );
  AOI21_X1 U21115 ( .B1(n18267), .B2(n17921), .A(n17920), .ZN(n17922) );
  AOI21_X1 U21116 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17923), .A(
        n17922), .ZN(n17924) );
  OAI211_X1 U21117 ( .C1(n18272), .C2(n18170), .A(n17925), .B(n17924), .ZN(
        P3_U2803) );
  INV_X1 U21118 ( .A(n17926), .ZN(n17942) );
  XNOR2_X1 U21119 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n17927), .ZN(
        n18278) );
  INV_X1 U21120 ( .A(n18012), .ZN(n17932) );
  INV_X2 U21121 ( .A(n18843), .ZN(n18982) );
  AOI21_X1 U21122 ( .B1(n18982), .B2(n17928), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17929) );
  OAI22_X1 U21123 ( .A1(n17930), .A2(n17929), .B1(n18476), .B2(n19175), .ZN(
        n17931) );
  AOI221_X1 U21124 ( .B1(n18093), .B2(n17933), .C1(n17932), .C2(n17933), .A(
        n17931), .ZN(n17938) );
  AND3_X1 U21125 ( .A1(n17935), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n17934), .ZN(n18274) );
  AOI22_X1 U21126 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17936), .B1(
        n17961), .B2(n18274), .ZN(n17937) );
  OAI211_X1 U21127 ( .C1(n18170), .C2(n18278), .A(n17938), .B(n17937), .ZN(
        P3_U2804) );
  AND2_X1 U21128 ( .A1(n17947), .A2(n18982), .ZN(n17966) );
  AOI211_X1 U21129 ( .C1(n17985), .C2(n17939), .A(n18251), .B(n17966), .ZN(
        n17974) );
  OAI21_X1 U21130 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18012), .A(
        n17974), .ZN(n17953) );
  AOI22_X1 U21131 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17953), .B1(
        n18093), .B2(n17940), .ZN(n17951) );
  AOI21_X1 U21132 ( .B1(n18052), .B2(n17942), .A(n17941), .ZN(n17943) );
  XNOR2_X1 U21133 ( .A(n17943), .B(n18286), .ZN(n18291) );
  XNOR2_X1 U21134 ( .A(n17944), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18288) );
  XNOR2_X1 U21135 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17945), .ZN(
        n18287) );
  OAI22_X1 U21136 ( .A1(n18238), .A2(n18288), .B1(n18169), .B2(n18287), .ZN(
        n17946) );
  AOI21_X1 U21137 ( .B1(n18156), .B2(n18291), .A(n17946), .ZN(n17950) );
  NAND2_X1 U21138 ( .A1(n18481), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18285) );
  NOR2_X1 U21139 ( .A1(n18101), .A2(n17947), .ZN(n17955) );
  OAI211_X1 U21140 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17955), .B(n17948), .ZN(n17949) );
  NAND4_X1 U21141 ( .A1(n17951), .A2(n17950), .A3(n18285), .A4(n17949), .ZN(
        P3_U2805) );
  INV_X1 U21142 ( .A(n18093), .ZN(n18115) );
  INV_X1 U21143 ( .A(n17952), .ZN(n17960) );
  NOR2_X1 U21144 ( .A1(n18476), .A2(n19171), .ZN(n18305) );
  AOI221_X1 U21145 ( .B1(n17955), .B2(n17954), .C1(n17953), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18305), .ZN(n17959) );
  NOR2_X1 U21146 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18316), .ZN(
        n18307) );
  AOI22_X1 U21147 ( .A1(n18254), .A2(n18294), .B1(n18123), .B2(n18293), .ZN(
        n17977) );
  AOI21_X1 U21148 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17956), .A(
        n16136), .ZN(n18309) );
  OAI22_X1 U21149 ( .A1(n17977), .A2(n18302), .B1(n18309), .B2(n18170), .ZN(
        n17957) );
  AOI21_X1 U21150 ( .B1(n17961), .B2(n18307), .A(n17957), .ZN(n17958) );
  OAI211_X1 U21151 ( .C1(n18115), .C2(n17960), .A(n17959), .B(n17958), .ZN(
        P3_U2806) );
  INV_X1 U21152 ( .A(n17961), .ZN(n17978) );
  AOI22_X1 U21153 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18168), .B1(
        n17979), .B2(n17963), .ZN(n17964) );
  NAND2_X1 U21154 ( .A1(n17962), .A2(n17964), .ZN(n17965) );
  XNOR2_X1 U21155 ( .A(n17965), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18313) );
  AOI22_X1 U21156 ( .A1(n18481), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17967), 
        .B2(n17966), .ZN(n17972) );
  NOR2_X1 U21157 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18012), .ZN(
        n17969) );
  AOI22_X1 U21158 ( .A1(n18093), .A2(n17970), .B1(n17969), .B2(n17968), .ZN(
        n17971) );
  OAI211_X1 U21159 ( .C1(n17974), .C2(n17973), .A(n17972), .B(n17971), .ZN(
        n17975) );
  AOI21_X1 U21160 ( .B1(n18156), .B2(n18313), .A(n17975), .ZN(n17976) );
  OAI221_X1 U21161 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17978), 
        .C1(n18316), .C2(n17977), .A(n17976), .ZN(P3_U2807) );
  INV_X1 U21162 ( .A(n17979), .ZN(n17980) );
  INV_X1 U21163 ( .A(n18323), .ZN(n18325) );
  NOR2_X1 U21164 ( .A1(n18318), .A2(n18325), .ZN(n18326) );
  OAI221_X1 U21165 ( .B1(n17980), .B2(n18326), .C1(n17980), .C2(n18051), .A(
        n17962), .ZN(n17981) );
  XNOR2_X1 U21166 ( .A(n18327), .B(n17981), .ZN(n18335) );
  NOR2_X1 U21167 ( .A1(n18396), .A2(n18238), .ZN(n18074) );
  NOR2_X1 U21168 ( .A1(n18397), .A2(n18169), .ZN(n18073) );
  NOR2_X1 U21169 ( .A1(n18074), .A2(n18073), .ZN(n18062) );
  OAI21_X1 U21170 ( .B1(n18006), .B2(n18326), .A(n18062), .ZN(n18003) );
  OR2_X1 U21171 ( .A1(n17983), .A2(n18101), .ZN(n17997) );
  AOI211_X1 U21172 ( .C1(n17996), .C2(n17990), .A(n17982), .B(n17997), .ZN(
        n17992) );
  AOI22_X1 U21173 ( .A1(n17985), .A2(n17984), .B1(n19107), .B2(n17983), .ZN(
        n17986) );
  NAND2_X1 U21174 ( .A1(n17986), .A2(n18242), .ZN(n18010) );
  AOI21_X1 U21175 ( .B1(n17932), .B2(n17987), .A(n18010), .ZN(n17995) );
  AOI22_X1 U21176 ( .A1(n18481), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18093), 
        .B2(n17988), .ZN(n17989) );
  OAI21_X1 U21177 ( .B1(n17995), .B2(n17990), .A(n17989), .ZN(n17991) );
  AOI211_X1 U21178 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18003), .A(
        n17992), .B(n17991), .ZN(n17994) );
  INV_X1 U21179 ( .A(n18063), .ZN(n18047) );
  NAND3_X1 U21180 ( .A1(n18047), .A2(n18326), .A3(n18327), .ZN(n17993) );
  OAI211_X1 U21181 ( .C1(n18170), .C2(n18335), .A(n17994), .B(n17993), .ZN(
        P3_U2808) );
  NAND2_X1 U21182 ( .A1(n18336), .A2(n18341), .ZN(n18347) );
  NAND2_X1 U21183 ( .A1(n18047), .A2(n18323), .ZN(n18029) );
  NAND2_X1 U21184 ( .A1(n18481), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18345) );
  OAI221_X1 U21185 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17997), .C1(
        n17996), .C2(n17995), .A(n18345), .ZN(n17998) );
  AOI21_X1 U21186 ( .B1(n18093), .B2(n17999), .A(n17998), .ZN(n18005) );
  NOR3_X1 U21187 ( .A1(n18030), .A2(n18168), .A3(n18000), .ZN(n18023) );
  INV_X1 U21188 ( .A(n18037), .ZN(n18024) );
  AOI22_X1 U21189 ( .A1(n18336), .A2(n18023), .B1(n18001), .B2(n18024), .ZN(
        n18002) );
  XNOR2_X1 U21190 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18002), .ZN(
        n18344) );
  AOI22_X1 U21191 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18003), .B1(
        n18156), .B2(n18344), .ZN(n18004) );
  OAI211_X1 U21192 ( .C1(n18347), .C2(n18029), .A(n18005), .B(n18004), .ZN(
        P3_U2809) );
  NOR2_X1 U21193 ( .A1(n18364), .A2(n18325), .ZN(n18321) );
  OAI21_X1 U21194 ( .B1(n18006), .B2(n18321), .A(n18062), .ZN(n18026) );
  OAI221_X1 U21195 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18036), 
        .C1(n18364), .C2(n18023), .A(n17962), .ZN(n18007) );
  XOR2_X1 U21196 ( .A(n18351), .B(n18007), .Z(n18354) );
  INV_X1 U21197 ( .A(n18354), .ZN(n18008) );
  NAND2_X1 U21198 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18351), .ZN(
        n18357) );
  OAI22_X1 U21199 ( .A1(n18170), .A2(n18008), .B1(n18029), .B2(n18357), .ZN(
        n18009) );
  AOI21_X1 U21200 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n18026), .A(
        n18009), .ZN(n18016) );
  NAND2_X1 U21201 ( .A1(n18481), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18355) );
  OAI221_X1 U21202 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18982), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18011), .A(n18010), .ZN(
        n18015) );
  OAI21_X1 U21203 ( .B1(n18093), .B2(n17932), .A(n18013), .ZN(n18014) );
  NAND4_X1 U21204 ( .A1(n18016), .A2(n18355), .A3(n18015), .A4(n18014), .ZN(
        P3_U2810) );
  AOI21_X1 U21205 ( .B1(n19107), .B2(n18018), .A(n18251), .ZN(n18044) );
  OAI21_X1 U21206 ( .B1(n18017), .B2(n18090), .A(n18044), .ZN(n18033) );
  NOR2_X1 U21207 ( .A1(n18101), .A2(n18018), .ZN(n18035) );
  OAI211_X1 U21208 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18035), .B(n18019), .ZN(n18020) );
  NAND2_X1 U21209 ( .A1(n18481), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18361) );
  OAI211_X1 U21210 ( .C1(n18115), .C2(n18021), .A(n18020), .B(n18361), .ZN(
        n18022) );
  AOI21_X1 U21211 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18033), .A(
        n18022), .ZN(n18028) );
  AOI21_X1 U21212 ( .B1(n18024), .B2(n18036), .A(n18023), .ZN(n18025) );
  XNOR2_X1 U21213 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n18025), .ZN(
        n18360) );
  AOI22_X1 U21214 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18026), .B1(
        n18156), .B2(n18360), .ZN(n18027) );
  OAI211_X1 U21215 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18029), .A(
        n18028), .B(n18027), .ZN(P3_U2811) );
  NAND2_X1 U21216 ( .A1(n18370), .A2(n18030), .ZN(n18377) );
  OAI22_X1 U21217 ( .A1(n18476), .A2(n19159), .B1(n18115), .B2(n18031), .ZN(
        n18032) );
  AOI221_X1 U21218 ( .B1(n18035), .B2(n18034), .C1(n18033), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18032), .ZN(n18040) );
  OAI21_X1 U21219 ( .B1(n18370), .B2(n18063), .A(n18062), .ZN(n18046) );
  AOI21_X1 U21220 ( .B1(n18052), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n18036), .ZN(n18038) );
  XNOR2_X1 U21221 ( .A(n18038), .B(n18037), .ZN(n18373) );
  AOI22_X1 U21222 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18046), .B1(
        n18156), .B2(n18373), .ZN(n18039) );
  OAI211_X1 U21223 ( .C1(n18063), .C2(n18377), .A(n18040), .B(n18039), .ZN(
        P3_U2812) );
  OAI21_X1 U21224 ( .B1(n18042), .B2(n18378), .A(n18041), .ZN(n18383) );
  AOI21_X1 U21225 ( .B1(n18982), .B2(n9785), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18043) );
  INV_X1 U21226 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19157) );
  OAI22_X1 U21227 ( .A1(n18044), .A2(n18043), .B1(n18476), .B2(n19157), .ZN(
        n18045) );
  AOI21_X1 U21228 ( .B1(n18156), .B2(n18383), .A(n18045), .ZN(n18049) );
  OAI221_X1 U21229 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18047), .A(n18046), .ZN(
        n18048) );
  OAI211_X1 U21230 ( .C1(n18250), .C2(n18050), .A(n18049), .B(n18048), .ZN(
        P3_U2813) );
  NAND2_X1 U21231 ( .A1(n18052), .A2(n18453), .ZN(n18149) );
  OAI22_X1 U21232 ( .A1(n18052), .A2(n18051), .B1(n18149), .B2(n18320), .ZN(
        n18053) );
  XNOR2_X1 U21233 ( .A(n18380), .B(n18053), .ZN(n18391) );
  AOI21_X1 U21234 ( .B1(n19107), .B2(n18055), .A(n18251), .ZN(n18079) );
  OAI21_X1 U21235 ( .B1(n18054), .B2(n18090), .A(n18079), .ZN(n18070) );
  AOI22_X1 U21236 ( .A1(n18481), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18070), .ZN(n18058) );
  NOR2_X1 U21237 ( .A1(n18101), .A2(n18055), .ZN(n18072) );
  OAI211_X1 U21238 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18072), .B(n18056), .ZN(n18057) );
  OAI211_X1 U21239 ( .C1(n18115), .C2(n18059), .A(n18058), .B(n18057), .ZN(
        n18060) );
  AOI21_X1 U21240 ( .B1(n18156), .B2(n18391), .A(n18060), .ZN(n18061) );
  OAI221_X1 U21241 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18063), 
        .C1(n18380), .C2(n18062), .A(n18061), .ZN(P3_U2814) );
  NAND2_X1 U21242 ( .A1(n18411), .A2(n18095), .ZN(n18064) );
  NOR3_X1 U21243 ( .A1(n18420), .A2(n18168), .A3(n18064), .ZN(n18065) );
  NAND2_X1 U21244 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18098), .ZN(
        n18442) );
  OAI21_X1 U21245 ( .B1(n18066), .B2(n18065), .A(n18442), .ZN(n18067) );
  XNOR2_X1 U21246 ( .A(n18067), .B(n18410), .ZN(n18403) );
  OAI22_X1 U21247 ( .A1(n18476), .A2(n19153), .B1(n18115), .B2(n18068), .ZN(
        n18069) );
  AOI221_X1 U21248 ( .B1(n18072), .B2(n18071), .C1(n18070), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18069), .ZN(n18076) );
  NAND2_X1 U21249 ( .A1(n18077), .A2(n18410), .ZN(n18406) );
  NAND2_X1 U21250 ( .A1(n18410), .A2(n18082), .ZN(n18401) );
  AOI22_X1 U21251 ( .A1(n18074), .A2(n18406), .B1(n18073), .B2(n18401), .ZN(
        n18075) );
  OAI211_X1 U21252 ( .C1(n18170), .C2(n18403), .A(n18076), .B(n18075), .ZN(
        P3_U2815) );
  INV_X1 U21253 ( .A(n18417), .ZN(n18083) );
  OAI221_X1 U21254 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18083), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18450), .A(n18077), .ZN(
        n18428) );
  INV_X1 U21255 ( .A(n18250), .ZN(n18217) );
  NOR3_X1 U21256 ( .A1(n18843), .A2(n18192), .A3(n18193), .ZN(n18181) );
  NAND2_X1 U21257 ( .A1(n18078), .A2(n18181), .ZN(n18128) );
  AOI221_X1 U21258 ( .B1(n18102), .B2(n9967), .C1(n18128), .C2(n9967), .A(
        n18079), .ZN(n18080) );
  NOR2_X1 U21259 ( .A1(n18476), .A2(n19152), .ZN(n18422) );
  AOI211_X1 U21260 ( .C1(n18081), .C2(n18217), .A(n18080), .B(n18422), .ZN(
        n18088) );
  OAI221_X1 U21261 ( .B1(n18083), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n18453), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n18082), .ZN(
        n18084) );
  INV_X1 U21262 ( .A(n18084), .ZN(n18424) );
  OAI22_X1 U21263 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18085), .B1(
        n18149), .B2(n18417), .ZN(n18086) );
  XNOR2_X1 U21264 ( .A(n18420), .B(n18086), .ZN(n18423) );
  AOI22_X1 U21265 ( .A1(n18123), .A2(n18424), .B1(n18156), .B2(n18423), .ZN(
        n18087) );
  OAI211_X1 U21266 ( .C1(n18238), .C2(n18428), .A(n18088), .B(n18087), .ZN(
        P3_U2816) );
  AOI21_X1 U21267 ( .B1(n19107), .B2(n18100), .A(n18251), .ZN(n18089) );
  OAI21_X1 U21268 ( .B1(n18091), .B2(n18090), .A(n18089), .ZN(n18110) );
  AOI22_X1 U21269 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18110), .B1(
        n18093), .B2(n18092), .ZN(n18106) );
  INV_X1 U21270 ( .A(n18094), .ZN(n18107) );
  AOI22_X1 U21271 ( .A1(n18095), .A2(n18411), .B1(n21047), .B2(n18168), .ZN(
        n18096) );
  AOI21_X1 U21272 ( .B1(n18107), .B2(n18168), .A(n18096), .ZN(n18097) );
  XNOR2_X1 U21273 ( .A(n18097), .B(n18098), .ZN(n18430) );
  NAND2_X1 U21274 ( .A1(n18411), .A2(n18450), .ZN(n18433) );
  NAND2_X1 U21275 ( .A1(n18411), .A2(n18453), .ZN(n18431) );
  AOI22_X1 U21276 ( .A1(n18254), .A2(n18433), .B1(n18123), .B2(n18431), .ZN(
        n18118) );
  INV_X1 U21277 ( .A(n18444), .ZN(n18429) );
  NAND2_X1 U21278 ( .A1(n18429), .A2(n18125), .ZN(n18119) );
  OAI22_X1 U21279 ( .A1(n18118), .A2(n18098), .B1(n18442), .B2(n18119), .ZN(
        n18099) );
  AOI21_X1 U21280 ( .B1(n18156), .B2(n18430), .A(n18099), .ZN(n18105) );
  NAND2_X1 U21281 ( .A1(n18481), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18104) );
  NOR2_X1 U21282 ( .A1(n18101), .A2(n18100), .ZN(n18112) );
  OAI211_X1 U21283 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18112), .B(n18102), .ZN(n18103) );
  NAND4_X1 U21284 ( .A1(n18106), .A2(n18105), .A3(n18104), .A4(n18103), .ZN(
        P3_U2817) );
  OAI21_X1 U21285 ( .B1(n18444), .B2(n18149), .A(n18107), .ZN(n18108) );
  XNOR2_X1 U21286 ( .A(n18108), .B(n21047), .ZN(n18443) );
  INV_X1 U21287 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18111) );
  NOR2_X1 U21288 ( .A1(n18476), .A2(n19147), .ZN(n18109) );
  AOI221_X1 U21289 ( .B1(n18112), .B2(n18111), .C1(n18110), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18109), .ZN(n18113) );
  OAI21_X1 U21290 ( .B1(n18115), .B2(n18114), .A(n18113), .ZN(n18116) );
  AOI21_X1 U21291 ( .B1(n18156), .B2(n18443), .A(n18116), .ZN(n18117) );
  OAI221_X1 U21292 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18119), 
        .C1(n21047), .C2(n18118), .A(n18117), .ZN(P3_U2818) );
  INV_X1 U21293 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18126) );
  NAND2_X1 U21294 ( .A1(n18456), .A2(n18126), .ZN(n18463) );
  INV_X1 U21295 ( .A(n18456), .ZN(n18141) );
  OAI21_X1 U21296 ( .B1(n18141), .B2(n18149), .A(n18120), .ZN(n18121) );
  XOR2_X1 U21297 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18121), .Z(
        n18449) );
  INV_X1 U21298 ( .A(n18450), .ZN(n18124) );
  AOI22_X1 U21299 ( .A1(n18254), .A2(n18124), .B1(n18123), .B2(n18122), .ZN(
        n18158) );
  NAND2_X1 U21300 ( .A1(n18141), .A2(n18125), .ZN(n18147) );
  AOI21_X1 U21301 ( .B1(n18158), .B2(n18147), .A(n18126), .ZN(n18133) );
  NAND3_X1 U21302 ( .A1(n18162), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18181), .ZN(n18135) );
  NOR2_X1 U21303 ( .A1(n18127), .A2(n18135), .ZN(n18137) );
  NAND2_X1 U21304 ( .A1(n18242), .A2(n18160), .ZN(n18247) );
  OAI211_X1 U21305 ( .C1(n18137), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n18247), .B(n18128), .ZN(n18130) );
  NAND2_X1 U21306 ( .A1(n18481), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18129) );
  OAI211_X1 U21307 ( .C1(n18250), .C2(n18131), .A(n18130), .B(n18129), .ZN(
        n18132) );
  AOI211_X1 U21308 ( .C1(n18156), .C2(n18449), .A(n18133), .B(n18132), .ZN(
        n18134) );
  OAI21_X1 U21309 ( .B1(n18159), .B2(n18463), .A(n18134), .ZN(P3_U2819) );
  INV_X1 U21310 ( .A(n18135), .ZN(n18153) );
  AOI21_X1 U21311 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18247), .A(
        n18153), .ZN(n18136) );
  NAND2_X1 U21312 ( .A1(n18481), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18469) );
  OAI21_X1 U21313 ( .B1(n18137), .B2(n18136), .A(n18469), .ZN(n18144) );
  OAI221_X1 U21314 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n9700), .C1(
        n18484), .C2(n18149), .A(n18142), .ZN(n18140) );
  NAND4_X1 U21315 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18138), .A3(
        n18484), .A4(n18168), .ZN(n18139) );
  OAI211_X1 U21316 ( .C1(n18149), .C2(n18141), .A(n18140), .B(n18139), .ZN(
        n18471) );
  OAI22_X1 U21317 ( .A1(n18158), .A2(n18142), .B1(n18170), .B2(n18471), .ZN(
        n18143) );
  AOI211_X1 U21318 ( .C1(n18145), .C2(n18217), .A(n18144), .B(n18143), .ZN(
        n18146) );
  OAI21_X1 U21319 ( .B1(n18148), .B2(n18147), .A(n18146), .ZN(P3_U2820) );
  NAND2_X1 U21320 ( .A1(n18149), .A2(n9700), .ZN(n18150) );
  XNOR2_X1 U21321 ( .A(n18150), .B(n18484), .ZN(n18479) );
  NOR2_X1 U21322 ( .A1(n18476), .A2(n19141), .ZN(n18155) );
  AOI22_X1 U21323 ( .A1(n18162), .A2(n18181), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18247), .ZN(n18152) );
  OAI22_X1 U21324 ( .A1(n18153), .A2(n18152), .B1(n18250), .B2(n18151), .ZN(
        n18154) );
  AOI211_X1 U21325 ( .C1(n18156), .C2(n18479), .A(n18155), .B(n18154), .ZN(
        n18157) );
  OAI221_X1 U21326 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18159), .C1(
        n18484), .C2(n18158), .A(n18157), .ZN(P3_U2821) );
  OAI21_X1 U21327 ( .B1(n18161), .B2(n18160), .A(n18242), .ZN(n18179) );
  INV_X1 U21328 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18164) );
  AOI211_X1 U21329 ( .C1(n18164), .C2(n18163), .A(n18162), .B(n18843), .ZN(
        n18165) );
  NOR2_X1 U21330 ( .A1(n18476), .A2(n19139), .ZN(n18501) );
  AOI211_X1 U21331 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18179), .A(
        n18165), .B(n18501), .ZN(n18173) );
  XNOR2_X1 U21332 ( .A(n21015), .B(n18166), .ZN(n18495) );
  AOI21_X1 U21333 ( .B1(n18168), .B2(n18497), .A(n18167), .ZN(n18505) );
  OAI22_X1 U21334 ( .A1(n18505), .A2(n18170), .B1(n18169), .B2(n18497), .ZN(
        n18171) );
  AOI21_X1 U21335 ( .B1(n18254), .B2(n18495), .A(n18171), .ZN(n18172) );
  OAI211_X1 U21336 ( .C1(n18250), .C2(n18174), .A(n18173), .B(n18172), .ZN(
        P3_U2822) );
  OAI21_X1 U21337 ( .B1(n18177), .B2(n18176), .A(n18175), .ZN(n18178) );
  XNOR2_X1 U21338 ( .A(n18178), .B(n18514), .ZN(n18509) );
  INV_X1 U21339 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19137) );
  NOR2_X1 U21340 ( .A1(n18476), .A2(n19137), .ZN(n18511) );
  AOI221_X1 U21341 ( .B1(n18181), .B2(n18180), .C1(n18179), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18511), .ZN(n18186) );
  AOI21_X1 U21342 ( .B1(n18514), .B2(n18183), .A(n18182), .ZN(n18506) );
  AOI22_X1 U21343 ( .A1(n18255), .A2(n18506), .B1(n18184), .B2(n18217), .ZN(
        n18185) );
  OAI211_X1 U21344 ( .C1(n18238), .C2(n18509), .A(n18186), .B(n18185), .ZN(
        P3_U2823) );
  NOR2_X1 U21345 ( .A1(n18843), .A2(n18192), .ZN(n18187) );
  AOI22_X1 U21346 ( .A1(n18481), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18187), 
        .B2(n18193), .ZN(n18196) );
  AOI21_X1 U21347 ( .B1(n9782), .B2(n18189), .A(n18188), .ZN(n18521) );
  OAI21_X1 U21348 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18191), .A(
        n18190), .ZN(n18523) );
  OAI21_X1 U21349 ( .B1(n18192), .B2(n18843), .A(n18247), .ZN(n18204) );
  OAI22_X1 U21350 ( .A1(n18238), .A2(n18523), .B1(n18193), .B2(n18204), .ZN(
        n18194) );
  AOI21_X1 U21351 ( .B1(n18255), .B2(n18521), .A(n18194), .ZN(n18195) );
  OAI211_X1 U21352 ( .C1(n18250), .C2(n18197), .A(n18196), .B(n18195), .ZN(
        P3_U2824) );
  OAI21_X1 U21353 ( .B1(n18200), .B2(n18199), .A(n18198), .ZN(n18532) );
  AOI21_X1 U21354 ( .B1(n18526), .B2(n18202), .A(n18201), .ZN(n18530) );
  AOI21_X1 U21355 ( .B1(n18203), .B2(n18242), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18205) );
  OAI22_X1 U21356 ( .A1(n18250), .A2(n18206), .B1(n18205), .B2(n18204), .ZN(
        n18207) );
  AOI21_X1 U21357 ( .B1(n18255), .B2(n18530), .A(n18207), .ZN(n18208) );
  NAND2_X1 U21358 ( .A1(n18481), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18525) );
  OAI211_X1 U21359 ( .C1(n18238), .C2(n18532), .A(n18208), .B(n18525), .ZN(
        P3_U2825) );
  AOI21_X1 U21360 ( .B1(n19107), .B2(n18209), .A(n18251), .ZN(n18229) );
  AOI21_X1 U21361 ( .B1(n18212), .B2(n18211), .A(n18210), .ZN(n18546) );
  OAI22_X1 U21362 ( .A1(n18546), .A2(n18238), .B1(n18476), .B2(n19131), .ZN(
        n18213) );
  AOI21_X1 U21363 ( .B1(n18982), .B2(n18214), .A(n18213), .ZN(n18220) );
  AOI21_X1 U21364 ( .B1(n9784), .B2(n18216), .A(n18215), .ZN(n18544) );
  AOI22_X1 U21365 ( .A1(n18255), .A2(n18544), .B1(n18218), .B2(n18217), .ZN(
        n18219) );
  OAI211_X1 U21366 ( .C1(n18229), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        P3_U2826) );
  OAI21_X1 U21367 ( .B1(n18224), .B2(n18223), .A(n18222), .ZN(n18548) );
  AOI21_X1 U21368 ( .B1(n18549), .B2(n18226), .A(n18225), .ZN(n18552) );
  AOI21_X1 U21369 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18242), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18228) );
  OAI22_X1 U21370 ( .A1(n18229), .A2(n18228), .B1(n18250), .B2(n18227), .ZN(
        n18230) );
  AOI21_X1 U21371 ( .B1(n18255), .B2(n18552), .A(n18230), .ZN(n18231) );
  NAND2_X1 U21372 ( .A1(n18481), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18547) );
  OAI211_X1 U21373 ( .C1(n18238), .C2(n18548), .A(n18231), .B(n18547), .ZN(
        P3_U2827) );
  AOI21_X1 U21374 ( .B1(n18234), .B2(n18233), .A(n18232), .ZN(n18567) );
  INV_X1 U21375 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19127) );
  NOR2_X1 U21376 ( .A1(n18476), .A2(n19127), .ZN(n18557) );
  OAI21_X1 U21377 ( .B1(n18237), .B2(n18236), .A(n18235), .ZN(n18571) );
  OAI22_X1 U21378 ( .A1(n18250), .A2(n18239), .B1(n18238), .B2(n18571), .ZN(
        n18240) );
  AOI211_X1 U21379 ( .C1(n18255), .C2(n18567), .A(n18557), .B(n18240), .ZN(
        n18241) );
  OAI221_X1 U21380 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18843), .C1(
        n18243), .C2(n18242), .A(n18241), .ZN(P3_U2828) );
  NOR2_X1 U21381 ( .A1(n18253), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18244) );
  XNOR2_X1 U21382 ( .A(n18244), .B(n18246), .ZN(n18579) );
  AOI22_X1 U21383 ( .A1(n18254), .A2(n18579), .B1(n18481), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18249) );
  AOI21_X1 U21384 ( .B1(n18246), .B2(n18252), .A(n18245), .ZN(n18573) );
  AOI22_X1 U21385 ( .A1(n18255), .A2(n18573), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18247), .ZN(n18248) );
  OAI211_X1 U21386 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18250), .A(
        n18249), .B(n18248), .ZN(P3_U2829) );
  AOI21_X1 U21387 ( .B1(n19102), .B2(n19248), .A(n18251), .ZN(n18258) );
  OAI21_X1 U21388 ( .B1(n18253), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18252), .ZN(n18589) );
  INV_X1 U21389 ( .A(n18589), .ZN(n18591) );
  AOI22_X1 U21390 ( .A1(n18591), .A2(n18255), .B1(n18254), .B2(n18589), .ZN(
        n18256) );
  NAND2_X1 U21391 ( .A1(n18481), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18587) );
  OAI211_X1 U21392 ( .C1(n18258), .C2(n18257), .A(n18256), .B(n18587), .ZN(
        P3_U2830) );
  AOI21_X1 U21393 ( .B1(n18584), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18259), .ZN(n18271) );
  NOR2_X1 U21394 ( .A1(n18585), .A2(n19068), .ZN(n18487) );
  NOR2_X1 U21395 ( .A1(n18260), .A2(n18487), .ZN(n18262) );
  AOI211_X1 U21396 ( .C1(n18432), .C2(n18263), .A(n18262), .B(n18261), .ZN(
        n18265) );
  NOR2_X1 U21397 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n9660), .ZN(
        n18561) );
  OAI21_X1 U21398 ( .B1(n18561), .B2(n18264), .A(n18560), .ZN(n18280) );
  OAI211_X1 U21399 ( .C1(n18266), .C2(n18451), .A(n18265), .B(n18280), .ZN(
        n18275) );
  OAI22_X1 U21400 ( .A1(n18269), .A2(n18268), .B1(n18267), .B2(n18275), .ZN(
        n18270) );
  OAI211_X1 U21401 ( .C1(n18272), .C2(n18504), .A(n18271), .B(n18270), .ZN(
        P3_U2835) );
  INV_X1 U21402 ( .A(n18273), .ZN(n18306) );
  AOI22_X1 U21403 ( .A1(n18481), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18306), 
        .B2(n18274), .ZN(n18277) );
  OAI211_X1 U21404 ( .C1(n18498), .C2(n18275), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18476), .ZN(n18276) );
  OAI211_X1 U21405 ( .C1(n18278), .C2(n18504), .A(n18277), .B(n18276), .ZN(
        P3_U2836) );
  INV_X1 U21406 ( .A(n18279), .ZN(n18281) );
  OAI21_X1 U21407 ( .B1(n18281), .B2(n18537), .A(n18280), .ZN(n18282) );
  OAI221_X1 U21408 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18283), 
        .C1(n18286), .C2(n18282), .A(n18586), .ZN(n18284) );
  OAI211_X1 U21409 ( .C1(n18575), .C2(n18286), .A(n18285), .B(n18284), .ZN(
        n18290) );
  INV_X1 U21410 ( .A(n18425), .ZN(n18496) );
  OAI22_X1 U21411 ( .A1(n18572), .A2(n18288), .B1(n18496), .B2(n18287), .ZN(
        n18289) );
  AOI211_X1 U21412 ( .C1(n18480), .C2(n18291), .A(n18290), .B(n18289), .ZN(
        n18292) );
  INV_X1 U21413 ( .A(n18292), .ZN(P3_U2837) );
  AOI22_X1 U21414 ( .A1(n19037), .A2(n18294), .B1(n18432), .B2(n18293), .ZN(
        n18298) );
  INV_X1 U21415 ( .A(n18295), .ZN(n18296) );
  OAI21_X1 U21416 ( .B1(n18561), .B2(n18296), .A(n18560), .ZN(n18297) );
  NAND3_X1 U21417 ( .A1(n18298), .A2(n18575), .A3(n18297), .ZN(n18301) );
  INV_X1 U21418 ( .A(n18301), .ZN(n18303) );
  OAI21_X1 U21419 ( .B1(n18299), .B2(n18537), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18300) );
  OAI21_X1 U21420 ( .B1(n18301), .B2(n18300), .A(n18476), .ZN(n18317) );
  AOI211_X1 U21421 ( .C1(n18491), .C2(n18303), .A(n18302), .B(n18317), .ZN(
        n18304) );
  AOI211_X1 U21422 ( .C1(n18307), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        n18308) );
  OAI21_X1 U21423 ( .B1(n18309), .B2(n18504), .A(n18308), .ZN(P3_U2838) );
  INV_X1 U21424 ( .A(n18310), .ZN(n18312) );
  NAND3_X1 U21425 ( .A1(n18312), .A2(n18311), .A3(n18575), .ZN(n18315) );
  AOI22_X1 U21426 ( .A1(n18481), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18480), 
        .B2(n18313), .ZN(n18314) );
  OAI221_X1 U21427 ( .B1(n18317), .B2(n18316), .C1(n18317), .C2(n18315), .A(
        n18314), .ZN(P3_U2839) );
  AOI22_X1 U21428 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18584), .B1(
        n18481), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n18334) );
  NOR2_X1 U21429 ( .A1(n18327), .A2(n18498), .ZN(n18331) );
  INV_X1 U21430 ( .A(n18318), .ZN(n18329) );
  NAND2_X1 U21431 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18319), .ZN(
        n18472) );
  NOR2_X1 U21432 ( .A1(n18320), .A2(n18472), .ZN(n18385) );
  INV_X1 U21433 ( .A(n18321), .ZN(n18349) );
  OAI21_X1 U21434 ( .B1(n18372), .B2(n18349), .A(n18585), .ZN(n18322) );
  OAI221_X1 U21435 ( .B1(n9660), .B2(n18323), .C1(n9660), .C2(n18385), .A(
        n18322), .ZN(n18324) );
  AOI221_X1 U21436 ( .B1(n18367), .B2(n19066), .C1(n18325), .C2(n19066), .A(
        n18324), .ZN(n18338) );
  NOR2_X1 U21437 ( .A1(n19037), .A2(n18432), .ZN(n18455) );
  OAI22_X1 U21438 ( .A1(n18465), .A2(n18336), .B1(n18326), .B2(n18455), .ZN(
        n18339) );
  AOI211_X1 U21439 ( .C1(n18434), .C2(n18341), .A(n18327), .B(n18339), .ZN(
        n18328) );
  OAI211_X1 U21440 ( .C1(n9660), .C2(n18329), .A(n18338), .B(n18328), .ZN(
        n18330) );
  OAI22_X1 U21441 ( .A1(n18396), .A2(n18451), .B1(n18397), .B2(n18452), .ZN(
        n18337) );
  OAI22_X1 U21442 ( .A1(n18332), .A2(n18331), .B1(n18330), .B2(n18337), .ZN(
        n18333) );
  OAI211_X1 U21443 ( .C1(n18335), .C2(n18504), .A(n18334), .B(n18333), .ZN(
        P3_U2840) );
  INV_X1 U21444 ( .A(n18336), .ZN(n18340) );
  NOR2_X1 U21445 ( .A1(n18498), .A2(n18337), .ZN(n18390) );
  NAND2_X1 U21446 ( .A1(n18390), .A2(n18338), .ZN(n18350) );
  AOI211_X1 U21447 ( .C1(n19068), .C2(n18340), .A(n18350), .B(n18339), .ZN(
        n18342) );
  NOR3_X1 U21448 ( .A1(n18481), .A2(n18342), .A3(n18341), .ZN(n18343) );
  AOI21_X1 U21449 ( .B1(n18480), .B2(n18344), .A(n18343), .ZN(n18346) );
  OAI211_X1 U21450 ( .C1(n18347), .C2(n18358), .A(n18346), .B(n18345), .ZN(
        P3_U2841) );
  INV_X1 U21451 ( .A(n18455), .ZN(n18348) );
  OAI221_X1 U21452 ( .B1(n18350), .B2(n18349), .C1(n18350), .C2(n18348), .A(
        n18476), .ZN(n18363) );
  NAND2_X1 U21453 ( .A1(n9660), .A2(n18537), .ZN(n18574) );
  NAND3_X1 U21454 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18364), .A3(n18574), 
        .ZN(n18352) );
  AOI21_X1 U21455 ( .B1(n18363), .B2(n18352), .A(n18351), .ZN(n18353) );
  AOI21_X1 U21456 ( .B1(n18354), .B2(n18480), .A(n18353), .ZN(n18356) );
  OAI211_X1 U21457 ( .C1(n18357), .C2(n18358), .A(n18356), .B(n18355), .ZN(
        P3_U2842) );
  INV_X1 U21458 ( .A(n18358), .ZN(n18359) );
  AOI22_X1 U21459 ( .A1(n18480), .A2(n18360), .B1(n18359), .B2(n18364), .ZN(
        n18362) );
  OAI211_X1 U21460 ( .C1(n18364), .C2(n18363), .A(n18362), .B(n18361), .ZN(
        P3_U2843) );
  AOI21_X1 U21461 ( .B1(n18365), .B2(n18416), .A(n18498), .ZN(n18467) );
  NAND2_X1 U21462 ( .A1(n18366), .A2(n18467), .ZN(n18395) );
  AOI221_X1 U21463 ( .B1(n18368), .B2(n19066), .C1(n18367), .C2(n19066), .A(
        n18561), .ZN(n18369) );
  OAI211_X1 U21464 ( .C1(n18370), .C2(n18455), .A(n18390), .B(n18369), .ZN(
        n18371) );
  AOI221_X1 U21465 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18379), 
        .C1(n18487), .C2(n18379), .A(n18481), .ZN(n18374) );
  AOI22_X1 U21466 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18374), .B1(
        n18480), .B2(n18373), .ZN(n18376) );
  NAND2_X1 U21467 ( .A1(n18481), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18375) );
  OAI211_X1 U21468 ( .C1(n18377), .C2(n18395), .A(n18376), .B(n18375), .ZN(
        P3_U2844) );
  NOR3_X1 U21469 ( .A1(n18481), .A2(n18379), .A3(n18378), .ZN(n18382) );
  NOR3_X1 U21470 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18380), .A3(
        n18395), .ZN(n18381) );
  AOI211_X1 U21471 ( .C1(n18480), .C2(n18383), .A(n18382), .B(n18381), .ZN(
        n18384) );
  OAI21_X1 U21472 ( .B1(n18476), .B2(n19157), .A(n18384), .ZN(P3_U2845) );
  AOI21_X1 U21473 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n9660), .A(
        n18385), .ZN(n18389) );
  INV_X1 U21474 ( .A(n18585), .ZN(n19070) );
  INV_X1 U21475 ( .A(n18386), .ZN(n18388) );
  AOI22_X1 U21476 ( .A1(n19066), .A2(n18388), .B1(n18585), .B2(n18387), .ZN(
        n18473) );
  OAI21_X1 U21477 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19070), .A(
        n18473), .ZN(n18458) );
  AOI211_X1 U21478 ( .C1(n18434), .C2(n18399), .A(n18389), .B(n18458), .ZN(
        n18398) );
  AOI221_X1 U21479 ( .B1(n18491), .B2(n18390), .C1(n18398), .C2(n18390), .A(
        n18481), .ZN(n18392) );
  AOI22_X1 U21480 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18392), .B1(
        n18480), .B2(n18391), .ZN(n18394) );
  NAND2_X1 U21481 ( .A1(n18481), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18393) );
  OAI211_X1 U21482 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18395), .A(
        n18394), .B(n18393), .ZN(P3_U2846) );
  NOR2_X1 U21483 ( .A1(n18396), .A2(n18572), .ZN(n18407) );
  NOR2_X1 U21484 ( .A1(n18397), .A2(n18452), .ZN(n18402) );
  AOI221_X1 U21485 ( .B1(n18399), .B2(n18410), .C1(n18416), .C2(n18410), .A(
        n18398), .ZN(n18400) );
  AOI21_X1 U21486 ( .B1(n18402), .B2(n18401), .A(n18400), .ZN(n18404) );
  OAI22_X1 U21487 ( .A1(n18404), .A2(n18498), .B1(n18504), .B2(n18403), .ZN(
        n18405) );
  AOI21_X1 U21488 ( .B1(n18407), .B2(n18406), .A(n18405), .ZN(n18409) );
  NAND2_X1 U21489 ( .A1(n18481), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18408) );
  OAI211_X1 U21490 ( .C1(n18575), .C2(n18410), .A(n18409), .B(n18408), .ZN(
        P3_U2847) );
  INV_X1 U21491 ( .A(n18574), .ZN(n18414) );
  AOI211_X1 U21492 ( .C1(n18434), .C2(n18417), .A(n18420), .B(n18458), .ZN(
        n18413) );
  INV_X1 U21493 ( .A(n18411), .ZN(n18412) );
  OAI21_X1 U21494 ( .B1(n18412), .B2(n18472), .A(n19068), .ZN(n18435) );
  OAI211_X1 U21495 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18414), .A(
        n18413), .B(n18435), .ZN(n18415) );
  NAND2_X1 U21496 ( .A1(n18586), .A2(n18415), .ZN(n18419) );
  OR2_X1 U21497 ( .A1(n18417), .A2(n18416), .ZN(n18418) );
  AOI222_X1 U21498 ( .A1(n18420), .A2(n18419), .B1(n18420), .B2(n18418), .C1(
        n18419), .C2(n18575), .ZN(n18421) );
  AOI211_X1 U21499 ( .C1(n18480), .C2(n18423), .A(n18422), .B(n18421), .ZN(
        n18427) );
  NAND2_X1 U21500 ( .A1(n18425), .A2(n18424), .ZN(n18426) );
  OAI211_X1 U21501 ( .C1(n18428), .C2(n18572), .A(n18427), .B(n18426), .ZN(
        P3_U2848) );
  NAND2_X1 U21502 ( .A1(n18429), .A2(n18467), .ZN(n18441) );
  AOI22_X1 U21503 ( .A1(n18481), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18480), 
        .B2(n18430), .ZN(n18440) );
  INV_X1 U21504 ( .A(n18458), .ZN(n18437) );
  AOI22_X1 U21505 ( .A1(n19037), .A2(n18433), .B1(n18432), .B2(n18431), .ZN(
        n18436) );
  NAND2_X1 U21506 ( .A1(n18434), .A2(n18444), .ZN(n18459) );
  NAND4_X1 U21507 ( .A1(n18437), .A2(n18436), .A3(n18435), .A4(n18459), .ZN(
        n18446) );
  OAI21_X1 U21508 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18465), .A(
        n18575), .ZN(n18438) );
  OAI211_X1 U21509 ( .C1(n18446), .C2(n18438), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18476), .ZN(n18439) );
  OAI211_X1 U21510 ( .C1(n18442), .C2(n18441), .A(n18440), .B(n18439), .ZN(
        P3_U2849) );
  AOI22_X1 U21511 ( .A1(n18481), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18480), 
        .B2(n18443), .ZN(n18448) );
  INV_X1 U21512 ( .A(n18467), .ZN(n18485) );
  OAI22_X1 U21513 ( .A1(n21047), .A2(n18498), .B1(n18444), .B2(n18485), .ZN(
        n18445) );
  OAI21_X1 U21514 ( .B1(n18446), .B2(n21047), .A(n18445), .ZN(n18447) );
  OAI211_X1 U21515 ( .C1(n18575), .C2(n21047), .A(n18448), .B(n18447), .ZN(
        P3_U2850) );
  AOI22_X1 U21516 ( .A1(n18481), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18480), 
        .B2(n18449), .ZN(n18462) );
  OAI22_X1 U21517 ( .A1(n18453), .A2(n18452), .B1(n18451), .B2(n18450), .ZN(
        n18478) );
  OAI21_X1 U21518 ( .B1(n18484), .B2(n18472), .A(n19068), .ZN(n18454) );
  OAI211_X1 U21519 ( .C1(n18456), .C2(n18455), .A(n18454), .B(n18575), .ZN(
        n18457) );
  NOR3_X1 U21520 ( .A1(n18458), .A2(n18478), .A3(n18457), .ZN(n18464) );
  OAI211_X1 U21521 ( .C1(n9660), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18464), .B(n18459), .ZN(n18460) );
  NAND3_X1 U21522 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18476), .A3(
        n18460), .ZN(n18461) );
  OAI211_X1 U21523 ( .C1(n18463), .C2(n18485), .A(n18462), .B(n18461), .ZN(
        P3_U2851) );
  AOI221_X1 U21524 ( .B1(n18465), .B2(n18464), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18464), .A(n18481), .ZN(
        n18468) );
  NOR2_X1 U21525 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18484), .ZN(
        n18466) );
  AOI22_X1 U21526 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18468), .B1(
        n18467), .B2(n18466), .ZN(n18470) );
  OAI211_X1 U21527 ( .C1(n18504), .C2(n18471), .A(n18470), .B(n18469), .ZN(
        P3_U2852) );
  INV_X1 U21528 ( .A(n18472), .ZN(n18475) );
  AOI21_X1 U21529 ( .B1(n21015), .B2(n18585), .A(n19068), .ZN(n18474) );
  OAI211_X1 U21530 ( .C1(n18475), .C2(n18474), .A(n18473), .B(n18575), .ZN(
        n18477) );
  OAI21_X1 U21531 ( .B1(n18478), .B2(n18477), .A(n18476), .ZN(n18483) );
  AOI22_X1 U21532 ( .A1(n18481), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18480), 
        .B2(n18479), .ZN(n18482) );
  OAI221_X1 U21533 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18485), .C1(
        n18484), .C2(n18483), .A(n18482), .ZN(P3_U2853) );
  OAI21_X1 U21534 ( .B1(n18491), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18490) );
  AOI21_X1 U21535 ( .B1(n19066), .B2(n18486), .A(n18561), .ZN(n18488) );
  AOI221_X1 U21536 ( .B1(n18489), .B2(n18488), .C1(n18487), .C2(n18488), .A(
        n18498), .ZN(n18517) );
  AOI21_X1 U21537 ( .B1(n18586), .B2(n18490), .A(n18517), .ZN(n18515) );
  OAI21_X1 U21538 ( .B1(n18491), .B2(n18515), .A(n18575), .ZN(n18502) );
  INV_X1 U21539 ( .A(n18536), .ZN(n18559) );
  OAI22_X1 U21540 ( .A1(n18559), .A2(n18537), .B1(n18534), .B2(n18492), .ZN(
        n18554) );
  NAND3_X1 U21541 ( .A1(n18493), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18554), .ZN(n18513) );
  NOR2_X1 U21542 ( .A1(n18514), .A2(n18513), .ZN(n18494) );
  AOI22_X1 U21543 ( .A1(n18495), .A2(n19037), .B1(n18494), .B2(n21015), .ZN(
        n18499) );
  OAI22_X1 U21544 ( .A1(n18499), .A2(n18498), .B1(n18497), .B2(n18496), .ZN(
        n18500) );
  AOI211_X1 U21545 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n18502), .A(
        n18501), .B(n18500), .ZN(n18503) );
  OAI21_X1 U21546 ( .B1(n18505), .B2(n18504), .A(n18503), .ZN(P3_U2854) );
  INV_X1 U21547 ( .A(n18506), .ZN(n18508) );
  NAND2_X1 U21548 ( .A1(n18507), .A2(n18586), .ZN(n18582) );
  OAI22_X1 U21549 ( .A1(n18572), .A2(n18509), .B1(n18508), .B2(n18582), .ZN(
        n18510) );
  AOI211_X1 U21550 ( .C1(n18584), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18511), .B(n18510), .ZN(n18512) );
  OAI221_X1 U21551 ( .B1(n18515), .B2(n18514), .C1(n18515), .C2(n18513), .A(
        n18512), .ZN(P3_U2855) );
  NAND2_X1 U21552 ( .A1(n18586), .A2(n18554), .ZN(n18533) );
  NOR3_X1 U21553 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18516), .A3(
        n18533), .ZN(n18520) );
  NOR2_X1 U21554 ( .A1(n18584), .A2(n18517), .ZN(n18527) );
  OAI22_X1 U21555 ( .A1(n18527), .A2(n18518), .B1(n18476), .B2(n19135), .ZN(
        n18519) );
  AOI211_X1 U21556 ( .C1(n18521), .C2(n18592), .A(n18520), .B(n18519), .ZN(
        n18522) );
  OAI21_X1 U21557 ( .B1(n18572), .B2(n18523), .A(n18522), .ZN(P3_U2856) );
  NOR4_X1 U21558 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18524), .A3(
        n18549), .A4(n18533), .ZN(n18529) );
  OAI21_X1 U21559 ( .B1(n18527), .B2(n18526), .A(n18525), .ZN(n18528) );
  AOI211_X1 U21560 ( .C1(n18530), .C2(n18592), .A(n18529), .B(n18528), .ZN(
        n18531) );
  OAI21_X1 U21561 ( .B1(n18572), .B2(n18532), .A(n18531), .ZN(P3_U2857) );
  NOR2_X1 U21562 ( .A1(n18476), .A2(n19131), .ZN(n18543) );
  NOR2_X1 U21563 ( .A1(n18549), .A2(n18533), .ZN(n18541) );
  AOI211_X1 U21564 ( .C1(n18534), .C2(n18560), .A(n18561), .B(n18549), .ZN(
        n18535) );
  OAI21_X1 U21565 ( .B1(n18537), .B2(n18536), .A(n18535), .ZN(n18553) );
  AOI21_X1 U21566 ( .B1(n18538), .B2(n18553), .A(n18584), .ZN(n18539) );
  INV_X1 U21567 ( .A(n18539), .ZN(n18540) );
  MUX2_X1 U21568 ( .A(n18541), .B(n18540), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n18542) );
  AOI211_X1 U21569 ( .C1(n18544), .C2(n18592), .A(n18543), .B(n18542), .ZN(
        n18545) );
  OAI21_X1 U21570 ( .B1(n18546), .B2(n18572), .A(n18545), .ZN(P3_U2858) );
  INV_X1 U21571 ( .A(n18547), .ZN(n18551) );
  OAI22_X1 U21572 ( .A1(n18549), .A2(n18575), .B1(n18572), .B2(n18548), .ZN(
        n18550) );
  AOI211_X1 U21573 ( .C1(n18552), .C2(n18592), .A(n18551), .B(n18550), .ZN(
        n18556) );
  OAI211_X1 U21574 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18554), .A(
        n18586), .B(n18553), .ZN(n18555) );
  NAND2_X1 U21575 ( .A1(n18556), .A2(n18555), .ZN(P3_U2859) );
  AOI21_X1 U21576 ( .B1(n18584), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18557), .ZN(n18570) );
  NOR2_X1 U21577 ( .A1(n20997), .A2(n19211), .ZN(n18558) );
  OAI221_X1 U21578 ( .B1(n18559), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18559), .C2(n18558), .A(n19066), .ZN(n18566) );
  OAI211_X1 U21579 ( .C1(n18561), .C2(n19211), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n18560), .ZN(n18565) );
  NAND3_X1 U21580 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18563), .A3(
        n18562), .ZN(n18564) );
  NAND3_X1 U21581 ( .A1(n18566), .A2(n18565), .A3(n18564), .ZN(n18568) );
  AOI22_X1 U21582 ( .A1(n18586), .A2(n18568), .B1(n18592), .B2(n18567), .ZN(
        n18569) );
  OAI211_X1 U21583 ( .C1(n18572), .C2(n18571), .A(n18570), .B(n18569), .ZN(
        P3_U2860) );
  INV_X1 U21584 ( .A(n18573), .ZN(n18583) );
  NAND3_X1 U21585 ( .A1(n18586), .A2(n20997), .A3(n18574), .ZN(n18593) );
  AOI21_X1 U21586 ( .B1(n18575), .B2(n18593), .A(n19211), .ZN(n18578) );
  AOI211_X1 U21587 ( .C1(n19070), .C2(n20997), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18576), .ZN(n18577) );
  AOI211_X1 U21588 ( .C1(n18590), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        n18581) );
  NAND2_X1 U21589 ( .A1(n18481), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18580) );
  OAI211_X1 U21590 ( .C1(n18583), .C2(n18582), .A(n18581), .B(n18580), .ZN(
        P3_U2861) );
  AOI21_X1 U21591 ( .B1(n18586), .B2(n18585), .A(n18584), .ZN(n18595) );
  INV_X1 U21592 ( .A(n18587), .ZN(n18588) );
  AOI221_X1 U21593 ( .B1(n18592), .B2(n18591), .C1(n18590), .C2(n18589), .A(
        n18588), .ZN(n18594) );
  OAI211_X1 U21594 ( .C1(n18595), .C2(n20997), .A(n18594), .B(n18593), .ZN(
        P3_U2862) );
  AOI21_X1 U21595 ( .B1(n18598), .B2(n18597), .A(n18596), .ZN(n19095) );
  OAI21_X1 U21596 ( .B1(n19095), .B2(n18643), .A(n18604), .ZN(n18599) );
  OAI221_X1 U21597 ( .B1(n18841), .B2(n18600), .C1(n18841), .C2(n18604), .A(
        n18599), .ZN(P3_U2863) );
  NAND2_X1 U21598 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19082), .ZN(
        n18772) );
  INV_X1 U21599 ( .A(n18772), .ZN(n18773) );
  NAND2_X1 U21600 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19079), .ZN(
        n18867) );
  INV_X1 U21601 ( .A(n18867), .ZN(n18866) );
  NOR2_X1 U21602 ( .A1(n18773), .A2(n18866), .ZN(n18602) );
  OAI22_X1 U21603 ( .A1(n18603), .A2(n19082), .B1(n18602), .B2(n18601), .ZN(
        P3_U2866) );
  INV_X1 U21604 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19083) );
  NOR2_X1 U21605 ( .A1(n19083), .A2(n18604), .ZN(P3_U2867) );
  NOR2_X1 U21606 ( .A1(n19079), .A2(n19082), .ZN(n18917) );
  INV_X1 U21607 ( .A(n18917), .ZN(n18915) );
  NAND2_X1 U21608 ( .A1(n19074), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18819) );
  NOR2_X2 U21609 ( .A1(n18915), .A2(n18819), .ZN(n19014) );
  INV_X1 U21610 ( .A(n19014), .ZN(n19036) );
  NAND2_X1 U21611 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18982), .ZN(n18951) );
  NOR2_X1 U21612 ( .A1(n19082), .A2(n18749), .ZN(n18980) );
  NAND2_X1 U21613 ( .A1(n18841), .A2(n18980), .ZN(n18954) );
  INV_X1 U21614 ( .A(n18954), .ZN(n18970) );
  AND2_X1 U21615 ( .A1(n18982), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18978) );
  AND2_X1 U21616 ( .A1(n18947), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18977) );
  INV_X1 U21617 ( .A(n18976), .ZN(n19100) );
  NAND2_X1 U21618 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19073) );
  NOR2_X2 U21619 ( .A1(n19073), .A2(n18915), .ZN(n19031) );
  NAND2_X1 U21620 ( .A1(n19074), .A2(n18841), .ZN(n19075) );
  NAND2_X1 U21621 ( .A1(n19079), .A2(n19082), .ZN(n18683) );
  NOR2_X2 U21622 ( .A1(n19075), .A2(n18683), .ZN(n18702) );
  NOR2_X1 U21623 ( .A1(n19031), .A2(n18702), .ZN(n18663) );
  NOR2_X1 U21624 ( .A1(n19100), .A2(n18663), .ZN(n18637) );
  AOI22_X1 U21625 ( .A1(n18970), .A2(n18978), .B1(n18977), .B2(n18637), .ZN(
        n18611) );
  AOI21_X1 U21626 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18663), .ZN(n18605) );
  NAND2_X1 U21627 ( .A1(n19036), .A2(n18954), .ZN(n18942) );
  AOI22_X1 U21628 ( .A1(n18947), .A2(n18605), .B1(n18982), .B2(n18942), .ZN(
        n18640) );
  INV_X1 U21629 ( .A(n18606), .ZN(n18607) );
  NAND2_X1 U21630 ( .A1(n18608), .A2(n18607), .ZN(n18638) );
  NOR2_X1 U21631 ( .A1(n18609), .A2(n18638), .ZN(n18948) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n18948), .ZN(n18610) );
  OAI211_X1 U21633 ( .C1(n19036), .C2(n18951), .A(n18611), .B(n18610), .ZN(
        P3_U2868) );
  NAND2_X1 U21634 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18982), .ZN(n18895) );
  AND2_X1 U21635 ( .A1(n18982), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18988) );
  NOR2_X2 U21636 ( .A1(n18842), .A2(n18612), .ZN(n18987) );
  AOI22_X1 U21637 ( .A1(n18970), .A2(n18988), .B1(n18637), .B2(n18987), .ZN(
        n18615) );
  NOR2_X1 U21638 ( .A1(n18613), .A2(n18638), .ZN(n18892) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n18892), .ZN(n18614) );
  OAI211_X1 U21640 ( .C1(n19036), .C2(n18895), .A(n18615), .B(n18614), .ZN(
        P3_U2869) );
  NAND2_X1 U21641 ( .A1(n18982), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18899) );
  NAND2_X1 U21642 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18982), .ZN(n18999) );
  INV_X1 U21643 ( .A(n18999), .ZN(n18896) );
  NOR2_X2 U21644 ( .A1(n18842), .A2(n18616), .ZN(n18994) );
  AOI22_X1 U21645 ( .A1(n19014), .A2(n18896), .B1(n18637), .B2(n18994), .ZN(
        n18619) );
  NOR2_X2 U21646 ( .A1(n18617), .A2(n18638), .ZN(n18996) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n18996), .ZN(n18618) );
  OAI211_X1 U21648 ( .C1(n18954), .C2(n18899), .A(n18619), .B(n18618), .ZN(
        P3_U2870) );
  NAND2_X1 U21649 ( .A1(n18982), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18929) );
  NAND2_X1 U21650 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18982), .ZN(n19005) );
  INV_X1 U21651 ( .A(n19005), .ZN(n18926) );
  NOR2_X2 U21652 ( .A1(n18842), .A2(n18620), .ZN(n19000) );
  AOI22_X1 U21653 ( .A1(n19014), .A2(n18926), .B1(n18637), .B2(n19000), .ZN(
        n18623) );
  NOR2_X2 U21654 ( .A1(n18621), .A2(n18638), .ZN(n19002) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n19002), .ZN(n18622) );
  OAI211_X1 U21656 ( .C1(n18954), .C2(n18929), .A(n18623), .B(n18622), .ZN(
        P3_U2871) );
  NAND2_X1 U21657 ( .A1(n18982), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18962) );
  NOR2_X1 U21658 ( .A1(n19573), .A2(n18843), .ZN(n18959) );
  NOR2_X2 U21659 ( .A1(n18842), .A2(n18624), .ZN(n19006) );
  AOI22_X1 U21660 ( .A1(n19014), .A2(n18959), .B1(n18637), .B2(n19006), .ZN(
        n18627) );
  NOR2_X2 U21661 ( .A1(n18625), .A2(n18638), .ZN(n19008) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n19008), .ZN(n18626) );
  OAI211_X1 U21663 ( .C1(n18954), .C2(n18962), .A(n18627), .B(n18626), .ZN(
        P3_U2872) );
  NAND2_X1 U21664 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18982), .ZN(n19019) );
  NAND2_X1 U21665 ( .A1(n18982), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18935) );
  INV_X1 U21666 ( .A(n18935), .ZN(n19013) );
  NOR2_X2 U21667 ( .A1(n18842), .A2(n18628), .ZN(n19012) );
  AOI22_X1 U21668 ( .A1(n18970), .A2(n19013), .B1(n18637), .B2(n19012), .ZN(
        n18631) );
  NOR2_X2 U21669 ( .A1(n18629), .A2(n18638), .ZN(n19015) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n19015), .ZN(n18630) );
  OAI211_X1 U21671 ( .C1(n19036), .C2(n19019), .A(n18631), .B(n18630), .ZN(
        P3_U2873) );
  NAND2_X1 U21672 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18982), .ZN(n19025) );
  NAND2_X1 U21673 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18982), .ZN(n18813) );
  INV_X1 U21674 ( .A(n18813), .ZN(n19021) );
  NOR2_X2 U21675 ( .A1(n18632), .A2(n18842), .ZN(n19020) );
  AOI22_X1 U21676 ( .A1(n19014), .A2(n19021), .B1(n18637), .B2(n19020), .ZN(
        n18635) );
  NOR2_X2 U21677 ( .A1(n18633), .A2(n18638), .ZN(n19022) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n19022), .ZN(n18634) );
  OAI211_X1 U21679 ( .C1(n18954), .C2(n19025), .A(n18635), .B(n18634), .ZN(
        P3_U2874) );
  NAND2_X1 U21680 ( .A1(n18982), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18975) );
  NAND2_X1 U21681 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18982), .ZN(n19035) );
  INV_X1 U21682 ( .A(n19035), .ZN(n18969) );
  NOR2_X2 U21683 ( .A1(n18636), .A2(n18842), .ZN(n19027) );
  AOI22_X1 U21684 ( .A1(n18970), .A2(n18969), .B1(n18637), .B2(n19027), .ZN(
        n18642) );
  NOR2_X2 U21685 ( .A1(n18639), .A2(n18638), .ZN(n19030) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18640), .B1(
        n18702), .B2(n19030), .ZN(n18641) );
  OAI211_X1 U21687 ( .C1(n19036), .C2(n18975), .A(n18642), .B(n18641), .ZN(
        P3_U2875) );
  NAND2_X1 U21688 ( .A1(n19074), .A2(n18976), .ZN(n18914) );
  NOR2_X1 U21689 ( .A1(n18683), .A2(n18914), .ZN(n18658) );
  AOI22_X1 U21690 ( .A1(n19031), .A2(n18978), .B1(n18977), .B2(n18658), .ZN(
        n18645) );
  INV_X1 U21691 ( .A(n18683), .ZN(n18685) );
  NOR2_X1 U21692 ( .A1(n18842), .A2(n18643), .ZN(n18979) );
  INV_X1 U21693 ( .A(n18979), .ZN(n18684) );
  NOR2_X1 U21694 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18684), .ZN(
        n18916) );
  AOI22_X1 U21695 ( .A1(n18982), .A2(n18980), .B1(n18685), .B2(n18916), .ZN(
        n18659) );
  NOR2_X2 U21696 ( .A1(n18819), .A2(n18683), .ZN(n18712) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18659), .B1(
        n18948), .B2(n18712), .ZN(n18644) );
  OAI211_X1 U21698 ( .C1(n18951), .C2(n18954), .A(n18645), .B(n18644), .ZN(
        P3_U2876) );
  INV_X1 U21699 ( .A(n18895), .ZN(n18989) );
  AOI22_X1 U21700 ( .A1(n18970), .A2(n18989), .B1(n18987), .B2(n18658), .ZN(
        n18647) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18659), .B1(
        n19031), .B2(n18988), .ZN(n18646) );
  OAI211_X1 U21702 ( .C1(n18992), .C2(n18727), .A(n18647), .B(n18646), .ZN(
        P3_U2877) );
  INV_X1 U21703 ( .A(n18899), .ZN(n18995) );
  AOI22_X1 U21704 ( .A1(n19031), .A2(n18995), .B1(n18994), .B2(n18658), .ZN(
        n18649) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18659), .B1(
        n18996), .B2(n18712), .ZN(n18648) );
  OAI211_X1 U21706 ( .C1(n18954), .C2(n18999), .A(n18649), .B(n18648), .ZN(
        P3_U2878) );
  INV_X1 U21707 ( .A(n19031), .ZN(n18993) );
  AOI22_X1 U21708 ( .A1(n18970), .A2(n18926), .B1(n19000), .B2(n18658), .ZN(
        n18651) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18659), .B1(
        n19002), .B2(n18712), .ZN(n18650) );
  OAI211_X1 U21710 ( .C1(n18993), .C2(n18929), .A(n18651), .B(n18650), .ZN(
        P3_U2879) );
  INV_X1 U21711 ( .A(n18959), .ZN(n19011) );
  INV_X1 U21712 ( .A(n18962), .ZN(n19007) );
  AOI22_X1 U21713 ( .A1(n19031), .A2(n19007), .B1(n19006), .B2(n18658), .ZN(
        n18653) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18659), .B1(
        n19008), .B2(n18712), .ZN(n18652) );
  OAI211_X1 U21715 ( .C1(n18954), .C2(n19011), .A(n18653), .B(n18652), .ZN(
        P3_U2880) );
  INV_X1 U21716 ( .A(n19019), .ZN(n18932) );
  AOI22_X1 U21717 ( .A1(n18970), .A2(n18932), .B1(n19012), .B2(n18658), .ZN(
        n18655) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18659), .B1(
        n19015), .B2(n18712), .ZN(n18654) );
  OAI211_X1 U21719 ( .C1(n18993), .C2(n18935), .A(n18655), .B(n18654), .ZN(
        P3_U2881) );
  AOI22_X1 U21720 ( .A1(n18970), .A2(n19021), .B1(n19020), .B2(n18658), .ZN(
        n18657) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18659), .B1(
        n19022), .B2(n18712), .ZN(n18656) );
  OAI211_X1 U21722 ( .C1(n18993), .C2(n19025), .A(n18657), .B(n18656), .ZN(
        P3_U2882) );
  INV_X1 U21723 ( .A(n18975), .ZN(n19029) );
  AOI22_X1 U21724 ( .A1(n18970), .A2(n19029), .B1(n19027), .B2(n18658), .ZN(
        n18661) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18659), .B1(
        n19030), .B2(n18712), .ZN(n18660) );
  OAI211_X1 U21726 ( .C1(n18993), .C2(n19035), .A(n18661), .B(n18660), .ZN(
        P3_U2883) );
  INV_X1 U21727 ( .A(n18948), .ZN(n18986) );
  NOR2_X1 U21728 ( .A1(n19074), .A2(n18683), .ZN(n18728) );
  NAND2_X1 U21729 ( .A1(n18728), .A2(n18841), .ZN(n18739) );
  INV_X1 U21730 ( .A(n18951), .ZN(n18983) );
  AOI21_X1 U21731 ( .B1(n18727), .B2(n18739), .A(n19100), .ZN(n18679) );
  AOI22_X1 U21732 ( .A1(n18983), .A2(n19031), .B1(n18977), .B2(n18679), .ZN(
        n18666) );
  INV_X1 U21733 ( .A(n18662), .ZN(n18944) );
  AOI221_X1 U21734 ( .B1(n18663), .B2(n18727), .C1(n18944), .C2(n18727), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18664) );
  OAI21_X1 U21735 ( .B1(n18745), .B2(n18664), .A(n18947), .ZN(n18680) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18680), .B1(
        n18702), .B2(n18978), .ZN(n18665) );
  OAI211_X1 U21737 ( .C1(n18986), .C2(n18739), .A(n18666), .B(n18665), .ZN(
        P3_U2884) );
  AOI22_X1 U21738 ( .A1(n19031), .A2(n18989), .B1(n18987), .B2(n18679), .ZN(
        n18668) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18680), .B1(
        n18702), .B2(n18988), .ZN(n18667) );
  OAI211_X1 U21740 ( .C1(n18992), .C2(n18739), .A(n18668), .B(n18667), .ZN(
        P3_U2885) );
  INV_X1 U21741 ( .A(n18702), .ZN(n18700) );
  AOI22_X1 U21742 ( .A1(n19031), .A2(n18896), .B1(n18994), .B2(n18679), .ZN(
        n18670) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18680), .B1(
        n18996), .B2(n18745), .ZN(n18669) );
  OAI211_X1 U21744 ( .C1(n18700), .C2(n18899), .A(n18670), .B(n18669), .ZN(
        P3_U2886) );
  AOI22_X1 U21745 ( .A1(n19031), .A2(n18926), .B1(n19000), .B2(n18679), .ZN(
        n18672) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18680), .B1(
        n19002), .B2(n18745), .ZN(n18671) );
  OAI211_X1 U21747 ( .C1(n18700), .C2(n18929), .A(n18672), .B(n18671), .ZN(
        P3_U2887) );
  AOI22_X1 U21748 ( .A1(n19031), .A2(n18959), .B1(n19006), .B2(n18679), .ZN(
        n18674) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18680), .B1(
        n19008), .B2(n18745), .ZN(n18673) );
  OAI211_X1 U21750 ( .C1(n18700), .C2(n18962), .A(n18674), .B(n18673), .ZN(
        P3_U2888) );
  AOI22_X1 U21751 ( .A1(n19031), .A2(n18932), .B1(n19012), .B2(n18679), .ZN(
        n18676) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18680), .B1(
        n19015), .B2(n18745), .ZN(n18675) );
  OAI211_X1 U21753 ( .C1(n18700), .C2(n18935), .A(n18676), .B(n18675), .ZN(
        P3_U2889) );
  INV_X1 U21754 ( .A(n19025), .ZN(n18809) );
  AOI22_X1 U21755 ( .A1(n18702), .A2(n18809), .B1(n19020), .B2(n18679), .ZN(
        n18678) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18680), .B1(
        n19022), .B2(n18745), .ZN(n18677) );
  OAI211_X1 U21757 ( .C1(n18993), .C2(n18813), .A(n18678), .B(n18677), .ZN(
        P3_U2890) );
  AOI22_X1 U21758 ( .A1(n19031), .A2(n19029), .B1(n19027), .B2(n18679), .ZN(
        n18682) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18680), .B1(
        n19030), .B2(n18745), .ZN(n18681) );
  OAI211_X1 U21760 ( .C1(n18700), .C2(n19035), .A(n18682), .B(n18681), .ZN(
        P3_U2891) );
  NOR2_X2 U21761 ( .A1(n19073), .A2(n18683), .ZN(n18768) );
  INV_X1 U21762 ( .A(n18768), .ZN(n18766) );
  AND2_X1 U21763 ( .A1(n18976), .A2(n18728), .ZN(n18701) );
  AOI22_X1 U21764 ( .A1(n18983), .A2(n18702), .B1(n18977), .B2(n18701), .ZN(
        n18687) );
  AOI21_X1 U21765 ( .B1(n19074), .B2(n18944), .A(n18684), .ZN(n18774) );
  NAND2_X1 U21766 ( .A1(n18685), .A2(n18774), .ZN(n18703) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18703), .B1(
        n18978), .B2(n18712), .ZN(n18686) );
  OAI211_X1 U21768 ( .C1(n18986), .C2(n18766), .A(n18687), .B(n18686), .ZN(
        P3_U2892) );
  AOI22_X1 U21769 ( .A1(n18702), .A2(n18989), .B1(n18987), .B2(n18701), .ZN(
        n18689) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18703), .B1(
        n18988), .B2(n18712), .ZN(n18688) );
  OAI211_X1 U21771 ( .C1(n18992), .C2(n18766), .A(n18689), .B(n18688), .ZN(
        P3_U2893) );
  AOI22_X1 U21772 ( .A1(n18702), .A2(n18896), .B1(n18994), .B2(n18701), .ZN(
        n18691) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18703), .B1(
        n18996), .B2(n18768), .ZN(n18690) );
  OAI211_X1 U21774 ( .C1(n18899), .C2(n18727), .A(n18691), .B(n18690), .ZN(
        P3_U2894) );
  AOI22_X1 U21775 ( .A1(n18702), .A2(n18926), .B1(n19000), .B2(n18701), .ZN(
        n18693) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18703), .B1(
        n19002), .B2(n18768), .ZN(n18692) );
  OAI211_X1 U21777 ( .C1(n18929), .C2(n18727), .A(n18693), .B(n18692), .ZN(
        P3_U2895) );
  AOI22_X1 U21778 ( .A1(n19007), .A2(n18712), .B1(n19006), .B2(n18701), .ZN(
        n18695) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18703), .B1(
        n19008), .B2(n18768), .ZN(n18694) );
  OAI211_X1 U21780 ( .C1(n18700), .C2(n19011), .A(n18695), .B(n18694), .ZN(
        P3_U2896) );
  AOI22_X1 U21781 ( .A1(n19012), .A2(n18701), .B1(n19013), .B2(n18712), .ZN(
        n18697) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18703), .B1(
        n19015), .B2(n18768), .ZN(n18696) );
  OAI211_X1 U21783 ( .C1(n18700), .C2(n19019), .A(n18697), .B(n18696), .ZN(
        P3_U2897) );
  AOI22_X1 U21784 ( .A1(n18809), .A2(n18712), .B1(n19020), .B2(n18701), .ZN(
        n18699) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18703), .B1(
        n19022), .B2(n18768), .ZN(n18698) );
  OAI211_X1 U21786 ( .C1(n18700), .C2(n18813), .A(n18699), .B(n18698), .ZN(
        P3_U2898) );
  AOI22_X1 U21787 ( .A1(n18702), .A2(n19029), .B1(n19027), .B2(n18701), .ZN(
        n18705) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18703), .B1(
        n19030), .B2(n18768), .ZN(n18704) );
  OAI211_X1 U21789 ( .C1(n19035), .C2(n18727), .A(n18705), .B(n18704), .ZN(
        P3_U2899) );
  NOR2_X1 U21790 ( .A1(n18768), .A2(n9655), .ZN(n18750) );
  NOR2_X1 U21791 ( .A1(n19100), .A2(n18750), .ZN(n18723) );
  AOI22_X1 U21792 ( .A1(n18977), .A2(n18723), .B1(n18978), .B2(n18745), .ZN(
        n18709) );
  NOR2_X1 U21793 ( .A1(n18712), .A2(n18745), .ZN(n18706) );
  OAI21_X1 U21794 ( .B1(n18706), .B2(n18944), .A(n18750), .ZN(n18707) );
  OAI211_X1 U21795 ( .C1(n9655), .C2(n19202), .A(n18947), .B(n18707), .ZN(
        n18724) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18724), .B1(
        n18948), .B2(n9655), .ZN(n18708) );
  OAI211_X1 U21797 ( .C1(n18951), .C2(n18727), .A(n18709), .B(n18708), .ZN(
        P3_U2900) );
  AOI22_X1 U21798 ( .A1(n18988), .A2(n18745), .B1(n18987), .B2(n18723), .ZN(
        n18711) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18724), .B1(
        n18892), .B2(n9655), .ZN(n18710) );
  OAI211_X1 U21800 ( .C1(n18895), .C2(n18727), .A(n18711), .B(n18710), .ZN(
        P3_U2901) );
  AOI22_X1 U21801 ( .A1(n18896), .A2(n18712), .B1(n18994), .B2(n18723), .ZN(
        n18714) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18724), .B1(
        n18996), .B2(n9655), .ZN(n18713) );
  OAI211_X1 U21803 ( .C1(n18899), .C2(n18739), .A(n18714), .B(n18713), .ZN(
        P3_U2902) );
  INV_X1 U21804 ( .A(n18929), .ZN(n19001) );
  AOI22_X1 U21805 ( .A1(n19001), .A2(n18745), .B1(n19000), .B2(n18723), .ZN(
        n18716) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18724), .B1(
        n19002), .B2(n9655), .ZN(n18715) );
  OAI211_X1 U21807 ( .C1(n19005), .C2(n18727), .A(n18716), .B(n18715), .ZN(
        P3_U2903) );
  AOI22_X1 U21808 ( .A1(n19007), .A2(n18745), .B1(n19006), .B2(n18723), .ZN(
        n18718) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18724), .B1(
        n19008), .B2(n9655), .ZN(n18717) );
  OAI211_X1 U21810 ( .C1(n19011), .C2(n18727), .A(n18718), .B(n18717), .ZN(
        P3_U2904) );
  AOI22_X1 U21811 ( .A1(n19012), .A2(n18723), .B1(n19013), .B2(n18745), .ZN(
        n18720) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18724), .B1(
        n19015), .B2(n9655), .ZN(n18719) );
  OAI211_X1 U21813 ( .C1(n19019), .C2(n18727), .A(n18720), .B(n18719), .ZN(
        P3_U2905) );
  AOI22_X1 U21814 ( .A1(n18809), .A2(n18745), .B1(n19020), .B2(n18723), .ZN(
        n18722) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18724), .B1(
        n19022), .B2(n9655), .ZN(n18721) );
  OAI211_X1 U21816 ( .C1(n18813), .C2(n18727), .A(n18722), .B(n18721), .ZN(
        P3_U2906) );
  AOI22_X1 U21817 ( .A1(n18969), .A2(n18745), .B1(n19027), .B2(n18723), .ZN(
        n18726) );
  AOI22_X1 U21818 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18724), .B1(
        n19030), .B2(n9655), .ZN(n18725) );
  OAI211_X1 U21819 ( .C1(n18975), .C2(n18727), .A(n18726), .B(n18725), .ZN(
        P3_U2907) );
  NOR2_X2 U21820 ( .A1(n18819), .A2(n18772), .ZN(n18815) );
  INV_X1 U21821 ( .A(n18815), .ZN(n18812) );
  NOR2_X1 U21822 ( .A1(n18914), .A2(n18772), .ZN(n18744) );
  AOI22_X1 U21823 ( .A1(n18983), .A2(n18745), .B1(n18977), .B2(n18744), .ZN(
        n18730) );
  AOI22_X1 U21824 ( .A1(n18982), .A2(n18728), .B1(n18916), .B2(n18773), .ZN(
        n18746) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18746), .B1(
        n18978), .B2(n18768), .ZN(n18729) );
  OAI211_X1 U21826 ( .C1(n18986), .C2(n18812), .A(n18730), .B(n18729), .ZN(
        P3_U2908) );
  AOI22_X1 U21827 ( .A1(n18989), .A2(n18745), .B1(n18987), .B2(n18744), .ZN(
        n18732) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18746), .B1(
        n18988), .B2(n18768), .ZN(n18731) );
  OAI211_X1 U21829 ( .C1(n18992), .C2(n18812), .A(n18732), .B(n18731), .ZN(
        P3_U2909) );
  AOI22_X1 U21830 ( .A1(n18896), .A2(n18745), .B1(n18994), .B2(n18744), .ZN(
        n18734) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18746), .B1(
        n18996), .B2(n18815), .ZN(n18733) );
  OAI211_X1 U21832 ( .C1(n18899), .C2(n18766), .A(n18734), .B(n18733), .ZN(
        P3_U2910) );
  AOI22_X1 U21833 ( .A1(n19001), .A2(n18768), .B1(n19000), .B2(n18744), .ZN(
        n18736) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18746), .B1(
        n19002), .B2(n18815), .ZN(n18735) );
  OAI211_X1 U21835 ( .C1(n19005), .C2(n18739), .A(n18736), .B(n18735), .ZN(
        P3_U2911) );
  AOI22_X1 U21836 ( .A1(n19007), .A2(n18768), .B1(n19006), .B2(n18744), .ZN(
        n18738) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18746), .B1(
        n19008), .B2(n18815), .ZN(n18737) );
  OAI211_X1 U21838 ( .C1(n19011), .C2(n18739), .A(n18738), .B(n18737), .ZN(
        P3_U2912) );
  AOI22_X1 U21839 ( .A1(n18932), .A2(n18745), .B1(n19012), .B2(n18744), .ZN(
        n18741) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18746), .B1(
        n19015), .B2(n18815), .ZN(n18740) );
  OAI211_X1 U21841 ( .C1(n18935), .C2(n18766), .A(n18741), .B(n18740), .ZN(
        P3_U2913) );
  AOI22_X1 U21842 ( .A1(n19021), .A2(n18745), .B1(n19020), .B2(n18744), .ZN(
        n18743) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18746), .B1(
        n19022), .B2(n18815), .ZN(n18742) );
  OAI211_X1 U21844 ( .C1(n19025), .C2(n18766), .A(n18743), .B(n18742), .ZN(
        P3_U2914) );
  AOI22_X1 U21845 ( .A1(n19029), .A2(n18745), .B1(n19027), .B2(n18744), .ZN(
        n18748) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18746), .B1(
        n19030), .B2(n18815), .ZN(n18747) );
  OAI211_X1 U21847 ( .C1(n19035), .C2(n18766), .A(n18748), .B(n18747), .ZN(
        P3_U2915) );
  NOR2_X1 U21848 ( .A1(n18749), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18820) );
  NAND2_X1 U21849 ( .A1(n18841), .A2(n18820), .ZN(n18840) );
  NOR2_X1 U21850 ( .A1(n18815), .A2(n18833), .ZN(n18795) );
  NOR2_X1 U21851 ( .A1(n19100), .A2(n18795), .ZN(n18767) );
  AOI22_X1 U21852 ( .A1(n18977), .A2(n18767), .B1(n18978), .B2(n9655), .ZN(
        n18753) );
  OAI21_X1 U21853 ( .B1(n18750), .B2(n18944), .A(n18795), .ZN(n18751) );
  OAI211_X1 U21854 ( .C1(n18833), .C2(n19202), .A(n18947), .B(n18751), .ZN(
        n18769) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18769), .B1(
        n18948), .B2(n18833), .ZN(n18752) );
  OAI211_X1 U21856 ( .C1(n18951), .C2(n18766), .A(n18753), .B(n18752), .ZN(
        P3_U2916) );
  AOI22_X1 U21857 ( .A1(n18989), .A2(n18768), .B1(n18987), .B2(n18767), .ZN(
        n18755) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18769), .B1(
        n18988), .B2(n9655), .ZN(n18754) );
  OAI211_X1 U21859 ( .C1(n18992), .C2(n18840), .A(n18755), .B(n18754), .ZN(
        P3_U2917) );
  INV_X1 U21860 ( .A(n9655), .ZN(n18794) );
  AOI22_X1 U21861 ( .A1(n18896), .A2(n18768), .B1(n18994), .B2(n18767), .ZN(
        n18757) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18769), .B1(
        n18996), .B2(n18833), .ZN(n18756) );
  OAI211_X1 U21863 ( .C1(n18899), .C2(n18794), .A(n18757), .B(n18756), .ZN(
        P3_U2918) );
  AOI22_X1 U21864 ( .A1(n19001), .A2(n9655), .B1(n19000), .B2(n18767), .ZN(
        n18759) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18769), .B1(
        n19002), .B2(n18833), .ZN(n18758) );
  OAI211_X1 U21866 ( .C1(n19005), .C2(n18766), .A(n18759), .B(n18758), .ZN(
        P3_U2919) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18769), .B1(
        n19006), .B2(n18767), .ZN(n18761) );
  AOI22_X1 U21868 ( .A1(n19007), .A2(n9655), .B1(n19008), .B2(n18833), .ZN(
        n18760) );
  OAI211_X1 U21869 ( .C1(n19011), .C2(n18766), .A(n18761), .B(n18760), .ZN(
        P3_U2920) );
  AOI22_X1 U21870 ( .A1(n18932), .A2(n18768), .B1(n19012), .B2(n18767), .ZN(
        n18763) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18769), .B1(
        n19015), .B2(n18833), .ZN(n18762) );
  OAI211_X1 U21872 ( .C1(n18935), .C2(n18794), .A(n18763), .B(n18762), .ZN(
        P3_U2921) );
  AOI22_X1 U21873 ( .A1(n18809), .A2(n9655), .B1(n19020), .B2(n18767), .ZN(
        n18765) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18769), .B1(
        n19022), .B2(n18833), .ZN(n18764) );
  OAI211_X1 U21875 ( .C1(n18813), .C2(n18766), .A(n18765), .B(n18764), .ZN(
        P3_U2922) );
  AOI22_X1 U21876 ( .A1(n19029), .A2(n18768), .B1(n19027), .B2(n18767), .ZN(
        n18771) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18769), .B1(
        n19030), .B2(n18833), .ZN(n18770) );
  OAI211_X1 U21878 ( .C1(n19035), .C2(n18794), .A(n18771), .B(n18770), .ZN(
        P3_U2923) );
  NOR2_X2 U21879 ( .A1(n19073), .A2(n18772), .ZN(n18862) );
  INV_X1 U21880 ( .A(n18862), .ZN(n18858) );
  AND2_X1 U21881 ( .A1(n18976), .A2(n18820), .ZN(n18790) );
  AOI22_X1 U21882 ( .A1(n18977), .A2(n18790), .B1(n18978), .B2(n18815), .ZN(
        n18776) );
  NAND2_X1 U21883 ( .A1(n18774), .A2(n18773), .ZN(n18791) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18791), .B1(
        n18983), .B2(n9655), .ZN(n18775) );
  OAI211_X1 U21885 ( .C1(n18986), .C2(n18858), .A(n18776), .B(n18775), .ZN(
        P3_U2924) );
  AOI22_X1 U21886 ( .A1(n18988), .A2(n18815), .B1(n18987), .B2(n18790), .ZN(
        n18778) );
  AOI22_X1 U21887 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18791), .B1(
        n18989), .B2(n9655), .ZN(n18777) );
  OAI211_X1 U21888 ( .C1(n18992), .C2(n18858), .A(n18778), .B(n18777), .ZN(
        P3_U2925) );
  AOI22_X1 U21889 ( .A1(n18896), .A2(n9655), .B1(n18994), .B2(n18790), .ZN(
        n18780) );
  AOI22_X1 U21890 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18791), .B1(
        n18996), .B2(n18862), .ZN(n18779) );
  OAI211_X1 U21891 ( .C1(n18899), .C2(n18812), .A(n18780), .B(n18779), .ZN(
        P3_U2926) );
  AOI22_X1 U21892 ( .A1(n18926), .A2(n9655), .B1(n19000), .B2(n18790), .ZN(
        n18782) );
  AOI22_X1 U21893 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18791), .B1(
        n19002), .B2(n18862), .ZN(n18781) );
  OAI211_X1 U21894 ( .C1(n18929), .C2(n18812), .A(n18782), .B(n18781), .ZN(
        P3_U2927) );
  AOI22_X1 U21895 ( .A1(n19007), .A2(n18815), .B1(n19006), .B2(n18790), .ZN(
        n18784) );
  AOI22_X1 U21896 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18791), .B1(
        n19008), .B2(n18862), .ZN(n18783) );
  OAI211_X1 U21897 ( .C1(n19011), .C2(n18794), .A(n18784), .B(n18783), .ZN(
        P3_U2928) );
  AOI22_X1 U21898 ( .A1(n18932), .A2(n9655), .B1(n19012), .B2(n18790), .ZN(
        n18787) );
  AOI22_X1 U21899 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18791), .B1(
        n19015), .B2(n18862), .ZN(n18786) );
  OAI211_X1 U21900 ( .C1(n18935), .C2(n18812), .A(n18787), .B(n18786), .ZN(
        P3_U2929) );
  AOI22_X1 U21901 ( .A1(n19021), .A2(n9655), .B1(n19020), .B2(n18790), .ZN(
        n18789) );
  AOI22_X1 U21902 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18791), .B1(
        n19022), .B2(n18862), .ZN(n18788) );
  OAI211_X1 U21903 ( .C1(n19025), .C2(n18812), .A(n18789), .B(n18788), .ZN(
        P3_U2930) );
  AOI22_X1 U21904 ( .A1(n18969), .A2(n18815), .B1(n19027), .B2(n18790), .ZN(
        n18793) );
  AOI22_X1 U21905 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18791), .B1(
        n19030), .B2(n18862), .ZN(n18792) );
  OAI211_X1 U21906 ( .C1(n18975), .C2(n18794), .A(n18793), .B(n18792), .ZN(
        P3_U2931) );
  NOR2_X2 U21907 ( .A1(n19075), .A2(n18867), .ZN(n18884) );
  NOR2_X1 U21908 ( .A1(n18862), .A2(n18884), .ZN(n18844) );
  NOR2_X1 U21909 ( .A1(n19100), .A2(n18844), .ZN(n18814) );
  AOI22_X1 U21910 ( .A1(n18977), .A2(n18814), .B1(n18978), .B2(n18833), .ZN(
        n18798) );
  OAI21_X1 U21911 ( .B1(n18795), .B2(n18944), .A(n18844), .ZN(n18796) );
  OAI211_X1 U21912 ( .C1(n18884), .C2(n19202), .A(n18947), .B(n18796), .ZN(
        n18816) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18816), .B1(
        n18948), .B2(n18884), .ZN(n18797) );
  OAI211_X1 U21914 ( .C1(n18951), .C2(n18812), .A(n18798), .B(n18797), .ZN(
        P3_U2932) );
  INV_X1 U21915 ( .A(n18884), .ZN(n18876) );
  AOI22_X1 U21916 ( .A1(n18989), .A2(n18815), .B1(n18987), .B2(n18814), .ZN(
        n18800) );
  AOI22_X1 U21917 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18816), .B1(
        n18988), .B2(n18833), .ZN(n18799) );
  OAI211_X1 U21918 ( .C1(n18992), .C2(n18876), .A(n18800), .B(n18799), .ZN(
        P3_U2933) );
  AOI22_X1 U21919 ( .A1(n18995), .A2(n18833), .B1(n18994), .B2(n18814), .ZN(
        n18802) );
  AOI22_X1 U21920 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18816), .B1(
        n18996), .B2(n18884), .ZN(n18801) );
  OAI211_X1 U21921 ( .C1(n18999), .C2(n18812), .A(n18802), .B(n18801), .ZN(
        P3_U2934) );
  AOI22_X1 U21922 ( .A1(n19001), .A2(n18833), .B1(n19000), .B2(n18814), .ZN(
        n18804) );
  AOI22_X1 U21923 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18816), .B1(
        n19002), .B2(n18884), .ZN(n18803) );
  OAI211_X1 U21924 ( .C1(n19005), .C2(n18812), .A(n18804), .B(n18803), .ZN(
        P3_U2935) );
  AOI22_X1 U21925 ( .A1(n18959), .A2(n18815), .B1(n19006), .B2(n18814), .ZN(
        n18806) );
  AOI22_X1 U21926 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18816), .B1(
        n19008), .B2(n18884), .ZN(n18805) );
  OAI211_X1 U21927 ( .C1(n18962), .C2(n18840), .A(n18806), .B(n18805), .ZN(
        P3_U2936) );
  AOI22_X1 U21928 ( .A1(n19012), .A2(n18814), .B1(n19013), .B2(n18833), .ZN(
        n18808) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18816), .B1(
        n19015), .B2(n18884), .ZN(n18807) );
  OAI211_X1 U21930 ( .C1(n19019), .C2(n18812), .A(n18808), .B(n18807), .ZN(
        P3_U2937) );
  AOI22_X1 U21931 ( .A1(n18809), .A2(n18833), .B1(n19020), .B2(n18814), .ZN(
        n18811) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18816), .B1(
        n19022), .B2(n18884), .ZN(n18810) );
  OAI211_X1 U21933 ( .C1(n18813), .C2(n18812), .A(n18811), .B(n18810), .ZN(
        P3_U2938) );
  AOI22_X1 U21934 ( .A1(n19029), .A2(n18815), .B1(n19027), .B2(n18814), .ZN(
        n18818) );
  AOI22_X1 U21935 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18816), .B1(
        n19030), .B2(n18884), .ZN(n18817) );
  OAI211_X1 U21936 ( .C1(n19035), .C2(n18840), .A(n18818), .B(n18817), .ZN(
        P3_U2939) );
  NOR2_X2 U21937 ( .A1(n18819), .A2(n18867), .ZN(n18906) );
  INV_X1 U21938 ( .A(n18906), .ZN(n18913) );
  NOR2_X1 U21939 ( .A1(n18914), .A2(n18867), .ZN(n18836) );
  AOI22_X1 U21940 ( .A1(n18983), .A2(n18833), .B1(n18977), .B2(n18836), .ZN(
        n18822) );
  AOI22_X1 U21941 ( .A1(n18982), .A2(n18820), .B1(n18916), .B2(n18866), .ZN(
        n18837) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18837), .B1(
        n18978), .B2(n18862), .ZN(n18821) );
  OAI211_X1 U21943 ( .C1(n18986), .C2(n18913), .A(n18822), .B(n18821), .ZN(
        P3_U2940) );
  AOI22_X1 U21944 ( .A1(n18989), .A2(n18833), .B1(n18987), .B2(n18836), .ZN(
        n18824) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18837), .B1(
        n18988), .B2(n18862), .ZN(n18823) );
  OAI211_X1 U21946 ( .C1(n18992), .C2(n18913), .A(n18824), .B(n18823), .ZN(
        P3_U2941) );
  AOI22_X1 U21947 ( .A1(n18995), .A2(n18862), .B1(n18994), .B2(n18836), .ZN(
        n18826) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18837), .B1(
        n18996), .B2(n18906), .ZN(n18825) );
  OAI211_X1 U21949 ( .C1(n18999), .C2(n18840), .A(n18826), .B(n18825), .ZN(
        P3_U2942) );
  AOI22_X1 U21950 ( .A1(n19001), .A2(n18862), .B1(n19000), .B2(n18836), .ZN(
        n18828) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18837), .B1(
        n19002), .B2(n18906), .ZN(n18827) );
  OAI211_X1 U21952 ( .C1(n19005), .C2(n18840), .A(n18828), .B(n18827), .ZN(
        P3_U2943) );
  AOI22_X1 U21953 ( .A1(n18959), .A2(n18833), .B1(n19006), .B2(n18836), .ZN(
        n18830) );
  AOI22_X1 U21954 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18837), .B1(
        n19008), .B2(n18906), .ZN(n18829) );
  OAI211_X1 U21955 ( .C1(n18962), .C2(n18858), .A(n18830), .B(n18829), .ZN(
        P3_U2944) );
  AOI22_X1 U21956 ( .A1(n19012), .A2(n18836), .B1(n19013), .B2(n18862), .ZN(
        n18832) );
  AOI22_X1 U21957 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18837), .B1(
        n19015), .B2(n18906), .ZN(n18831) );
  OAI211_X1 U21958 ( .C1(n19019), .C2(n18840), .A(n18832), .B(n18831), .ZN(
        P3_U2945) );
  AOI22_X1 U21959 ( .A1(n19021), .A2(n18833), .B1(n19020), .B2(n18836), .ZN(
        n18835) );
  AOI22_X1 U21960 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18837), .B1(
        n19022), .B2(n18906), .ZN(n18834) );
  OAI211_X1 U21961 ( .C1(n19025), .C2(n18858), .A(n18835), .B(n18834), .ZN(
        P3_U2946) );
  AOI22_X1 U21962 ( .A1(n18969), .A2(n18862), .B1(n19027), .B2(n18836), .ZN(
        n18839) );
  AOI22_X1 U21963 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18837), .B1(
        n19030), .B2(n18906), .ZN(n18838) );
  OAI211_X1 U21964 ( .C1(n18975), .C2(n18840), .A(n18839), .B(n18838), .ZN(
        P3_U2947) );
  NOR2_X1 U21965 ( .A1(n19074), .A2(n18867), .ZN(n18918) );
  NAND2_X1 U21966 ( .A1(n18841), .A2(n18918), .ZN(n18925) );
  NOR2_X1 U21967 ( .A1(n18906), .A2(n18938), .ZN(n18888) );
  NOR2_X1 U21968 ( .A1(n19100), .A2(n18888), .ZN(n18861) );
  AOI22_X1 U21969 ( .A1(n18977), .A2(n18861), .B1(n18978), .B2(n18884), .ZN(
        n18847) );
  OAI22_X1 U21970 ( .A1(n18844), .A2(n18843), .B1(n18888), .B2(n18842), .ZN(
        n18845) );
  OAI21_X1 U21971 ( .B1(n18938), .B2(n19202), .A(n18845), .ZN(n18863) );
  AOI22_X1 U21972 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18863), .B1(
        n18948), .B2(n18938), .ZN(n18846) );
  OAI211_X1 U21973 ( .C1(n18951), .C2(n18858), .A(n18847), .B(n18846), .ZN(
        P3_U2948) );
  AOI22_X1 U21974 ( .A1(n18988), .A2(n18884), .B1(n18987), .B2(n18861), .ZN(
        n18849) );
  AOI22_X1 U21975 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18863), .B1(
        n18892), .B2(n18938), .ZN(n18848) );
  OAI211_X1 U21976 ( .C1(n18895), .C2(n18858), .A(n18849), .B(n18848), .ZN(
        P3_U2949) );
  AOI22_X1 U21977 ( .A1(n18995), .A2(n18884), .B1(n18994), .B2(n18861), .ZN(
        n18851) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18863), .B1(
        n18996), .B2(n18938), .ZN(n18850) );
  OAI211_X1 U21979 ( .C1(n18999), .C2(n18858), .A(n18851), .B(n18850), .ZN(
        P3_U2950) );
  AOI22_X1 U21980 ( .A1(n18926), .A2(n18862), .B1(n19000), .B2(n18861), .ZN(
        n18853) );
  AOI22_X1 U21981 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18863), .B1(
        n19002), .B2(n18938), .ZN(n18852) );
  OAI211_X1 U21982 ( .C1(n18929), .C2(n18876), .A(n18853), .B(n18852), .ZN(
        P3_U2951) );
  AOI22_X1 U21983 ( .A1(n19007), .A2(n18884), .B1(n19006), .B2(n18861), .ZN(
        n18855) );
  AOI22_X1 U21984 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18863), .B1(
        n19008), .B2(n18938), .ZN(n18854) );
  OAI211_X1 U21985 ( .C1(n19011), .C2(n18858), .A(n18855), .B(n18854), .ZN(
        P3_U2952) );
  AOI22_X1 U21986 ( .A1(n19012), .A2(n18861), .B1(n19013), .B2(n18884), .ZN(
        n18857) );
  AOI22_X1 U21987 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18863), .B1(
        n19015), .B2(n18938), .ZN(n18856) );
  OAI211_X1 U21988 ( .C1(n19019), .C2(n18858), .A(n18857), .B(n18856), .ZN(
        P3_U2953) );
  AOI22_X1 U21989 ( .A1(n19021), .A2(n18862), .B1(n19020), .B2(n18861), .ZN(
        n18860) );
  AOI22_X1 U21990 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18863), .B1(
        n19022), .B2(n18938), .ZN(n18859) );
  OAI211_X1 U21991 ( .C1(n19025), .C2(n18876), .A(n18860), .B(n18859), .ZN(
        P3_U2954) );
  AOI22_X1 U21992 ( .A1(n19029), .A2(n18862), .B1(n19027), .B2(n18861), .ZN(
        n18865) );
  AOI22_X1 U21993 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18863), .B1(
        n19030), .B2(n18938), .ZN(n18864) );
  OAI211_X1 U21994 ( .C1(n19035), .C2(n18876), .A(n18865), .B(n18864), .ZN(
        P3_U2955) );
  AND2_X1 U21995 ( .A1(n18976), .A2(n18918), .ZN(n18883) );
  AOI22_X1 U21996 ( .A1(n18977), .A2(n18883), .B1(n18978), .B2(n18906), .ZN(
        n18869) );
  AOI22_X1 U21997 ( .A1(n18982), .A2(n18866), .B1(n18979), .B2(n18918), .ZN(
        n18885) );
  NOR2_X2 U21998 ( .A1(n19073), .A2(n18867), .ZN(n18965) );
  AOI22_X1 U21999 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18885), .B1(
        n18948), .B2(n18965), .ZN(n18868) );
  OAI211_X1 U22000 ( .C1(n18951), .C2(n18876), .A(n18869), .B(n18868), .ZN(
        P3_U2956) );
  INV_X1 U22001 ( .A(n18965), .ZN(n18974) );
  AOI22_X1 U22002 ( .A1(n18989), .A2(n18884), .B1(n18987), .B2(n18883), .ZN(
        n18871) );
  AOI22_X1 U22003 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18885), .B1(
        n18988), .B2(n18906), .ZN(n18870) );
  OAI211_X1 U22004 ( .C1(n18992), .C2(n18974), .A(n18871), .B(n18870), .ZN(
        P3_U2957) );
  AOI22_X1 U22005 ( .A1(n18896), .A2(n18884), .B1(n18994), .B2(n18883), .ZN(
        n18873) );
  AOI22_X1 U22006 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18885), .B1(
        n18996), .B2(n18965), .ZN(n18872) );
  OAI211_X1 U22007 ( .C1(n18899), .C2(n18913), .A(n18873), .B(n18872), .ZN(
        P3_U2958) );
  AOI22_X1 U22008 ( .A1(n19001), .A2(n18906), .B1(n19000), .B2(n18883), .ZN(
        n18875) );
  AOI22_X1 U22009 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18885), .B1(
        n19002), .B2(n18965), .ZN(n18874) );
  OAI211_X1 U22010 ( .C1(n19005), .C2(n18876), .A(n18875), .B(n18874), .ZN(
        P3_U2959) );
  AOI22_X1 U22011 ( .A1(n18959), .A2(n18884), .B1(n19006), .B2(n18883), .ZN(
        n18878) );
  AOI22_X1 U22012 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18885), .B1(
        n19008), .B2(n18965), .ZN(n18877) );
  OAI211_X1 U22013 ( .C1(n18962), .C2(n18913), .A(n18878), .B(n18877), .ZN(
        P3_U2960) );
  AOI22_X1 U22014 ( .A1(n18932), .A2(n18884), .B1(n19012), .B2(n18883), .ZN(
        n18880) );
  AOI22_X1 U22015 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18885), .B1(
        n19015), .B2(n18965), .ZN(n18879) );
  OAI211_X1 U22016 ( .C1(n18935), .C2(n18913), .A(n18880), .B(n18879), .ZN(
        P3_U2961) );
  AOI22_X1 U22017 ( .A1(n19021), .A2(n18884), .B1(n19020), .B2(n18883), .ZN(
        n18882) );
  AOI22_X1 U22018 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18885), .B1(
        n19022), .B2(n18965), .ZN(n18881) );
  OAI211_X1 U22019 ( .C1(n19025), .C2(n18913), .A(n18882), .B(n18881), .ZN(
        P3_U2962) );
  AOI22_X1 U22020 ( .A1(n19029), .A2(n18884), .B1(n19027), .B2(n18883), .ZN(
        n18887) );
  AOI22_X1 U22021 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18885), .B1(
        n19030), .B2(n18965), .ZN(n18886) );
  OAI211_X1 U22022 ( .C1(n19035), .C2(n18913), .A(n18887), .B(n18886), .ZN(
        P3_U2963) );
  NOR2_X2 U22023 ( .A1(n19075), .A2(n18915), .ZN(n19028) );
  NOR2_X1 U22024 ( .A1(n18965), .A2(n19028), .ZN(n18945) );
  NOR2_X1 U22025 ( .A1(n19100), .A2(n18945), .ZN(n18909) );
  AOI22_X1 U22026 ( .A1(n18977), .A2(n18909), .B1(n18978), .B2(n18938), .ZN(
        n18891) );
  OAI21_X1 U22027 ( .B1(n18888), .B2(n18944), .A(n18945), .ZN(n18889) );
  OAI211_X1 U22028 ( .C1(n19028), .C2(n19202), .A(n18947), .B(n18889), .ZN(
        n18910) );
  AOI22_X1 U22029 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18910), .B1(
        n18948), .B2(n19028), .ZN(n18890) );
  OAI211_X1 U22030 ( .C1(n18951), .C2(n18913), .A(n18891), .B(n18890), .ZN(
        P3_U2964) );
  AOI22_X1 U22031 ( .A1(n18988), .A2(n18938), .B1(n18987), .B2(n18909), .ZN(
        n18894) );
  AOI22_X1 U22032 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18910), .B1(
        n18892), .B2(n19028), .ZN(n18893) );
  OAI211_X1 U22033 ( .C1(n18895), .C2(n18913), .A(n18894), .B(n18893), .ZN(
        P3_U2965) );
  AOI22_X1 U22034 ( .A1(n18896), .A2(n18906), .B1(n18994), .B2(n18909), .ZN(
        n18898) );
  AOI22_X1 U22035 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18910), .B1(
        n18996), .B2(n19028), .ZN(n18897) );
  OAI211_X1 U22036 ( .C1(n18899), .C2(n18925), .A(n18898), .B(n18897), .ZN(
        P3_U2966) );
  AOI22_X1 U22037 ( .A1(n18926), .A2(n18906), .B1(n19000), .B2(n18909), .ZN(
        n18901) );
  AOI22_X1 U22038 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18910), .B1(
        n19002), .B2(n19028), .ZN(n18900) );
  OAI211_X1 U22039 ( .C1(n18929), .C2(n18925), .A(n18901), .B(n18900), .ZN(
        P3_U2967) );
  AOI22_X1 U22040 ( .A1(n19007), .A2(n18938), .B1(n19006), .B2(n18909), .ZN(
        n18903) );
  AOI22_X1 U22041 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18910), .B1(
        n19008), .B2(n19028), .ZN(n18902) );
  OAI211_X1 U22042 ( .C1(n19011), .C2(n18913), .A(n18903), .B(n18902), .ZN(
        P3_U2968) );
  AOI22_X1 U22043 ( .A1(n19012), .A2(n18909), .B1(n19013), .B2(n18938), .ZN(
        n18905) );
  AOI22_X1 U22044 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18910), .B1(
        n19015), .B2(n19028), .ZN(n18904) );
  OAI211_X1 U22045 ( .C1(n19019), .C2(n18913), .A(n18905), .B(n18904), .ZN(
        P3_U2969) );
  AOI22_X1 U22046 ( .A1(n19021), .A2(n18906), .B1(n19020), .B2(n18909), .ZN(
        n18908) );
  AOI22_X1 U22047 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18910), .B1(
        n19022), .B2(n19028), .ZN(n18907) );
  OAI211_X1 U22048 ( .C1(n19025), .C2(n18925), .A(n18908), .B(n18907), .ZN(
        P3_U2970) );
  AOI22_X1 U22049 ( .A1(n18969), .A2(n18938), .B1(n19027), .B2(n18909), .ZN(
        n18912) );
  AOI22_X1 U22050 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18910), .B1(
        n19030), .B2(n19028), .ZN(n18911) );
  OAI211_X1 U22051 ( .C1(n18975), .C2(n18913), .A(n18912), .B(n18911), .ZN(
        P3_U2971) );
  NOR2_X1 U22052 ( .A1(n18915), .A2(n18914), .ZN(n18981) );
  AOI22_X1 U22053 ( .A1(n18977), .A2(n18981), .B1(n18978), .B2(n18965), .ZN(
        n18920) );
  AOI22_X1 U22054 ( .A1(n18982), .A2(n18918), .B1(n18917), .B2(n18916), .ZN(
        n18939) );
  AOI22_X1 U22055 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18939), .B1(
        n19014), .B2(n18948), .ZN(n18919) );
  OAI211_X1 U22056 ( .C1(n18951), .C2(n18925), .A(n18920), .B(n18919), .ZN(
        P3_U2972) );
  AOI22_X1 U22057 ( .A1(n18989), .A2(n18938), .B1(n18987), .B2(n18981), .ZN(
        n18922) );
  AOI22_X1 U22058 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18939), .B1(
        n18988), .B2(n18965), .ZN(n18921) );
  OAI211_X1 U22059 ( .C1(n19036), .C2(n18992), .A(n18922), .B(n18921), .ZN(
        P3_U2973) );
  AOI22_X1 U22060 ( .A1(n18995), .A2(n18965), .B1(n18994), .B2(n18981), .ZN(
        n18924) );
  AOI22_X1 U22061 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18939), .B1(
        n19014), .B2(n18996), .ZN(n18923) );
  OAI211_X1 U22062 ( .C1(n18999), .C2(n18925), .A(n18924), .B(n18923), .ZN(
        P3_U2974) );
  AOI22_X1 U22063 ( .A1(n18926), .A2(n18938), .B1(n19000), .B2(n18981), .ZN(
        n18928) );
  AOI22_X1 U22064 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18939), .B1(
        n19014), .B2(n19002), .ZN(n18927) );
  OAI211_X1 U22065 ( .C1(n18929), .C2(n18974), .A(n18928), .B(n18927), .ZN(
        P3_U2975) );
  AOI22_X1 U22066 ( .A1(n18959), .A2(n18938), .B1(n19006), .B2(n18981), .ZN(
        n18931) );
  AOI22_X1 U22067 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18939), .B1(
        n19014), .B2(n19008), .ZN(n18930) );
  OAI211_X1 U22068 ( .C1(n18962), .C2(n18974), .A(n18931), .B(n18930), .ZN(
        P3_U2976) );
  AOI22_X1 U22069 ( .A1(n18932), .A2(n18938), .B1(n19012), .B2(n18981), .ZN(
        n18934) );
  AOI22_X1 U22070 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18939), .B1(
        n19014), .B2(n19015), .ZN(n18933) );
  OAI211_X1 U22071 ( .C1(n18935), .C2(n18974), .A(n18934), .B(n18933), .ZN(
        P3_U2977) );
  AOI22_X1 U22072 ( .A1(n19021), .A2(n18938), .B1(n19020), .B2(n18981), .ZN(
        n18937) );
  AOI22_X1 U22073 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18939), .B1(
        n19014), .B2(n19022), .ZN(n18936) );
  OAI211_X1 U22074 ( .C1(n19025), .C2(n18974), .A(n18937), .B(n18936), .ZN(
        P3_U2978) );
  AOI22_X1 U22075 ( .A1(n19029), .A2(n18938), .B1(n19027), .B2(n18981), .ZN(
        n18941) );
  AOI22_X1 U22076 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18939), .B1(
        n19014), .B2(n19030), .ZN(n18940) );
  OAI211_X1 U22077 ( .C1(n19035), .C2(n18974), .A(n18941), .B(n18940), .ZN(
        P3_U2979) );
  INV_X1 U22078 ( .A(n18942), .ZN(n18943) );
  NOR2_X1 U22079 ( .A1(n19100), .A2(n18943), .ZN(n18968) );
  AOI22_X1 U22080 ( .A1(n18977), .A2(n18968), .B1(n18978), .B2(n19028), .ZN(
        n18950) );
  OAI21_X1 U22081 ( .B1(n18945), .B2(n18944), .A(n18943), .ZN(n18946) );
  OAI211_X1 U22082 ( .C1(n18970), .C2(n19202), .A(n18947), .B(n18946), .ZN(
        n18971) );
  AOI22_X1 U22083 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18948), .ZN(n18949) );
  OAI211_X1 U22084 ( .C1(n18951), .C2(n18974), .A(n18950), .B(n18949), .ZN(
        P3_U2980) );
  AOI22_X1 U22085 ( .A1(n18989), .A2(n18965), .B1(n18987), .B2(n18968), .ZN(
        n18953) );
  AOI22_X1 U22086 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18971), .B1(
        n18988), .B2(n19028), .ZN(n18952) );
  OAI211_X1 U22087 ( .C1(n18954), .C2(n18992), .A(n18953), .B(n18952), .ZN(
        P3_U2981) );
  AOI22_X1 U22088 ( .A1(n18995), .A2(n19028), .B1(n18994), .B2(n18968), .ZN(
        n18956) );
  AOI22_X1 U22089 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18996), .ZN(n18955) );
  OAI211_X1 U22090 ( .C1(n18999), .C2(n18974), .A(n18956), .B(n18955), .ZN(
        P3_U2982) );
  AOI22_X1 U22091 ( .A1(n19001), .A2(n19028), .B1(n19000), .B2(n18968), .ZN(
        n18958) );
  AOI22_X1 U22092 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n19002), .ZN(n18957) );
  OAI211_X1 U22093 ( .C1(n19005), .C2(n18974), .A(n18958), .B(n18957), .ZN(
        P3_U2983) );
  INV_X1 U22094 ( .A(n19028), .ZN(n19018) );
  AOI22_X1 U22095 ( .A1(n18959), .A2(n18965), .B1(n19006), .B2(n18968), .ZN(
        n18961) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n19008), .ZN(n18960) );
  OAI211_X1 U22097 ( .C1(n18962), .C2(n19018), .A(n18961), .B(n18960), .ZN(
        P3_U2984) );
  AOI22_X1 U22098 ( .A1(n19012), .A2(n18968), .B1(n19013), .B2(n19028), .ZN(
        n18964) );
  AOI22_X1 U22099 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n19015), .ZN(n18963) );
  OAI211_X1 U22100 ( .C1(n19019), .C2(n18974), .A(n18964), .B(n18963), .ZN(
        P3_U2985) );
  AOI22_X1 U22101 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18971), .B1(
        n19020), .B2(n18968), .ZN(n18967) );
  AOI22_X1 U22102 ( .A1(n18970), .A2(n19022), .B1(n19021), .B2(n18965), .ZN(
        n18966) );
  OAI211_X1 U22103 ( .C1(n19025), .C2(n19018), .A(n18967), .B(n18966), .ZN(
        P3_U2986) );
  AOI22_X1 U22104 ( .A1(n18969), .A2(n19028), .B1(n19027), .B2(n18968), .ZN(
        n18973) );
  AOI22_X1 U22105 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n19030), .ZN(n18972) );
  OAI211_X1 U22106 ( .C1(n18975), .C2(n18974), .A(n18973), .B(n18972), .ZN(
        P3_U2987) );
  AND2_X1 U22107 ( .A1(n18976), .A2(n18980), .ZN(n19026) );
  AOI22_X1 U22108 ( .A1(n19014), .A2(n18978), .B1(n18977), .B2(n19026), .ZN(
        n18985) );
  AOI22_X1 U22109 ( .A1(n18982), .A2(n18981), .B1(n18980), .B2(n18979), .ZN(
        n19032) );
  AOI22_X1 U22110 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19032), .B1(
        n18983), .B2(n19028), .ZN(n18984) );
  OAI211_X1 U22111 ( .C1(n18993), .C2(n18986), .A(n18985), .B(n18984), .ZN(
        P3_U2988) );
  AOI22_X1 U22112 ( .A1(n19014), .A2(n18988), .B1(n18987), .B2(n19026), .ZN(
        n18991) );
  AOI22_X1 U22113 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19032), .B1(
        n18989), .B2(n19028), .ZN(n18990) );
  OAI211_X1 U22114 ( .C1(n18993), .C2(n18992), .A(n18991), .B(n18990), .ZN(
        P3_U2989) );
  AOI22_X1 U22115 ( .A1(n19014), .A2(n18995), .B1(n18994), .B2(n19026), .ZN(
        n18998) );
  AOI22_X1 U22116 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19032), .B1(
        n19031), .B2(n18996), .ZN(n18997) );
  OAI211_X1 U22117 ( .C1(n18999), .C2(n19018), .A(n18998), .B(n18997), .ZN(
        P3_U2990) );
  AOI22_X1 U22118 ( .A1(n19014), .A2(n19001), .B1(n19000), .B2(n19026), .ZN(
        n19004) );
  AOI22_X1 U22119 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19032), .B1(
        n19031), .B2(n19002), .ZN(n19003) );
  OAI211_X1 U22120 ( .C1(n19005), .C2(n19018), .A(n19004), .B(n19003), .ZN(
        P3_U2991) );
  AOI22_X1 U22121 ( .A1(n19014), .A2(n19007), .B1(n19006), .B2(n19026), .ZN(
        n19010) );
  AOI22_X1 U22122 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19032), .B1(
        n19031), .B2(n19008), .ZN(n19009) );
  OAI211_X1 U22123 ( .C1(n19011), .C2(n19018), .A(n19010), .B(n19009), .ZN(
        P3_U2992) );
  AOI22_X1 U22124 ( .A1(n19014), .A2(n19013), .B1(n19012), .B2(n19026), .ZN(
        n19017) );
  AOI22_X1 U22125 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19032), .B1(
        n19031), .B2(n19015), .ZN(n19016) );
  OAI211_X1 U22126 ( .C1(n19019), .C2(n19018), .A(n19017), .B(n19016), .ZN(
        P3_U2993) );
  AOI22_X1 U22127 ( .A1(n19021), .A2(n19028), .B1(n19020), .B2(n19026), .ZN(
        n19024) );
  AOI22_X1 U22128 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19032), .B1(
        n19031), .B2(n19022), .ZN(n19023) );
  OAI211_X1 U22129 ( .C1(n19036), .C2(n19025), .A(n19024), .B(n19023), .ZN(
        P3_U2994) );
  AOI22_X1 U22130 ( .A1(n19029), .A2(n19028), .B1(n19027), .B2(n19026), .ZN(
        n19034) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19032), .B1(
        n19031), .B2(n19030), .ZN(n19033) );
  OAI211_X1 U22132 ( .C1(n19036), .C2(n19035), .A(n19034), .B(n19033), .ZN(
        P3_U2995) );
  NOR2_X1 U22133 ( .A1(n19066), .A2(n19037), .ZN(n19039) );
  OAI222_X1 U22134 ( .A1(n19043), .A2(n19042), .B1(n19041), .B2(n19040), .C1(
        n19039), .C2(n19038), .ZN(n19244) );
  OAI21_X1 U22135 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19044), .ZN(n19045) );
  OAI211_X1 U22136 ( .C1(n21004), .C2(n19067), .A(n19046), .B(n19045), .ZN(
        n19088) );
  OAI21_X1 U22137 ( .B1(n9660), .B2(n19232), .A(n19070), .ZN(n19059) );
  AOI22_X1 U22138 ( .A1(n19066), .A2(n19048), .B1(n19060), .B2(n19059), .ZN(
        n19049) );
  NOR2_X1 U22139 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19049), .ZN(
        n19204) );
  INV_X1 U22140 ( .A(n19050), .ZN(n19054) );
  AOI21_X1 U22141 ( .B1(n19053), .B2(n19052), .A(n19051), .ZN(n19062) );
  OAI221_X1 U22142 ( .B1(n19060), .B2(n19055), .C1(n19060), .C2(n19054), .A(
        n19062), .ZN(n19056) );
  AOI22_X1 U22143 ( .A1(n19219), .A2(n19061), .B1(n19057), .B2(n19056), .ZN(
        n19205) );
  AOI21_X1 U22144 ( .B1(n19205), .B2(n19067), .A(n19207), .ZN(n19058) );
  AOI21_X1 U22145 ( .B1(n19067), .B2(n19204), .A(n19058), .ZN(n19086) );
  INV_X1 U22146 ( .A(n19067), .ZN(n19077) );
  INV_X1 U22147 ( .A(n19059), .ZN(n19071) );
  AOI211_X1 U22148 ( .C1(n19219), .C2(n19227), .A(n19071), .B(n19060), .ZN(
        n19065) );
  INV_X1 U22149 ( .A(n19061), .ZN(n19063) );
  NOR3_X1 U22150 ( .A1(n19063), .A2(n19062), .A3(n19219), .ZN(n19064) );
  AOI211_X1 U22151 ( .C1(n19066), .C2(n19213), .A(n19065), .B(n19064), .ZN(
        n19216) );
  AOI22_X1 U22152 ( .A1(n19077), .A2(n19219), .B1(n19216), .B2(n19067), .ZN(
        n19081) );
  NOR2_X1 U22153 ( .A1(n19069), .A2(n19068), .ZN(n19072) );
  AOI22_X1 U22154 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19070), .B1(
        n19072), .B2(n19232), .ZN(n19229) );
  OAI22_X1 U22155 ( .A1(n19072), .A2(n19220), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19071), .ZN(n19225) );
  AOI222_X1 U22156 ( .A1(n19229), .A2(n19225), .B1(n19229), .B2(n19074), .C1(
        n19225), .C2(n19073), .ZN(n19076) );
  OAI21_X1 U22157 ( .B1(n19077), .B2(n19076), .A(n19075), .ZN(n19080) );
  AND2_X1 U22158 ( .A1(n19081), .A2(n19080), .ZN(n19078) );
  OAI221_X1 U22159 ( .B1(n19081), .B2(n19080), .C1(n19079), .C2(n19078), .A(
        n19083), .ZN(n19085) );
  AOI21_X1 U22160 ( .B1(n19083), .B2(n19082), .A(n19081), .ZN(n19084) );
  AOI222_X1 U22161 ( .A1(n19086), .A2(n19085), .B1(n19086), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19085), .C2(n19084), .ZN(
        n19087) );
  NOR4_X1 U22162 ( .A1(n19089), .A2(n19244), .A3(n19088), .A4(n19087), .ZN(
        n19099) );
  OAI211_X1 U22163 ( .C1(n19092), .C2(n19091), .A(n19090), .B(n19099), .ZN(
        n19201) );
  OAI21_X1 U22164 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19093), .A(n19201), 
        .ZN(n19101) );
  AOI221_X1 U22165 ( .B1(n19095), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19101), 
        .C2(P3_STATE2_REG_0__SCAN_IN), .A(n19094), .ZN(n19098) );
  INV_X1 U22166 ( .A(n19228), .ZN(n19214) );
  NAND2_X1 U22167 ( .A1(n19252), .A2(n19096), .ZN(n19104) );
  OAI211_X1 U22168 ( .C1(n19214), .C2(n19248), .A(n19249), .B(n19104), .ZN(
        n19097) );
  OAI211_X1 U22169 ( .C1(n19099), .C2(n19254), .A(n19098), .B(n19097), .ZN(
        P3_U2996) );
  NAND3_X1 U22170 ( .A1(n19252), .A2(n19106), .A3(n19261), .ZN(n19109) );
  OR3_X1 U22171 ( .A1(n19102), .A2(n19101), .A3(n19100), .ZN(n19103) );
  NAND4_X1 U22172 ( .A1(n19105), .A2(n19104), .A3(n19109), .A4(n19103), .ZN(
        P3_U2997) );
  OR3_X1 U22173 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19107), .A3(n19106), 
        .ZN(n19108) );
  AND3_X1 U22174 ( .A1(n19109), .A2(n19200), .A3(n19108), .ZN(P3_U2998) );
  AND2_X1 U22175 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19196), .ZN(
        P3_U2999) );
  AND2_X1 U22176 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19196), .ZN(
        P3_U3000) );
  AND2_X1 U22177 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19196), .ZN(
        P3_U3001) );
  AND2_X1 U22178 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19196), .ZN(
        P3_U3002) );
  AND2_X1 U22179 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19196), .ZN(
        P3_U3003) );
  AND2_X1 U22180 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19196), .ZN(
        P3_U3004) );
  AND2_X1 U22181 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19196), .ZN(
        P3_U3005) );
  AND2_X1 U22182 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19196), .ZN(
        P3_U3006) );
  AND2_X1 U22183 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19196), .ZN(
        P3_U3007) );
  AND2_X1 U22184 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19196), .ZN(
        P3_U3008) );
  AND2_X1 U22185 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19196), .ZN(
        P3_U3009) );
  AND2_X1 U22186 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19196), .ZN(
        P3_U3010) );
  AND2_X1 U22187 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19196), .ZN(
        P3_U3011) );
  AND2_X1 U22188 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19196), .ZN(
        P3_U3012) );
  AND2_X1 U22189 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19196), .ZN(
        P3_U3013) );
  AND2_X1 U22190 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19196), .ZN(
        P3_U3014) );
  AND2_X1 U22191 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19196), .ZN(
        P3_U3015) );
  AND2_X1 U22192 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19196), .ZN(
        P3_U3016) );
  AND2_X1 U22193 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19196), .ZN(
        P3_U3017) );
  AND2_X1 U22194 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19196), .ZN(
        P3_U3018) );
  AND2_X1 U22195 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19196), .ZN(
        P3_U3019) );
  AND2_X1 U22196 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19196), .ZN(
        P3_U3020) );
  AND2_X1 U22197 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19196), .ZN(P3_U3021) );
  AND2_X1 U22198 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19196), .ZN(P3_U3022) );
  AND2_X1 U22199 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19196), .ZN(P3_U3023) );
  AND2_X1 U22200 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19196), .ZN(P3_U3024) );
  AND2_X1 U22201 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19196), .ZN(P3_U3025) );
  AND2_X1 U22202 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19196), .ZN(P3_U3026) );
  AND2_X1 U22203 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19196), .ZN(P3_U3027) );
  AND2_X1 U22204 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19196), .ZN(P3_U3028) );
  NOR2_X1 U22205 ( .A1(n19110), .A2(n20769), .ZN(n19114) );
  NAND2_X1 U22206 ( .A1(HOLD), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19115) );
  INV_X1 U22207 ( .A(n19115), .ZN(n19120) );
  INV_X1 U22208 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19111) );
  NOR3_X1 U22209 ( .A1(n19114), .A2(n19120), .A3(n19111), .ZN(n19113) );
  NAND2_X1 U22210 ( .A1(n19252), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19118) );
  AND2_X1 U22211 ( .A1(n19118), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19124) );
  INV_X1 U22212 ( .A(NA), .ZN(n20775) );
  OAI21_X1 U22213 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n20775), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n19123) );
  INV_X1 U22214 ( .A(n19123), .ZN(n19112) );
  OAI22_X1 U22215 ( .A1(n19260), .A2(n19113), .B1(n19124), .B2(n19112), .ZN(
        P3_U3029) );
  AOI22_X1 U22216 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n19125), .ZN(n19117) );
  OAI211_X1 U22217 ( .C1(n19117), .C2(n19122), .A(n19118), .B(n19116), .ZN(
        P3_U3030) );
  OAI22_X1 U22218 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19118), .ZN(n19119) );
  OAI22_X1 U22219 ( .A1(n19120), .A2(n19119), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19121) );
  OAI22_X1 U22220 ( .A1(n19124), .A2(n19123), .B1(n19122), .B2(n19121), .ZN(
        P3_U3031) );
  OAI222_X1 U22221 ( .A1(n19234), .A2(n19187), .B1(n19126), .B2(n19260), .C1(
        n19127), .C2(n19183), .ZN(P3_U3032) );
  INV_X1 U22222 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19129) );
  OAI222_X1 U22223 ( .A1(n19183), .A2(n19129), .B1(n19128), .B2(n19260), .C1(
        n19127), .C2(n19187), .ZN(P3_U3033) );
  OAI222_X1 U22224 ( .A1(n19183), .A2(n19131), .B1(n19130), .B2(n19260), .C1(
        n19129), .C2(n19187), .ZN(P3_U3034) );
  INV_X1 U22225 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19134) );
  OAI222_X1 U22226 ( .A1(n19183), .A2(n19134), .B1(n19132), .B2(n19260), .C1(
        n19131), .C2(n19187), .ZN(P3_U3035) );
  OAI222_X1 U22227 ( .A1(n19134), .A2(n19187), .B1(n19133), .B2(n19260), .C1(
        n19135), .C2(n19183), .ZN(P3_U3036) );
  OAI222_X1 U22228 ( .A1(n19183), .A2(n19137), .B1(n19136), .B2(n19260), .C1(
        n19135), .C2(n19187), .ZN(P3_U3037) );
  OAI222_X1 U22229 ( .A1(n19183), .A2(n19139), .B1(n19138), .B2(n19260), .C1(
        n19137), .C2(n19187), .ZN(P3_U3038) );
  OAI222_X1 U22230 ( .A1(n19183), .A2(n19141), .B1(n19140), .B2(n19260), .C1(
        n19139), .C2(n19187), .ZN(P3_U3039) );
  OAI222_X1 U22231 ( .A1(n19183), .A2(n19143), .B1(n19142), .B2(n19260), .C1(
        n19141), .C2(n19187), .ZN(P3_U3040) );
  INV_X1 U22232 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19145) );
  OAI222_X1 U22233 ( .A1(n19183), .A2(n19145), .B1(n19144), .B2(n19260), .C1(
        n19143), .C2(n19187), .ZN(P3_U3041) );
  OAI222_X1 U22234 ( .A1(n19183), .A2(n19147), .B1(n19146), .B2(n19260), .C1(
        n19145), .C2(n19187), .ZN(P3_U3042) );
  INV_X1 U22235 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19149) );
  OAI222_X1 U22236 ( .A1(n19183), .A2(n19149), .B1(n19148), .B2(n19260), .C1(
        n19147), .C2(n19187), .ZN(P3_U3043) );
  OAI222_X1 U22237 ( .A1(n19183), .A2(n19152), .B1(n19150), .B2(n19260), .C1(
        n19149), .C2(n19187), .ZN(P3_U3044) );
  OAI222_X1 U22238 ( .A1(n19152), .A2(n19187), .B1(n19151), .B2(n19260), .C1(
        n19153), .C2(n19183), .ZN(P3_U3045) );
  OAI222_X1 U22239 ( .A1(n19183), .A2(n19155), .B1(n19154), .B2(n19260), .C1(
        n19153), .C2(n19187), .ZN(P3_U3046) );
  OAI222_X1 U22240 ( .A1(n19183), .A2(n19157), .B1(n19156), .B2(n19260), .C1(
        n19155), .C2(n19187), .ZN(P3_U3047) );
  OAI222_X1 U22241 ( .A1(n19183), .A2(n19159), .B1(n19158), .B2(n19260), .C1(
        n19157), .C2(n19187), .ZN(P3_U3048) );
  OAI222_X1 U22242 ( .A1(n19183), .A2(n19161), .B1(n19160), .B2(n19260), .C1(
        n19159), .C2(n19187), .ZN(P3_U3049) );
  INV_X1 U22243 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19164) );
  OAI222_X1 U22244 ( .A1(n19183), .A2(n19164), .B1(n19162), .B2(n19260), .C1(
        n19161), .C2(n19187), .ZN(P3_U3050) );
  INV_X1 U22245 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19165) );
  OAI222_X1 U22246 ( .A1(n19164), .A2(n19187), .B1(n19163), .B2(n19260), .C1(
        n19165), .C2(n19183), .ZN(P3_U3051) );
  INV_X1 U22247 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19167) );
  OAI222_X1 U22248 ( .A1(n19183), .A2(n19167), .B1(n19166), .B2(n19260), .C1(
        n19165), .C2(n19187), .ZN(P3_U3052) );
  OAI222_X1 U22249 ( .A1(n19183), .A2(n19170), .B1(n19168), .B2(n19260), .C1(
        n19167), .C2(n19187), .ZN(P3_U3053) );
  OAI222_X1 U22250 ( .A1(n19170), .A2(n19187), .B1(n19169), .B2(n19260), .C1(
        n19171), .C2(n19183), .ZN(P3_U3054) );
  INV_X1 U22251 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19173) );
  OAI222_X1 U22252 ( .A1(n19183), .A2(n19173), .B1(n19172), .B2(n19260), .C1(
        n19171), .C2(n19187), .ZN(P3_U3055) );
  OAI222_X1 U22253 ( .A1(n19183), .A2(n19175), .B1(n19174), .B2(n19260), .C1(
        n19173), .C2(n19187), .ZN(P3_U3056) );
  OAI222_X1 U22254 ( .A1(n19183), .A2(n19177), .B1(n19176), .B2(n19260), .C1(
        n19175), .C2(n19187), .ZN(P3_U3057) );
  OAI222_X1 U22255 ( .A1(n19183), .A2(n19180), .B1(n19178), .B2(n19260), .C1(
        n19177), .C2(n19187), .ZN(P3_U3058) );
  OAI222_X1 U22256 ( .A1(n19187), .A2(n19180), .B1(n19179), .B2(n19260), .C1(
        n19181), .C2(n19183), .ZN(P3_U3059) );
  OAI222_X1 U22257 ( .A1(n19183), .A2(n19186), .B1(n19182), .B2(n19260), .C1(
        n19181), .C2(n19187), .ZN(P3_U3060) );
  OAI222_X1 U22258 ( .A1(n19187), .A2(n19186), .B1(n19185), .B2(n19260), .C1(
        n19184), .C2(n19183), .ZN(P3_U3061) );
  INV_X1 U22259 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19188) );
  AOI22_X1 U22260 ( .A1(n19260), .A2(n19189), .B1(n19188), .B2(n19258), .ZN(
        P3_U3274) );
  INV_X1 U22261 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19237) );
  INV_X1 U22262 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19190) );
  AOI22_X1 U22263 ( .A1(n19260), .A2(n19237), .B1(n19190), .B2(n19258), .ZN(
        P3_U3275) );
  INV_X1 U22264 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19191) );
  AOI22_X1 U22265 ( .A1(n19260), .A2(n19192), .B1(n19191), .B2(n19258), .ZN(
        P3_U3276) );
  INV_X1 U22266 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19240) );
  INV_X1 U22267 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19193) );
  AOI22_X1 U22268 ( .A1(n19260), .A2(n19240), .B1(n19193), .B2(n19258), .ZN(
        P3_U3277) );
  INV_X1 U22269 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19195) );
  INV_X1 U22270 ( .A(n19197), .ZN(n19194) );
  AOI21_X1 U22271 ( .B1(n19196), .B2(n19195), .A(n19194), .ZN(P3_U3280) );
  OAI21_X1 U22272 ( .B1(n19199), .B2(n19198), .A(n19197), .ZN(P3_U3281) );
  OAI221_X1 U22273 ( .B1(n19202), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19202), 
        .C2(n19201), .A(n19200), .ZN(P3_U3282) );
  AOI22_X1 U22274 ( .A1(n19262), .A2(n19204), .B1(n19228), .B2(n19203), .ZN(
        n19209) );
  INV_X1 U22275 ( .A(n19205), .ZN(n19206) );
  AOI21_X1 U22276 ( .B1(n19262), .B2(n19206), .A(n19233), .ZN(n19208) );
  OAI22_X1 U22277 ( .A1(n19233), .A2(n19209), .B1(n19208), .B2(n19207), .ZN(
        P3_U3285) );
  AOI22_X1 U22278 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19211), .B2(n19210), .ZN(
        n19221) );
  NOR2_X1 U22279 ( .A1(n20997), .A2(n19212), .ZN(n19222) );
  INV_X1 U22280 ( .A(n19262), .ZN(n19215) );
  OAI22_X1 U22281 ( .A1(n19216), .A2(n19215), .B1(n19214), .B2(n19213), .ZN(
        n19217) );
  AOI21_X1 U22282 ( .B1(n19221), .B2(n19222), .A(n19217), .ZN(n19218) );
  AOI22_X1 U22283 ( .A1(n19233), .A2(n19219), .B1(n19218), .B2(n19230), .ZN(
        P3_U3288) );
  INV_X1 U22284 ( .A(n19220), .ZN(n19224) );
  INV_X1 U22285 ( .A(n19221), .ZN(n19223) );
  AOI222_X1 U22286 ( .A1(n19225), .A2(n19262), .B1(n19228), .B2(n19224), .C1(
        n19223), .C2(n19222), .ZN(n19226) );
  AOI22_X1 U22287 ( .A1(n19233), .A2(n19227), .B1(n19226), .B2(n19230), .ZN(
        P3_U3289) );
  AOI222_X1 U22288 ( .A1(n20997), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19229), 
        .B2(n19262), .C1(n19232), .C2(n19228), .ZN(n19231) );
  AOI22_X1 U22289 ( .A1(n19233), .A2(n19232), .B1(n19231), .B2(n19230), .ZN(
        P3_U3290) );
  AOI21_X1 U22290 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19235) );
  AOI22_X1 U22291 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19235), .B2(n19234), .ZN(n19238) );
  AOI22_X1 U22292 ( .A1(n19241), .A2(n19238), .B1(n19237), .B2(n19236), .ZN(
        P3_U3292) );
  OAI21_X1 U22293 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19241), .ZN(n19239) );
  OAI21_X1 U22294 ( .B1(n19241), .B2(n19240), .A(n19239), .ZN(P3_U3293) );
  INV_X1 U22295 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19242) );
  AOI22_X1 U22296 ( .A1(n19260), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19242), 
        .B2(n19258), .ZN(P3_U3294) );
  MUX2_X1 U22297 ( .A(P3_MORE_REG_SCAN_IN), .B(n19244), .S(n19243), .Z(
        P3_U3295) );
  OAI21_X1 U22298 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19246), .A(n19245), 
        .ZN(n19247) );
  AOI211_X1 U22299 ( .C1(n19265), .C2(n19247), .A(n19252), .B(n19261), .ZN(
        n19250) );
  OAI21_X1 U22300 ( .B1(n19250), .B2(n19249), .A(n19248), .ZN(n19257) );
  NOR2_X1 U22301 ( .A1(n19252), .A2(n19251), .ZN(n19253) );
  AOI211_X1 U22302 ( .C1(n19255), .C2(n19254), .A(n19253), .B(n19264), .ZN(
        n19256) );
  MUX2_X1 U22303 ( .A(n19257), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n19256), 
        .Z(P3_U3296) );
  INV_X1 U22304 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19267) );
  INV_X1 U22305 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19259) );
  AOI22_X1 U22306 ( .A1(n19260), .A2(n19267), .B1(n19259), .B2(n19258), .ZN(
        P3_U3297) );
  AOI21_X1 U22307 ( .B1(n19262), .B2(n19261), .A(n19264), .ZN(n19268) );
  INV_X1 U22308 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19263) );
  AOI22_X1 U22309 ( .A1(n19265), .A2(n19264), .B1(n19268), .B2(n19263), .ZN(
        P3_U3298) );
  AOI21_X1 U22310 ( .B1(n19268), .B2(n19267), .A(n19266), .ZN(P3_U3299) );
  INV_X1 U22311 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20131) );
  INV_X1 U22312 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19269) );
  NAND2_X1 U22313 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20149), .ZN(n20139) );
  NAND2_X1 U22314 ( .A1(n20131), .A2(n20130), .ZN(n20135) );
  OAI21_X1 U22315 ( .B1(n20131), .B2(n20139), .A(n20135), .ZN(n20217) );
  OAI21_X1 U22316 ( .B1(n20131), .B2(n19269), .A(n20129), .ZN(P2_U2815) );
  INV_X1 U22317 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19271) );
  OAI22_X1 U22318 ( .A1(n19272), .A2(n19271), .B1(n20278), .B2(n19270), .ZN(
        P2_U2816) );
  NAND2_X1 U22319 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20131), .ZN(n20289) );
  AOI21_X1 U22320 ( .B1(n20131), .B2(n20149), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19273) );
  AOI22_X1 U22321 ( .A1(n20197), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19273), 
        .B2(n20289), .ZN(P2_U2817) );
  OAI21_X1 U22322 ( .B1(n20143), .B2(BS16), .A(n20217), .ZN(n20215) );
  OAI21_X1 U22323 ( .B1(n20217), .B2(n19952), .A(n20215), .ZN(P2_U2818) );
  AND2_X1 U22324 ( .A1(n20122), .A2(n19274), .ZN(n20266) );
  OAI21_X1 U22325 ( .B1(n20266), .B2(n19276), .A(n19275), .ZN(P2_U2819) );
  NOR4_X1 U22326 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19286) );
  NOR4_X1 U22327 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19285) );
  NOR4_X1 U22328 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19277) );
  INV_X1 U22329 ( .A(P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21025) );
  INV_X1 U22330 ( .A(P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20872) );
  NAND3_X1 U22331 ( .A1(n19277), .A2(n21025), .A3(n20872), .ZN(n19283) );
  NOR4_X1 U22332 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19281) );
  NOR4_X1 U22333 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19280) );
  NOR4_X1 U22334 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19279) );
  NOR4_X1 U22335 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19278) );
  NAND4_X1 U22336 ( .A1(n19281), .A2(n19280), .A3(n19279), .A4(n19278), .ZN(
        n19282) );
  AOI211_X1 U22337 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19283), .B(n19282), .ZN(n19284) );
  NAND3_X1 U22338 ( .A1(n19286), .A2(n19285), .A3(n19284), .ZN(n19292) );
  NOR2_X1 U22339 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19292), .ZN(n19287) );
  INV_X1 U22340 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20213) );
  AOI22_X1 U22341 ( .A1(n19287), .A2(n19406), .B1(n19292), .B2(n20213), .ZN(
        P2_U2820) );
  OR3_X1 U22342 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19291) );
  INV_X1 U22343 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20211) );
  AOI22_X1 U22344 ( .A1(n19287), .A2(n19291), .B1(n19292), .B2(n20211), .ZN(
        P2_U2821) );
  INV_X1 U22345 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20216) );
  NAND2_X1 U22346 ( .A1(n19287), .A2(n20216), .ZN(n19290) );
  INV_X1 U22347 ( .A(n19292), .ZN(n19293) );
  INV_X1 U22348 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20996) );
  OAI21_X1 U22349 ( .B1(n19406), .B2(n20996), .A(n19293), .ZN(n19288) );
  OAI21_X1 U22350 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19293), .A(n19288), 
        .ZN(n19289) );
  OAI221_X1 U22351 ( .B1(n19290), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19290), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19289), .ZN(P2_U2822) );
  INV_X1 U22352 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20209) );
  OAI221_X1 U22353 ( .B1(n19293), .B2(n20209), .C1(n19292), .C2(n19291), .A(
        n19290), .ZN(P2_U2823) );
  AOI22_X1 U22354 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19417), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19392), .ZN(n19304) );
  AOI22_X1 U22355 ( .A1(n19295), .A2(n19294), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19411), .ZN(n19303) );
  AOI22_X1 U22356 ( .A1(n19297), .A2(n19396), .B1(n19296), .B2(n19377), .ZN(
        n19302) );
  OAI211_X1 U22357 ( .C1(n19300), .C2(n19299), .A(n9671), .B(n19298), .ZN(
        n19301) );
  NAND4_X1 U22358 ( .A1(n19304), .A2(n19303), .A3(n19302), .A4(n19301), .ZN(
        P2_U2835) );
  OAI21_X1 U22359 ( .B1(n20180), .B2(n19405), .A(n19363), .ZN(n19307) );
  OAI22_X1 U22360 ( .A1(n19305), .A2(n19404), .B1(n10945), .B2(n19352), .ZN(
        n19306) );
  AOI211_X1 U22361 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19417), .A(
        n19307), .B(n19306), .ZN(n19314) );
  NOR2_X1 U22362 ( .A1(n19379), .A2(n19308), .ZN(n19310) );
  XNOR2_X1 U22363 ( .A(n19310), .B(n19309), .ZN(n19312) );
  AOI22_X1 U22364 ( .A1(n19312), .A2(n9671), .B1(n19311), .B2(n19396), .ZN(
        n19313) );
  OAI211_X1 U22365 ( .C1(n19315), .C2(n19408), .A(n19314), .B(n19313), .ZN(
        P2_U2837) );
  INV_X1 U22366 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20176) );
  OAI21_X1 U22367 ( .B1(n20176), .B2(n19405), .A(n19363), .ZN(n19318) );
  OAI22_X1 U22368 ( .A1(n19316), .A2(n19404), .B1(n10936), .B2(n19352), .ZN(
        n19317) );
  AOI211_X1 U22369 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19417), .A(
        n19318), .B(n19317), .ZN(n19325) );
  INV_X1 U22370 ( .A(n19319), .ZN(n19323) );
  XOR2_X1 U22371 ( .A(n19321), .B(n19320), .Z(n19322) );
  AOI22_X1 U22372 ( .A1(n19323), .A2(n19396), .B1(n9671), .B2(n19322), .ZN(
        n19324) );
  OAI211_X1 U22373 ( .C1(n19326), .C2(n19408), .A(n19325), .B(n19324), .ZN(
        P2_U2839) );
  OAI21_X1 U22374 ( .B1(n19379), .B2(n19327), .A(n9671), .ZN(n19329) );
  OAI22_X1 U22375 ( .A1(n19334), .A2(n19329), .B1(n19328), .B2(n19389), .ZN(
        n19330) );
  AOI21_X1 U22376 ( .B1(n19411), .B2(P2_EBX_REG_14__SCAN_IN), .A(n19330), .ZN(
        n19331) );
  OAI21_X1 U22377 ( .B1(n19332), .B2(n19404), .A(n19331), .ZN(n19333) );
  AOI211_X1 U22378 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19392), .A(n19529), 
        .B(n19333), .ZN(n19338) );
  AOI22_X1 U22379 ( .A1(n19336), .A2(n19396), .B1(n19335), .B2(n19334), .ZN(
        n19337) );
  OAI211_X1 U22380 ( .C1(n19432), .C2(n19408), .A(n19338), .B(n19337), .ZN(
        P2_U2841) );
  OAI22_X1 U22381 ( .A1(n19340), .A2(n19404), .B1(n19352), .B2(n19339), .ZN(
        n19341) );
  INV_X1 U22382 ( .A(n19341), .ZN(n19342) );
  OAI211_X1 U22383 ( .C1(n20166), .C2(n19405), .A(n19342), .B(n19363), .ZN(
        n19343) );
  AOI21_X1 U22384 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19417), .A(
        n19343), .ZN(n19350) );
  NOR2_X1 U22385 ( .A1(n19379), .A2(n19344), .ZN(n19346) );
  XNOR2_X1 U22386 ( .A(n19346), .B(n19345), .ZN(n19348) );
  AOI22_X1 U22387 ( .A1(n19348), .A2(n9671), .B1(n19347), .B2(n19396), .ZN(
        n19349) );
  OAI211_X1 U22388 ( .C1(n19444), .C2(n19408), .A(n19350), .B(n19349), .ZN(
        P2_U2845) );
  INV_X1 U22389 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19351) );
  OAI222_X1 U22390 ( .A1(n19404), .A2(n19354), .B1(n19353), .B2(n19352), .C1(
        n19351), .C2(n19389), .ZN(n19355) );
  AOI211_X1 U22391 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19392), .A(n19529), .B(
        n19355), .ZN(n19362) );
  NOR2_X1 U22392 ( .A1(n19379), .A2(n19356), .ZN(n19358) );
  XNOR2_X1 U22393 ( .A(n19358), .B(n19357), .ZN(n19360) );
  AOI22_X1 U22394 ( .A1(n19360), .A2(n9671), .B1(n19359), .B2(n19396), .ZN(
        n19361) );
  OAI211_X1 U22395 ( .C1(n19451), .C2(n19408), .A(n19362), .B(n19361), .ZN(
        P2_U2847) );
  OAI21_X1 U22396 ( .B1(n20159), .B2(n19405), .A(n19363), .ZN(n19366) );
  OAI22_X1 U22397 ( .A1(n19364), .A2(n19404), .B1(n10046), .B2(n19389), .ZN(
        n19365) );
  AOI211_X1 U22398 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19411), .A(n19366), .B(
        n19365), .ZN(n19373) );
  NOR2_X1 U22399 ( .A1(n19379), .A2(n19367), .ZN(n19369) );
  XNOR2_X1 U22400 ( .A(n19369), .B(n19368), .ZN(n19371) );
  AOI22_X1 U22401 ( .A1(n19371), .A2(n9671), .B1(n19370), .B2(n19396), .ZN(
        n19372) );
  OAI211_X1 U22402 ( .C1(n19408), .C2(n19453), .A(n19373), .B(n19372), .ZN(
        P2_U2849) );
  AOI21_X1 U22403 ( .B1(P2_REIP_REG_4__SCAN_IN), .B2(n19392), .A(n19529), .ZN(
        n19388) );
  INV_X1 U22404 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19374) );
  OAI22_X1 U22405 ( .A1(n19404), .A2(n19375), .B1(n19389), .B2(n19374), .ZN(
        n19376) );
  INV_X1 U22406 ( .A(n19376), .ZN(n19387) );
  AOI22_X1 U22407 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19411), .B1(n19377), .B2(
        n19464), .ZN(n19386) );
  NOR2_X1 U22408 ( .A1(n19379), .A2(n19378), .ZN(n19380) );
  XNOR2_X1 U22409 ( .A(n19541), .B(n19380), .ZN(n19384) );
  OAI22_X1 U22410 ( .A1(n19466), .A2(n19382), .B1(n19381), .B2(n19413), .ZN(
        n19383) );
  AOI21_X1 U22411 ( .B1(n19384), .B2(n9671), .A(n19383), .ZN(n19385) );
  NAND4_X1 U22412 ( .A1(n19388), .A2(n19387), .A3(n19386), .A4(n19385), .ZN(
        P2_U2851) );
  OAI22_X1 U22413 ( .A1(n19404), .A2(n19390), .B1(n12092), .B2(n19389), .ZN(
        n19391) );
  AOI21_X1 U22414 ( .B1(P2_REIP_REG_1__SCAN_IN), .B2(n19392), .A(n19391), .ZN(
        n19394) );
  NAND2_X1 U22415 ( .A1(n19411), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19393) );
  OAI211_X1 U22416 ( .C1(n19455), .C2(n19408), .A(n19394), .B(n19393), .ZN(
        n19395) );
  AOI21_X1 U22417 ( .B1(n10437), .B2(n19396), .A(n19395), .ZN(n19399) );
  AOI22_X1 U22418 ( .A1(n20248), .A2(n19416), .B1(n12092), .B2(n19397), .ZN(
        n19398) );
  OAI211_X1 U22419 ( .C1(n20126), .C2(n19400), .A(n19399), .B(n19398), .ZN(
        P2_U2854) );
  INV_X1 U22420 ( .A(n19402), .ZN(n19403) );
  OAI22_X1 U22421 ( .A1(n19406), .A2(n19405), .B1(n19404), .B2(n19403), .ZN(
        n19410) );
  NOR2_X1 U22422 ( .A1(n19408), .A2(n19407), .ZN(n19409) );
  AOI211_X1 U22423 ( .C1(P2_EBX_REG_0__SCAN_IN), .C2(n19411), .A(n19410), .B(
        n19409), .ZN(n19412) );
  OAI21_X1 U22424 ( .B1(n19414), .B2(n19413), .A(n19412), .ZN(n19415) );
  AOI21_X1 U22425 ( .B1(n19827), .B2(n19416), .A(n19415), .ZN(n19419) );
  NAND2_X1 U22426 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19417), .ZN(
        n19418) );
  OAI211_X1 U22427 ( .C1(n15875), .C2(n20126), .A(n19419), .B(n19418), .ZN(
        P2_U2855) );
  AOI22_X1 U22428 ( .A1(n19421), .A2(n19486), .B1(n19420), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19424) );
  AOI22_X1 U22429 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n19422), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19485), .ZN(n19423) );
  NAND2_X1 U22430 ( .A1(n19424), .A2(n19423), .ZN(P2_U2888) );
  INV_X1 U22431 ( .A(n19425), .ZN(n19430) );
  INV_X1 U22432 ( .A(n19426), .ZN(n19428) );
  OAI222_X1 U22433 ( .A1(n12130), .A2(n19463), .B1(n19430), .B2(n19462), .C1(
        n19429), .C2(n19492), .ZN(P2_U2904) );
  INV_X1 U22434 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19497) );
  OAI222_X1 U22435 ( .A1(n19497), .A2(n19463), .B1(n19432), .B2(n19462), .C1(
        n19492), .C2(n19431), .ZN(P2_U2905) );
  INV_X1 U22436 ( .A(n19492), .ZN(n19446) );
  AOI22_X1 U22437 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n19485), .B1(n19433), 
        .B2(n19446), .ZN(n19434) );
  OAI21_X1 U22438 ( .B1(n19462), .B2(n19435), .A(n19434), .ZN(P2_U2906) );
  INV_X1 U22439 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19501) );
  INV_X1 U22440 ( .A(n19436), .ZN(n19438) );
  OAI222_X1 U22441 ( .A1(n19501), .A2(n19463), .B1(n19438), .B2(n19462), .C1(
        n19492), .C2(n19437), .ZN(P2_U2907) );
  INV_X1 U22442 ( .A(n19439), .ZN(n19442) );
  AOI22_X1 U22443 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(n19485), .B1(n19440), 
        .B2(n19446), .ZN(n19441) );
  OAI21_X1 U22444 ( .B1(n19462), .B2(n19442), .A(n19441), .ZN(P2_U2908) );
  INV_X1 U22445 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19505) );
  OAI222_X1 U22446 ( .A1(n19505), .A2(n19463), .B1(n19444), .B2(n19462), .C1(
        n19492), .C2(n19443), .ZN(P2_U2909) );
  INV_X1 U22447 ( .A(n19445), .ZN(n19449) );
  AOI22_X1 U22448 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19485), .B1(n19447), .B2(
        n19446), .ZN(n19448) );
  OAI21_X1 U22449 ( .B1(n19462), .B2(n19449), .A(n19448), .ZN(P2_U2910) );
  INV_X1 U22450 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19510) );
  OAI222_X1 U22451 ( .A1(n19510), .A2(n19463), .B1(n19451), .B2(n19462), .C1(
        n19492), .C2(n19450), .ZN(P2_U2911) );
  INV_X1 U22452 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19512) );
  OAI222_X1 U22453 ( .A1(n19512), .A2(n19463), .B1(n19452), .B2(n19462), .C1(
        n19492), .C2(n19592), .ZN(P2_U2912) );
  OAI222_X1 U22454 ( .A1(n11136), .A2(n19463), .B1(n19453), .B2(n19462), .C1(
        n19492), .C2(n19580), .ZN(P2_U2913) );
  INV_X1 U22455 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19515) );
  NAND2_X1 U22456 ( .A1(n19860), .A2(n19454), .ZN(n19457) );
  XNOR2_X1 U22457 ( .A(n19860), .B(n20228), .ZN(n19471) );
  XOR2_X1 U22458 ( .A(n20241), .B(n20239), .Z(n19477) );
  XNOR2_X1 U22459 ( .A(n20227), .B(n20250), .ZN(n19481) );
  NAND2_X1 U22460 ( .A1(n19827), .A2(n19489), .ZN(n19488) );
  AOI22_X1 U22461 ( .A1(n19481), .A2(n19488), .B1(n20227), .B2(n19455), .ZN(
        n19476) );
  INV_X1 U22462 ( .A(n20239), .ZN(n19456) );
  OAI22_X1 U22463 ( .A1(n19477), .A2(n19476), .B1(n19456), .B2(n20241), .ZN(
        n19472) );
  NAND2_X1 U22464 ( .A1(n19471), .A2(n19472), .ZN(n19470) );
  AOI21_X1 U22465 ( .B1(n19457), .B2(n19470), .A(n19464), .ZN(n19465) );
  NOR3_X1 U22466 ( .A1(n19465), .A2(n19466), .A3(n19458), .ZN(n19460) );
  NOR2_X1 U22467 ( .A1(n19460), .A2(n19459), .ZN(n19461) );
  OAI222_X1 U22468 ( .A1(n19515), .A2(n19463), .B1(n19577), .B2(n19492), .C1(
        n19462), .C2(n19461), .ZN(P2_U2914) );
  AOI22_X1 U22469 ( .A1(n19464), .A2(n19486), .B1(n19485), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19469) );
  XOR2_X1 U22470 ( .A(n19466), .B(n19465), .Z(n19467) );
  NAND2_X1 U22471 ( .A1(n19467), .A2(n19487), .ZN(n19468) );
  OAI211_X1 U22472 ( .C1(n19574), .C2(n19492), .A(n19469), .B(n19468), .ZN(
        P2_U2915) );
  AOI22_X1 U22473 ( .A1(n19486), .A2(n20228), .B1(n19485), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19475) );
  OAI21_X1 U22474 ( .B1(n19472), .B2(n19471), .A(n19470), .ZN(n19473) );
  NAND2_X1 U22475 ( .A1(n19473), .A2(n19487), .ZN(n19474) );
  OAI211_X1 U22476 ( .C1(n19570), .C2(n19492), .A(n19475), .B(n19474), .ZN(
        P2_U2916) );
  AOI22_X1 U22477 ( .A1(n19486), .A2(n20241), .B1(n19485), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19480) );
  XNOR2_X1 U22478 ( .A(n19477), .B(n19476), .ZN(n19478) );
  NAND2_X1 U22479 ( .A1(n19478), .A2(n19487), .ZN(n19479) );
  OAI211_X1 U22480 ( .C1(n19565), .C2(n19492), .A(n19480), .B(n19479), .ZN(
        P2_U2917) );
  AOI22_X1 U22481 ( .A1(n19486), .A2(n20250), .B1(n19485), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19484) );
  XNOR2_X1 U22482 ( .A(n19481), .B(n19488), .ZN(n19482) );
  NAND2_X1 U22483 ( .A1(n19482), .A2(n19487), .ZN(n19483) );
  OAI211_X1 U22484 ( .C1(n19560), .C2(n19492), .A(n19484), .B(n19483), .ZN(
        P2_U2918) );
  AOI22_X1 U22485 ( .A1(n19486), .A2(n19489), .B1(n19485), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19491) );
  OAI211_X1 U22486 ( .C1(n19827), .C2(n19489), .A(n19488), .B(n19487), .ZN(
        n19490) );
  OAI211_X1 U22487 ( .C1(n19553), .C2(n19492), .A(n19491), .B(n19490), .ZN(
        P2_U2919) );
  NOR2_X1 U22488 ( .A1(n19509), .A2(n19493), .ZN(P2_U2920) );
  AOI22_X1 U22489 ( .A1(n19521), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19495) );
  OAI21_X1 U22490 ( .B1(n12130), .B2(n19527), .A(n19495), .ZN(P2_U2936) );
  AOI22_X1 U22491 ( .A1(n19521), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19496) );
  OAI21_X1 U22492 ( .B1(n19497), .B2(n19527), .A(n19496), .ZN(P2_U2937) );
  AOI22_X1 U22493 ( .A1(n19525), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19498) );
  OAI21_X1 U22494 ( .B1(n19499), .B2(n19527), .A(n19498), .ZN(P2_U2938) );
  AOI22_X1 U22495 ( .A1(n19525), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19500) );
  OAI21_X1 U22496 ( .B1(n19501), .B2(n19527), .A(n19500), .ZN(P2_U2939) );
  AOI22_X1 U22497 ( .A1(n19525), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19502) );
  OAI21_X1 U22498 ( .B1(n19503), .B2(n19527), .A(n19502), .ZN(P2_U2940) );
  AOI22_X1 U22499 ( .A1(n19525), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19504) );
  OAI21_X1 U22500 ( .B1(n19505), .B2(n19527), .A(n19504), .ZN(P2_U2941) );
  AOI22_X1 U22501 ( .A1(n19525), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19506) );
  OAI21_X1 U22502 ( .B1(n19507), .B2(n19527), .A(n19506), .ZN(P2_U2942) );
  INV_X1 U22503 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n21030) );
  OAI222_X1 U22504 ( .A1(n20273), .A2(n21030), .B1(n19527), .B2(n19510), .C1(
        n19509), .C2(n19508), .ZN(P2_U2943) );
  AOI22_X1 U22505 ( .A1(n19525), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19511) );
  OAI21_X1 U22506 ( .B1(n19512), .B2(n19527), .A(n19511), .ZN(P2_U2944) );
  AOI22_X1 U22507 ( .A1(n19521), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19513) );
  OAI21_X1 U22508 ( .B1(n11136), .B2(n19527), .A(n19513), .ZN(P2_U2945) );
  AOI22_X1 U22509 ( .A1(n19521), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19514) );
  OAI21_X1 U22510 ( .B1(n19515), .B2(n19527), .A(n19514), .ZN(P2_U2946) );
  INV_X1 U22511 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U22512 ( .A1(n19521), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19516) );
  OAI21_X1 U22513 ( .B1(n20896), .B2(n19527), .A(n19516), .ZN(P2_U2947) );
  INV_X1 U22514 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19518) );
  AOI22_X1 U22515 ( .A1(n19521), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19517) );
  OAI21_X1 U22516 ( .B1(n19518), .B2(n19527), .A(n19517), .ZN(P2_U2948) );
  INV_X1 U22517 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19520) );
  AOI22_X1 U22518 ( .A1(n19521), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19519) );
  OAI21_X1 U22519 ( .B1(n19520), .B2(n19527), .A(n19519), .ZN(P2_U2949) );
  INV_X1 U22520 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19523) );
  AOI22_X1 U22521 ( .A1(n19521), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19524), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19522) );
  OAI21_X1 U22522 ( .B1(n19523), .B2(n19527), .A(n19522), .ZN(P2_U2950) );
  INV_X1 U22523 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U22524 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n19525), .B1(n19524), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19526) );
  OAI21_X1 U22525 ( .B1(n19528), .B2(n19527), .A(n19526), .ZN(P2_U2951) );
  AOI22_X1 U22526 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19530), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19529), .ZN(n19540) );
  INV_X1 U22527 ( .A(n19531), .ZN(n19535) );
  OAI22_X1 U22528 ( .A1(n19535), .A2(n19534), .B1(n19533), .B2(n19532), .ZN(
        n19536) );
  AOI21_X1 U22529 ( .B1(n19538), .B2(n19537), .A(n19536), .ZN(n19539) );
  OAI211_X1 U22530 ( .C1(n19542), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3010) );
  AOI22_X1 U22531 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19583), .ZN(n20072) );
  INV_X1 U22532 ( .A(n19589), .ZN(n19568) );
  AND2_X1 U22533 ( .A1(n20279), .A2(n19568), .ZN(n20060) );
  NAND2_X1 U22534 ( .A1(n20236), .A2(n20243), .ZN(n19677) );
  NOR2_X1 U22535 ( .A1(n19829), .A2(n19677), .ZN(n19591) );
  AOI22_X1 U22536 ( .A1(n20069), .A2(n20116), .B1(n20060), .B2(n19591), .ZN(
        n19559) );
  INV_X1 U22537 ( .A(n19647), .ZN(n19546) );
  OAI21_X1 U22538 ( .B1(n20116), .B2(n19546), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19547) );
  NAND2_X1 U22539 ( .A1(n19547), .A2(n20223), .ZN(n19557) );
  NOR2_X1 U22540 ( .A1(n20236), .A2(n19548), .ZN(n20111) );
  NOR2_X1 U22541 ( .A1(n20111), .A2(n19591), .ZN(n19556) );
  INV_X1 U22542 ( .A(n19556), .ZN(n19552) );
  INV_X1 U22543 ( .A(n19554), .ZN(n19550) );
  INV_X1 U22544 ( .A(n20223), .ZN(n20232) );
  INV_X1 U22545 ( .A(n19591), .ZN(n19549) );
  OAI211_X1 U22546 ( .C1(n19550), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20232), 
        .B(n19549), .ZN(n19551) );
  OAI211_X1 U22547 ( .C1(n19557), .C2(n19552), .A(n20067), .B(n19551), .ZN(
        n19594) );
  NOR2_X2 U22548 ( .A1(n19553), .A2(n19775), .ZN(n20061) );
  OAI21_X1 U22549 ( .B1(n19554), .B2(n19591), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19555) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19594), .B1(
        n20061), .B2(n19593), .ZN(n19558) );
  OAI211_X1 U22551 ( .C1(n20072), .C2(n19647), .A(n19559), .B(n19558), .ZN(
        P2_U3048) );
  AOI22_X1 U22552 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19583), .ZN(n20035) );
  NOR2_X2 U22553 ( .A1(n16723), .A2(n19589), .ZN(n20073) );
  AOI22_X1 U22554 ( .A1(n20032), .A2(n20116), .B1(n20073), .B2(n19591), .ZN(
        n19562) );
  NOR2_X2 U22555 ( .A1(n19560), .A2(n19775), .ZN(n20074) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19594), .B1(
        n20074), .B2(n19593), .ZN(n19561) );
  OAI211_X1 U22557 ( .C1(n20035), .C2(n19647), .A(n19562), .B(n19561), .ZN(
        P2_U3049) );
  AOI22_X1 U22558 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19583), .ZN(n20084) );
  NOR2_X2 U22559 ( .A1(n19564), .A2(n19589), .ZN(n20079) );
  AOI22_X1 U22560 ( .A1(n20036), .A2(n20116), .B1(n20079), .B2(n19591), .ZN(
        n19567) );
  NOR2_X2 U22561 ( .A1(n19565), .A2(n19775), .ZN(n20080) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19594), .B1(
        n20080), .B2(n19593), .ZN(n19566) );
  OAI211_X1 U22563 ( .C1(n20039), .C2(n19647), .A(n19567), .B(n19566), .ZN(
        P2_U3050) );
  AOI22_X1 U22564 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19583), .ZN(n19968) );
  AOI22_X1 U22565 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19583), .ZN(n20090) );
  AOI22_X1 U22566 ( .A1(n19965), .A2(n20116), .B1(n20085), .B2(n19591), .ZN(
        n19572) );
  NOR2_X2 U22567 ( .A1(n19570), .A2(n19775), .ZN(n20086) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19594), .B1(
        n20086), .B2(n19593), .ZN(n19571) );
  OAI211_X1 U22569 ( .C1(n19968), .C2(n19647), .A(n19572), .B(n19571), .ZN(
        P2_U3051) );
  AOI22_X1 U22570 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19583), .ZN(n20096) );
  OAI22_X2 U22571 ( .A1(n14485), .A2(n19584), .B1(n19573), .B2(n19585), .ZN(
        n20093) );
  NOR2_X2 U22572 ( .A1(n11352), .A2(n19589), .ZN(n20091) );
  AOI22_X1 U22573 ( .A1(n20093), .A2(n20116), .B1(n20091), .B2(n19591), .ZN(
        n19576) );
  NOR2_X2 U22574 ( .A1(n19574), .A2(n19775), .ZN(n20092) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19594), .B1(
        n20092), .B2(n19593), .ZN(n19575) );
  OAI211_X1 U22576 ( .C1(n20096), .C2(n19647), .A(n19576), .B(n19575), .ZN(
        P2_U3052) );
  AOI22_X1 U22577 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19583), .ZN(n20102) );
  AOI22_X1 U22578 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19583), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n9657), .ZN(n20009) );
  INV_X1 U22579 ( .A(n20009), .ZN(n20099) );
  NOR2_X2 U22580 ( .A1(n11007), .A2(n19589), .ZN(n20097) );
  AOI22_X1 U22581 ( .A1(n20099), .A2(n20116), .B1(n20097), .B2(n19591), .ZN(
        n19579) );
  NOR2_X2 U22582 ( .A1(n19577), .A2(n19775), .ZN(n20098) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19594), .B1(
        n20098), .B2(n19593), .ZN(n19578) );
  OAI211_X1 U22584 ( .C1(n20102), .C2(n19647), .A(n19579), .B(n19578), .ZN(
        P2_U3053) );
  AOI22_X1 U22585 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19583), .ZN(n20110) );
  AOI22_X1 U22586 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19583), .ZN(n20013) );
  NOR2_X2 U22587 ( .A1(n10372), .A2(n19589), .ZN(n20103) );
  AOI22_X1 U22588 ( .A1(n20105), .A2(n20116), .B1(n20103), .B2(n19591), .ZN(
        n19582) );
  NOR2_X2 U22589 ( .A1(n19580), .A2(n19775), .ZN(n20104) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19594), .B1(
        n20104), .B2(n19593), .ZN(n19581) );
  OAI211_X1 U22591 ( .C1(n20110), .C2(n19647), .A(n19582), .B(n19581), .ZN(
        P2_U3054) );
  AOI22_X1 U22592 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9657), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19583), .ZN(n20056) );
  OAI22_X2 U22593 ( .A1(n19588), .A2(n19584), .B1(n19586), .B2(n19585), .ZN(
        n20050) );
  NOR2_X2 U22594 ( .A1(n19590), .A2(n19589), .ZN(n20112) );
  AOI22_X1 U22595 ( .A1(n20050), .A2(n20116), .B1(n20112), .B2(n19591), .ZN(
        n19596) );
  NOR2_X2 U22596 ( .A1(n19592), .A2(n19775), .ZN(n20113) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19594), .B1(
        n20113), .B2(n19593), .ZN(n19595) );
  OAI211_X1 U22598 ( .C1(n20056), .C2(n19647), .A(n19596), .B(n19595), .ZN(
        P2_U3055) );
  NOR3_X1 U22599 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20263), .A3(
        n19677), .ZN(n19606) );
  INV_X1 U22600 ( .A(n19606), .ZN(n19639) );
  AND2_X1 U22601 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19639), .ZN(n19597) );
  NAND2_X1 U22602 ( .A1(n10682), .A2(n19597), .ZN(n19603) );
  OR2_X1 U22603 ( .A1(n19677), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19602) );
  AOI21_X1 U22604 ( .B1(n20269), .B2(n19602), .A(n19800), .ZN(n19598) );
  NAND2_X1 U22605 ( .A1(n19603), .A2(n19598), .ZN(n19642) );
  INV_X1 U22606 ( .A(n20061), .ZN(n19600) );
  INV_X1 U22607 ( .A(n20060), .ZN(n19599) );
  OAI22_X1 U22608 ( .A1(n19642), .A2(n19600), .B1(n19599), .B2(n19639), .ZN(
        n19601) );
  INV_X1 U22609 ( .A(n19601), .ZN(n19608) );
  NAND2_X1 U22610 ( .A1(n19860), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19801) );
  OAI21_X1 U22611 ( .B1(n19801), .B2(n19861), .A(n19602), .ZN(n19604) );
  AND2_X1 U22612 ( .A1(n19604), .A2(n19603), .ZN(n19605) );
  OAI211_X1 U22613 ( .C1(n19606), .C2(n20268), .A(n19605), .B(n20067), .ZN(
        n19644) );
  NAND2_X1 U22614 ( .A1(n19828), .A2(n19807), .ZN(n19650) );
  INV_X1 U22615 ( .A(n20072), .ZN(n19992) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n19992), .ZN(n19607) );
  OAI211_X1 U22617 ( .C1(n19995), .C2(n19647), .A(n19608), .B(n19607), .ZN(
        P2_U3056) );
  INV_X1 U22618 ( .A(n20074), .ZN(n19610) );
  INV_X1 U22619 ( .A(n20073), .ZN(n19609) );
  OAI22_X1 U22620 ( .A1(n19642), .A2(n19610), .B1(n19609), .B2(n19639), .ZN(
        n19611) );
  INV_X1 U22621 ( .A(n19611), .ZN(n19613) );
  INV_X1 U22622 ( .A(n20035), .ZN(n20075) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n20075), .ZN(n19612) );
  OAI211_X1 U22624 ( .C1(n20078), .C2(n19647), .A(n19613), .B(n19612), .ZN(
        P2_U3057) );
  INV_X1 U22625 ( .A(n20080), .ZN(n19615) );
  INV_X1 U22626 ( .A(n20079), .ZN(n19614) );
  OAI22_X1 U22627 ( .A1(n19642), .A2(n19615), .B1(n19614), .B2(n19639), .ZN(
        n19616) );
  INV_X1 U22628 ( .A(n19616), .ZN(n19618) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n20081), .ZN(n19617) );
  OAI211_X1 U22630 ( .C1(n20084), .C2(n19647), .A(n19618), .B(n19617), .ZN(
        P2_U3058) );
  INV_X1 U22631 ( .A(n20086), .ZN(n19620) );
  INV_X1 U22632 ( .A(n20085), .ZN(n19619) );
  OAI22_X1 U22633 ( .A1(n19642), .A2(n19620), .B1(n19619), .B2(n19639), .ZN(
        n19621) );
  INV_X1 U22634 ( .A(n19621), .ZN(n19623) );
  INV_X1 U22635 ( .A(n19968), .ZN(n20087) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n20087), .ZN(n19622) );
  OAI211_X1 U22637 ( .C1(n20090), .C2(n19647), .A(n19623), .B(n19622), .ZN(
        P2_U3059) );
  INV_X1 U22638 ( .A(n20092), .ZN(n19625) );
  INV_X1 U22639 ( .A(n20091), .ZN(n19624) );
  OAI22_X1 U22640 ( .A1(n19642), .A2(n19625), .B1(n19624), .B2(n19639), .ZN(
        n19626) );
  INV_X1 U22641 ( .A(n19626), .ZN(n19628) );
  INV_X1 U22642 ( .A(n20096), .ZN(n20002) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n20002), .ZN(n19627) );
  OAI211_X1 U22644 ( .C1(n20005), .C2(n19647), .A(n19628), .B(n19627), .ZN(
        P2_U3060) );
  INV_X1 U22645 ( .A(n20098), .ZN(n19630) );
  INV_X1 U22646 ( .A(n20097), .ZN(n19629) );
  OAI22_X1 U22647 ( .A1(n19642), .A2(n19630), .B1(n19629), .B2(n19639), .ZN(
        n19631) );
  INV_X1 U22648 ( .A(n19631), .ZN(n19633) );
  INV_X1 U22649 ( .A(n20102), .ZN(n20006) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n20006), .ZN(n19632) );
  OAI211_X1 U22651 ( .C1(n20009), .C2(n19647), .A(n19633), .B(n19632), .ZN(
        P2_U3061) );
  INV_X1 U22652 ( .A(n20104), .ZN(n19635) );
  INV_X1 U22653 ( .A(n20103), .ZN(n19634) );
  OAI22_X1 U22654 ( .A1(n19642), .A2(n19635), .B1(n19634), .B2(n19639), .ZN(
        n19636) );
  INV_X1 U22655 ( .A(n19636), .ZN(n19638) );
  INV_X1 U22656 ( .A(n20110), .ZN(n20010) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n20010), .ZN(n19637) );
  OAI211_X1 U22658 ( .C1(n20013), .C2(n19647), .A(n19638), .B(n19637), .ZN(
        P2_U3062) );
  INV_X1 U22659 ( .A(n20050), .ZN(n20121) );
  INV_X1 U22660 ( .A(n20113), .ZN(n19641) );
  INV_X1 U22661 ( .A(n20112), .ZN(n19640) );
  OAI22_X1 U22662 ( .A1(n19642), .A2(n19641), .B1(n19640), .B2(n19639), .ZN(
        n19643) );
  INV_X1 U22663 ( .A(n19643), .ZN(n19646) );
  INV_X1 U22664 ( .A(n20056), .ZN(n20115) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19644), .B1(
        n19672), .B2(n20115), .ZN(n19645) );
  OAI211_X1 U22666 ( .C1(n20121), .C2(n19647), .A(n19646), .B(n19645), .ZN(
        P2_U3063) );
  NOR3_X2 U22667 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20252), .A3(
        n19677), .ZN(n19670) );
  OAI21_X1 U22668 ( .B1(n10620), .B2(n19670), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19649) );
  NOR2_X1 U22669 ( .A1(n19892), .A2(n19677), .ZN(n19651) );
  INV_X1 U22670 ( .A(n19651), .ZN(n19648) );
  NAND2_X1 U22671 ( .A1(n19649), .A2(n19648), .ZN(n19671) );
  AOI22_X1 U22672 ( .A1(n19671), .A2(n20061), .B1(n20060), .B2(n19670), .ZN(
        n19657) );
  AOI21_X1 U22673 ( .B1(n10620), .B2(n20268), .A(n19670), .ZN(n19654) );
  AOI21_X1 U22674 ( .B1(n19706), .B2(n19650), .A(n19952), .ZN(n19652) );
  NOR2_X1 U22675 ( .A1(n19652), .A2(n19651), .ZN(n19653) );
  MUX2_X1 U22676 ( .A(n19654), .B(n19653), .S(n20223), .Z(n19655) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n20069), .ZN(n19656) );
  OAI211_X1 U22678 ( .C1(n20072), .C2(n19706), .A(n19657), .B(n19656), .ZN(
        P2_U3064) );
  AOI22_X1 U22679 ( .A1(n19671), .A2(n20074), .B1(n20073), .B2(n19670), .ZN(
        n19659) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n20032), .ZN(n19658) );
  OAI211_X1 U22681 ( .C1(n20035), .C2(n19706), .A(n19659), .B(n19658), .ZN(
        P2_U3065) );
  AOI22_X1 U22682 ( .A1(n19671), .A2(n20080), .B1(n20079), .B2(n19670), .ZN(
        n19661) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n20036), .ZN(n19660) );
  OAI211_X1 U22684 ( .C1(n20039), .C2(n19706), .A(n19661), .B(n19660), .ZN(
        P2_U3066) );
  AOI22_X1 U22685 ( .A1(n19671), .A2(n20086), .B1(n20085), .B2(n19670), .ZN(
        n19663) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n19965), .ZN(n19662) );
  OAI211_X1 U22687 ( .C1(n19968), .C2(n19706), .A(n19663), .B(n19662), .ZN(
        P2_U3067) );
  AOI22_X1 U22688 ( .A1(n19671), .A2(n20092), .B1(n20091), .B2(n19670), .ZN(
        n19665) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n20093), .ZN(n19664) );
  OAI211_X1 U22690 ( .C1(n20096), .C2(n19706), .A(n19665), .B(n19664), .ZN(
        P2_U3068) );
  AOI22_X1 U22691 ( .A1(n19671), .A2(n20098), .B1(n20097), .B2(n19670), .ZN(
        n19667) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n20099), .ZN(n19666) );
  OAI211_X1 U22693 ( .C1(n20102), .C2(n19706), .A(n19667), .B(n19666), .ZN(
        P2_U3069) );
  AOI22_X1 U22694 ( .A1(n19671), .A2(n20104), .B1(n20103), .B2(n19670), .ZN(
        n19669) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n20105), .ZN(n19668) );
  OAI211_X1 U22696 ( .C1(n20110), .C2(n19706), .A(n19669), .B(n19668), .ZN(
        P2_U3070) );
  AOI22_X1 U22697 ( .A1(n19671), .A2(n20113), .B1(n20112), .B2(n19670), .ZN(
        n19675) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19673), .B1(
        n19672), .B2(n20050), .ZN(n19674) );
  OAI211_X1 U22699 ( .C1(n20056), .C2(n19706), .A(n19675), .B(n19674), .ZN(
        P2_U3071) );
  NOR2_X1 U22700 ( .A1(n19920), .A2(n19677), .ZN(n19701) );
  AOI22_X1 U22701 ( .A1(n19992), .A2(n19734), .B1(n19701), .B2(n20060), .ZN(
        n19687) );
  INV_X1 U22702 ( .A(n20224), .ZN(n19676) );
  OAI21_X1 U22703 ( .B1(n19801), .B2(n19676), .A(n20223), .ZN(n19685) );
  NOR2_X1 U22704 ( .A1(n20252), .A2(n19677), .ZN(n19682) );
  OAI21_X1 U22705 ( .B1(n19678), .B2(n20269), .A(n20268), .ZN(n19680) );
  INV_X1 U22706 ( .A(n19701), .ZN(n19679) );
  AOI21_X1 U22707 ( .B1(n19680), .B2(n19679), .A(n19775), .ZN(n19681) );
  OAI21_X1 U22708 ( .B1(n19685), .B2(n19682), .A(n19681), .ZN(n19703) );
  INV_X1 U22709 ( .A(n19682), .ZN(n19684) );
  NOR2_X1 U22710 ( .A1(n19678), .A2(n19701), .ZN(n19683) );
  OAI22_X1 U22711 ( .A1(n19685), .A2(n19684), .B1(n19683), .B2(n20269), .ZN(
        n19702) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19703), .B1(
        n20061), .B2(n19702), .ZN(n19686) );
  OAI211_X1 U22713 ( .C1(n19995), .C2(n19706), .A(n19687), .B(n19686), .ZN(
        P2_U3072) );
  AOI22_X1 U22714 ( .A1(n20075), .A2(n19734), .B1(n19701), .B2(n20073), .ZN(
        n19689) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19703), .B1(
        n20074), .B2(n19702), .ZN(n19688) );
  OAI211_X1 U22716 ( .C1(n20078), .C2(n19706), .A(n19689), .B(n19688), .ZN(
        P2_U3073) );
  INV_X1 U22717 ( .A(n19706), .ZN(n19692) );
  AOI22_X1 U22718 ( .A1(n20036), .A2(n19692), .B1(n19701), .B2(n20079), .ZN(
        n19691) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19703), .B1(
        n20080), .B2(n19702), .ZN(n19690) );
  OAI211_X1 U22720 ( .C1(n20039), .C2(n19732), .A(n19691), .B(n19690), .ZN(
        P2_U3074) );
  AOI22_X1 U22721 ( .A1(n19965), .A2(n19692), .B1(n19701), .B2(n20085), .ZN(
        n19694) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19703), .B1(
        n20086), .B2(n19702), .ZN(n19693) );
  OAI211_X1 U22723 ( .C1(n19968), .C2(n19732), .A(n19694), .B(n19693), .ZN(
        P2_U3075) );
  AOI22_X1 U22724 ( .A1(n20002), .A2(n19734), .B1(n19701), .B2(n20091), .ZN(
        n19696) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19703), .B1(
        n20092), .B2(n19702), .ZN(n19695) );
  OAI211_X1 U22726 ( .C1(n20005), .C2(n19706), .A(n19696), .B(n19695), .ZN(
        P2_U3076) );
  AOI22_X1 U22727 ( .A1(n20006), .A2(n19734), .B1(n19701), .B2(n20097), .ZN(
        n19698) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19703), .B1(
        n20098), .B2(n19702), .ZN(n19697) );
  OAI211_X1 U22729 ( .C1(n20009), .C2(n19706), .A(n19698), .B(n19697), .ZN(
        P2_U3077) );
  AOI22_X1 U22730 ( .A1(n20010), .A2(n19734), .B1(n19701), .B2(n20103), .ZN(
        n19700) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19703), .B1(
        n20104), .B2(n19702), .ZN(n19699) );
  OAI211_X1 U22732 ( .C1(n20013), .C2(n19706), .A(n19700), .B(n19699), .ZN(
        P2_U3078) );
  AOI22_X1 U22733 ( .A1(n20115), .A2(n19734), .B1(n19701), .B2(n20112), .ZN(
        n19705) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19703), .B1(
        n20113), .B2(n19702), .ZN(n19704) );
  OAI211_X1 U22735 ( .C1(n20121), .C2(n19706), .A(n19705), .B(n19704), .ZN(
        P2_U3079) );
  NOR2_X1 U22736 ( .A1(n19769), .A2(n19829), .ZN(n19733) );
  AOI22_X1 U22737 ( .A1(n19992), .A2(n19758), .B1(n20060), .B2(n19733), .ZN(
        n19719) );
  OAI21_X1 U22738 ( .B1(n19758), .B2(n19734), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19707) );
  NAND2_X1 U22739 ( .A1(n19707), .A2(n20223), .ZN(n19717) );
  NAND2_X1 U22740 ( .A1(n19709), .A2(n19708), .ZN(n19949) );
  NOR2_X1 U22741 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19949), .ZN(
        n19713) );
  OAI21_X1 U22742 ( .B1(n19714), .B2(n20269), .A(n20268), .ZN(n19711) );
  INV_X1 U22743 ( .A(n19733), .ZN(n19710) );
  AOI21_X1 U22744 ( .B1(n19711), .B2(n19710), .A(n19775), .ZN(n19712) );
  INV_X1 U22745 ( .A(n19713), .ZN(n19716) );
  OAI21_X1 U22746 ( .B1(n19714), .B2(n19733), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19715) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19736), .B1(
        n20061), .B2(n19735), .ZN(n19718) );
  OAI211_X1 U22748 ( .C1(n19995), .C2(n19732), .A(n19719), .B(n19718), .ZN(
        P2_U3080) );
  AOI22_X1 U22749 ( .A1(n20032), .A2(n19734), .B1(n20073), .B2(n19733), .ZN(
        n19721) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19736), .B1(
        n20074), .B2(n19735), .ZN(n19720) );
  OAI211_X1 U22751 ( .C1(n20035), .C2(n19766), .A(n19721), .B(n19720), .ZN(
        P2_U3081) );
  AOI22_X1 U22752 ( .A1(n20081), .A2(n19758), .B1(n19733), .B2(n20079), .ZN(
        n19723) );
  AOI22_X1 U22753 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19736), .B1(
        n20080), .B2(n19735), .ZN(n19722) );
  OAI211_X1 U22754 ( .C1(n20084), .C2(n19732), .A(n19723), .B(n19722), .ZN(
        P2_U3082) );
  AOI22_X1 U22755 ( .A1(n19965), .A2(n19734), .B1(n20085), .B2(n19733), .ZN(
        n19725) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19736), .B1(
        n20086), .B2(n19735), .ZN(n19724) );
  OAI211_X1 U22757 ( .C1(n19968), .C2(n19766), .A(n19725), .B(n19724), .ZN(
        P2_U3083) );
  AOI22_X1 U22758 ( .A1(n20093), .A2(n19734), .B1(n20091), .B2(n19733), .ZN(
        n19727) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19736), .B1(
        n20092), .B2(n19735), .ZN(n19726) );
  OAI211_X1 U22760 ( .C1(n20096), .C2(n19766), .A(n19727), .B(n19726), .ZN(
        P2_U3084) );
  AOI22_X1 U22761 ( .A1(n20006), .A2(n19758), .B1(n20097), .B2(n19733), .ZN(
        n19729) );
  AOI22_X1 U22762 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19736), .B1(
        n20098), .B2(n19735), .ZN(n19728) );
  OAI211_X1 U22763 ( .C1(n20009), .C2(n19732), .A(n19729), .B(n19728), .ZN(
        P2_U3085) );
  AOI22_X1 U22764 ( .A1(n20010), .A2(n19758), .B1(n20103), .B2(n19733), .ZN(
        n19731) );
  AOI22_X1 U22765 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19736), .B1(
        n20104), .B2(n19735), .ZN(n19730) );
  OAI211_X1 U22766 ( .C1(n20013), .C2(n19732), .A(n19731), .B(n19730), .ZN(
        P2_U3086) );
  AOI22_X1 U22767 ( .A1(n20050), .A2(n19734), .B1(n20112), .B2(n19733), .ZN(
        n19738) );
  AOI22_X1 U22768 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19736), .B1(
        n20113), .B2(n19735), .ZN(n19737) );
  OAI211_X1 U22769 ( .C1(n20056), .C2(n19766), .A(n19738), .B(n19737), .ZN(
        P2_U3087) );
  NOR2_X1 U22770 ( .A1(n19769), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19741) );
  INV_X1 U22771 ( .A(n19741), .ZN(n19744) );
  NOR2_X1 U22772 ( .A1(n20263), .A2(n19744), .ZN(n19761) );
  AOI22_X1 U22773 ( .A1(n19992), .A2(n19793), .B1(n20060), .B2(n19761), .ZN(
        n19747) );
  OAI21_X1 U22774 ( .B1(n19801), .B2(n19990), .A(n20223), .ZN(n19745) );
  INV_X1 U22775 ( .A(n19761), .ZN(n19739) );
  OAI211_X1 U22776 ( .C1(n10631), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20232), 
        .B(n19739), .ZN(n19740) );
  OAI211_X1 U22777 ( .C1(n19745), .C2(n19741), .A(n20067), .B(n19740), .ZN(
        n19763) );
  OAI21_X1 U22778 ( .B1(n19742), .B2(n19761), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19743) );
  OAI21_X1 U22779 ( .B1(n19745), .B2(n19744), .A(n19743), .ZN(n19762) );
  AOI22_X1 U22780 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19763), .B1(
        n20061), .B2(n19762), .ZN(n19746) );
  OAI211_X1 U22781 ( .C1(n19995), .C2(n19766), .A(n19747), .B(n19746), .ZN(
        P2_U3088) );
  AOI22_X1 U22782 ( .A1(n20075), .A2(n19793), .B1(n20073), .B2(n19761), .ZN(
        n19749) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19763), .B1(
        n20074), .B2(n19762), .ZN(n19748) );
  OAI211_X1 U22784 ( .C1(n20078), .C2(n19766), .A(n19749), .B(n19748), .ZN(
        P2_U3089) );
  AOI22_X1 U22785 ( .A1(n20036), .A2(n19758), .B1(n20079), .B2(n19761), .ZN(
        n19751) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19763), .B1(
        n20080), .B2(n19762), .ZN(n19750) );
  OAI211_X1 U22787 ( .C1(n20039), .C2(n19770), .A(n19751), .B(n19750), .ZN(
        P2_U3090) );
  AOI22_X1 U22788 ( .A1(n19965), .A2(n19758), .B1(n20085), .B2(n19761), .ZN(
        n19753) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19763), .B1(
        n20086), .B2(n19762), .ZN(n19752) );
  OAI211_X1 U22790 ( .C1(n19968), .C2(n19770), .A(n19753), .B(n19752), .ZN(
        P2_U3091) );
  AOI22_X1 U22791 ( .A1(n20002), .A2(n19793), .B1(n20091), .B2(n19761), .ZN(
        n19755) );
  AOI22_X1 U22792 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19763), .B1(
        n20092), .B2(n19762), .ZN(n19754) );
  OAI211_X1 U22793 ( .C1(n20005), .C2(n19766), .A(n19755), .B(n19754), .ZN(
        P2_U3092) );
  AOI22_X1 U22794 ( .A1(n20006), .A2(n19793), .B1(n20097), .B2(n19761), .ZN(
        n19757) );
  AOI22_X1 U22795 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19763), .B1(
        n20098), .B2(n19762), .ZN(n19756) );
  OAI211_X1 U22796 ( .C1(n20009), .C2(n19766), .A(n19757), .B(n19756), .ZN(
        P2_U3093) );
  AOI22_X1 U22797 ( .A1(n20105), .A2(n19758), .B1(n20103), .B2(n19761), .ZN(
        n19760) );
  AOI22_X1 U22798 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19763), .B1(
        n20104), .B2(n19762), .ZN(n19759) );
  OAI211_X1 U22799 ( .C1(n20110), .C2(n19770), .A(n19760), .B(n19759), .ZN(
        P2_U3094) );
  AOI22_X1 U22800 ( .A1(n20115), .A2(n19793), .B1(n20112), .B2(n19761), .ZN(
        n19765) );
  AOI22_X1 U22801 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19763), .B1(
        n20113), .B2(n19762), .ZN(n19764) );
  OAI211_X1 U22802 ( .C1(n20121), .C2(n19766), .A(n19765), .B(n19764), .ZN(
        P2_U3095) );
  NOR3_X2 U22803 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20057), .ZN(n19791) );
  OAI21_X1 U22804 ( .B1(n10622), .B2(n19791), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19768) );
  OAI21_X1 U22805 ( .B1(n19769), .B2(n19892), .A(n19768), .ZN(n19792) );
  AOI22_X1 U22806 ( .A1(n19792), .A2(n20061), .B1(n20060), .B2(n19791), .ZN(
        n19778) );
  AOI21_X1 U22807 ( .B1(n19770), .B2(n19826), .A(n19952), .ZN(n19771) );
  AOI21_X1 U22808 ( .B1(n19773), .B2(n19772), .A(n19771), .ZN(n19776) );
  AOI211_X1 U22809 ( .C1(n10622), .C2(n20268), .A(n20223), .B(n19791), .ZN(
        n19774) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n20069), .ZN(n19777) );
  OAI211_X1 U22811 ( .C1(n20072), .C2(n19826), .A(n19778), .B(n19777), .ZN(
        P2_U3096) );
  AOI22_X1 U22812 ( .A1(n19792), .A2(n20074), .B1(n20073), .B2(n19791), .ZN(
        n19780) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n20032), .ZN(n19779) );
  OAI211_X1 U22814 ( .C1(n20035), .C2(n19826), .A(n19780), .B(n19779), .ZN(
        P2_U3097) );
  AOI22_X1 U22815 ( .A1(n19792), .A2(n20080), .B1(n20079), .B2(n19791), .ZN(
        n19782) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n20036), .ZN(n19781) );
  OAI211_X1 U22817 ( .C1(n20039), .C2(n19826), .A(n19782), .B(n19781), .ZN(
        P2_U3098) );
  AOI22_X1 U22818 ( .A1(n19792), .A2(n20086), .B1(n20085), .B2(n19791), .ZN(
        n19784) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n19965), .ZN(n19783) );
  OAI211_X1 U22820 ( .C1(n19968), .C2(n19826), .A(n19784), .B(n19783), .ZN(
        P2_U3099) );
  AOI22_X1 U22821 ( .A1(n19792), .A2(n20092), .B1(n20091), .B2(n19791), .ZN(
        n19786) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n20093), .ZN(n19785) );
  OAI211_X1 U22823 ( .C1(n20096), .C2(n19826), .A(n19786), .B(n19785), .ZN(
        P2_U3100) );
  AOI22_X1 U22824 ( .A1(n19792), .A2(n20098), .B1(n20097), .B2(n19791), .ZN(
        n19788) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n20099), .ZN(n19787) );
  OAI211_X1 U22826 ( .C1(n20102), .C2(n19826), .A(n19788), .B(n19787), .ZN(
        P2_U3101) );
  AOI22_X1 U22827 ( .A1(n19792), .A2(n20104), .B1(n20103), .B2(n19791), .ZN(
        n19790) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n20105), .ZN(n19789) );
  OAI211_X1 U22829 ( .C1(n20110), .C2(n19826), .A(n19790), .B(n19789), .ZN(
        P2_U3102) );
  AOI22_X1 U22830 ( .A1(n19792), .A2(n20113), .B1(n20112), .B2(n19791), .ZN(
        n19796) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19794), .B1(
        n19793), .B2(n20050), .ZN(n19795) );
  OAI211_X1 U22832 ( .C1(n20056), .C2(n19826), .A(n19796), .B(n19795), .ZN(
        P2_U3103) );
  OR2_X1 U22833 ( .A1(n20057), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19803) );
  AND2_X1 U22834 ( .A1(n19832), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19797) );
  NAND2_X1 U22835 ( .A1(n19798), .A2(n19797), .ZN(n19805) );
  INV_X1 U22836 ( .A(n19805), .ZN(n19799) );
  AOI211_X2 U22837 ( .C1(n19803), .C2(n20269), .A(n19800), .B(n19799), .ZN(
        n19822) );
  INV_X1 U22838 ( .A(n19832), .ZN(n19835) );
  AOI22_X1 U22839 ( .A1(n19822), .A2(n20061), .B1(n19835), .B2(n20060), .ZN(
        n19809) );
  OR2_X1 U22840 ( .A1(n19802), .A2(n19801), .ZN(n20233) );
  NAND2_X1 U22841 ( .A1(n20233), .A2(n19803), .ZN(n19806) );
  NAND2_X1 U22842 ( .A1(n19832), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19804) );
  NAND4_X1 U22843 ( .A1(n19806), .A2(n20067), .A3(n19805), .A4(n19804), .ZN(
        n19823) );
  NAND2_X1 U22844 ( .A1(n19807), .A2(n20062), .ZN(n19851) );
  AOI22_X1 U22845 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n19992), .ZN(n19808) );
  OAI211_X1 U22846 ( .C1(n19995), .C2(n19826), .A(n19809), .B(n19808), .ZN(
        P2_U3104) );
  AOI22_X1 U22847 ( .A1(n19822), .A2(n20074), .B1(n19835), .B2(n20073), .ZN(
        n19811) );
  AOI22_X1 U22848 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n20075), .ZN(n19810) );
  OAI211_X1 U22849 ( .C1(n20078), .C2(n19826), .A(n19811), .B(n19810), .ZN(
        P2_U3105) );
  AOI22_X1 U22850 ( .A1(n19822), .A2(n20080), .B1(n19835), .B2(n20079), .ZN(
        n19813) );
  AOI22_X1 U22851 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n20081), .ZN(n19812) );
  OAI211_X1 U22852 ( .C1(n20084), .C2(n19826), .A(n19813), .B(n19812), .ZN(
        P2_U3106) );
  AOI22_X1 U22853 ( .A1(n19822), .A2(n20086), .B1(n19835), .B2(n20085), .ZN(
        n19815) );
  AOI22_X1 U22854 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n20087), .ZN(n19814) );
  OAI211_X1 U22855 ( .C1(n20090), .C2(n19826), .A(n19815), .B(n19814), .ZN(
        P2_U3107) );
  AOI22_X1 U22856 ( .A1(n19822), .A2(n20092), .B1(n19835), .B2(n20091), .ZN(
        n19817) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n20002), .ZN(n19816) );
  OAI211_X1 U22858 ( .C1(n20005), .C2(n19826), .A(n19817), .B(n19816), .ZN(
        P2_U3108) );
  AOI22_X1 U22859 ( .A1(n19822), .A2(n20098), .B1(n19835), .B2(n20097), .ZN(
        n19819) );
  AOI22_X1 U22860 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n20006), .ZN(n19818) );
  OAI211_X1 U22861 ( .C1(n20009), .C2(n19826), .A(n19819), .B(n19818), .ZN(
        P2_U3109) );
  AOI22_X1 U22862 ( .A1(n19822), .A2(n20104), .B1(n19835), .B2(n20103), .ZN(
        n19821) );
  AOI22_X1 U22863 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n20010), .ZN(n19820) );
  OAI211_X1 U22864 ( .C1(n20013), .C2(n19826), .A(n19821), .B(n19820), .ZN(
        P2_U3110) );
  AOI22_X1 U22865 ( .A1(n19822), .A2(n20113), .B1(n19835), .B2(n20112), .ZN(
        n19825) );
  AOI22_X1 U22866 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19823), .B1(
        n19855), .B2(n20115), .ZN(n19824) );
  OAI211_X1 U22867 ( .C1(n20121), .C2(n19826), .A(n19825), .B(n19824), .ZN(
        P2_U3111) );
  NAND2_X1 U22868 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20243), .ZN(
        n19919) );
  NOR2_X1 U22869 ( .A1(n19829), .A2(n19919), .ZN(n19854) );
  AOI22_X1 U22870 ( .A1(n20069), .A2(n19855), .B1(n20060), .B2(n19854), .ZN(
        n19840) );
  NAND2_X1 U22871 ( .A1(n19882), .A2(n19851), .ZN(n19830) );
  AOI21_X1 U22872 ( .B1(n19830), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20232), 
        .ZN(n19834) );
  OAI21_X1 U22873 ( .B1(n19836), .B2(n20269), .A(n20268), .ZN(n19831) );
  AOI21_X1 U22874 ( .B1(n19834), .B2(n19832), .A(n19831), .ZN(n19833) );
  OAI21_X1 U22875 ( .B1(n19854), .B2(n19833), .A(n20067), .ZN(n19857) );
  OAI21_X1 U22876 ( .B1(n19835), .B2(n19854), .A(n19834), .ZN(n19838) );
  OAI21_X1 U22877 ( .B1(n19836), .B2(n19854), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19837) );
  NAND2_X1 U22878 ( .A1(n19838), .A2(n19837), .ZN(n19856) );
  AOI22_X1 U22879 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19857), .B1(
        n20061), .B2(n19856), .ZN(n19839) );
  OAI211_X1 U22880 ( .C1(n20072), .C2(n19882), .A(n19840), .B(n19839), .ZN(
        P2_U3112) );
  AOI22_X1 U22881 ( .A1(n20032), .A2(n19855), .B1(n20073), .B2(n19854), .ZN(
        n19842) );
  AOI22_X1 U22882 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19857), .B1(
        n20074), .B2(n19856), .ZN(n19841) );
  OAI211_X1 U22883 ( .C1(n20035), .C2(n19882), .A(n19842), .B(n19841), .ZN(
        P2_U3113) );
  INV_X1 U22884 ( .A(n19882), .ZN(n19885) );
  AOI22_X1 U22885 ( .A1(n20081), .A2(n19885), .B1(n20079), .B2(n19854), .ZN(
        n19844) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19857), .B1(
        n20080), .B2(n19856), .ZN(n19843) );
  OAI211_X1 U22887 ( .C1(n20084), .C2(n19851), .A(n19844), .B(n19843), .ZN(
        P2_U3114) );
  AOI22_X1 U22888 ( .A1(n19965), .A2(n19855), .B1(n20085), .B2(n19854), .ZN(
        n19846) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19857), .B1(
        n20086), .B2(n19856), .ZN(n19845) );
  OAI211_X1 U22890 ( .C1(n19968), .C2(n19882), .A(n19846), .B(n19845), .ZN(
        P2_U3115) );
  AOI22_X1 U22891 ( .A1(n20093), .A2(n19855), .B1(n20091), .B2(n19854), .ZN(
        n19848) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19857), .B1(
        n20092), .B2(n19856), .ZN(n19847) );
  OAI211_X1 U22893 ( .C1(n20096), .C2(n19882), .A(n19848), .B(n19847), .ZN(
        P2_U3116) );
  AOI22_X1 U22894 ( .A1(n20006), .A2(n19885), .B1(n20097), .B2(n19854), .ZN(
        n19850) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19857), .B1(
        n20098), .B2(n19856), .ZN(n19849) );
  OAI211_X1 U22896 ( .C1(n20009), .C2(n19851), .A(n19850), .B(n19849), .ZN(
        P2_U3117) );
  AOI22_X1 U22897 ( .A1(n20105), .A2(n19855), .B1(n20103), .B2(n19854), .ZN(
        n19853) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19857), .B1(
        n20104), .B2(n19856), .ZN(n19852) );
  OAI211_X1 U22899 ( .C1(n20110), .C2(n19882), .A(n19853), .B(n19852), .ZN(
        P2_U3118) );
  AOI22_X1 U22900 ( .A1(n20050), .A2(n19855), .B1(n20112), .B2(n19854), .ZN(
        n19859) );
  AOI22_X1 U22901 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19857), .B1(
        n20113), .B2(n19856), .ZN(n19858) );
  OAI211_X1 U22902 ( .C1(n20056), .C2(n19882), .A(n19859), .B(n19858), .ZN(
        P2_U3119) );
  INV_X1 U22903 ( .A(n19915), .ZN(n19890) );
  NOR3_X2 U22904 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20263), .A3(
        n19919), .ZN(n19893) );
  AOI22_X1 U22905 ( .A1(n20069), .A2(n19885), .B1(n20060), .B2(n19893), .ZN(
        n19871) );
  INV_X1 U22906 ( .A(n19860), .ZN(n20229) );
  NAND2_X1 U22907 ( .A1(n20229), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19987) );
  OAI21_X1 U22908 ( .B1(n19987), .B2(n19861), .A(n20223), .ZN(n19869) );
  NOR2_X1 U22909 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19919), .ZN(
        n19864) );
  INV_X1 U22910 ( .A(n19893), .ZN(n19862) );
  OAI211_X1 U22911 ( .C1(n19865), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20232), 
        .B(n19862), .ZN(n19863) );
  OAI211_X1 U22912 ( .C1(n19869), .C2(n19864), .A(n20067), .B(n19863), .ZN(
        n19887) );
  INV_X1 U22913 ( .A(n19864), .ZN(n19868) );
  INV_X1 U22914 ( .A(n19865), .ZN(n19866) );
  OAI21_X1 U22915 ( .B1(n19866), .B2(n19893), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19867) );
  OAI21_X1 U22916 ( .B1(n19869), .B2(n19868), .A(n19867), .ZN(n19886) );
  AOI22_X1 U22917 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19887), .B1(
        n20061), .B2(n19886), .ZN(n19870) );
  OAI211_X1 U22918 ( .C1(n20072), .C2(n19890), .A(n19871), .B(n19870), .ZN(
        P2_U3120) );
  AOI22_X1 U22919 ( .A1(n19915), .A2(n20075), .B1(n20073), .B2(n19893), .ZN(
        n19873) );
  AOI22_X1 U22920 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19887), .B1(
        n20074), .B2(n19886), .ZN(n19872) );
  OAI211_X1 U22921 ( .C1(n20078), .C2(n19882), .A(n19873), .B(n19872), .ZN(
        P2_U3121) );
  AOI22_X1 U22922 ( .A1(n20036), .A2(n19885), .B1(n20079), .B2(n19893), .ZN(
        n19875) );
  AOI22_X1 U22923 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19887), .B1(
        n20080), .B2(n19886), .ZN(n19874) );
  OAI211_X1 U22924 ( .C1(n20039), .C2(n19890), .A(n19875), .B(n19874), .ZN(
        P2_U3122) );
  AOI22_X1 U22925 ( .A1(n19965), .A2(n19885), .B1(n20085), .B2(n19893), .ZN(
        n19877) );
  AOI22_X1 U22926 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19887), .B1(
        n20086), .B2(n19886), .ZN(n19876) );
  OAI211_X1 U22927 ( .C1(n19968), .C2(n19890), .A(n19877), .B(n19876), .ZN(
        P2_U3123) );
  AOI22_X1 U22928 ( .A1(n19915), .A2(n20002), .B1(n20091), .B2(n19893), .ZN(
        n19879) );
  AOI22_X1 U22929 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19887), .B1(
        n20092), .B2(n19886), .ZN(n19878) );
  OAI211_X1 U22930 ( .C1(n20005), .C2(n19882), .A(n19879), .B(n19878), .ZN(
        P2_U3124) );
  AOI22_X1 U22931 ( .A1(n19915), .A2(n20006), .B1(n20097), .B2(n19893), .ZN(
        n19881) );
  AOI22_X1 U22932 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19887), .B1(
        n20098), .B2(n19886), .ZN(n19880) );
  OAI211_X1 U22933 ( .C1(n20009), .C2(n19882), .A(n19881), .B(n19880), .ZN(
        P2_U3125) );
  AOI22_X1 U22934 ( .A1(n20105), .A2(n19885), .B1(n20103), .B2(n19893), .ZN(
        n19884) );
  AOI22_X1 U22935 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19887), .B1(
        n20104), .B2(n19886), .ZN(n19883) );
  OAI211_X1 U22936 ( .C1(n20110), .C2(n19890), .A(n19884), .B(n19883), .ZN(
        P2_U3126) );
  AOI22_X1 U22937 ( .A1(n20050), .A2(n19885), .B1(n20112), .B2(n19893), .ZN(
        n19889) );
  AOI22_X1 U22938 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19887), .B1(
        n20113), .B2(n19886), .ZN(n19888) );
  OAI211_X1 U22939 ( .C1(n20056), .C2(n19890), .A(n19889), .B(n19888), .ZN(
        P2_U3127) );
  NOR3_X2 U22940 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20252), .A3(
        n19919), .ZN(n19913) );
  OAI21_X1 U22941 ( .B1(n19894), .B2(n19913), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19891) );
  OAI21_X1 U22942 ( .B1(n19919), .B2(n19892), .A(n19891), .ZN(n19914) );
  AOI22_X1 U22943 ( .A1(n19914), .A2(n20061), .B1(n20060), .B2(n19913), .ZN(
        n19900) );
  INV_X1 U22944 ( .A(n19942), .ZN(n19945) );
  AOI221_X1 U22945 ( .B1(n19915), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19945), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19893), .ZN(n19896) );
  INV_X1 U22946 ( .A(n19894), .ZN(n19895) );
  MUX2_X1 U22947 ( .A(n19896), .B(n19895), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19897) );
  NOR2_X1 U22948 ( .A1(n19897), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19898) );
  AOI22_X1 U22949 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n20069), .ZN(n19899) );
  OAI211_X1 U22950 ( .C1(n20072), .C2(n19942), .A(n19900), .B(n19899), .ZN(
        P2_U3128) );
  AOI22_X1 U22951 ( .A1(n19914), .A2(n20074), .B1(n20073), .B2(n19913), .ZN(
        n19902) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n20032), .ZN(n19901) );
  OAI211_X1 U22953 ( .C1(n20035), .C2(n19942), .A(n19902), .B(n19901), .ZN(
        P2_U3129) );
  AOI22_X1 U22954 ( .A1(n19914), .A2(n20080), .B1(n20079), .B2(n19913), .ZN(
        n19904) );
  AOI22_X1 U22955 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n20036), .ZN(n19903) );
  OAI211_X1 U22956 ( .C1(n20039), .C2(n19942), .A(n19904), .B(n19903), .ZN(
        P2_U3130) );
  AOI22_X1 U22957 ( .A1(n19914), .A2(n20086), .B1(n20085), .B2(n19913), .ZN(
        n19906) );
  AOI22_X1 U22958 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19965), .ZN(n19905) );
  OAI211_X1 U22959 ( .C1(n19968), .C2(n19942), .A(n19906), .B(n19905), .ZN(
        P2_U3131) );
  AOI22_X1 U22960 ( .A1(n19914), .A2(n20092), .B1(n20091), .B2(n19913), .ZN(
        n19908) );
  AOI22_X1 U22961 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n20093), .ZN(n19907) );
  OAI211_X1 U22962 ( .C1(n20096), .C2(n19942), .A(n19908), .B(n19907), .ZN(
        P2_U3132) );
  AOI22_X1 U22963 ( .A1(n19914), .A2(n20098), .B1(n20097), .B2(n19913), .ZN(
        n19910) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n20099), .ZN(n19909) );
  OAI211_X1 U22965 ( .C1(n20102), .C2(n19942), .A(n19910), .B(n19909), .ZN(
        P2_U3133) );
  AOI22_X1 U22966 ( .A1(n19914), .A2(n20104), .B1(n20103), .B2(n19913), .ZN(
        n19912) );
  AOI22_X1 U22967 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n20105), .ZN(n19911) );
  OAI211_X1 U22968 ( .C1(n20110), .C2(n19942), .A(n19912), .B(n19911), .ZN(
        P2_U3134) );
  AOI22_X1 U22969 ( .A1(n19914), .A2(n20113), .B1(n20112), .B2(n19913), .ZN(
        n19918) );
  AOI22_X1 U22970 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n20050), .ZN(n19917) );
  OAI211_X1 U22971 ( .C1(n20056), .C2(n19942), .A(n19918), .B(n19917), .ZN(
        P2_U3135) );
  OR2_X1 U22972 ( .A1(n20252), .A2(n19919), .ZN(n19924) );
  OR2_X1 U22973 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19924), .ZN(n19922) );
  INV_X1 U22974 ( .A(n10628), .ZN(n19921) );
  NOR2_X1 U22975 ( .A1(n19920), .A2(n19919), .ZN(n19943) );
  NOR3_X1 U22976 ( .A1(n19921), .A2(n19943), .A3(n20269), .ZN(n19923) );
  AOI21_X1 U22977 ( .B1(n20269), .B2(n19922), .A(n19923), .ZN(n19944) );
  AOI22_X1 U22978 ( .A1(n19944), .A2(n20061), .B1(n20060), .B2(n19943), .ZN(
        n19929) );
  INV_X1 U22979 ( .A(n19987), .ZN(n20063) );
  NAND2_X1 U22980 ( .A1(n20063), .A2(n20224), .ZN(n19925) );
  AOI21_X1 U22981 ( .B1(n19925), .B2(n19924), .A(n19923), .ZN(n19926) );
  OAI211_X1 U22982 ( .C1(n19943), .C2(n20268), .A(n19926), .B(n20067), .ZN(
        n19946) );
  NAND2_X1 U22983 ( .A1(n19927), .A2(n20224), .ZN(n19953) );
  AOI22_X1 U22984 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19946), .B1(
        n19977), .B2(n19992), .ZN(n19928) );
  OAI211_X1 U22985 ( .C1(n19995), .C2(n19942), .A(n19929), .B(n19928), .ZN(
        P2_U3136) );
  AOI22_X1 U22986 ( .A1(n19944), .A2(n20074), .B1(n20073), .B2(n19943), .ZN(
        n19931) );
  AOI22_X1 U22987 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n20032), .ZN(n19930) );
  OAI211_X1 U22988 ( .C1(n20035), .C2(n19953), .A(n19931), .B(n19930), .ZN(
        P2_U3137) );
  AOI22_X1 U22989 ( .A1(n19944), .A2(n20080), .B1(n20079), .B2(n19943), .ZN(
        n19933) );
  AOI22_X1 U22990 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19946), .B1(
        n19977), .B2(n20081), .ZN(n19932) );
  OAI211_X1 U22991 ( .C1(n20084), .C2(n19942), .A(n19933), .B(n19932), .ZN(
        P2_U3138) );
  AOI22_X1 U22992 ( .A1(n19944), .A2(n20086), .B1(n20085), .B2(n19943), .ZN(
        n19935) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19946), .B1(
        n19977), .B2(n20087), .ZN(n19934) );
  OAI211_X1 U22994 ( .C1(n20090), .C2(n19942), .A(n19935), .B(n19934), .ZN(
        P2_U3139) );
  AOI22_X1 U22995 ( .A1(n19944), .A2(n20092), .B1(n20091), .B2(n19943), .ZN(
        n19937) );
  AOI22_X1 U22996 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n20093), .ZN(n19936) );
  OAI211_X1 U22997 ( .C1(n20096), .C2(n19953), .A(n19937), .B(n19936), .ZN(
        P2_U3140) );
  AOI22_X1 U22998 ( .A1(n19944), .A2(n20098), .B1(n20097), .B2(n19943), .ZN(
        n19939) );
  AOI22_X1 U22999 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19946), .B1(
        n19977), .B2(n20006), .ZN(n19938) );
  OAI211_X1 U23000 ( .C1(n20009), .C2(n19942), .A(n19939), .B(n19938), .ZN(
        P2_U3141) );
  AOI22_X1 U23001 ( .A1(n19944), .A2(n20104), .B1(n20103), .B2(n19943), .ZN(
        n19941) );
  AOI22_X1 U23002 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19946), .B1(
        n19977), .B2(n20010), .ZN(n19940) );
  OAI211_X1 U23003 ( .C1(n20013), .C2(n19942), .A(n19941), .B(n19940), .ZN(
        P2_U3142) );
  AOI22_X1 U23004 ( .A1(n19944), .A2(n20113), .B1(n20112), .B2(n19943), .ZN(
        n19948) );
  AOI22_X1 U23005 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n20050), .ZN(n19947) );
  OAI211_X1 U23006 ( .C1(n20056), .C2(n19953), .A(n19948), .B(n19947), .ZN(
        P2_U3143) );
  NOR2_X1 U23007 ( .A1(n20236), .A2(n19949), .ZN(n19957) );
  INV_X1 U23008 ( .A(n19957), .ZN(n19951) );
  NAND3_X1 U23009 ( .A1(n20252), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19985) );
  NOR2_X1 U23010 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19985), .ZN(
        n19975) );
  OAI21_X1 U23011 ( .B1(n10636), .B2(n19975), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19950) );
  OAI21_X1 U23012 ( .B1(n19951), .B2(n20232), .A(n19950), .ZN(n19976) );
  AOI22_X1 U23013 ( .A1(n19976), .A2(n20061), .B1(n20060), .B2(n19975), .ZN(
        n19960) );
  AOI21_X1 U23014 ( .B1(n20018), .B2(n19953), .A(n19952), .ZN(n19958) );
  INV_X1 U23015 ( .A(n19975), .ZN(n19954) );
  OAI211_X1 U23016 ( .C1(n19955), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20232), 
        .B(n19954), .ZN(n19956) );
  OAI211_X1 U23017 ( .C1(n19958), .C2(n19957), .A(n20067), .B(n19956), .ZN(
        n19978) );
  AOI22_X1 U23018 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n20069), .ZN(n19959) );
  OAI211_X1 U23019 ( .C1(n20072), .C2(n20018), .A(n19960), .B(n19959), .ZN(
        P2_U3144) );
  AOI22_X1 U23020 ( .A1(n19976), .A2(n20074), .B1(n20073), .B2(n19975), .ZN(
        n19962) );
  AOI22_X1 U23021 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n20032), .ZN(n19961) );
  OAI211_X1 U23022 ( .C1(n20035), .C2(n20018), .A(n19962), .B(n19961), .ZN(
        P2_U3145) );
  AOI22_X1 U23023 ( .A1(n19976), .A2(n20080), .B1(n20079), .B2(n19975), .ZN(
        n19964) );
  AOI22_X1 U23024 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n20036), .ZN(n19963) );
  OAI211_X1 U23025 ( .C1(n20039), .C2(n20018), .A(n19964), .B(n19963), .ZN(
        P2_U3146) );
  AOI22_X1 U23026 ( .A1(n19976), .A2(n20086), .B1(n20085), .B2(n19975), .ZN(
        n19967) );
  AOI22_X1 U23027 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n19965), .ZN(n19966) );
  OAI211_X1 U23028 ( .C1(n19968), .C2(n20018), .A(n19967), .B(n19966), .ZN(
        P2_U3147) );
  AOI22_X1 U23029 ( .A1(n19976), .A2(n20092), .B1(n20091), .B2(n19975), .ZN(
        n19970) );
  AOI22_X1 U23030 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n20093), .ZN(n19969) );
  OAI211_X1 U23031 ( .C1(n20096), .C2(n20018), .A(n19970), .B(n19969), .ZN(
        P2_U3148) );
  AOI22_X1 U23032 ( .A1(n19976), .A2(n20098), .B1(n20097), .B2(n19975), .ZN(
        n19972) );
  AOI22_X1 U23033 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n20099), .ZN(n19971) );
  OAI211_X1 U23034 ( .C1(n20102), .C2(n20018), .A(n19972), .B(n19971), .ZN(
        P2_U3149) );
  AOI22_X1 U23035 ( .A1(n19976), .A2(n20104), .B1(n20103), .B2(n19975), .ZN(
        n19974) );
  AOI22_X1 U23036 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n20105), .ZN(n19973) );
  OAI211_X1 U23037 ( .C1(n20110), .C2(n20018), .A(n19974), .B(n19973), .ZN(
        P2_U3150) );
  AOI22_X1 U23038 ( .A1(n19976), .A2(n20113), .B1(n20112), .B2(n19975), .ZN(
        n19980) );
  AOI22_X1 U23039 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19978), .B1(
        n19977), .B2(n20050), .ZN(n19979) );
  OAI211_X1 U23040 ( .C1(n20056), .C2(n20018), .A(n19980), .B(n19979), .ZN(
        P2_U3151) );
  NOR2_X1 U23041 ( .A1(n20263), .A2(n19985), .ZN(n20021) );
  INV_X1 U23042 ( .A(n20021), .ZN(n19981) );
  NAND3_X1 U23043 ( .A1(n19982), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19981), 
        .ZN(n19988) );
  OAI21_X1 U23044 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19985), .A(n20269), 
        .ZN(n19983) );
  AOI22_X1 U23045 ( .A1(n20014), .A2(n20061), .B1(n20060), .B2(n20021), .ZN(
        n19994) );
  NAND2_X1 U23046 ( .A1(n19984), .A2(n20268), .ZN(n19986) );
  NOR2_X1 U23047 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20268), .ZN(
        n20258) );
  OAI22_X1 U23048 ( .A1(n19987), .A2(n19986), .B1(n20258), .B2(n19985), .ZN(
        n19989) );
  NAND3_X1 U23049 ( .A1(n19989), .A2(n20067), .A3(n19988), .ZN(n20015) );
  AOI22_X1 U23050 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n19992), .ZN(n19993) );
  OAI211_X1 U23051 ( .C1(n19995), .C2(n20018), .A(n19994), .B(n19993), .ZN(
        P2_U3152) );
  AOI22_X1 U23052 ( .A1(n20014), .A2(n20074), .B1(n20073), .B2(n20021), .ZN(
        n19997) );
  AOI22_X1 U23053 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n20075), .ZN(n19996) );
  OAI211_X1 U23054 ( .C1(n20078), .C2(n20018), .A(n19997), .B(n19996), .ZN(
        P2_U3153) );
  AOI22_X1 U23055 ( .A1(n20014), .A2(n20080), .B1(n20079), .B2(n20021), .ZN(
        n19999) );
  AOI22_X1 U23056 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n20081), .ZN(n19998) );
  OAI211_X1 U23057 ( .C1(n20084), .C2(n20018), .A(n19999), .B(n19998), .ZN(
        P2_U3154) );
  AOI22_X1 U23058 ( .A1(n20014), .A2(n20086), .B1(n20085), .B2(n20021), .ZN(
        n20001) );
  AOI22_X1 U23059 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n20087), .ZN(n20000) );
  OAI211_X1 U23060 ( .C1(n20090), .C2(n20018), .A(n20001), .B(n20000), .ZN(
        P2_U3155) );
  AOI22_X1 U23061 ( .A1(n20014), .A2(n20092), .B1(n20091), .B2(n20021), .ZN(
        n20004) );
  AOI22_X1 U23062 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n20002), .ZN(n20003) );
  OAI211_X1 U23063 ( .C1(n20005), .C2(n20018), .A(n20004), .B(n20003), .ZN(
        P2_U3156) );
  AOI22_X1 U23064 ( .A1(n20014), .A2(n20098), .B1(n20097), .B2(n20021), .ZN(
        n20008) );
  AOI22_X1 U23065 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n20006), .ZN(n20007) );
  OAI211_X1 U23066 ( .C1(n20009), .C2(n20018), .A(n20008), .B(n20007), .ZN(
        P2_U3157) );
  AOI22_X1 U23067 ( .A1(n20014), .A2(n20104), .B1(n20103), .B2(n20021), .ZN(
        n20012) );
  AOI22_X1 U23068 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n20010), .ZN(n20011) );
  OAI211_X1 U23069 ( .C1(n20013), .C2(n20018), .A(n20012), .B(n20011), .ZN(
        P2_U3158) );
  AOI22_X1 U23070 ( .A1(n20014), .A2(n20113), .B1(n20112), .B2(n20021), .ZN(
        n20017) );
  AOI22_X1 U23071 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20015), .B1(
        n20051), .B2(n20115), .ZN(n20016) );
  OAI211_X1 U23072 ( .C1(n20121), .C2(n20018), .A(n20017), .B(n20016), .ZN(
        P2_U3159) );
  NOR3_X2 U23073 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20236), .A3(
        n20057), .ZN(n20049) );
  AOI22_X1 U23074 ( .A1(n20051), .A2(n20069), .B1(n20060), .B2(n20049), .ZN(
        n20031) );
  OAI21_X1 U23075 ( .B1(n20051), .B2(n20106), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20020) );
  NAND2_X1 U23076 ( .A1(n20020), .A2(n20223), .ZN(n20029) );
  NOR2_X1 U23077 ( .A1(n20049), .A2(n20021), .ZN(n20028) );
  INV_X1 U23078 ( .A(n20028), .ZN(n20025) );
  INV_X1 U23079 ( .A(n20026), .ZN(n20023) );
  INV_X1 U23080 ( .A(n20049), .ZN(n20022) );
  OAI211_X1 U23081 ( .C1(n20023), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20232), 
        .B(n20022), .ZN(n20024) );
  OAI211_X1 U23082 ( .C1(n20029), .C2(n20025), .A(n20067), .B(n20024), .ZN(
        n20053) );
  OAI21_X1 U23083 ( .B1(n20026), .B2(n20049), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20027) );
  AOI22_X1 U23084 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20053), .B1(
        n20061), .B2(n20052), .ZN(n20030) );
  OAI211_X1 U23085 ( .C1(n20072), .C2(n20120), .A(n20031), .B(n20030), .ZN(
        P2_U3160) );
  AOI22_X1 U23086 ( .A1(n20051), .A2(n20032), .B1(n20073), .B2(n20049), .ZN(
        n20034) );
  AOI22_X1 U23087 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20053), .B1(
        n20074), .B2(n20052), .ZN(n20033) );
  OAI211_X1 U23088 ( .C1(n20035), .C2(n20120), .A(n20034), .B(n20033), .ZN(
        P2_U3161) );
  AOI22_X1 U23089 ( .A1(n20051), .A2(n20036), .B1(n20079), .B2(n20049), .ZN(
        n20038) );
  AOI22_X1 U23090 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20053), .B1(
        n20080), .B2(n20052), .ZN(n20037) );
  OAI211_X1 U23091 ( .C1(n20039), .C2(n20120), .A(n20038), .B(n20037), .ZN(
        P2_U3162) );
  INV_X1 U23092 ( .A(n20051), .ZN(n20042) );
  AOI22_X1 U23093 ( .A1(n20087), .A2(n20106), .B1(n20085), .B2(n20049), .ZN(
        n20041) );
  AOI22_X1 U23094 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20053), .B1(
        n20086), .B2(n20052), .ZN(n20040) );
  OAI211_X1 U23095 ( .C1(n20090), .C2(n20042), .A(n20041), .B(n20040), .ZN(
        P2_U3163) );
  AOI22_X1 U23096 ( .A1(n20051), .A2(n20093), .B1(n20091), .B2(n20049), .ZN(
        n20044) );
  AOI22_X1 U23097 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20053), .B1(
        n20092), .B2(n20052), .ZN(n20043) );
  OAI211_X1 U23098 ( .C1(n20096), .C2(n20120), .A(n20044), .B(n20043), .ZN(
        P2_U3164) );
  AOI22_X1 U23099 ( .A1(n20051), .A2(n20099), .B1(n20097), .B2(n20049), .ZN(
        n20046) );
  AOI22_X1 U23100 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20053), .B1(
        n20098), .B2(n20052), .ZN(n20045) );
  OAI211_X1 U23101 ( .C1(n20102), .C2(n20120), .A(n20046), .B(n20045), .ZN(
        P2_U3165) );
  AOI22_X1 U23102 ( .A1(n20051), .A2(n20105), .B1(n20103), .B2(n20049), .ZN(
        n20048) );
  AOI22_X1 U23103 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20053), .B1(
        n20104), .B2(n20052), .ZN(n20047) );
  OAI211_X1 U23104 ( .C1(n20110), .C2(n20120), .A(n20048), .B(n20047), .ZN(
        P2_U3166) );
  AOI22_X1 U23105 ( .A1(n20051), .A2(n20050), .B1(n20112), .B2(n20049), .ZN(
        n20055) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20053), .B1(
        n20113), .B2(n20052), .ZN(n20054) );
  OAI211_X1 U23107 ( .C1(n20056), .C2(n20120), .A(n20055), .B(n20054), .ZN(
        P2_U3167) );
  INV_X1 U23108 ( .A(n20116), .ZN(n20109) );
  OR2_X1 U23109 ( .A1(n20236), .A2(n20057), .ZN(n20065) );
  OR2_X1 U23110 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20065), .ZN(n20059) );
  NOR3_X1 U23111 ( .A1(n20058), .A2(n20111), .A3(n20269), .ZN(n20064) );
  AOI21_X1 U23112 ( .B1(n20269), .B2(n20059), .A(n20064), .ZN(n20114) );
  AOI22_X1 U23113 ( .A1(n20114), .A2(n20061), .B1(n20060), .B2(n20111), .ZN(
        n20071) );
  NAND2_X1 U23114 ( .A1(n20063), .A2(n20062), .ZN(n20066) );
  AOI21_X1 U23115 ( .B1(n20066), .B2(n20065), .A(n20064), .ZN(n20068) );
  OAI211_X1 U23116 ( .C1(n20111), .C2(n20268), .A(n20068), .B(n20067), .ZN(
        n20117) );
  AOI22_X1 U23117 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20117), .B1(
        n20106), .B2(n20069), .ZN(n20070) );
  OAI211_X1 U23118 ( .C1(n20072), .C2(n20109), .A(n20071), .B(n20070), .ZN(
        P2_U3168) );
  AOI22_X1 U23119 ( .A1(n20114), .A2(n20074), .B1(n20073), .B2(n20111), .ZN(
        n20077) );
  AOI22_X1 U23120 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20075), .ZN(n20076) );
  OAI211_X1 U23121 ( .C1(n20078), .C2(n20120), .A(n20077), .B(n20076), .ZN(
        P2_U3169) );
  AOI22_X1 U23122 ( .A1(n20114), .A2(n20080), .B1(n20079), .B2(n20111), .ZN(
        n20083) );
  AOI22_X1 U23123 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20081), .ZN(n20082) );
  OAI211_X1 U23124 ( .C1(n20084), .C2(n20120), .A(n20083), .B(n20082), .ZN(
        P2_U3170) );
  AOI22_X1 U23125 ( .A1(n20114), .A2(n20086), .B1(n20085), .B2(n20111), .ZN(
        n20089) );
  AOI22_X1 U23126 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20087), .ZN(n20088) );
  OAI211_X1 U23127 ( .C1(n20090), .C2(n20120), .A(n20089), .B(n20088), .ZN(
        P2_U3171) );
  AOI22_X1 U23128 ( .A1(n20114), .A2(n20092), .B1(n20091), .B2(n20111), .ZN(
        n20095) );
  AOI22_X1 U23129 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20117), .B1(
        n20106), .B2(n20093), .ZN(n20094) );
  OAI211_X1 U23130 ( .C1(n20096), .C2(n20109), .A(n20095), .B(n20094), .ZN(
        P2_U3172) );
  AOI22_X1 U23131 ( .A1(n20114), .A2(n20098), .B1(n20097), .B2(n20111), .ZN(
        n20101) );
  AOI22_X1 U23132 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20117), .B1(
        n20106), .B2(n20099), .ZN(n20100) );
  OAI211_X1 U23133 ( .C1(n20102), .C2(n20109), .A(n20101), .B(n20100), .ZN(
        P2_U3173) );
  AOI22_X1 U23134 ( .A1(n20114), .A2(n20104), .B1(n20103), .B2(n20111), .ZN(
        n20108) );
  AOI22_X1 U23135 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20117), .B1(
        n20106), .B2(n20105), .ZN(n20107) );
  OAI211_X1 U23136 ( .C1(n20110), .C2(n20109), .A(n20108), .B(n20107), .ZN(
        P2_U3174) );
  AOI22_X1 U23137 ( .A1(n20114), .A2(n20113), .B1(n20112), .B2(n20111), .ZN(
        n20119) );
  AOI22_X1 U23138 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20115), .ZN(n20118) );
  OAI211_X1 U23139 ( .C1(n20121), .C2(n20120), .A(n20119), .B(n20118), .ZN(
        P2_U3175) );
  AOI21_X1 U23140 ( .B1(n20219), .B2(n20123), .A(n20122), .ZN(n20127) );
  OAI211_X1 U23141 ( .C1(n20128), .C2(n20124), .A(n20274), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20125) );
  OAI211_X1 U23142 ( .C1(n20128), .C2(n20127), .A(n20126), .B(n20125), .ZN(
        P2_U3177) );
  AND2_X1 U23143 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20129), .ZN(
        P2_U3179) );
  AND2_X1 U23144 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20129), .ZN(
        P2_U3180) );
  AND2_X1 U23145 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20129), .ZN(
        P2_U3181) );
  AND2_X1 U23146 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20129), .ZN(
        P2_U3182) );
  NOR2_X1 U23147 ( .A1(n20872), .A2(n20217), .ZN(P2_U3183) );
  AND2_X1 U23148 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20129), .ZN(
        P2_U3184) );
  AND2_X1 U23149 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20129), .ZN(
        P2_U3185) );
  AND2_X1 U23150 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20129), .ZN(
        P2_U3186) );
  AND2_X1 U23151 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20129), .ZN(
        P2_U3187) );
  AND2_X1 U23152 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20129), .ZN(
        P2_U3188) );
  AND2_X1 U23153 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20129), .ZN(
        P2_U3189) );
  AND2_X1 U23154 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20129), .ZN(
        P2_U3190) );
  AND2_X1 U23155 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20129), .ZN(
        P2_U3191) );
  AND2_X1 U23156 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20129), .ZN(
        P2_U3192) );
  AND2_X1 U23157 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20129), .ZN(
        P2_U3193) );
  AND2_X1 U23158 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20129), .ZN(
        P2_U3194) );
  AND2_X1 U23159 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20129), .ZN(
        P2_U3195) );
  AND2_X1 U23160 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20129), .ZN(
        P2_U3196) );
  AND2_X1 U23161 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20129), .ZN(
        P2_U3197) );
  AND2_X1 U23162 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20129), .ZN(
        P2_U3198) );
  AND2_X1 U23163 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20129), .ZN(
        P2_U3199) );
  AND2_X1 U23164 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20129), .ZN(
        P2_U3200) );
  AND2_X1 U23165 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20129), .ZN(P2_U3201) );
  AND2_X1 U23166 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20129), .ZN(P2_U3202) );
  AND2_X1 U23167 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20129), .ZN(P2_U3203) );
  AND2_X1 U23168 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20129), .ZN(P2_U3204) );
  NOR2_X1 U23169 ( .A1(n21025), .A2(n20217), .ZN(P2_U3205) );
  AND2_X1 U23170 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20129), .ZN(P2_U3206) );
  AND2_X1 U23171 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20129), .ZN(P2_U3207) );
  AND2_X1 U23172 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20129), .ZN(P2_U3208) );
  NOR2_X1 U23173 ( .A1(n20276), .A2(n20130), .ZN(n20142) );
  INV_X1 U23174 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20287) );
  OR3_X1 U23175 ( .A1(n20142), .A2(n20287), .A3(n20131), .ZN(n20133) );
  AOI211_X1 U23176 ( .C1(n20769), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n20143), .B(n20197), .ZN(n20132) );
  NOR2_X1 U23177 ( .A1(n20775), .A2(n20135), .ZN(n20148) );
  AOI211_X1 U23178 ( .C1(n20149), .C2(n20133), .A(n20132), .B(n20148), .ZN(
        n20134) );
  INV_X1 U23179 ( .A(n20134), .ZN(P2_U3209) );
  AOI21_X1 U23180 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20769), .A(n20149), 
        .ZN(n20140) );
  NOR2_X1 U23181 ( .A1(n20287), .A2(n20140), .ZN(n20136) );
  AOI21_X1 U23182 ( .B1(n20136), .B2(n20135), .A(n20142), .ZN(n20138) );
  INV_X1 U23183 ( .A(n20280), .ZN(n20137) );
  OAI211_X1 U23184 ( .C1(n20769), .C2(n20139), .A(n20138), .B(n20137), .ZN(
        P2_U3210) );
  AOI21_X1 U23185 ( .B1(n20141), .B2(n20274), .A(n20140), .ZN(n20147) );
  AOI22_X1 U23186 ( .A1(n20287), .A2(n20143), .B1(n20775), .B2(n20142), .ZN(
        n20144) );
  INV_X1 U23187 ( .A(n20144), .ZN(n20145) );
  OAI211_X1 U23188 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20145), .ZN(n20146) );
  OAI21_X1 U23189 ( .B1(n20148), .B2(n20147), .A(n20146), .ZN(P2_U3211) );
  NAND2_X1 U23190 ( .A1(n20197), .A2(n20149), .ZN(n20207) );
  CLKBUF_X1 U23191 ( .A(n20207), .Z(n20202) );
  OAI222_X1 U23192 ( .A1(n20203), .A2(n20996), .B1(n20150), .B2(n20197), .C1(
        n20152), .C2(n20202), .ZN(P2_U3212) );
  OAI222_X1 U23193 ( .A1(n20203), .A2(n20152), .B1(n20151), .B2(n20197), .C1(
        n20154), .C2(n20202), .ZN(P2_U3213) );
  INV_X1 U23194 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20155) );
  OAI222_X1 U23195 ( .A1(n20203), .A2(n20154), .B1(n20153), .B2(n20197), .C1(
        n20155), .C2(n20202), .ZN(P2_U3214) );
  OAI222_X1 U23196 ( .A1(n20202), .A2(n20157), .B1(n20156), .B2(n20197), .C1(
        n20155), .C2(n20203), .ZN(P2_U3215) );
  OAI222_X1 U23197 ( .A1(n20207), .A2(n20159), .B1(n20158), .B2(n20197), .C1(
        n20157), .C2(n20203), .ZN(P2_U3216) );
  OAI222_X1 U23198 ( .A1(n20207), .A2(n13312), .B1(n20160), .B2(n20197), .C1(
        n20159), .C2(n20203), .ZN(P2_U3217) );
  OAI222_X1 U23199 ( .A1(n20207), .A2(n20162), .B1(n20161), .B2(n20197), .C1(
        n13312), .C2(n20203), .ZN(P2_U3218) );
  INV_X1 U23200 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20164) );
  OAI222_X1 U23201 ( .A1(n20207), .A2(n20164), .B1(n20163), .B2(n20197), .C1(
        n20162), .C2(n20203), .ZN(P2_U3219) );
  OAI222_X1 U23202 ( .A1(n20207), .A2(n20166), .B1(n20165), .B2(n20197), .C1(
        n20164), .C2(n20203), .ZN(P2_U3220) );
  OAI222_X1 U23203 ( .A1(n20202), .A2(n15205), .B1(n20167), .B2(n20197), .C1(
        n20166), .C2(n20203), .ZN(P2_U3221) );
  OAI222_X1 U23204 ( .A1(n20202), .A2(n13260), .B1(n20168), .B2(n20197), .C1(
        n15205), .C2(n20203), .ZN(P2_U3222) );
  OAI222_X1 U23205 ( .A1(n20202), .A2(n20170), .B1(n20169), .B2(n20197), .C1(
        n13260), .C2(n20203), .ZN(P2_U3223) );
  INV_X1 U23206 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20172) );
  OAI222_X1 U23207 ( .A1(n20202), .A2(n20172), .B1(n20171), .B2(n20197), .C1(
        n20170), .C2(n20203), .ZN(P2_U3224) );
  OAI222_X1 U23208 ( .A1(n20202), .A2(n20174), .B1(n20173), .B2(n20197), .C1(
        n20172), .C2(n20203), .ZN(P2_U3225) );
  OAI222_X1 U23209 ( .A1(n20202), .A2(n20176), .B1(n20175), .B2(n20197), .C1(
        n20174), .C2(n20203), .ZN(P2_U3226) );
  OAI222_X1 U23210 ( .A1(n20207), .A2(n20178), .B1(n20177), .B2(n20197), .C1(
        n20176), .C2(n20203), .ZN(P2_U3227) );
  OAI222_X1 U23211 ( .A1(n20207), .A2(n20180), .B1(n20179), .B2(n20197), .C1(
        n20178), .C2(n20203), .ZN(P2_U3228) );
  OAI222_X1 U23212 ( .A1(n20207), .A2(n15493), .B1(n20181), .B2(n20197), .C1(
        n20180), .C2(n20203), .ZN(P2_U3229) );
  OAI222_X1 U23213 ( .A1(n20207), .A2(n20183), .B1(n20182), .B2(n20197), .C1(
        n15493), .C2(n20203), .ZN(P2_U3230) );
  OAI222_X1 U23214 ( .A1(n20207), .A2(n20185), .B1(n20184), .B2(n20197), .C1(
        n20183), .C2(n20203), .ZN(P2_U3231) );
  OAI222_X1 U23215 ( .A1(n20207), .A2(n20187), .B1(n20186), .B2(n20197), .C1(
        n20185), .C2(n20203), .ZN(P2_U3232) );
  OAI222_X1 U23216 ( .A1(n20202), .A2(n20189), .B1(n20188), .B2(n20197), .C1(
        n20187), .C2(n20203), .ZN(P2_U3233) );
  OAI222_X1 U23217 ( .A1(n20202), .A2(n20191), .B1(n20190), .B2(n20197), .C1(
        n20189), .C2(n20203), .ZN(P2_U3234) );
  INV_X1 U23218 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20193) );
  OAI222_X1 U23219 ( .A1(n20202), .A2(n20193), .B1(n20192), .B2(n20197), .C1(
        n20191), .C2(n20203), .ZN(P2_U3235) );
  OAI222_X1 U23220 ( .A1(n20202), .A2(n20195), .B1(n20194), .B2(n20197), .C1(
        n20193), .C2(n20203), .ZN(P2_U3236) );
  OAI222_X1 U23221 ( .A1(n20202), .A2(n15394), .B1(n20196), .B2(n20197), .C1(
        n20195), .C2(n20203), .ZN(P2_U3237) );
  OAI222_X1 U23222 ( .A1(n20203), .A2(n15394), .B1(n20198), .B2(n20197), .C1(
        n20199), .C2(n20202), .ZN(P2_U3238) );
  OAI222_X1 U23223 ( .A1(n20202), .A2(n15383), .B1(n20200), .B2(n20197), .C1(
        n20199), .C2(n20203), .ZN(P2_U3239) );
  INV_X1 U23224 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20204) );
  OAI222_X1 U23225 ( .A1(n20202), .A2(n20204), .B1(n20201), .B2(n20197), .C1(
        n15383), .C2(n20203), .ZN(P2_U3240) );
  INV_X1 U23226 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20206) );
  OAI222_X1 U23227 ( .A1(n20207), .A2(n20206), .B1(n20205), .B2(n20197), .C1(
        n20204), .C2(n20203), .ZN(P2_U3241) );
  INV_X1 U23228 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U23229 ( .A1(n20197), .A2(n20209), .B1(n20208), .B2(n20289), .ZN(
        P2_U3585) );
  MUX2_X1 U23230 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20197), .Z(P2_U3586) );
  INV_X1 U23231 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20210) );
  AOI22_X1 U23232 ( .A1(n20197), .A2(n20211), .B1(n20210), .B2(n20289), .ZN(
        P2_U3587) );
  INV_X1 U23233 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20212) );
  AOI22_X1 U23234 ( .A1(n20197), .A2(n20213), .B1(n20212), .B2(n20289), .ZN(
        P2_U3588) );
  OAI21_X1 U23235 ( .B1(n20217), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20215), 
        .ZN(n20214) );
  INV_X1 U23236 ( .A(n20214), .ZN(P2_U3591) );
  OAI21_X1 U23237 ( .B1(n20217), .B2(n20216), .A(n20215), .ZN(P2_U3592) );
  NAND3_X1 U23238 ( .A1(n20222), .A2(n20219), .A3(n20218), .ZN(n20220) );
  OAI21_X1 U23239 ( .B1(n20222), .B2(n20221), .A(n20220), .ZN(P2_U3595) );
  AND2_X1 U23240 ( .A1(n20223), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20244) );
  NAND2_X1 U23241 ( .A1(n20224), .A2(n20244), .ZN(n20237) );
  NAND2_X1 U23242 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20225), .ZN(n20226) );
  OAI21_X1 U23243 ( .B1(n20227), .B2(n20226), .A(n20254), .ZN(n20238) );
  NAND2_X1 U23244 ( .A1(n20237), .A2(n20238), .ZN(n20230) );
  AOI22_X1 U23245 ( .A1(n20230), .A2(n20229), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20228), .ZN(n20231) );
  OAI21_X1 U23246 ( .B1(n20233), .B2(n20232), .A(n20231), .ZN(n20234) );
  INV_X1 U23247 ( .A(n20234), .ZN(n20235) );
  AOI22_X1 U23248 ( .A1(n20264), .A2(n20236), .B1(n20235), .B2(n20261), .ZN(
        P2_U3602) );
  OAI21_X1 U23249 ( .B1(n20239), .B2(n20238), .A(n20237), .ZN(n20240) );
  AOI21_X1 U23250 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20241), .A(n20240), 
        .ZN(n20242) );
  AOI22_X1 U23251 ( .A1(n20264), .A2(n20243), .B1(n20242), .B2(n20261), .ZN(
        P2_U3603) );
  INV_X1 U23252 ( .A(n20244), .ZN(n20247) );
  NAND3_X1 U23253 ( .A1(n20248), .A2(n20254), .A3(n20245), .ZN(n20246) );
  OAI21_X1 U23254 ( .B1(n20248), .B2(n20247), .A(n20246), .ZN(n20249) );
  AOI21_X1 U23255 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20250), .A(n20249), 
        .ZN(n20251) );
  AOI22_X1 U23256 ( .A1(n20264), .A2(n20252), .B1(n20251), .B2(n20261), .ZN(
        P2_U3604) );
  INV_X1 U23257 ( .A(n20253), .ZN(n20260) );
  INV_X1 U23258 ( .A(n20254), .ZN(n20255) );
  NOR2_X1 U23259 ( .A1(n20256), .A2(n20255), .ZN(n20257) );
  AOI211_X1 U23260 ( .C1(n20260), .C2(n20259), .A(n20258), .B(n20257), .ZN(
        n20262) );
  AOI22_X1 U23261 ( .A1(n20264), .A2(n20263), .B1(n20262), .B2(n20261), .ZN(
        P2_U3605) );
  INV_X1 U23262 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20265) );
  AOI22_X1 U23263 ( .A1(n20197), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20265), 
        .B2(n20289), .ZN(P2_U3608) );
  MUX2_X1 U23264 ( .A(P2_MORE_REG_SCAN_IN), .B(n20267), .S(n20266), .Z(
        P2_U3609) );
  OAI21_X1 U23265 ( .B1(n20270), .B2(n20269), .A(n20268), .ZN(n20271) );
  OAI211_X1 U23266 ( .C1(n20274), .C2(n20273), .A(n20272), .B(n20271), .ZN(
        n20288) );
  AOI21_X1 U23267 ( .B1(n20276), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n20275), 
        .ZN(n20285) );
  AOI21_X1 U23268 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20280), .A(n20277), 
        .ZN(n20283) );
  NOR3_X1 U23269 ( .A1(n20280), .A2(n20279), .A3(n20278), .ZN(n20282) );
  MUX2_X1 U23270 ( .A(n20283), .B(n20282), .S(n20281), .Z(n20284) );
  OAI21_X1 U23271 ( .B1(n20285), .B2(n20284), .A(n20288), .ZN(n20286) );
  OAI21_X1 U23272 ( .B1(n20288), .B2(n20287), .A(n20286), .ZN(P2_U3610) );
  INV_X1 U23273 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20290) );
  AOI22_X1 U23274 ( .A1(n20197), .A2(n20291), .B1(n20290), .B2(n20289), .ZN(
        P2_U3611) );
  OAI21_X1 U23275 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20763), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20778) );
  NOR2_X2 U23276 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20763), .ZN(n20866) );
  OAI21_X1 U23277 ( .B1(n20778), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20867), .ZN(
        n20292) );
  INV_X1 U23278 ( .A(n20292), .ZN(P1_U2802) );
  OAI21_X1 U23279 ( .B1(n20294), .B2(n20293), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20295) );
  OAI21_X1 U23280 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20296), .A(n20295), 
        .ZN(P1_U2803) );
  NOR2_X1 U23281 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20298) );
  OAI21_X1 U23282 ( .B1(n20298), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20867), .ZN(
        n20297) );
  OAI21_X1 U23283 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20867), .A(n20297), 
        .ZN(P1_U2804) );
  OAI21_X1 U23284 ( .B1(BS16), .B2(n20298), .A(n20845), .ZN(n20843) );
  OAI21_X1 U23285 ( .B1(n20845), .B2(n20702), .A(n20843), .ZN(P1_U2805) );
  OAI21_X1 U23286 ( .B1(n20301), .B2(n20300), .A(n20299), .ZN(P1_U2806) );
  NOR4_X1 U23287 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20305) );
  NOR4_X1 U23288 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20304) );
  NOR4_X1 U23289 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20303) );
  NOR4_X1 U23290 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20302) );
  NAND4_X1 U23291 ( .A1(n20305), .A2(n20304), .A3(n20303), .A4(n20302), .ZN(
        n20311) );
  NOR4_X1 U23292 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20309) );
  AOI211_X1 U23293 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20308) );
  NOR4_X1 U23294 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20307) );
  NOR4_X1 U23295 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20306) );
  NAND4_X1 U23296 ( .A1(n20309), .A2(n20308), .A3(n20307), .A4(n20306), .ZN(
        n20310) );
  NOR2_X1 U23297 ( .A1(n20311), .A2(n20310), .ZN(n20850) );
  INV_X1 U23298 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20838) );
  NOR3_X1 U23299 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20313) );
  OAI21_X1 U23300 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20313), .A(n20850), .ZN(
        n20312) );
  OAI21_X1 U23301 ( .B1(n20850), .B2(n20838), .A(n20312), .ZN(P1_U2807) );
  INV_X1 U23302 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20844) );
  AOI21_X1 U23303 ( .B1(n20846), .B2(n20844), .A(n20313), .ZN(n20314) );
  INV_X1 U23304 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20835) );
  INV_X1 U23305 ( .A(n20850), .ZN(n20852) );
  AOI22_X1 U23306 ( .A1(n20850), .A2(n20314), .B1(n20835), .B2(n20852), .ZN(
        P1_U2808) );
  OAI21_X1 U23307 ( .B1(n20316), .B2(n20315), .A(n16489), .ZN(n20319) );
  NOR2_X1 U23308 ( .A1(n20317), .A2(n20376), .ZN(n20318) );
  AOI211_X1 U23309 ( .C1(P1_EBX_REG_9__SCAN_IN), .C2(n20354), .A(n20319), .B(
        n20318), .ZN(n20328) );
  INV_X1 U23310 ( .A(n20320), .ZN(n20323) );
  AOI22_X1 U23311 ( .A1(n20323), .A2(n20348), .B1(n20322), .B2(n20321), .ZN(
        n20327) );
  OAI21_X1 U23312 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20325), .A(n20324), .ZN(
        n20326) );
  NAND3_X1 U23313 ( .A1(n20328), .A2(n20327), .A3(n20326), .ZN(P1_U2831) );
  NAND2_X1 U23314 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20330) );
  AOI21_X1 U23315 ( .B1(n20381), .B2(P1_REIP_REG_4__SCAN_IN), .A(n20329), .ZN(
        n20380) );
  AOI21_X1 U23316 ( .B1(n20331), .B2(n20330), .A(n20380), .ZN(n20344) );
  AOI22_X1 U23317 ( .A1(n20332), .A2(n20356), .B1(n20354), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20333) );
  OAI21_X1 U23318 ( .B1(n20334), .B2(n20384), .A(n20333), .ZN(n20335) );
  AOI211_X1 U23319 ( .C1(n20374), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16482), .B(n20335), .ZN(n20340) );
  NOR2_X1 U23320 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20336), .ZN(n20337) );
  AOI22_X1 U23321 ( .A1(n20338), .A2(n20348), .B1(n20381), .B2(n20337), .ZN(
        n20339) );
  OAI211_X1 U23322 ( .C1(n20344), .C2(n20790), .A(n20340), .B(n20339), .ZN(
        P1_U2833) );
  OAI22_X1 U23323 ( .A1(n20342), .A2(n20376), .B1(n20341), .B2(n20372), .ZN(
        n20343) );
  AOI211_X1 U23324 ( .C1(n20374), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16482), .B(n20343), .ZN(n20352) );
  INV_X1 U23325 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20788) );
  NAND2_X1 U23326 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20381), .ZN(n20363) );
  NOR2_X1 U23327 ( .A1(n20788), .A2(n20363), .ZN(n20346) );
  INV_X1 U23328 ( .A(n20344), .ZN(n20345) );
  MUX2_X1 U23329 ( .A(n20346), .B(n20345), .S(P1_REIP_REG_6__SCAN_IN), .Z(
        n20350) );
  AND2_X1 U23330 ( .A1(n20348), .A2(n20347), .ZN(n20349) );
  NOR2_X1 U23331 ( .A1(n20350), .A2(n20349), .ZN(n20351) );
  OAI211_X1 U23332 ( .C1(n20353), .C2(n20384), .A(n20352), .B(n20351), .ZN(
        P1_U2834) );
  AOI22_X1 U23333 ( .A1(n20356), .A2(n20355), .B1(n20354), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20357) );
  OAI21_X1 U23334 ( .B1(n20358), .B2(n20384), .A(n20357), .ZN(n20359) );
  AOI211_X1 U23335 ( .C1(n20374), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16482), .B(n20359), .ZN(n20362) );
  AOI22_X1 U23336 ( .A1(n20379), .A2(n20360), .B1(n20380), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20361) );
  OAI211_X1 U23337 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n20363), .A(n20362), .B(
        n20361), .ZN(P1_U2835) );
  NOR2_X1 U23338 ( .A1(n20365), .A2(n20364), .ZN(n20378) );
  INV_X1 U23339 ( .A(n20366), .ZN(n20367) );
  OAI21_X1 U23340 ( .B1(n20369), .B2(n20368), .A(n20367), .ZN(n20371) );
  NAND2_X1 U23341 ( .A1(n20371), .A2(n20370), .ZN(n20463) );
  NOR2_X1 U23342 ( .A1(n20372), .A2(n20389), .ZN(n20373) );
  AOI211_X1 U23343 ( .C1(n20374), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16482), .B(n20373), .ZN(n20375) );
  OAI21_X1 U23344 ( .B1(n20376), .B2(n20463), .A(n20375), .ZN(n20377) );
  AOI211_X1 U23345 ( .C1(n20379), .C2(n20455), .A(n20378), .B(n20377), .ZN(
        n20383) );
  OAI21_X1 U23346 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n20381), .A(n20380), .ZN(
        n20382) );
  OAI211_X1 U23347 ( .C1(n20384), .C2(n20460), .A(n20383), .B(n20382), .ZN(
        P1_U2836) );
  NOR2_X1 U23348 ( .A1(n20385), .A2(n20463), .ZN(n20386) );
  AOI21_X1 U23349 ( .B1(n20455), .B2(n20387), .A(n20386), .ZN(n20388) );
  OAI21_X1 U23350 ( .B1(n20390), .B2(n20389), .A(n20388), .ZN(P1_U2868) );
  INV_X1 U23351 ( .A(n20391), .ZN(n20393) );
  AOI22_X1 U23352 ( .A1(n20393), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20858), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20392) );
  OAI21_X1 U23353 ( .B1(n21046), .B2(n20395), .A(n20392), .ZN(P1_U2911) );
  AOI22_X1 U23354 ( .A1(n20393), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20858), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n20394) );
  OAI21_X1 U23355 ( .B1(n21011), .B2(n20395), .A(n20394), .ZN(P1_U2917) );
  AOI22_X1 U23356 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20397) );
  OAI21_X1 U23357 ( .B1(n12397), .B2(n20418), .A(n20397), .ZN(P1_U2921) );
  AOI22_X1 U23358 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20398) );
  OAI21_X1 U23359 ( .B1(n13805), .B2(n20418), .A(n20398), .ZN(P1_U2922) );
  AOI22_X1 U23360 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20399) );
  OAI21_X1 U23361 ( .B1(n13845), .B2(n20418), .A(n20399), .ZN(P1_U2923) );
  AOI22_X1 U23362 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20400) );
  OAI21_X1 U23363 ( .B1(n14746), .B2(n20418), .A(n20400), .ZN(P1_U2924) );
  AOI22_X1 U23364 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20401) );
  OAI21_X1 U23365 ( .B1(n13841), .B2(n20418), .A(n20401), .ZN(P1_U2925) );
  INV_X1 U23366 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20403) );
  AOI22_X1 U23367 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20402) );
  OAI21_X1 U23368 ( .B1(n20403), .B2(n20418), .A(n20402), .ZN(P1_U2926) );
  INV_X1 U23369 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20405) );
  AOI22_X1 U23370 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20404) );
  OAI21_X1 U23371 ( .B1(n20405), .B2(n20418), .A(n20404), .ZN(P1_U2927) );
  AOI22_X1 U23372 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20406) );
  OAI21_X1 U23373 ( .B1(n13373), .B2(n20418), .A(n20406), .ZN(P1_U2928) );
  AOI22_X1 U23374 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20407) );
  OAI21_X1 U23375 ( .B1(n13175), .B2(n20418), .A(n20407), .ZN(P1_U2929) );
  AOI22_X1 U23376 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20408) );
  OAI21_X1 U23377 ( .B1(n13048), .B2(n20418), .A(n20408), .ZN(P1_U2930) );
  AOI22_X1 U23378 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20409) );
  OAI21_X1 U23379 ( .B1(n12890), .B2(n20418), .A(n20409), .ZN(P1_U2931) );
  AOI22_X1 U23380 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20410) );
  OAI21_X1 U23381 ( .B1(n20411), .B2(n20418), .A(n20410), .ZN(P1_U2932) );
  AOI22_X1 U23382 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20412) );
  OAI21_X1 U23383 ( .B1(n12748), .B2(n20418), .A(n20412), .ZN(P1_U2933) );
  AOI22_X1 U23384 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20413), .B1(n20415), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20414) );
  OAI21_X1 U23385 ( .B1(n12602), .B2(n20418), .A(n20414), .ZN(P1_U2934) );
  AOI22_X1 U23386 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20416) );
  OAI21_X1 U23387 ( .B1(n12503), .B2(n20418), .A(n20416), .ZN(P1_U2935) );
  AOI22_X1 U23388 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20858), .B1(n20415), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20417) );
  OAI21_X1 U23389 ( .B1(n12234), .B2(n20418), .A(n20417), .ZN(P1_U2936) );
  AOI22_X1 U23390 ( .A1(n20447), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20442), .ZN(n20420) );
  NAND2_X1 U23391 ( .A1(n20432), .A2(n20419), .ZN(n20434) );
  NAND2_X1 U23392 ( .A1(n20420), .A2(n20434), .ZN(P1_U2945) );
  AOI22_X1 U23393 ( .A1(n20447), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20442), .ZN(n20422) );
  NAND2_X1 U23394 ( .A1(n20432), .A2(n20421), .ZN(n20436) );
  NAND2_X1 U23395 ( .A1(n20422), .A2(n20436), .ZN(P1_U2946) );
  AOI22_X1 U23396 ( .A1(n20447), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20442), .ZN(n20424) );
  NAND2_X1 U23397 ( .A1(n20432), .A2(n20423), .ZN(n20438) );
  NAND2_X1 U23398 ( .A1(n20424), .A2(n20438), .ZN(P1_U2947) );
  AOI22_X1 U23399 ( .A1(n20447), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20442), .ZN(n20426) );
  NAND2_X1 U23400 ( .A1(n20432), .A2(n20425), .ZN(n20440) );
  NAND2_X1 U23401 ( .A1(n20426), .A2(n20440), .ZN(P1_U2948) );
  AOI22_X1 U23402 ( .A1(n20447), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20442), .ZN(n20428) );
  NAND2_X1 U23403 ( .A1(n20432), .A2(n20427), .ZN(n20443) );
  NAND2_X1 U23404 ( .A1(n20428), .A2(n20443), .ZN(P1_U2949) );
  AOI22_X1 U23405 ( .A1(n20447), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20442), .ZN(n20430) );
  NAND2_X1 U23406 ( .A1(n20432), .A2(n20429), .ZN(n20445) );
  NAND2_X1 U23407 ( .A1(n20430), .A2(n20445), .ZN(P1_U2950) );
  AOI22_X1 U23408 ( .A1(n20447), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20442), .ZN(n20433) );
  NAND2_X1 U23409 ( .A1(n20432), .A2(n20431), .ZN(n20448) );
  NAND2_X1 U23410 ( .A1(n20433), .A2(n20448), .ZN(P1_U2951) );
  AOI22_X1 U23411 ( .A1(n20447), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20442), .ZN(n20435) );
  NAND2_X1 U23412 ( .A1(n20435), .A2(n20434), .ZN(P1_U2960) );
  AOI22_X1 U23413 ( .A1(n20447), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20442), .ZN(n20437) );
  NAND2_X1 U23414 ( .A1(n20437), .A2(n20436), .ZN(P1_U2961) );
  AOI22_X1 U23415 ( .A1(n20447), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20442), .ZN(n20439) );
  NAND2_X1 U23416 ( .A1(n20439), .A2(n20438), .ZN(P1_U2962) );
  AOI22_X1 U23417 ( .A1(n20447), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20442), .ZN(n20441) );
  NAND2_X1 U23418 ( .A1(n20441), .A2(n20440), .ZN(P1_U2963) );
  AOI22_X1 U23419 ( .A1(n20447), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20442), .ZN(n20444) );
  NAND2_X1 U23420 ( .A1(n20444), .A2(n20443), .ZN(P1_U2964) );
  AOI22_X1 U23421 ( .A1(n20447), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20442), .ZN(n20446) );
  NAND2_X1 U23422 ( .A1(n20446), .A2(n20445), .ZN(P1_U2965) );
  AOI22_X1 U23423 ( .A1(n20447), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20442), .ZN(n20449) );
  NAND2_X1 U23424 ( .A1(n20449), .A2(n20448), .ZN(P1_U2966) );
  AOI22_X1 U23425 ( .A1(n20450), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n16482), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20459) );
  OAI21_X1 U23426 ( .B1(n20453), .B2(n20452), .A(n20451), .ZN(n20454) );
  INV_X1 U23427 ( .A(n20454), .ZN(n20467) );
  AOI22_X1 U23428 ( .A1(n20467), .A2(n20457), .B1(n20456), .B2(n20455), .ZN(
        n20458) );
  OAI211_X1 U23429 ( .C1(n20461), .C2(n20460), .A(n20459), .B(n20458), .ZN(
        P1_U2995) );
  OAI21_X1 U23430 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20462), .ZN(n20470) );
  INV_X1 U23431 ( .A(n20463), .ZN(n20464) );
  AOI22_X1 U23432 ( .A1(n20464), .A2(n20481), .B1(n16482), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20469) );
  NAND2_X1 U23433 ( .A1(n20483), .A2(n20465), .ZN(n20466) );
  OAI211_X1 U23434 ( .C1(n20497), .C2(n20498), .A(n20466), .B(n20487), .ZN(
        n20474) );
  AOI22_X1 U23435 ( .A1(n20467), .A2(n20509), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20474), .ZN(n20468) );
  OAI211_X1 U23436 ( .C1(n20478), .C2(n20470), .A(n20469), .B(n20468), .ZN(
        P1_U3027) );
  INV_X1 U23437 ( .A(n20471), .ZN(n20473) );
  AOI21_X1 U23438 ( .B1(n20473), .B2(n20481), .A(n20472), .ZN(n20477) );
  AOI22_X1 U23439 ( .A1(n20475), .A2(n20509), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20474), .ZN(n20476) );
  OAI211_X1 U23440 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20478), .A(
        n20477), .B(n20476), .ZN(P1_U3028) );
  INV_X1 U23441 ( .A(n20479), .ZN(n20482) );
  AOI21_X1 U23442 ( .B1(n20482), .B2(n20481), .A(n20480), .ZN(n20496) );
  NAND2_X1 U23443 ( .A1(n20870), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20492) );
  NOR2_X1 U23444 ( .A1(n9985), .A2(n20500), .ZN(n20485) );
  AOI22_X1 U23445 ( .A1(n20485), .A2(n20484), .B1(n20500), .B2(n20483), .ZN(
        n20486) );
  AOI21_X1 U23446 ( .B1(n20487), .B2(n20486), .A(n20870), .ZN(n20488) );
  INV_X1 U23447 ( .A(n20488), .ZN(n20491) );
  NAND3_X1 U23448 ( .A1(n12986), .A2(n20489), .A3(n20509), .ZN(n20490) );
  OAI211_X1 U23449 ( .C1(n20493), .C2(n20492), .A(n20491), .B(n20490), .ZN(
        n20494) );
  INV_X1 U23450 ( .A(n20494), .ZN(n20495) );
  OAI211_X1 U23451 ( .C1(n20498), .C2(n20497), .A(n20496), .B(n20495), .ZN(
        P1_U3029) );
  NAND2_X1 U23452 ( .A1(n20500), .A2(n20499), .ZN(n20513) );
  OAI21_X1 U23453 ( .B1(n20503), .B2(n20502), .A(n20501), .ZN(n20504) );
  INV_X1 U23454 ( .A(n20504), .ZN(n20512) );
  INV_X1 U23455 ( .A(n20505), .ZN(n20510) );
  OAI21_X1 U23456 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20507), .A(
        n20506), .ZN(n20508) );
  AOI22_X1 U23457 ( .A1(n20510), .A2(n20509), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20508), .ZN(n20511) );
  OAI211_X1 U23458 ( .C1(n20514), .C2(n20513), .A(n20512), .B(n20511), .ZN(
        P1_U3030) );
  NOR2_X1 U23459 ( .A1(n20516), .A2(n20515), .ZN(P1_U3032) );
  INV_X1 U23460 ( .A(n20585), .ZN(n20518) );
  NAND2_X1 U23461 ( .A1(n20555), .A2(n20518), .ZN(n20525) );
  INV_X1 U23462 ( .A(n20525), .ZN(n20547) );
  AOI22_X1 U23463 ( .A1(n20548), .A2(n20708), .B1(n20547), .B2(n20701), .ZN(
        n20534) );
  INV_X1 U23464 ( .A(n20582), .ZN(n20519) );
  OAI21_X1 U23465 ( .B1(n20519), .B2(n20548), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20520) );
  NAND2_X1 U23466 ( .A1(n20520), .A2(n20622), .ZN(n20532) );
  NOR2_X1 U23467 ( .A1(n20522), .A2(n20521), .ZN(n20528) );
  OR2_X1 U23468 ( .A1(n20524), .A2(n20523), .ZN(n20588) );
  AOI22_X1 U23469 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20588), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20525), .ZN(n20526) );
  OAI211_X1 U23470 ( .C1(n20532), .C2(n20528), .A(n20527), .B(n20526), .ZN(
        n20550) );
  INV_X1 U23471 ( .A(n20528), .ZN(n20531) );
  INV_X1 U23472 ( .A(n20529), .ZN(n20530) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20550), .B1(
        n20700), .B2(n20549), .ZN(n20533) );
  OAI211_X1 U23474 ( .C1(n20711), .C2(n20582), .A(n20534), .B(n20533), .ZN(
        P1_U3033) );
  AOI22_X1 U23475 ( .A1(n20548), .A2(n20714), .B1(n20547), .B2(n20713), .ZN(
        n20536) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20550), .B1(
        n20712), .B2(n20549), .ZN(n20535) );
  OAI211_X1 U23477 ( .C1(n20717), .C2(n20582), .A(n20536), .B(n20535), .ZN(
        P1_U3034) );
  AOI22_X1 U23478 ( .A1(n20548), .A2(n20720), .B1(n20547), .B2(n20719), .ZN(
        n20538) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20550), .B1(
        n20718), .B2(n20549), .ZN(n20537) );
  OAI211_X1 U23480 ( .C1(n20723), .C2(n20582), .A(n20538), .B(n20537), .ZN(
        P1_U3035) );
  AOI22_X1 U23481 ( .A1(n20548), .A2(n20726), .B1(n20547), .B2(n20725), .ZN(
        n20540) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20550), .B1(
        n20724), .B2(n20549), .ZN(n20539) );
  OAI211_X1 U23483 ( .C1(n20729), .C2(n20582), .A(n20540), .B(n20539), .ZN(
        P1_U3036) );
  AOI22_X1 U23484 ( .A1(n20548), .A2(n20732), .B1(n20547), .B2(n20731), .ZN(
        n20542) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20550), .B1(
        n20730), .B2(n20549), .ZN(n20541) );
  OAI211_X1 U23486 ( .C1(n20735), .C2(n20582), .A(n20542), .B(n20541), .ZN(
        P1_U3037) );
  AOI22_X1 U23487 ( .A1(n20548), .A2(n20738), .B1(n20547), .B2(n20737), .ZN(
        n20544) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20550), .B1(
        n20736), .B2(n20549), .ZN(n20543) );
  OAI211_X1 U23489 ( .C1(n20741), .C2(n20582), .A(n20544), .B(n20543), .ZN(
        P1_U3038) );
  AOI22_X1 U23490 ( .A1(n20548), .A2(n20744), .B1(n20547), .B2(n21074), .ZN(
        n20546) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20550), .B1(
        n20742), .B2(n20549), .ZN(n20545) );
  OAI211_X1 U23492 ( .C1(n20747), .C2(n20582), .A(n20546), .B(n20545), .ZN(
        P1_U3039) );
  AOI22_X1 U23493 ( .A1(n20548), .A2(n20752), .B1(n20547), .B2(n20751), .ZN(
        n20552) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20550), .B1(
        n20749), .B2(n20549), .ZN(n20551) );
  OAI211_X1 U23495 ( .C1(n20758), .C2(n20582), .A(n20552), .B(n20551), .ZN(
        P1_U3040) );
  INV_X1 U23496 ( .A(n20553), .ZN(n20695) );
  NAND2_X1 U23497 ( .A1(n20555), .A2(n20554), .ZN(n20557) );
  NOR2_X1 U23498 ( .A1(n20693), .A2(n20557), .ZN(n20576) );
  AOI21_X1 U23499 ( .B1(n20556), .B2(n20695), .A(n20576), .ZN(n20558) );
  OAI22_X1 U23500 ( .A1(n20558), .A2(n20703), .B1(n20557), .B2(n20697), .ZN(
        n20577) );
  AOI22_X1 U23501 ( .A1(n20577), .A2(n20700), .B1(n20701), .B2(n20576), .ZN(
        n20563) );
  INV_X1 U23502 ( .A(n20557), .ZN(n20561) );
  OAI21_X1 U23503 ( .B1(n20559), .B2(n20702), .A(n20558), .ZN(n20560) );
  OAI221_X1 U23504 ( .B1(n20658), .B2(n20561), .C1(n20703), .C2(n20560), .A(
        n20705), .ZN(n20579) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20623), .ZN(n20562) );
  OAI211_X1 U23506 ( .C1(n20626), .C2(n20582), .A(n20563), .B(n20562), .ZN(
        P1_U3041) );
  AOI22_X1 U23507 ( .A1(n20577), .A2(n20712), .B1(n20713), .B2(n20576), .ZN(
        n20565) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20661), .ZN(n20564) );
  OAI211_X1 U23509 ( .C1(n20664), .C2(n20582), .A(n20565), .B(n20564), .ZN(
        P1_U3042) );
  AOI22_X1 U23510 ( .A1(n20577), .A2(n20718), .B1(n20719), .B2(n20576), .ZN(
        n20567) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20665), .ZN(n20566) );
  OAI211_X1 U23512 ( .C1(n20668), .C2(n20582), .A(n20567), .B(n20566), .ZN(
        P1_U3043) );
  AOI22_X1 U23513 ( .A1(n20577), .A2(n20724), .B1(n20725), .B2(n20576), .ZN(
        n20569) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20669), .ZN(n20568) );
  OAI211_X1 U23515 ( .C1(n20672), .C2(n20582), .A(n20569), .B(n20568), .ZN(
        P1_U3044) );
  AOI22_X1 U23516 ( .A1(n20577), .A2(n20730), .B1(n20731), .B2(n20576), .ZN(
        n20571) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20633), .ZN(n20570) );
  OAI211_X1 U23518 ( .C1(n20636), .C2(n20582), .A(n20571), .B(n20570), .ZN(
        P1_U3045) );
  AOI22_X1 U23519 ( .A1(n20577), .A2(n20736), .B1(n20737), .B2(n20576), .ZN(
        n20573) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20637), .ZN(n20572) );
  OAI211_X1 U23521 ( .C1(n20640), .C2(n20582), .A(n20573), .B(n20572), .ZN(
        P1_U3046) );
  AOI22_X1 U23522 ( .A1(n20577), .A2(n20742), .B1(n21074), .B2(n20576), .ZN(
        n20575) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20679), .ZN(n20574) );
  OAI211_X1 U23524 ( .C1(n20682), .C2(n20582), .A(n20575), .B(n20574), .ZN(
        P1_U3047) );
  AOI22_X1 U23525 ( .A1(n20577), .A2(n20749), .B1(n20751), .B2(n20576), .ZN(
        n20581) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20579), .B1(
        n20578), .B2(n20685), .ZN(n20580) );
  OAI211_X1 U23527 ( .C1(n20691), .C2(n20582), .A(n20581), .B(n20580), .ZN(
        P1_U3048) );
  NOR2_X1 U23528 ( .A1(n20585), .A2(n20615), .ZN(n20610) );
  NAND3_X1 U23529 ( .A1(n20616), .A2(n20622), .A3(n20591), .ZN(n20586) );
  OAI21_X1 U23530 ( .B1(n20588), .B2(n20587), .A(n20586), .ZN(n20609) );
  AOI22_X1 U23531 ( .A1(n20701), .A2(n20610), .B1(n20700), .B2(n20609), .ZN(
        n20596) );
  INV_X1 U23532 ( .A(n20611), .ZN(n20589) );
  AOI21_X1 U23533 ( .B1(n20589), .B2(n20649), .A(n20702), .ZN(n20590) );
  AOI21_X1 U23534 ( .B1(n20616), .B2(n20591), .A(n20590), .ZN(n20592) );
  NOR2_X1 U23535 ( .A1(n20592), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20594) );
  AOI22_X1 U23536 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n20611), .B2(n20708), .ZN(n20595) );
  OAI211_X1 U23537 ( .C1(n20711), .C2(n20649), .A(n20596), .B(n20595), .ZN(
        P1_U3065) );
  AOI22_X1 U23538 ( .A1(n20713), .A2(n20610), .B1(n20712), .B2(n20609), .ZN(
        n20598) );
  AOI22_X1 U23539 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n20611), .B2(n20714), .ZN(n20597) );
  OAI211_X1 U23540 ( .C1(n20717), .C2(n20649), .A(n20598), .B(n20597), .ZN(
        P1_U3066) );
  AOI22_X1 U23541 ( .A1(n20719), .A2(n20610), .B1(n20718), .B2(n20609), .ZN(
        n20600) );
  AOI22_X1 U23542 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n20611), .B2(n20720), .ZN(n20599) );
  OAI211_X1 U23543 ( .C1(n20723), .C2(n20649), .A(n20600), .B(n20599), .ZN(
        P1_U3067) );
  AOI22_X1 U23544 ( .A1(n20725), .A2(n20610), .B1(n20724), .B2(n20609), .ZN(
        n20602) );
  AOI22_X1 U23545 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n20611), .B2(n20726), .ZN(n20601) );
  OAI211_X1 U23546 ( .C1(n20729), .C2(n20649), .A(n20602), .B(n20601), .ZN(
        P1_U3068) );
  AOI22_X1 U23547 ( .A1(n20731), .A2(n20610), .B1(n20730), .B2(n20609), .ZN(
        n20604) );
  AOI22_X1 U23548 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n20611), .B2(n20732), .ZN(n20603) );
  OAI211_X1 U23549 ( .C1(n20735), .C2(n20649), .A(n20604), .B(n20603), .ZN(
        P1_U3069) );
  AOI22_X1 U23550 ( .A1(n20737), .A2(n20610), .B1(n20736), .B2(n20609), .ZN(
        n20606) );
  AOI22_X1 U23551 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n20611), .B2(n20738), .ZN(n20605) );
  OAI211_X1 U23552 ( .C1(n20741), .C2(n20649), .A(n20606), .B(n20605), .ZN(
        P1_U3070) );
  AOI22_X1 U23553 ( .A1(n21074), .A2(n20610), .B1(n20742), .B2(n20609), .ZN(
        n20608) );
  AOI22_X1 U23554 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n20611), .B2(n20744), .ZN(n20607) );
  OAI211_X1 U23555 ( .C1(n20747), .C2(n20649), .A(n20608), .B(n20607), .ZN(
        P1_U3071) );
  AOI22_X1 U23556 ( .A1(n20751), .A2(n20610), .B1(n20749), .B2(n20609), .ZN(
        n20614) );
  AOI22_X1 U23557 ( .A1(n20612), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n20611), .B2(n20752), .ZN(n20613) );
  OAI211_X1 U23558 ( .C1(n20758), .C2(n20649), .A(n20614), .B(n20613), .ZN(
        P1_U3072) );
  NOR2_X1 U23559 ( .A1(n20615), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20621) );
  INV_X1 U23560 ( .A(n20621), .ZN(n20617) );
  NOR2_X1 U23561 ( .A1(n20693), .A2(n20617), .ZN(n20644) );
  AOI21_X1 U23562 ( .B1(n20616), .B2(n20695), .A(n20644), .ZN(n20618) );
  OAI22_X1 U23563 ( .A1(n20618), .A2(n20703), .B1(n20617), .B2(n20697), .ZN(
        n20643) );
  AOI22_X1 U23564 ( .A1(n20701), .A2(n20644), .B1(n20643), .B2(n20700), .ZN(
        n20625) );
  OAI211_X1 U23565 ( .C1(n20619), .C2(n20702), .A(n20622), .B(n20618), .ZN(
        n20620) );
  OAI211_X1 U23566 ( .C1(n20622), .C2(n20621), .A(n20705), .B(n20620), .ZN(
        n20646) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20623), .ZN(n20624) );
  OAI211_X1 U23568 ( .C1(n20626), .C2(n20649), .A(n20625), .B(n20624), .ZN(
        P1_U3073) );
  AOI22_X1 U23569 ( .A1(n20713), .A2(n20644), .B1(n20643), .B2(n20712), .ZN(
        n20628) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20661), .ZN(n20627) );
  OAI211_X1 U23571 ( .C1(n20664), .C2(n20649), .A(n20628), .B(n20627), .ZN(
        P1_U3074) );
  AOI22_X1 U23572 ( .A1(n20719), .A2(n20644), .B1(n20643), .B2(n20718), .ZN(
        n20630) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20665), .ZN(n20629) );
  OAI211_X1 U23574 ( .C1(n20668), .C2(n20649), .A(n20630), .B(n20629), .ZN(
        P1_U3075) );
  AOI22_X1 U23575 ( .A1(n20725), .A2(n20644), .B1(n20643), .B2(n20724), .ZN(
        n20632) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20669), .ZN(n20631) );
  OAI211_X1 U23577 ( .C1(n20672), .C2(n20649), .A(n20632), .B(n20631), .ZN(
        P1_U3076) );
  AOI22_X1 U23578 ( .A1(n20731), .A2(n20644), .B1(n20643), .B2(n20730), .ZN(
        n20635) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20633), .ZN(n20634) );
  OAI211_X1 U23580 ( .C1(n20636), .C2(n20649), .A(n20635), .B(n20634), .ZN(
        P1_U3077) );
  AOI22_X1 U23581 ( .A1(n20737), .A2(n20644), .B1(n20643), .B2(n20736), .ZN(
        n20639) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20637), .ZN(n20638) );
  OAI211_X1 U23583 ( .C1(n20640), .C2(n20649), .A(n20639), .B(n20638), .ZN(
        P1_U3078) );
  AOI22_X1 U23584 ( .A1(n21074), .A2(n20644), .B1(n20643), .B2(n20742), .ZN(
        n20642) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20679), .ZN(n20641) );
  OAI211_X1 U23586 ( .C1(n20682), .C2(n20649), .A(n20642), .B(n20641), .ZN(
        P1_U3079) );
  AOI22_X1 U23587 ( .A1(n20751), .A2(n20644), .B1(n20643), .B2(n20749), .ZN(
        n20648) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20685), .ZN(n20647) );
  OAI211_X1 U23589 ( .C1(n20691), .C2(n20649), .A(n20648), .B(n20647), .ZN(
        P1_U3080) );
  INV_X1 U23590 ( .A(n20650), .ZN(n20652) );
  NOR2_X1 U23591 ( .A1(n20651), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20657) );
  INV_X1 U23592 ( .A(n20657), .ZN(n20653) );
  NOR2_X1 U23593 ( .A1(n20693), .A2(n20653), .ZN(n20683) );
  AOI21_X1 U23594 ( .B1(n20652), .B2(n20695), .A(n20683), .ZN(n20654) );
  OAI22_X1 U23595 ( .A1(n20654), .A2(n20703), .B1(n20653), .B2(n20697), .ZN(
        n20684) );
  AOI22_X1 U23596 ( .A1(n20684), .A2(n20700), .B1(n20701), .B2(n20683), .ZN(
        n20660) );
  OAI21_X1 U23597 ( .B1(n20655), .B2(n20702), .A(n20654), .ZN(n20656) );
  OAI221_X1 U23598 ( .B1(n20658), .B2(n20657), .C1(n20703), .C2(n20656), .A(
        n20705), .ZN(n20687) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20687), .B1(
        n20675), .B2(n20708), .ZN(n20659) );
  OAI211_X1 U23600 ( .C1(n20711), .C2(n20678), .A(n20660), .B(n20659), .ZN(
        P1_U3105) );
  AOI22_X1 U23601 ( .A1(n20684), .A2(n20712), .B1(n20713), .B2(n20683), .ZN(
        n20663) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20661), .ZN(n20662) );
  OAI211_X1 U23603 ( .C1(n20664), .C2(n20690), .A(n20663), .B(n20662), .ZN(
        P1_U3106) );
  AOI22_X1 U23604 ( .A1(n20684), .A2(n20718), .B1(n20719), .B2(n20683), .ZN(
        n20667) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20665), .ZN(n20666) );
  OAI211_X1 U23606 ( .C1(n20668), .C2(n20690), .A(n20667), .B(n20666), .ZN(
        P1_U3107) );
  AOI22_X1 U23607 ( .A1(n20684), .A2(n20724), .B1(n20725), .B2(n20683), .ZN(
        n20671) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20669), .ZN(n20670) );
  OAI211_X1 U23609 ( .C1(n20672), .C2(n20690), .A(n20671), .B(n20670), .ZN(
        P1_U3108) );
  AOI22_X1 U23610 ( .A1(n20684), .A2(n20730), .B1(n20731), .B2(n20683), .ZN(
        n20674) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20687), .B1(
        n20675), .B2(n20732), .ZN(n20673) );
  OAI211_X1 U23612 ( .C1(n20735), .C2(n20678), .A(n20674), .B(n20673), .ZN(
        P1_U3109) );
  AOI22_X1 U23613 ( .A1(n20684), .A2(n20736), .B1(n20737), .B2(n20683), .ZN(
        n20677) );
  AOI22_X1 U23614 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20687), .B1(
        n20675), .B2(n20738), .ZN(n20676) );
  OAI211_X1 U23615 ( .C1(n20741), .C2(n20678), .A(n20677), .B(n20676), .ZN(
        P1_U3110) );
  AOI22_X1 U23616 ( .A1(n20684), .A2(n20742), .B1(n21074), .B2(n20683), .ZN(
        n20681) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20679), .ZN(n20680) );
  OAI211_X1 U23618 ( .C1(n20682), .C2(n20690), .A(n20681), .B(n20680), .ZN(
        P1_U3111) );
  AOI22_X1 U23619 ( .A1(n20684), .A2(n20749), .B1(n20751), .B2(n20683), .ZN(
        n20689) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20685), .ZN(n20688) );
  OAI211_X1 U23621 ( .C1(n20691), .C2(n20690), .A(n20689), .B(n20688), .ZN(
        P1_U3112) );
  NOR2_X1 U23622 ( .A1(n20692), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20706) );
  INV_X1 U23623 ( .A(n20706), .ZN(n20698) );
  NOR2_X1 U23624 ( .A1(n20693), .A2(n20698), .ZN(n20750) );
  INV_X1 U23625 ( .A(n20694), .ZN(n20696) );
  AOI21_X1 U23626 ( .B1(n20696), .B2(n20695), .A(n20750), .ZN(n20699) );
  OAI22_X1 U23627 ( .A1(n20699), .A2(n20703), .B1(n20698), .B2(n20697), .ZN(
        n20748) );
  AOI22_X1 U23628 ( .A1(n20701), .A2(n20750), .B1(n20700), .B2(n20748), .ZN(
        n20710) );
  NOR3_X1 U23629 ( .A1(n20704), .A2(n20703), .A3(n20702), .ZN(n20707) );
  OAI21_X1 U23630 ( .B1(n20707), .B2(n20706), .A(n20705), .ZN(n20754) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20708), .ZN(n20709) );
  OAI211_X1 U23632 ( .C1(n20711), .C2(n20757), .A(n20710), .B(n20709), .ZN(
        P1_U3137) );
  AOI22_X1 U23633 ( .A1(n20713), .A2(n20750), .B1(n20712), .B2(n20748), .ZN(
        n20716) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20714), .ZN(n20715) );
  OAI211_X1 U23635 ( .C1(n20717), .C2(n20757), .A(n20716), .B(n20715), .ZN(
        P1_U3138) );
  AOI22_X1 U23636 ( .A1(n20719), .A2(n20750), .B1(n20718), .B2(n20748), .ZN(
        n20722) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20720), .ZN(n20721) );
  OAI211_X1 U23638 ( .C1(n20723), .C2(n20757), .A(n20722), .B(n20721), .ZN(
        P1_U3139) );
  AOI22_X1 U23639 ( .A1(n20725), .A2(n20750), .B1(n20724), .B2(n20748), .ZN(
        n20728) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20726), .ZN(n20727) );
  OAI211_X1 U23641 ( .C1(n20729), .C2(n20757), .A(n20728), .B(n20727), .ZN(
        P1_U3140) );
  AOI22_X1 U23642 ( .A1(n20731), .A2(n20750), .B1(n20730), .B2(n20748), .ZN(
        n20734) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20732), .ZN(n20733) );
  OAI211_X1 U23644 ( .C1(n20735), .C2(n20757), .A(n20734), .B(n20733), .ZN(
        P1_U3141) );
  AOI22_X1 U23645 ( .A1(n20737), .A2(n20750), .B1(n20736), .B2(n20748), .ZN(
        n20740) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20738), .ZN(n20739) );
  OAI211_X1 U23647 ( .C1(n20741), .C2(n20757), .A(n20740), .B(n20739), .ZN(
        P1_U3142) );
  AOI22_X1 U23648 ( .A1(n21074), .A2(n20750), .B1(n20742), .B2(n20748), .ZN(
        n20746) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20744), .ZN(n20745) );
  OAI211_X1 U23650 ( .C1(n20747), .C2(n20757), .A(n20746), .B(n20745), .ZN(
        P1_U3143) );
  AOI22_X1 U23651 ( .A1(n20751), .A2(n20750), .B1(n20749), .B2(n20748), .ZN(
        n20756) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20754), .B1(
        n20753), .B2(n20752), .ZN(n20755) );
  OAI211_X1 U23653 ( .C1(n20758), .C2(n20757), .A(n20756), .B(n20755), .ZN(
        P1_U3144) );
  INV_X1 U23654 ( .A(n20759), .ZN(n20761) );
  NAND2_X1 U23655 ( .A1(n20761), .A2(n20760), .ZN(P1_U3163) );
  INV_X1 U23656 ( .A(n20845), .ZN(n20841) );
  AND2_X1 U23657 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20841), .ZN(
        P1_U3164) );
  AND2_X1 U23658 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20841), .ZN(
        P1_U3165) );
  AND2_X1 U23659 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20841), .ZN(
        P1_U3166) );
  AND2_X1 U23660 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20841), .ZN(
        P1_U3167) );
  AND2_X1 U23661 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20841), .ZN(
        P1_U3168) );
  AND2_X1 U23662 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20841), .ZN(
        P1_U3169) );
  AND2_X1 U23663 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20841), .ZN(
        P1_U3170) );
  AND2_X1 U23664 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20841), .ZN(
        P1_U3171) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20841), .ZN(
        P1_U3172) );
  AND2_X1 U23666 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20841), .ZN(
        P1_U3173) );
  AND2_X1 U23667 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20841), .ZN(
        P1_U3174) );
  AND2_X1 U23668 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20841), .ZN(
        P1_U3175) );
  AND2_X1 U23669 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20841), .ZN(
        P1_U3176) );
  AND2_X1 U23670 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20841), .ZN(
        P1_U3177) );
  AND2_X1 U23671 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20841), .ZN(
        P1_U3178) );
  AND2_X1 U23672 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20841), .ZN(
        P1_U3179) );
  AND2_X1 U23673 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20841), .ZN(
        P1_U3180) );
  AND2_X1 U23674 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20841), .ZN(
        P1_U3181) );
  AND2_X1 U23675 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20841), .ZN(
        P1_U3182) );
  AND2_X1 U23676 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20841), .ZN(
        P1_U3183) );
  AND2_X1 U23677 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20841), .ZN(
        P1_U3184) );
  AND2_X1 U23678 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20841), .ZN(
        P1_U3185) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20841), .ZN(P1_U3186) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20841), .ZN(P1_U3187) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20841), .ZN(P1_U3188) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20841), .ZN(P1_U3189) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20841), .ZN(P1_U3190) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20841), .ZN(P1_U3191) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20841), .ZN(P1_U3192) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20841), .ZN(P1_U3193) );
  NAND2_X1 U23687 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20762), .ZN(n20774) );
  INV_X1 U23688 ( .A(n20774), .ZN(n20767) );
  NAND2_X1 U23689 ( .A1(n20780), .A2(n20763), .ZN(n20765) );
  NAND2_X1 U23690 ( .A1(n20775), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20768) );
  AOI22_X1 U23691 ( .A1(HOLD), .A2(n20765), .B1(n20768), .B2(n20764), .ZN(
        n20766) );
  OAI22_X1 U23692 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20767), .B1(n20866), 
        .B2(n20766), .ZN(P1_U3194) );
  INV_X1 U23693 ( .A(n20768), .ZN(n20771) );
  AOI21_X1 U23694 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20780), .A(n20769), .ZN(n20770) );
  AOI21_X1 U23695 ( .B1(n20772), .B2(n20771), .A(n20770), .ZN(n20779) );
  NAND3_X1 U23696 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20773), .A3(n20775), 
        .ZN(n20777) );
  OAI211_X1 U23697 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20775), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20774), .ZN(n20776) );
  OAI221_X1 U23698 ( .B1(n20779), .B2(n20778), .C1(n20779), .C2(n20777), .A(
        n20776), .ZN(P1_U3196) );
  NAND2_X1 U23699 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20866), .ZN(n20828) );
  INV_X1 U23700 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20781) );
  NAND2_X1 U23701 ( .A1(n20866), .A2(n20780), .ZN(n20832) );
  OAI222_X1 U23702 ( .A1(n20828), .A2(n20846), .B1(n20782), .B2(n20866), .C1(
        n20781), .C2(n20832), .ZN(P1_U3197) );
  INV_X1 U23703 ( .A(n20828), .ZN(n20830) );
  INV_X1 U23704 ( .A(n20832), .ZN(n20826) );
  AOI222_X1 U23705 ( .A1(n20830), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20812), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20826), .ZN(n20783) );
  INV_X1 U23706 ( .A(n20783), .ZN(P1_U3198) );
  AOI22_X1 U23707 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(n20812), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n20826), .ZN(n20784) );
  OAI21_X1 U23708 ( .B1(n20785), .B2(n20828), .A(n20784), .ZN(P1_U3199) );
  AOI22_X1 U23709 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20812), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n20830), .ZN(n20786) );
  OAI21_X1 U23710 ( .B1(n20788), .B2(n20832), .A(n20786), .ZN(P1_U3200) );
  INV_X1 U23711 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20787) );
  OAI222_X1 U23712 ( .A1(n20828), .A2(n20788), .B1(n20787), .B2(n20866), .C1(
        n16488), .C2(n20832), .ZN(P1_U3201) );
  INV_X1 U23713 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20789) );
  OAI222_X1 U23714 ( .A1(n20828), .A2(n16488), .B1(n20789), .B2(n20866), .C1(
        n20790), .C2(n20832), .ZN(P1_U3202) );
  INV_X1 U23715 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20791) );
  OAI222_X1 U23716 ( .A1(n20832), .A2(n20793), .B1(n20791), .B2(n20866), .C1(
        n20790), .C2(n20828), .ZN(P1_U3203) );
  INV_X1 U23717 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20912) );
  INV_X1 U23718 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20792) );
  OAI222_X1 U23719 ( .A1(n20828), .A2(n20793), .B1(n20912), .B2(n20866), .C1(
        n20792), .C2(n20832), .ZN(P1_U3204) );
  AOI222_X1 U23720 ( .A1(n20826), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20867), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20830), .ZN(n20794) );
  INV_X1 U23721 ( .A(n20794), .ZN(P1_U3205) );
  AOI22_X1 U23722 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20812), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20826), .ZN(n20795) );
  OAI21_X1 U23723 ( .B1(n20796), .B2(n20828), .A(n20795), .ZN(P1_U3206) );
  INV_X1 U23724 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20800) );
  AOI22_X1 U23725 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20812), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20830), .ZN(n20797) );
  OAI21_X1 U23726 ( .B1(n20800), .B2(n20832), .A(n20797), .ZN(P1_U3207) );
  INV_X1 U23727 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20799) );
  OAI222_X1 U23728 ( .A1(n20828), .A2(n20800), .B1(n20799), .B2(n20866), .C1(
        n20798), .C2(n20832), .ZN(P1_U3208) );
  AOI222_X1 U23729 ( .A1(n20830), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20867), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20826), .ZN(n20801) );
  INV_X1 U23730 ( .A(n20801), .ZN(P1_U3209) );
  AOI222_X1 U23731 ( .A1(n20830), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20812), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20826), .ZN(n20802) );
  INV_X1 U23732 ( .A(n20802), .ZN(P1_U3210) );
  INV_X1 U23733 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20806) );
  INV_X1 U23734 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20804) );
  OAI222_X1 U23735 ( .A1(n20832), .A2(n20806), .B1(n20804), .B2(n20866), .C1(
        n20803), .C2(n20828), .ZN(P1_U3211) );
  INV_X1 U23736 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20805) );
  OAI222_X1 U23737 ( .A1(n20828), .A2(n20806), .B1(n20805), .B2(n20866), .C1(
        n20808), .C2(n20832), .ZN(P1_U3212) );
  AOI22_X1 U23738 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20812), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20826), .ZN(n20807) );
  OAI21_X1 U23739 ( .B1(n20808), .B2(n20828), .A(n20807), .ZN(P1_U3213) );
  AOI22_X1 U23740 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20867), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20830), .ZN(n20809) );
  OAI21_X1 U23741 ( .B1(n20811), .B2(n20832), .A(n20809), .ZN(P1_U3214) );
  AOI22_X1 U23742 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20867), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20826), .ZN(n20810) );
  OAI21_X1 U23743 ( .B1(n20811), .B2(n20828), .A(n20810), .ZN(P1_U3215) );
  AOI22_X1 U23744 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20812), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20830), .ZN(n20813) );
  OAI21_X1 U23745 ( .B1(n20814), .B2(n20832), .A(n20813), .ZN(P1_U3216) );
  INV_X1 U23746 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20877) );
  OAI222_X1 U23747 ( .A1(n20828), .A2(n20814), .B1(n20877), .B2(n20866), .C1(
        n14819), .C2(n20832), .ZN(P1_U3217) );
  AOI222_X1 U23748 ( .A1(n20830), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20867), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20826), .ZN(n20815) );
  INV_X1 U23749 ( .A(n20815), .ZN(P1_U3218) );
  AOI22_X1 U23750 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20867), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(n20826), .ZN(n20816) );
  OAI21_X1 U23751 ( .B1(n20817), .B2(n20828), .A(n20816), .ZN(P1_U3219) );
  AOI22_X1 U23752 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n20867), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(n20830), .ZN(n20818) );
  OAI21_X1 U23753 ( .B1(n20820), .B2(n20832), .A(n20818), .ZN(P1_U3220) );
  INV_X1 U23754 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20819) );
  INV_X1 U23755 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20822) );
  OAI222_X1 U23756 ( .A1(n20828), .A2(n20820), .B1(n20819), .B2(n20866), .C1(
        n20822), .C2(n20832), .ZN(P1_U3221) );
  INV_X1 U23757 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20821) );
  OAI222_X1 U23758 ( .A1(n20828), .A2(n20822), .B1(n20821), .B2(n20866), .C1(
        n20824), .C2(n20832), .ZN(P1_U3222) );
  AOI22_X1 U23759 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20826), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20867), .ZN(n20823) );
  OAI21_X1 U23760 ( .B1(n20824), .B2(n20828), .A(n20823), .ZN(P1_U3223) );
  AOI22_X1 U23761 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20830), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20867), .ZN(n20825) );
  OAI21_X1 U23762 ( .B1(n20829), .B2(n20832), .A(n20825), .ZN(P1_U3224) );
  AOI22_X1 U23763 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20826), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20867), .ZN(n20827) );
  OAI21_X1 U23764 ( .B1(n20829), .B2(n20828), .A(n20827), .ZN(P1_U3225) );
  AOI22_X1 U23765 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20830), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20867), .ZN(n20831) );
  OAI21_X1 U23766 ( .B1(n20833), .B2(n20832), .A(n20831), .ZN(P1_U3226) );
  INV_X1 U23767 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U23768 ( .A1(n20866), .A2(n20835), .B1(n20834), .B2(n20867), .ZN(
        P1_U3458) );
  INV_X1 U23769 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20848) );
  INV_X1 U23770 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U23771 ( .A1(n20866), .A2(n20848), .B1(n20836), .B2(n20867), .ZN(
        P1_U3459) );
  INV_X1 U23772 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20837) );
  AOI22_X1 U23773 ( .A1(n20866), .A2(n20838), .B1(n20837), .B2(n20867), .ZN(
        P1_U3460) );
  INV_X1 U23774 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20853) );
  INV_X1 U23775 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20839) );
  AOI22_X1 U23776 ( .A1(n20866), .A2(n20853), .B1(n20839), .B2(n20867), .ZN(
        P1_U3461) );
  INV_X1 U23777 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20842) );
  INV_X1 U23778 ( .A(n20843), .ZN(n20840) );
  AOI21_X1 U23779 ( .B1(n20842), .B2(n20841), .A(n20840), .ZN(P1_U3464) );
  OAI21_X1 U23780 ( .B1(n20845), .B2(n20844), .A(n20843), .ZN(P1_U3465) );
  AOI21_X1 U23781 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20847) );
  AOI22_X1 U23782 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20847), .B2(n20846), .ZN(n20849) );
  AOI22_X1 U23783 ( .A1(n20850), .A2(n20849), .B1(n20848), .B2(n20852), .ZN(
        P1_U3481) );
  NOR2_X1 U23784 ( .A1(n20852), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20851) );
  AOI22_X1 U23785 ( .A1(n20853), .A2(n20852), .B1(n12317), .B2(n20851), .ZN(
        P1_U3482) );
  AOI22_X1 U23786 ( .A1(n20866), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20854), 
        .B2(n20867), .ZN(P1_U3483) );
  AOI211_X1 U23787 ( .C1(n20858), .C2(n20857), .A(n20856), .B(n20855), .ZN(
        n20865) );
  OAI211_X1 U23788 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20860), .A(n20859), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20862) );
  AOI21_X1 U23789 ( .B1(n20862), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20861), 
        .ZN(n20864) );
  NAND2_X1 U23790 ( .A1(n20865), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20863) );
  OAI21_X1 U23791 ( .B1(n20865), .B2(n20864), .A(n20863), .ZN(P1_U3485) );
  OAI22_X1 U23792 ( .A1(n20867), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20866), .ZN(n20868) );
  INV_X1 U23793 ( .A(n20868), .ZN(P1_U3486) );
  AOI22_X1 U23794 ( .A1(n20871), .A2(keyinput120), .B1(n20870), .B2(keyinput79), .ZN(n20869) );
  OAI221_X1 U23795 ( .B1(n20871), .B2(keyinput120), .C1(n20870), .C2(
        keyinput79), .A(n20869), .ZN(n20875) );
  XOR2_X1 U23796 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B(keyinput115), .Z(
        n20874) );
  XNOR2_X1 U23797 ( .A(n20872), .B(keyinput113), .ZN(n20873) );
  OR3_X1 U23798 ( .A1(n20875), .A2(n20874), .A3(n20873), .ZN(n20882) );
  AOI22_X1 U23799 ( .A1(n20877), .A2(keyinput92), .B1(n21031), .B2(keyinput89), 
        .ZN(n20876) );
  OAI221_X1 U23800 ( .B1(n20877), .B2(keyinput92), .C1(n21031), .C2(keyinput89), .A(n20876), .ZN(n20881) );
  AOI22_X1 U23801 ( .A1(n20879), .A2(keyinput127), .B1(keyinput97), .B2(n11416), .ZN(n20878) );
  OAI221_X1 U23802 ( .B1(n20879), .B2(keyinput127), .C1(n11416), .C2(
        keyinput97), .A(n20878), .ZN(n20880) );
  NOR3_X1 U23803 ( .A1(n20882), .A2(n20881), .A3(n20880), .ZN(n20922) );
  AOI22_X1 U23804 ( .A1(n20999), .A2(keyinput93), .B1(keyinput101), .B2(n21027), .ZN(n20883) );
  OAI221_X1 U23805 ( .B1(n20999), .B2(keyinput93), .C1(n21027), .C2(
        keyinput101), .A(n20883), .ZN(n20892) );
  AOI22_X1 U23806 ( .A1(n12092), .A2(keyinput66), .B1(keyinput104), .B2(n20885), .ZN(n20884) );
  OAI221_X1 U23807 ( .B1(n12092), .B2(keyinput66), .C1(n20885), .C2(
        keyinput104), .A(n20884), .ZN(n20891) );
  AOI22_X1 U23808 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput69), 
        .B1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B2(keyinput117), .ZN(n20886) );
  OAI221_X1 U23809 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput69), 
        .C1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .C2(keyinput117), .A(n20886), 
        .ZN(n20890) );
  XOR2_X1 U23810 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(keyinput114), .Z(
        n20888) );
  XNOR2_X1 U23811 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B(keyinput68), .ZN(
        n20887) );
  NAND2_X1 U23812 ( .A1(n20888), .A2(n20887), .ZN(n20889) );
  NOR4_X1 U23813 ( .A1(n20892), .A2(n20891), .A3(n20890), .A4(n20889), .ZN(
        n20921) );
  AOI22_X1 U23814 ( .A1(n21046), .A2(keyinput70), .B1(keyinput122), .B2(n20997), .ZN(n20893) );
  OAI221_X1 U23815 ( .B1(n21046), .B2(keyinput70), .C1(n20997), .C2(
        keyinput122), .A(n20893), .ZN(n20903) );
  AOI22_X1 U23816 ( .A1(n20896), .A2(keyinput82), .B1(keyinput123), .B2(n20895), .ZN(n20894) );
  OAI221_X1 U23817 ( .B1(n20896), .B2(keyinput82), .C1(n20895), .C2(
        keyinput123), .A(n20894), .ZN(n20902) );
  AOI22_X1 U23818 ( .A1(n21041), .A2(keyinput118), .B1(keyinput110), .B2(
        n21040), .ZN(n20897) );
  OAI221_X1 U23819 ( .B1(n21041), .B2(keyinput118), .C1(n21040), .C2(
        keyinput110), .A(n20897), .ZN(n20901) );
  INV_X1 U23820 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n20899) );
  AOI22_X1 U23821 ( .A1(n21015), .A2(keyinput125), .B1(n20899), .B2(keyinput96), .ZN(n20898) );
  OAI221_X1 U23822 ( .B1(n21015), .B2(keyinput125), .C1(n20899), .C2(
        keyinput96), .A(n20898), .ZN(n20900) );
  NOR4_X1 U23823 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n20920) );
  AOI22_X1 U23824 ( .A1(n21001), .A2(keyinput74), .B1(keyinput94), .B2(n20905), 
        .ZN(n20904) );
  OAI221_X1 U23825 ( .B1(n21001), .B2(keyinput74), .C1(n20905), .C2(keyinput94), .A(n20904), .ZN(n20909) );
  XOR2_X1 U23826 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B(keyinput90), .Z(
        n20908) );
  XNOR2_X1 U23827 ( .A(n20906), .B(keyinput98), .ZN(n20907) );
  OR3_X1 U23828 ( .A1(n20909), .A2(n20908), .A3(n20907), .ZN(n20918) );
  AOI22_X1 U23829 ( .A1(n20912), .A2(keyinput76), .B1(keyinput116), .B2(n20911), .ZN(n20910) );
  OAI221_X1 U23830 ( .B1(n20912), .B2(keyinput76), .C1(n20911), .C2(
        keyinput116), .A(n20910), .ZN(n20917) );
  INV_X1 U23831 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20915) );
  AOI22_X1 U23832 ( .A1(n20915), .A2(keyinput112), .B1(keyinput91), .B2(n20914), .ZN(n20913) );
  OAI221_X1 U23833 ( .B1(n20915), .B2(keyinput112), .C1(n20914), .C2(
        keyinput91), .A(n20913), .ZN(n20916) );
  NOR3_X1 U23834 ( .A1(n20918), .A2(n20917), .A3(n20916), .ZN(n20919) );
  NAND4_X1 U23835 ( .A1(n20922), .A2(n20921), .A3(n20920), .A4(n20919), .ZN(
        n21061) );
  AOI22_X1 U23836 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput67), 
        .B1(P3_REIP_REG_29__SCAN_IN), .B2(keyinput106), .ZN(n20923) );
  OAI221_X1 U23837 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput67), 
        .C1(P3_REIP_REG_29__SCAN_IN), .C2(keyinput106), .A(n20923), .ZN(n20930) );
  AOI22_X1 U23838 ( .A1(BUF1_REG_7__SCAN_IN), .A2(keyinput84), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput83), .ZN(n20924) );
  OAI221_X1 U23839 ( .B1(BUF1_REG_7__SCAN_IN), .B2(keyinput84), .C1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(keyinput83), .A(n20924), .ZN(
        n20929) );
  AOI22_X1 U23840 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput87), .B1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .B2(keyinput80), .ZN(n20925) );
  OAI221_X1 U23841 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput87), .C1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .C2(keyinput80), .A(n20925), .ZN(
        n20928) );
  AOI22_X1 U23842 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput81), 
        .B1(P2_REIP_REG_1__SCAN_IN), .B2(keyinput77), .ZN(n20926) );
  OAI221_X1 U23843 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput81), 
        .C1(P2_REIP_REG_1__SCAN_IN), .C2(keyinput77), .A(n20926), .ZN(n20927)
         );
  NOR4_X1 U23844 ( .A1(n20930), .A2(n20929), .A3(n20928), .A4(n20927), .ZN(
        n20958) );
  AOI22_X1 U23845 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput72), .B1(
        P1_INSTQUEUE_REG_13__7__SCAN_IN), .B2(keyinput108), .ZN(n20931) );
  OAI221_X1 U23846 ( .B1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput72), 
        .C1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .C2(keyinput108), .A(n20931), 
        .ZN(n20938) );
  AOI22_X1 U23847 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput100), .B1(
        P1_INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput88), .ZN(n20932) );
  OAI221_X1 U23848 ( .B1(P2_DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput100), .C1(
        P1_INSTQUEUE_REG_2__1__SCAN_IN), .C2(keyinput88), .A(n20932), .ZN(
        n20937) );
  AOI22_X1 U23849 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(keyinput124), 
        .B1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B2(keyinput64), .ZN(n20933) );
  OAI221_X1 U23850 ( .B1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput124), 
        .C1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .C2(keyinput64), .A(n20933), .ZN(
        n20936) );
  AOI22_X1 U23851 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(keyinput99), 
        .B1(P3_EBX_REG_27__SCAN_IN), .B2(keyinput119), .ZN(n20934) );
  OAI221_X1 U23852 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput99), 
        .C1(P3_EBX_REG_27__SCAN_IN), .C2(keyinput119), .A(n20934), .ZN(n20935)
         );
  NOR4_X1 U23853 ( .A1(n20938), .A2(n20937), .A3(n20936), .A4(n20935), .ZN(
        n20957) );
  AOI22_X1 U23854 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput121), .B1(
        P2_INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput126), .ZN(n20939) );
  OAI221_X1 U23855 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput121), .C1(
        P2_INSTQUEUE_REG_8__5__SCAN_IN), .C2(keyinput126), .A(n20939), .ZN(
        n20946) );
  AOI22_X1 U23856 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(keyinput95), .B1(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput73), .ZN(n20940) );
  OAI221_X1 U23857 ( .B1(P1_ADDRESS_REG_12__SCAN_IN), .B2(keyinput95), .C1(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput73), .A(n20940), .ZN(
        n20945) );
  AOI22_X1 U23858 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput75), 
        .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput71), .ZN(n20941) );
  OAI221_X1 U23859 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput75), 
        .C1(P1_EBX_REG_1__SCAN_IN), .C2(keyinput71), .A(n20941), .ZN(n20944)
         );
  AOI22_X1 U23860 ( .A1(BUF1_REG_8__SCAN_IN), .A2(keyinput65), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput78), .ZN(n20942) );
  OAI221_X1 U23861 ( .B1(BUF1_REG_8__SCAN_IN), .B2(keyinput65), .C1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .C2(keyinput78), .A(n20942), .ZN(
        n20943) );
  NOR4_X1 U23862 ( .A1(n20946), .A2(n20945), .A3(n20944), .A4(n20943), .ZN(
        n20956) );
  AOI22_X1 U23863 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(keyinput85), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(keyinput86), .ZN(n20947) );
  OAI221_X1 U23864 ( .B1(P2_LWORD_REG_8__SCAN_IN), .B2(keyinput85), .C1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(keyinput86), .A(n20947), .ZN(
        n20954) );
  AOI22_X1 U23865 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(keyinput103), 
        .B1(P1_ADDRESS_REG_15__SCAN_IN), .B2(keyinput107), .ZN(n20948) );
  OAI221_X1 U23866 ( .B1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput103), 
        .C1(P1_ADDRESS_REG_15__SCAN_IN), .C2(keyinput107), .A(n20948), .ZN(
        n20953) );
  AOI22_X1 U23867 ( .A1(DATAI_16_), .A2(keyinput102), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(keyinput111), .ZN(n20949) );
  OAI221_X1 U23868 ( .B1(DATAI_16_), .B2(keyinput102), .C1(
        P2_EAX_REG_28__SCAN_IN), .C2(keyinput111), .A(n20949), .ZN(n20952) );
  AOI22_X1 U23869 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(keyinput109), .B1(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput105), .ZN(n20950) );
  OAI221_X1 U23870 ( .B1(P2_LWORD_REG_0__SCAN_IN), .B2(keyinput109), .C1(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .C2(keyinput105), .A(n20950), .ZN(
        n20951) );
  NOR4_X1 U23871 ( .A1(n20954), .A2(n20953), .A3(n20952), .A4(n20951), .ZN(
        n20955) );
  NAND4_X1 U23872 ( .A1(n20958), .A2(n20957), .A3(n20956), .A4(n20955), .ZN(
        n21060) );
  OAI22_X1 U23873 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(keyinput18), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(keyinput56), .ZN(n20959) );
  AOI221_X1 U23874 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(keyinput18), .C1(
        keyinput56), .C2(P3_EAX_REG_21__SCAN_IN), .A(n20959), .ZN(n20966) );
  OAI22_X1 U23875 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput33), 
        .B1(P1_ADDRESS_REG_12__SCAN_IN), .B2(keyinput31), .ZN(n20960) );
  AOI221_X1 U23876 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput33), 
        .C1(keyinput31), .C2(P1_ADDRESS_REG_12__SCAN_IN), .A(n20960), .ZN(
        n20965) );
  OAI22_X1 U23877 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(keyinput22), .B1(
        keyinput17), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20961) );
  AOI221_X1 U23878 ( .B1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(keyinput22), 
        .C1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(keyinput17), .A(n20961), 
        .ZN(n20964) );
  OAI22_X1 U23879 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(keyinput60), 
        .B1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput59), .ZN(n20962) );
  AOI221_X1 U23880 ( .B1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput60), 
        .C1(keyinput59), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(n20962), .ZN(
        n20963) );
  NAND4_X1 U23881 ( .A1(n20966), .A2(n20965), .A3(n20964), .A4(n20963), .ZN(
        n20994) );
  OAI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(keyinput48), .B1(
        keyinput27), .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n20967) );
  AOI221_X1 U23883 ( .B1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(keyinput48), 
        .C1(P3_DATAO_REG_8__SCAN_IN), .C2(keyinput27), .A(n20967), .ZN(n20974)
         );
  OAI22_X1 U23884 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(keyinput35), 
        .B1(keyinput49), .B2(P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20968) );
  AOI221_X1 U23885 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput35), 
        .C1(P2_DATAWIDTH_REG_27__SCAN_IN), .C2(keyinput49), .A(n20968), .ZN(
        n20973) );
  OAI22_X1 U23886 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(keyinput42), .B1(
        keyinput52), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n20969) );
  AOI221_X1 U23887 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(keyinput42), .C1(
        P3_EBX_REG_7__SCAN_IN), .C2(keyinput52), .A(n20969), .ZN(n20972) );
  OAI22_X1 U23888 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(keyinput19), .B1(
        keyinput45), .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n20970) );
  AOI221_X1 U23889 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput19), 
        .C1(P2_LWORD_REG_0__SCAN_IN), .C2(keyinput45), .A(n20970), .ZN(n20971)
         );
  NAND4_X1 U23890 ( .A1(n20974), .A2(n20973), .A3(n20972), .A4(n20971), .ZN(
        n20993) );
  OAI22_X1 U23891 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput15), 
        .B1(keyinput12), .B2(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20975) );
  AOI221_X1 U23892 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput15), 
        .C1(P1_ADDRESS_REG_7__SCAN_IN), .C2(keyinput12), .A(n20975), .ZN(
        n20982) );
  OAI22_X1 U23893 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(keyinput43), .B1(
        keyinput30), .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n20976) );
  AOI221_X1 U23894 ( .B1(P1_ADDRESS_REG_15__SCAN_IN), .B2(keyinput43), .C1(
        P3_DATAO_REG_26__SCAN_IN), .C2(keyinput30), .A(n20976), .ZN(n20981) );
  OAI22_X1 U23895 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(keyinput62), .B1(
        keyinput39), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n20977) );
  AOI221_X1 U23896 ( .B1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput62), 
        .C1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .C2(keyinput39), .A(n20977), .ZN(
        n20980) );
  OAI22_X1 U23897 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(keyinput4), .B1(
        keyinput34), .B2(P3_LWORD_REG_3__SCAN_IN), .ZN(n20978) );
  AOI221_X1 U23898 ( .B1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput4), .C1(
        P3_LWORD_REG_3__SCAN_IN), .C2(keyinput34), .A(n20978), .ZN(n20979) );
  NAND4_X1 U23899 ( .A1(n20982), .A2(n20981), .A3(n20980), .A4(n20979), .ZN(
        n20992) );
  OAI22_X1 U23900 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(keyinput55), .B1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput3), .ZN(n20983) );
  AOI221_X1 U23901 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(keyinput55), .C1(
        keyinput3), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(n20983), .ZN(
        n20990) );
  OAI22_X1 U23902 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(keyinput63), .B1(
        keyinput40), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20984) );
  AOI221_X1 U23903 ( .B1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(keyinput63), 
        .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(keyinput40), .A(n20984), 
        .ZN(n20989) );
  OAI22_X1 U23904 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(keyinput32), 
        .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput7), .ZN(n20985) );
  AOI221_X1 U23905 ( .B1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput32), 
        .C1(keyinput7), .C2(P1_EBX_REG_1__SCAN_IN), .A(n20985), .ZN(n20988) );
  OAI22_X1 U23906 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(keyinput28), .B1(
        keyinput38), .B2(DATAI_16_), .ZN(n20986) );
  AOI221_X1 U23907 ( .B1(P1_ADDRESS_REG_20__SCAN_IN), .B2(keyinput28), .C1(
        DATAI_16_), .C2(keyinput38), .A(n20986), .ZN(n20987) );
  NAND4_X1 U23908 ( .A1(n20990), .A2(n20989), .A3(n20988), .A4(n20987), .ZN(
        n20991) );
  NOR4_X1 U23909 ( .A1(n20994), .A2(n20993), .A3(n20992), .A4(n20991), .ZN(
        n21059) );
  AOI22_X1 U23910 ( .A1(n20997), .A2(keyinput58), .B1(n20996), .B2(keyinput13), 
        .ZN(n20995) );
  OAI221_X1 U23911 ( .B1(n20997), .B2(keyinput58), .C1(n20996), .C2(keyinput13), .A(n20995), .ZN(n21008) );
  AOI22_X1 U23912 ( .A1(n20999), .A2(keyinput29), .B1(n10046), .B2(keyinput9), 
        .ZN(n20998) );
  OAI221_X1 U23913 ( .B1(n20999), .B2(keyinput29), .C1(n10046), .C2(keyinput9), 
        .A(n20998), .ZN(n21007) );
  INV_X1 U23914 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n21002) );
  AOI22_X1 U23915 ( .A1(n21002), .A2(keyinput24), .B1(keyinput10), .B2(n21001), 
        .ZN(n21000) );
  OAI221_X1 U23916 ( .B1(n21002), .B2(keyinput24), .C1(n21001), .C2(keyinput10), .A(n21000), .ZN(n21006) );
  AOI22_X1 U23917 ( .A1(n12427), .A2(keyinput1), .B1(keyinput11), .B2(n21004), 
        .ZN(n21003) );
  OAI221_X1 U23918 ( .B1(n12427), .B2(keyinput1), .C1(n21004), .C2(keyinput11), 
        .A(n21003), .ZN(n21005) );
  NOR4_X1 U23919 ( .A1(n21008), .A2(n21007), .A3(n21006), .A4(n21005), .ZN(
        n21057) );
  AOI22_X1 U23920 ( .A1(n21011), .A2(keyinput23), .B1(keyinput50), .B2(n21010), 
        .ZN(n21009) );
  OAI221_X1 U23921 ( .B1(n21011), .B2(keyinput23), .C1(n21010), .C2(keyinput50), .A(n21009), .ZN(n21023) );
  INV_X1 U23922 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21013) );
  AOI22_X1 U23923 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(keyinput14), .B1(
        n21013), .B2(keyinput0), .ZN(n21012) );
  OAI221_X1 U23924 ( .B1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput14), 
        .C1(n21013), .C2(keyinput0), .A(n21012), .ZN(n21022) );
  AOI22_X1 U23925 ( .A1(n21016), .A2(keyinput57), .B1(keyinput61), .B2(n21015), 
        .ZN(n21014) );
  OAI221_X1 U23926 ( .B1(n21016), .B2(keyinput57), .C1(n21015), .C2(keyinput61), .A(n21014), .ZN(n21021) );
  INV_X1 U23927 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21019) );
  AOI22_X1 U23928 ( .A1(n21019), .A2(keyinput41), .B1(keyinput20), .B2(n21018), 
        .ZN(n21017) );
  OAI221_X1 U23929 ( .B1(n21019), .B2(keyinput41), .C1(n21018), .C2(keyinput20), .A(n21017), .ZN(n21020) );
  NOR4_X1 U23930 ( .A1(n21023), .A2(n21022), .A3(n21021), .A4(n21020), .ZN(
        n21056) );
  AOI22_X1 U23931 ( .A1(n12092), .A2(keyinput2), .B1(keyinput36), .B2(n21025), 
        .ZN(n21024) );
  OAI221_X1 U23932 ( .B1(n12092), .B2(keyinput2), .C1(n21025), .C2(keyinput36), 
        .A(n21024), .ZN(n21037) );
  INV_X1 U23933 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n21028) );
  AOI22_X1 U23934 ( .A1(n21028), .A2(keyinput53), .B1(keyinput37), .B2(n21027), 
        .ZN(n21026) );
  OAI221_X1 U23935 ( .B1(n21028), .B2(keyinput53), .C1(n21027), .C2(keyinput37), .A(n21026), .ZN(n21036) );
  AOI22_X1 U23936 ( .A1(n21031), .A2(keyinput25), .B1(keyinput21), .B2(n21030), 
        .ZN(n21029) );
  OAI221_X1 U23937 ( .B1(n21031), .B2(keyinput25), .C1(n21030), .C2(keyinput21), .A(n21029), .ZN(n21035) );
  XNOR2_X1 U23938 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B(keyinput26), .ZN(
        n21033) );
  XNOR2_X1 U23939 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B(keyinput16), .ZN(
        n21032) );
  NAND2_X1 U23940 ( .A1(n21033), .A2(n21032), .ZN(n21034) );
  NOR4_X1 U23941 ( .A1(n21037), .A2(n21036), .A3(n21035), .A4(n21034), .ZN(
        n21055) );
  AOI22_X1 U23942 ( .A1(n21040), .A2(keyinput46), .B1(n21039), .B2(keyinput47), 
        .ZN(n21038) );
  OAI221_X1 U23943 ( .B1(n21040), .B2(keyinput46), .C1(n21039), .C2(keyinput47), .A(n21038), .ZN(n21044) );
  XNOR2_X1 U23944 ( .A(n21041), .B(keyinput54), .ZN(n21043) );
  XOR2_X1 U23945 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B(keyinput51), .Z(
        n21042) );
  OR3_X1 U23946 ( .A1(n21044), .A2(n21043), .A3(n21042), .ZN(n21053) );
  AOI22_X1 U23947 ( .A1(n21047), .A2(keyinput5), .B1(keyinput6), .B2(n21046), 
        .ZN(n21045) );
  OAI221_X1 U23948 ( .B1(n21047), .B2(keyinput5), .C1(n21046), .C2(keyinput6), 
        .A(n21045), .ZN(n21052) );
  INV_X1 U23949 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21050) );
  INV_X1 U23950 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n21049) );
  AOI22_X1 U23951 ( .A1(n21050), .A2(keyinput8), .B1(n21049), .B2(keyinput44), 
        .ZN(n21048) );
  OAI221_X1 U23952 ( .B1(n21050), .B2(keyinput8), .C1(n21049), .C2(keyinput44), 
        .A(n21048), .ZN(n21051) );
  NOR3_X1 U23953 ( .A1(n21053), .A2(n21052), .A3(n21051), .ZN(n21054) );
  AND4_X1 U23954 ( .A1(n21057), .A2(n21056), .A3(n21055), .A4(n21054), .ZN(
        n21058) );
  OAI211_X1 U23955 ( .C1(n21061), .C2(n21060), .A(n21059), .B(n21058), .ZN(
        n21073) );
  NAND2_X1 U23956 ( .A1(n21062), .A2(DATAI_22_), .ZN(n21067) );
  AOI22_X1 U23957 ( .A1(n21065), .A2(n21064), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n21063), .ZN(n21066) );
  OAI211_X1 U23958 ( .C1(n16859), .C2(n21068), .A(n21067), .B(n21066), .ZN(
        n21069) );
  INV_X1 U23959 ( .A(n21069), .ZN(n21070) );
  OAI21_X1 U23960 ( .B1(n21071), .B2(n14717), .A(n21070), .ZN(n21072) );
  XNOR2_X1 U23961 ( .A(n21073), .B(n21072), .ZN(P1_U2882) );
  AND2_X1 U14887 ( .A1(n11878), .A2(n11882), .ZN(n11983) );
  BUF_X1 U11251 ( .A(n11674), .Z(n11778) );
  BUF_X1 U11101 ( .A(n10446), .Z(n10458) );
  INV_X1 U11108 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20268) );
  INV_X1 U12718 ( .A(n15894), .ZN(n9795) );
  CLKBUF_X2 U11131 ( .A(n13337), .Z(n9682) );
  NOR2_X1 U11135 ( .A1(n12911), .A2(n12905), .ZN(n21074) );
  CLKBUF_X1 U11136 ( .A(n11979), .Z(n12905) );
  CLKBUF_X3 U11137 ( .A(n13337), .Z(n9681) );
  INV_X1 U11138 ( .A(n9660), .ZN(n19068) );
  NAND2_X1 U11401 ( .A1(n16062), .A2(n18222), .ZN(n16064) );
  CLKBUF_X1 U11428 ( .A(n13184), .Z(n14456) );
  OR2_X1 U11430 ( .A1(n18481), .A2(n19264), .ZN(n21075) );
  OR2_X1 U11477 ( .A1(n17239), .A2(n19094), .ZN(n21076) );
  CLKBUF_X1 U12188 ( .A(n17883), .Z(n17891) );
endmodule

