

module b14_C_AntiSAT_k_256_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075;

  OAI21_X1 U2470 ( .B1(n2307), .B2(n2306), .A(n2304), .ZN(n3760) );
  INV_X2 U2471 ( .A(n2600), .ZN(n2972) );
  CLKBUF_X1 U2472 ( .A(n3150), .Z(n2232) );
  INV_X1 U2474 ( .A(n2600), .ZN(n2971) );
  INV_X1 U2475 ( .A(n2973), .ZN(n2984) );
  AND2_X1 U2476 ( .A1(n3905), .A2(n3902), .ZN(n3878) );
  NAND2_X1 U2477 ( .A1(n3269), .A2(n3005), .ZN(n2973) );
  NAND2_X1 U2478 ( .A1(n2558), .A2(IR_REG_31__SCAN_IN), .ZN(n2317) );
  NOR2_X1 U2479 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2449)
         );
  NAND4_X1 U2480 ( .A1(n2641), .A2(n2640), .A3(n2639), .A4(n2638), .ZN(n3449)
         );
  AND2_X1 U2481 ( .A1(n3106), .A2(n3105), .ZN(n2228) );
  INV_X1 U2482 ( .A(n3387), .ZN(n3394) );
  OAI21_X2 U2484 ( .B1(n4457), .B2(n2280), .A(n3181), .ZN(n4469) );
  INV_X1 U2485 ( .A(n2599), .ZN(n2229) );
  INV_X1 U2486 ( .A(n2229), .ZN(n2230) );
  INV_X1 U2487 ( .A(n2229), .ZN(n2231) );
  XNOR2_X1 U2488 ( .A(n2446), .B(IR_REG_1__SCAN_IN), .ZN(n3150) );
  AND2_X4 U2489 ( .A1(n4385), .A2(n2578), .ZN(n2603) );
  XNOR2_X2 U2490 ( .A(n2451), .B(IR_REG_2__SCAN_IN), .ZN(n3146) );
  BUF_X4 U2491 ( .A(n2650), .Z(n2977) );
  INV_X1 U2492 ( .A(n2742), .ZN(n2233) );
  INV_X1 U2493 ( .A(n2233), .ZN(n2234) );
  INV_X2 U2494 ( .A(n2233), .ZN(n2235) );
  XNOR2_X2 U2495 ( .A(n2317), .B(n2559), .ZN(n2595) );
  AOI21_X1 U2496 ( .B1(n3769), .B2(n3770), .A(n3772), .ZN(n3805) );
  AOI21_X1 U2497 ( .B1(n3228), .B2(n3229), .A(n2648), .ZN(n3239) );
  INV_X2 U2498 ( .A(n2629), .ZN(n2658) );
  INV_X2 U2499 ( .A(n3251), .ZN(n2598) );
  OAI21_X1 U2500 ( .B1(n3144), .B2(n3163), .A(n2453), .ZN(n3387) );
  BUF_X2 U2501 ( .A(n2521), .Z(n3144) );
  AND2_X1 U2502 ( .A1(n2567), .A2(n3869), .ZN(n4629) );
  MUX2_X1 U2503 ( .A(REG0_REG_28__SCAN_IN), .B(n3123), .S(n4673), .Z(n3124) );
  AOI21_X1 U2504 ( .B1(n4073), .B2(n4197), .A(n4072), .ZN(n4293) );
  NAND2_X1 U2505 ( .A1(n2326), .A2(n2323), .ZN(n3769) );
  AND2_X1 U2506 ( .A1(n4219), .A2(n4169), .ZN(n4190) );
  AND2_X1 U2507 ( .A1(n3797), .A2(n2938), .ZN(n3739) );
  NAND2_X1 U2508 ( .A1(n3798), .A2(n3799), .ZN(n3797) );
  AND2_X1 U2509 ( .A1(n3668), .A2(n3079), .ZN(n3684) );
  AND2_X1 U2510 ( .A1(n4044), .A2(n4543), .ZN(n4045) );
  NAND2_X1 U2511 ( .A1(n3075), .A2(n2293), .ZN(n3606) );
  OAI21_X1 U2512 ( .B1(n3437), .B2(n2784), .A(n2783), .ZN(n3534) );
  AOI21_X1 U2513 ( .B1(n4534), .B2(n4043), .A(n4042), .ZN(n4044) );
  OAI21_X1 U2514 ( .B1(n3494), .B2(n3581), .A(n3580), .ZN(n4039) );
  NAND2_X1 U2515 ( .A1(n2298), .A2(n3913), .ZN(n3273) );
  NAND2_X1 U2516 ( .A1(n4508), .A2(n3491), .ZN(n3492) );
  NAND2_X1 U2517 ( .A1(n3486), .A2(n3487), .ZN(n3488) );
  NAND2_X2 U2518 ( .A1(n2566), .A2(n4268), .ZN(n4273) );
  OAI21_X1 U2519 ( .B1(n3420), .B2(n3183), .A(n4470), .ZN(n3184) );
  INV_X2 U2520 ( .A(n4004), .ZN(U4043) );
  INV_X1 U2521 ( .A(n2578), .ZN(n3131) );
  OAI21_X1 U2522 ( .B1(n2521), .B2(n2448), .A(n2447), .ZN(n2599) );
  AND2_X2 U2523 ( .A1(n2579), .A2(n2578), .ZN(n2651) );
  NAND2_X1 U2524 ( .A1(n2595), .A2(n4390), .ZN(n3269) );
  NAND2_X2 U2525 ( .A1(n2445), .A2(n2444), .ZN(n2521) );
  INV_X1 U2526 ( .A(n3869), .ZN(n4390) );
  OR2_X1 U2527 ( .A1(n2527), .A2(n2553), .ZN(n2528) );
  AND2_X1 U2528 ( .A1(n2318), .A2(n2268), .ZN(n2558) );
  AND2_X1 U2529 ( .A1(n2454), .A2(n2430), .ZN(n2431) );
  AND2_X1 U2530 ( .A1(n2418), .A2(n2429), .ZN(n2346) );
  INV_X1 U2531 ( .A(IR_REG_17__SCAN_IN), .ZN(n2504) );
  INV_X1 U2532 ( .A(IR_REG_2__SCAN_IN), .ZN(n2429) );
  NOR2_X2 U2533 ( .A1(n4345), .A2(n3717), .ZN(n3705) );
  AND2_X4 U2534 ( .A1(n2596), .A2(n2597), .ZN(n2600) );
  OAI21_X1 U2535 ( .B1(n2583), .B2(n2585), .A(n2442), .ZN(n2445) );
  NAND2_X1 U2536 ( .A1(n2597), .A2(n3137), .ZN(n3140) );
  INV_X1 U2537 ( .A(IR_REG_19__SCAN_IN), .ZN(n2518) );
  XNOR2_X1 U2538 ( .A(n2299), .B(n2973), .ZN(n2621) );
  OAI22_X1 U2539 ( .A1(n3451), .A2(n2971), .B1(n3026), .B2(n2627), .ZN(n2299)
         );
  NAND2_X1 U2540 ( .A1(n2602), .A2(n2601), .ZN(n2620) );
  OR2_X1 U2541 ( .A1(n3451), .A2(n2629), .ZN(n2602) );
  AOI21_X1 U2542 ( .B1(n2413), .B2(n2415), .A(n2240), .ZN(n2411) );
  INV_X1 U2543 ( .A(n2413), .ZN(n2412) );
  INV_X1 U2544 ( .A(n3854), .ZN(n2416) );
  INV_X1 U2545 ( .A(n2406), .ZN(n2402) );
  NOR2_X1 U2546 ( .A1(n2256), .A2(n3055), .ZN(n2404) );
  OAI21_X1 U2547 ( .B1(n2378), .B2(n2375), .A(n2263), .ZN(n2374) );
  INV_X1 U2548 ( .A(n3053), .ZN(n2375) );
  INV_X1 U2549 ( .A(n3944), .ZN(n3825) );
  NAND2_X1 U2550 ( .A1(n3451), .A2(n2231), .ZN(n3901) );
  INV_X1 U2551 ( .A(IR_REG_5__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U2552 ( .A1(n4562), .A2(n4032), .ZN(n4574) );
  AOI21_X1 U2553 ( .B1(n4150), .B2(n3060), .A(n2253), .ZN(n4132) );
  OAI21_X1 U2554 ( .B1(n3273), .B2(n3069), .A(n3921), .ZN(n3375) );
  AND3_X1 U2555 ( .A1(n3115), .A2(n3114), .A3(n3113), .ZN(n3121) );
  NOR2_X1 U2556 ( .A1(n2438), .A2(n2437), .ZN(n2439) );
  NOR2_X1 U2557 ( .A1(n2570), .A2(IR_REG_28__SCAN_IN), .ZN(n2421) );
  INV_X1 U2558 ( .A(IR_REG_22__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U2559 ( .A1(n4574), .A2(n4575), .ZN(n4573) );
  INV_X1 U2560 ( .A(n4548), .ZN(n2363) );
  INV_X1 U2561 ( .A(n3532), .ZN(n2335) );
  AND2_X1 U2562 ( .A1(n2894), .A2(n2893), .ZN(n2896) );
  OAI21_X1 U2563 ( .B1(n3173), .B2(n2371), .A(n3191), .ZN(n2370) );
  NAND2_X1 U2564 ( .A1(n3576), .A2(n3575), .ZN(n3577) );
  NOR2_X1 U2565 ( .A1(n4530), .A2(REG2_REG_13__SCAN_IN), .ZN(n4042) );
  INV_X1 U2566 ( .A(n3951), .ZN(n2286) );
  AND2_X1 U2567 ( .A1(n3832), .A2(n2285), .ZN(n2284) );
  OR2_X1 U2568 ( .A1(n2286), .A2(n3946), .ZN(n2285) );
  NAND2_X1 U2569 ( .A1(n4222), .A2(n4239), .ZN(n2406) );
  NAND2_X1 U2570 ( .A1(n3684), .A2(n3081), .ZN(n4229) );
  NAND2_X1 U2571 ( .A1(n3606), .A2(n3936), .ZN(n2295) );
  NAND2_X1 U2572 ( .A1(n3988), .A2(n3285), .ZN(n3921) );
  NAND2_X1 U2573 ( .A1(n3447), .A2(n3878), .ZN(n2292) );
  NAND2_X1 U2574 ( .A1(n3025), .A2(n3026), .ZN(n3898) );
  AND2_X1 U2575 ( .A1(n4389), .A2(n4390), .ZN(n3141) );
  NOR2_X1 U2576 ( .A1(n3860), .A2(n2342), .ZN(n2341) );
  NAND2_X1 U2577 ( .A1(n2568), .A2(n2296), .ZN(n2570) );
  AND2_X1 U2578 ( .A1(n2443), .A2(n2569), .ZN(n2296) );
  NOR2_X1 U2579 ( .A1(n2676), .A2(n2322), .ZN(n2320) );
  OR2_X1 U2580 ( .A1(n3531), .A2(n2335), .ZN(n2333) );
  AND2_X1 U2581 ( .A1(n3531), .A2(n2335), .ZN(n2334) );
  OR2_X1 U2582 ( .A1(n2734), .A2(n2733), .ZN(n2735) );
  INV_X1 U2583 ( .A(n2314), .ZN(n2305) );
  AND2_X1 U2584 ( .A1(n2310), .A2(n2309), .ZN(n2308) );
  NAND2_X1 U2585 ( .A1(n3780), .A2(n2935), .ZN(n2327) );
  AND2_X1 U2586 ( .A1(n2933), .A2(n2934), .ZN(n2324) );
  NAND2_X1 U2587 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  NAND2_X1 U2588 ( .A1(n2911), .A2(REG3_REG_23__SCAN_IN), .ZN(n2940) );
  NOR2_X1 U2589 ( .A1(n3789), .A2(n2315), .ZN(n2314) );
  INV_X1 U2590 ( .A(n3723), .ZN(n2315) );
  NAND2_X1 U2591 ( .A1(n2312), .A2(n2311), .ZN(n2310) );
  INV_X1 U2592 ( .A(n3789), .ZN(n2312) );
  NAND2_X1 U2593 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  INV_X1 U2594 ( .A(n4413), .ZN(n2862) );
  INV_X1 U2595 ( .A(n4412), .ZN(n2863) );
  INV_X1 U2596 ( .A(n3988), .ZN(n3349) );
  CLKBUF_X1 U2597 ( .A(n2603), .Z(n3206) );
  AND2_X1 U2599 ( .A1(n4385), .A2(n3131), .ZN(n2650) );
  NAND2_X1 U2600 ( .A1(n2351), .A2(n2350), .ZN(n3171) );
  AOI21_X1 U2601 ( .B1(n2236), .B2(n3168), .A(n4475), .ZN(n2350) );
  NAND2_X1 U2602 ( .A1(n4469), .A2(n3182), .ZN(n4470) );
  XNOR2_X1 U2603 ( .A(n3172), .B(n4623), .ZN(n4486) );
  NAND2_X1 U2604 ( .A1(n4486), .A2(REG1_REG_6__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U2605 ( .A1(n3188), .A2(n3187), .ZN(n3486) );
  AOI21_X1 U2606 ( .B1(REG1_REG_9__SCAN_IN), .B2(n3501), .A(n4503), .ZN(n3502)
         );
  NAND2_X1 U2607 ( .A1(n2354), .A2(n2353), .ZN(n3576) );
  INV_X1 U2608 ( .A(n3506), .ZN(n2353) );
  XNOR2_X1 U2609 ( .A(n4039), .B(n2278), .ZN(n3582) );
  NAND2_X1 U2610 ( .A1(n3582), .A2(REG2_REG_12__SCAN_IN), .ZN(n4041) );
  OR2_X1 U2611 ( .A1(n4025), .A2(n4543), .ZN(n4026) );
  NOR2_X1 U2612 ( .A1(n4540), .A2(n4539), .ZN(n4538) );
  NOR2_X1 U2613 ( .A1(n2273), .A2(n4587), .ZN(n4586) );
  NOR2_X1 U2614 ( .A1(n2951), .A2(n5043), .ZN(n2965) );
  AND2_X1 U2615 ( .A1(n2965), .A2(REG3_REG_27__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U2616 ( .A1(n2265), .A2(n2416), .ZN(n2413) );
  AND2_X1 U2617 ( .A1(n3099), .A2(n3815), .ZN(n4103) );
  AOI21_X1 U2618 ( .B1(n4168), .B2(n3059), .A(n3058), .ZN(n4150) );
  NOR2_X1 U2619 ( .A1(n4191), .A2(n4179), .ZN(n3058) );
  OAI21_X1 U2620 ( .B1(n4248), .B2(n2396), .A(n2395), .ZN(n4188) );
  OR2_X1 U2621 ( .A1(n2401), .A2(n2254), .ZN(n2396) );
  OR2_X1 U2622 ( .A1(n2398), .A2(n2254), .ZN(n2395) );
  AND2_X1 U2623 ( .A1(n2406), .A2(n3056), .ZN(n2403) );
  AOI21_X1 U2624 ( .B1(n2380), .B2(n2379), .A(n2261), .ZN(n2378) );
  INV_X1 U2625 ( .A(n2252), .ZN(n2379) );
  NAND2_X1 U2626 ( .A1(n2252), .A2(n3052), .ZN(n2382) );
  OR2_X1 U2627 ( .A1(n3983), .A2(n3628), .ZN(n3051) );
  AND2_X1 U2628 ( .A1(n2785), .A2(REG3_REG_13__SCAN_IN), .ZN(n2794) );
  NAND2_X1 U2629 ( .A1(n3355), .A2(n2386), .ZN(n2385) );
  NOR2_X1 U2630 ( .A1(n2389), .A2(n2428), .ZN(n2386) );
  OR2_X1 U2631 ( .A1(n2387), .A2(n2428), .ZN(n2384) );
  AOI21_X1 U2632 ( .B1(n2390), .B2(n2388), .A(n2250), .ZN(n2387) );
  INV_X1 U2633 ( .A(n2245), .ZN(n2388) );
  INV_X1 U2634 ( .A(n3274), .ZN(n3430) );
  NAND2_X1 U2635 ( .A1(n3330), .A2(n3915), .ZN(n2298) );
  NAND2_X1 U2636 ( .A1(n2551), .A2(n2537), .ZN(n3134) );
  XNOR2_X1 U2637 ( .A(n2573), .B(n3127), .ZN(n2579) );
  NAND2_X1 U2638 ( .A1(n3130), .A2(IR_REG_31__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U2639 ( .A1(n2572), .A2(IR_REG_31__SCAN_IN), .ZN(n2575) );
  INV_X1 U2640 ( .A(n2522), .ZN(n2523) );
  OAI21_X1 U2641 ( .B1(n2557), .B2(n2556), .A(n2555), .ZN(n3142) );
  OR2_X1 U2642 ( .A1(n2554), .A2(n2553), .ZN(n2557) );
  NAND2_X1 U2643 ( .A1(n2466), .A2(n2436), .ZN(n2486) );
  AND4_X1 U2644 ( .A1(n2435), .A2(n2434), .A3(n2433), .A4(n2481), .ZN(n2436)
         );
  INV_X1 U2645 ( .A(IR_REG_8__SCAN_IN), .ZN(n2433) );
  INV_X1 U2646 ( .A(IR_REG_11__SCAN_IN), .ZN(n2481) );
  OR2_X1 U2647 ( .A1(n2477), .A2(IR_REG_9__SCAN_IN), .ZN(n2480) );
  INV_X1 U2648 ( .A(n4107), .ZN(n3736) );
  NAND2_X1 U2649 ( .A1(n3733), .A2(n3732), .ZN(n2301) );
  MUX2_X1 U2650 ( .A(n3146), .B(DATAI_2_), .S(n2521), .Z(n3448) );
  INV_X1 U2651 ( .A(n4234), .ZN(n4410) );
  INV_X1 U2652 ( .A(n4446), .ZN(n3812) );
  AND2_X1 U2653 ( .A1(n2994), .A2(n2993), .ZN(n4441) );
  NOR2_X1 U2654 ( .A1(n4536), .A2(n4537), .ZN(n4535) );
  INV_X1 U2655 ( .A(n4584), .ZN(n2360) );
  NOR2_X1 U2656 ( .A1(n4586), .A2(n2271), .ZN(n4589) );
  NAND2_X1 U2657 ( .A1(n2272), .A2(n4588), .ZN(n2271) );
  NAND2_X1 U2658 ( .A1(n2273), .A2(n4587), .ZN(n2272) );
  AOI21_X1 U2659 ( .B1(n4585), .B2(n4584), .A(n4583), .ZN(n4590) );
  INV_X1 U2660 ( .A(n4577), .ZN(n4583) );
  NAND2_X1 U2661 ( .A1(n4573), .A2(n2270), .ZN(n2357) );
  AND2_X1 U2662 ( .A1(n2975), .A2(REG3_REG_28__SCAN_IN), .ZN(n4075) );
  NAND2_X1 U2663 ( .A1(n2347), .A2(n4400), .ZN(n4345) );
  NAND2_X1 U2664 ( .A1(n2558), .A2(n2520), .ZN(n4058) );
  OR2_X1 U2665 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  INV_X1 U2666 ( .A(n4052), .ZN(n4608) );
  INV_X1 U2667 ( .A(n3590), .ZN(n2332) );
  INV_X1 U2668 ( .A(IR_REG_13__SCAN_IN), .ZN(n4781) );
  NOR2_X1 U2669 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2441)
         );
  OR2_X1 U2670 ( .A1(n2724), .A2(n3426), .ZN(n2726) );
  NAND2_X1 U2671 ( .A1(n2330), .A2(n2329), .ZN(n2831) );
  AOI21_X1 U2672 ( .B1(n2334), .B2(n2331), .A(n2269), .ZN(n2329) );
  NAND2_X1 U2673 ( .A1(n3534), .A2(n2331), .ZN(n2330) );
  AND2_X1 U2674 ( .A1(n2333), .A2(n2332), .ZN(n2331) );
  NAND2_X1 U2675 ( .A1(n4479), .A2(REG1_REG_5__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U2676 ( .A1(n2362), .A2(n2361), .ZN(n2364) );
  AOI21_X1 U2677 ( .B1(n4028), .B2(n2363), .A(n2426), .ZN(n2361) );
  NAND2_X1 U2678 ( .A1(n4538), .A2(n2363), .ZN(n2362) );
  AOI21_X1 U2679 ( .B1(n3088), .B2(n2284), .A(n2282), .ZN(n2281) );
  NAND2_X1 U2680 ( .A1(n2283), .A2(n3949), .ZN(n2282) );
  NAND2_X1 U2681 ( .A1(n2284), .A2(n2286), .ZN(n2283) );
  AOI21_X1 U2682 ( .B1(n2400), .B2(n2399), .A(n2262), .ZN(n2398) );
  INV_X1 U2683 ( .A(n2403), .ZN(n2399) );
  AND2_X1 U2684 ( .A1(n4170), .A2(n3089), .ZN(n3865) );
  NOR2_X1 U2685 ( .A1(n2294), .A2(n3892), .ZN(n2293) );
  NOR2_X1 U2686 ( .A1(n3040), .A2(n3372), .ZN(n3043) );
  NAND2_X1 U2687 ( .A1(n3349), .A2(n3322), .ZN(n3068) );
  NAND2_X1 U2688 ( .A1(n3911), .A2(n3908), .ZN(n3259) );
  OAI21_X1 U2689 ( .B1(n4118), .B2(n4195), .A(n3103), .ZN(n3104) );
  INV_X1 U2690 ( .A(n4126), .ZN(n3096) );
  NAND2_X1 U2691 ( .A1(n4318), .A2(n2242), .ZN(n4123) );
  NOR2_X1 U2692 ( .A1(n3094), .A2(n3095), .ZN(n2345) );
  INV_X1 U2693 ( .A(n3517), .ZN(n3523) );
  NOR2_X1 U2694 ( .A1(n2237), .A2(n3322), .ZN(n2338) );
  NAND2_X1 U2695 ( .A1(n3026), .A2(n2609), .ZN(n3315) );
  NAND4_X1 U2696 ( .A1(n4781), .A2(n2505), .A3(n2507), .A4(n2504), .ZN(n2437)
         );
  AND2_X1 U2697 ( .A1(n2421), .A2(n2420), .ZN(n2574) );
  NOR2_X1 U2698 ( .A1(n2522), .A2(IR_REG_26__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U2699 ( .A1(n2257), .A2(n2297), .ZN(n2522) );
  INV_X1 U2700 ( .A(IR_REG_20__SCAN_IN), .ZN(n2559) );
  AND2_X1 U2701 ( .A1(n2803), .A2(n2804), .ZN(n3590) );
  INV_X1 U2702 ( .A(n2627), .ZN(n2986) );
  AND2_X1 U2703 ( .A1(n3144), .A2(DATAI_24_), .ZN(n3095) );
  OR2_X1 U2704 ( .A1(n2712), .A2(n2701), .ZN(n2743) );
  AND2_X1 U2705 ( .A1(n2877), .A2(n2876), .ZN(n2311) );
  AND2_X1 U2706 ( .A1(n2766), .A2(n2765), .ZN(n3543) );
  AND2_X1 U2707 ( .A1(n2767), .A2(REG3_REG_12__SCAN_IN), .ZN(n2785) );
  NOR2_X1 U2708 ( .A1(n2901), .A2(n2900), .ZN(n2911) );
  NOR2_X1 U2709 ( .A1(n2758), .A2(n3439), .ZN(n2767) );
  INV_X1 U2710 ( .A(n2622), .ZN(n2303) );
  AND2_X1 U2711 ( .A1(n2600), .A2(n3006), .ZN(n3011) );
  INV_X1 U2712 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2280) );
  NAND2_X1 U2713 ( .A1(n4487), .A2(n3185), .ZN(n3188) );
  NAND2_X1 U2714 ( .A1(n2369), .A2(n2371), .ZN(n2368) );
  OR2_X1 U2715 ( .A1(n4513), .A2(n3503), .ZN(n2354) );
  INV_X1 U2716 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3439) );
  AND2_X1 U2717 ( .A1(n2244), .A2(n2349), .ZN(n4525) );
  NOR2_X1 U2718 ( .A1(n4525), .A2(n4524), .ZN(n4523) );
  XNOR2_X1 U2719 ( .A(n2364), .B(n4612), .ZN(n4564) );
  NAND2_X1 U2720 ( .A1(n4564), .A2(n4563), .ZN(n4562) );
  NOR2_X1 U2721 ( .A1(n4551), .A2(n4047), .ZN(n4048) );
  INV_X1 U2722 ( .A(n4046), .ZN(n4047) );
  NAND2_X1 U2723 ( .A1(n4570), .A2(n4051), .ZN(n2273) );
  NAND2_X1 U2724 ( .A1(n4083), .A2(n4082), .ZN(n4284) );
  NAND2_X1 U2725 ( .A1(n2409), .A2(n2408), .ZN(n4079) );
  AOI21_X1 U2726 ( .B1(n2411), .B2(n2412), .A(n2259), .ZN(n2408) );
  OAI21_X1 U2727 ( .B1(n3088), .B2(n2286), .A(n2284), .ZN(n4152) );
  NAND2_X1 U2728 ( .A1(n4188), .A2(n4189), .ZN(n4187) );
  NAND2_X1 U2729 ( .A1(n3088), .A2(n3946), .ZN(n4217) );
  AND2_X1 U2730 ( .A1(n3144), .A2(DATAI_21_), .ZN(n4210) );
  NOR2_X1 U2731 ( .A1(n4241), .A2(n4210), .ZN(n4209) );
  AND2_X1 U2732 ( .A1(n2865), .A2(REG3_REG_19__SCAN_IN), .ZN(n2878) );
  INV_X1 U2733 ( .A(n2372), .ZN(n3690) );
  NAND2_X1 U2734 ( .A1(n2380), .A2(n3053), .ZN(n2376) );
  INV_X1 U2735 ( .A(n2374), .ZN(n2373) );
  INV_X1 U2736 ( .A(n3684), .ZN(n3701) );
  NOR2_X1 U2737 ( .A1(n3636), .A2(n3077), .ZN(n2347) );
  NOR2_X1 U2738 ( .A1(n2817), .A2(n4398), .ZN(n2838) );
  NAND2_X1 U2739 ( .A1(n3669), .A2(n3851), .ZN(n3668) );
  INV_X1 U2740 ( .A(n2807), .ZN(n2808) );
  NAND2_X1 U2741 ( .A1(n2794), .A2(REG3_REG_14__SCAN_IN), .ZN(n2807) );
  AND4_X1 U2742 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(n3631)
         );
  NAND2_X1 U2743 ( .A1(n3075), .A2(n3891), .ZN(n3561) );
  NOR2_X1 U2744 ( .A1(n2394), .A2(n2248), .ZN(n2390) );
  INV_X1 U2745 ( .A(n3359), .ZN(n3519) );
  NAND2_X1 U2746 ( .A1(n3070), .A2(n3922), .ZN(n3357) );
  INV_X1 U2747 ( .A(n4195), .ZN(n4260) );
  AND3_X1 U2748 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U2749 ( .A1(n2510), .A2(n2316), .ZN(n2318) );
  AND2_X1 U2750 ( .A1(n2509), .A2(n2514), .ZN(n2316) );
  INV_X1 U2751 ( .A(IR_REG_18__SCAN_IN), .ZN(n2515) );
  AND2_X1 U2752 ( .A1(n2510), .A2(n2509), .ZN(n2516) );
  NAND2_X1 U2753 ( .A1(n4386), .A2(n3141), .ZN(n4195) );
  NAND2_X1 U2754 ( .A1(n3967), .A2(n3100), .ZN(n4197) );
  INV_X1 U2755 ( .A(n4197), .ZN(n4262) );
  NOR2_X1 U2756 ( .A1(n4284), .A2(n4288), .ZN(n4283) );
  AND2_X1 U2757 ( .A1(n4391), .A2(n4629), .ZN(n4287) );
  AND2_X1 U2758 ( .A1(n3116), .A2(n3118), .ZN(n4083) );
  NOR2_X1 U2759 ( .A1(n4123), .A2(n3096), .ZN(n4124) );
  NAND2_X1 U2760 ( .A1(n4318), .A2(n2345), .ZN(n4160) );
  NAND2_X1 U2761 ( .A1(n4318), .A2(n4179), .ZN(n4178) );
  AND2_X1 U2762 ( .A1(n4209), .A2(n4202), .ZN(n4318) );
  NAND2_X1 U2763 ( .A1(n3705), .A2(n2340), .ZN(n4241) );
  AND2_X1 U2764 ( .A1(n2341), .A2(n4226), .ZN(n2340) );
  INV_X1 U2765 ( .A(n2347), .ZN(n3673) );
  NOR2_X1 U2766 ( .A1(n3616), .A2(n3615), .ZN(n3638) );
  NAND2_X1 U2767 ( .A1(n3524), .A2(n3523), .ZN(n3568) );
  OR2_X1 U2768 ( .A1(n3568), .A2(n3567), .ZN(n3616) );
  NOR2_X1 U2769 ( .A1(n3369), .A2(n3432), .ZN(n3469) );
  AND2_X1 U2770 ( .A1(n3469), .A2(n3477), .ZN(n3524) );
  INV_X1 U2771 ( .A(n4656), .ZN(n4661) );
  NAND2_X1 U2772 ( .A1(n2337), .A2(n2338), .ZN(n3367) );
  INV_X1 U2773 ( .A(n3331), .ZN(n3329) );
  NOR2_X1 U2774 ( .A1(n3252), .A2(n3411), .ZN(n3416) );
  NOR2_X1 U2775 ( .A1(n3252), .A2(n2237), .ZN(n3327) );
  NAND2_X1 U2776 ( .A1(n3613), .A2(n4668), .ZN(n4656) );
  NOR2_X1 U2777 ( .A1(n3315), .A2(n3448), .ZN(n4636) );
  INV_X1 U2778 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4892) );
  AOI21_X1 U2779 ( .B1(n2533), .B2(IR_REG_25__SCAN_IN), .A(n2532), .ZN(n2534)
         );
  XOR2_X1 U2780 ( .A(n2562), .B(n2569), .Z(n3869) );
  INV_X1 U2781 ( .A(IR_REG_15__SCAN_IN), .ZN(n2506) );
  OR2_X1 U2782 ( .A1(n2494), .A2(n2553), .ZN(n2501) );
  AND2_X1 U2783 ( .A1(n2510), .A2(n2507), .ZN(n2494) );
  INV_X1 U2784 ( .A(n2510), .ZN(n2490) );
  AND2_X1 U2785 ( .A1(n2478), .A2(n2480), .ZN(n3501) );
  INV_X1 U2786 ( .A(IR_REG_6__SCAN_IN), .ZN(n2432) );
  INV_X1 U2787 ( .A(n2452), .ZN(n2417) );
  NOR2_X1 U2788 ( .A1(n3291), .A2(n3292), .ZN(n2321) );
  AOI21_X1 U2789 ( .B1(n2246), .B2(n3291), .A(n2320), .ZN(n2319) );
  INV_X1 U2790 ( .A(n3628), .ZN(n3637) );
  OR2_X1 U2791 ( .A1(n3534), .A2(n2334), .ZN(n2328) );
  NAND2_X1 U2792 ( .A1(n2741), .A2(n2740), .ZN(n3480) );
  AND4_X2 U2793 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(n3386)
         );
  NAND2_X1 U2794 ( .A1(n3144), .A2(DATAI_3_), .ZN(n2453) );
  NAND2_X1 U2795 ( .A1(n2308), .A2(n4417), .ZN(n2306) );
  NAND2_X1 U2796 ( .A1(n2308), .A2(n2305), .ZN(n2304) );
  INV_X1 U2797 ( .A(n4415), .ZN(n2307) );
  AOI21_X1 U2798 ( .B1(n2937), .B2(n2325), .A(n2324), .ZN(n2323) );
  NAND2_X1 U2799 ( .A1(n3797), .A2(n2258), .ZN(n2326) );
  INV_X1 U2800 ( .A(n3780), .ZN(n2325) );
  OAI21_X1 U2801 ( .B1(n3739), .B2(n2933), .A(n2934), .ZN(n3779) );
  OAI21_X1 U2802 ( .B1(n2521), .B2(n2459), .A(n2458), .ZN(n3261) );
  INV_X1 U2803 ( .A(n4461), .ZN(n2459) );
  AND4_X1 U2804 ( .A1(n2892), .A2(n2891), .A3(n2890), .A4(n2889), .ZN(n4227)
         );
  NAND2_X1 U2805 ( .A1(n3014), .A2(n4386), .ZN(n4430) );
  NAND2_X1 U2806 ( .A1(n2313), .A2(n2310), .ZN(n3787) );
  NAND2_X1 U2807 ( .A1(n3722), .A2(n2314), .ZN(n2313) );
  AOI21_X1 U2808 ( .B1(n3722), .B2(n3723), .A(n2311), .ZN(n3791) );
  INV_X1 U2809 ( .A(n3076), .ZN(n3615) );
  NAND2_X1 U2810 ( .A1(n3750), .A2(n2622), .ZN(n3224) );
  NAND2_X1 U2811 ( .A1(n3014), .A2(n3013), .ZN(n4429) );
  NAND2_X1 U2812 ( .A1(n3245), .A2(n2676), .ZN(n3294) );
  AND2_X1 U2813 ( .A1(n3007), .A2(n3197), .ZN(n4446) );
  AND4_X1 U2814 ( .A1(n2824), .A2(n2823), .A3(n2822), .A4(n2821), .ZN(n4428)
         );
  INV_X1 U2815 ( .A(n3631), .ZN(n3984) );
  NAND2_X1 U2816 ( .A1(n2697), .A2(n2696), .ZN(n3988) );
  AND2_X1 U2817 ( .A1(n2695), .A2(n2424), .ZN(n2697) );
  NAND4_X1 U2818 ( .A1(n2683), .A2(n2682), .A3(n2681), .A4(n2680), .ZN(n3989)
         );
  OR2_X1 U2819 ( .A1(n2597), .A2(n4606), .ZN(n4004) );
  NAND2_X1 U2820 ( .A1(n2656), .A2(n2655), .ZN(n3991) );
  AND3_X1 U2821 ( .A1(n2654), .A2(n2653), .A3(n2652), .ZN(n2655) );
  INV_X1 U2822 ( .A(n3386), .ZN(n3753) );
  NAND2_X1 U2823 ( .A1(n2650), .A2(REG3_REG_1__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U2824 ( .A1(n3148), .A2(n4015), .ZN(n4019) );
  INV_X1 U2825 ( .A(n2352), .ZN(n4476) );
  OAI21_X1 U2826 ( .B1(n4459), .B2(n3168), .A(n2236), .ZN(n2352) );
  XNOR2_X1 U2827 ( .A(n3184), .B(n4623), .ZN(n4488) );
  NAND2_X1 U2828 ( .A1(n4488), .A2(REG2_REG_6__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U2829 ( .A1(n4498), .A2(n3489), .ZN(n4509) );
  NAND2_X1 U2830 ( .A1(n4509), .A2(n4510), .ZN(n4508) );
  XNOR2_X1 U2831 ( .A(n3502), .B(n4522), .ZN(n4514) );
  NOR2_X1 U2832 ( .A1(n4514), .A2(n4515), .ZN(n4513) );
  INV_X1 U2833 ( .A(n2354), .ZN(n3507) );
  INV_X1 U2834 ( .A(n2349), .ZN(n2348) );
  NAND2_X1 U2835 ( .A1(n2244), .A2(n3578), .ZN(n3579) );
  NAND2_X1 U2836 ( .A1(n4041), .A2(n4040), .ZN(n4530) );
  NAND2_X1 U2837 ( .A1(n2277), .A2(n2274), .ZN(n4536) );
  NAND2_X1 U2838 ( .A1(n2276), .A2(n2275), .ZN(n2274) );
  INV_X1 U2839 ( .A(n4543), .ZN(n2275) );
  NOR2_X1 U2840 ( .A1(n4549), .A2(n4548), .ZN(n4547) );
  NOR2_X1 U2841 ( .A1(n4538), .A2(n4028), .ZN(n4549) );
  NOR2_X1 U2842 ( .A1(n4455), .A2(n4386), .ZN(n4556) );
  XNOR2_X1 U2843 ( .A(n4048), .B(n2498), .ZN(n2279) );
  NAND2_X1 U2844 ( .A1(n2279), .A2(n3674), .ZN(n4561) );
  NAND2_X1 U2845 ( .A1(n4037), .A2(n4036), .ZN(n2358) );
  OAI22_X1 U2846 ( .A1(n2243), .A2(n2358), .B1(n4036), .B2(n4037), .ZN(n2356)
         );
  OR2_X1 U2847 ( .A1(n4075), .A2(n2976), .ZN(n4090) );
  OR2_X1 U2848 ( .A1(n2975), .A2(n2966), .ZN(n4107) );
  NAND2_X1 U2849 ( .A1(n2410), .A2(n2413), .ZN(n4104) );
  NAND2_X1 U2850 ( .A1(n4132), .A2(n2414), .ZN(n2410) );
  NAND2_X1 U2851 ( .A1(n2397), .A2(n2400), .ZN(n4208) );
  NAND2_X1 U2852 ( .A1(n4248), .A2(n2403), .ZN(n2397) );
  AND2_X1 U2853 ( .A1(n2405), .A2(n2407), .ZN(n4236) );
  NAND2_X1 U2854 ( .A1(n4248), .A2(n3056), .ZN(n2405) );
  OAI21_X1 U2855 ( .B1(n3651), .B2(n2381), .A(n2378), .ZN(n3700) );
  NAND2_X1 U2856 ( .A1(n2377), .A2(n2380), .ZN(n3665) );
  NAND2_X1 U2857 ( .A1(n3651), .A2(n2252), .ZN(n2377) );
  NAND2_X1 U2858 ( .A1(n2385), .A2(n2384), .ZN(n3566) );
  NAND2_X1 U2859 ( .A1(n2391), .A2(n2393), .ZN(n3468) );
  INV_X1 U2860 ( .A(n2394), .ZN(n2393) );
  OR2_X1 U2861 ( .A1(n2564), .A2(n3120), .ZN(n2566) );
  OR2_X1 U2862 ( .A1(n3140), .A2(n3111), .ZN(n4268) );
  INV_X1 U2863 ( .A(n4598), .ZN(n4266) );
  AND2_X1 U2864 ( .A1(n3286), .A2(n2598), .ZN(n4598) );
  INV_X1 U2865 ( .A(n4268), .ZN(n4594) );
  INV_X1 U2866 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2290) );
  AND2_X2 U2867 ( .A1(n3121), .A2(n3120), .ZN(n4684) );
  XNOR2_X1 U2868 ( .A(n4283), .B(n2339), .ZN(n4278) );
  INV_X1 U2869 ( .A(n3965), .ZN(n2339) );
  NAND2_X1 U2870 ( .A1(n2228), .A2(n2291), .ZN(n3123) );
  OR2_X1 U2871 ( .A1(n4088), .A2(n4661), .ZN(n2291) );
  AND2_X1 U2872 ( .A1(n3705), .A2(n4420), .ZN(n4265) );
  AND2_X2 U2873 ( .A1(n3122), .A2(n3121), .ZN(n4673) );
  INV_X1 U2874 ( .A(n4606), .ZN(n3137) );
  AND2_X1 U2875 ( .A1(n2563), .A2(n2529), .ZN(n3135) );
  NAND2_X1 U2876 ( .A1(n3198), .A2(n3134), .ZN(n4685) );
  NOR2_X1 U2877 ( .A1(n2571), .A2(IR_REG_29__SCAN_IN), .ZN(n2419) );
  INV_X1 U2878 ( .A(IR_REG_30__SCAN_IN), .ZN(n3127) );
  INV_X1 U2879 ( .A(n3013), .ZN(n4386) );
  NAND2_X1 U2880 ( .A1(n2535), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  XNOR2_X1 U2881 ( .A(n2528), .B(IR_REG_24__SCAN_IN), .ZN(n4388) );
  INV_X1 U2882 ( .A(n2567), .ZN(n4389) );
  AND2_X1 U2883 ( .A1(n2483), .A2(n2484), .ZN(n4394) );
  NAND2_X1 U2884 ( .A1(n2450), .A2(IR_REG_31__SCAN_IN), .ZN(n2451) );
  INV_X1 U2885 ( .A(n2449), .ZN(n2450) );
  NAND2_X1 U2886 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2446)
         );
  NAND2_X1 U2887 ( .A1(n2301), .A2(n2427), .ZN(n2300) );
  AOI21_X1 U2888 ( .B1(n4582), .B2(n4590), .A(n4589), .ZN(n4591) );
  NAND2_X1 U2889 ( .A1(n4573), .A2(n2243), .ZN(n4582) );
  OAI211_X1 U2890 ( .C1(n4573), .C2(n2358), .A(n2357), .B(n2355), .ZN(n4062)
         );
  INV_X1 U2891 ( .A(n2356), .ZN(n2355) );
  INV_X1 U2892 ( .A(n2287), .ZN(U3546) );
  AOI21_X1 U2893 ( .B1(n3123), .B2(n4684), .A(n2288), .ZN(n2287) );
  NAND2_X1 U2894 ( .A1(n3119), .A2(n2289), .ZN(n2288) );
  OR2_X1 U2895 ( .A1(n4684), .A2(n2290), .ZN(n2289) );
  NAND2_X1 U2896 ( .A1(n3169), .A2(n4461), .ZN(n2236) );
  NAND2_X1 U2897 ( .A1(n3329), .A2(n3418), .ZN(n2237) );
  AND2_X1 U2898 ( .A1(n4410), .A2(n4264), .ZN(n3055) );
  INV_X1 U2899 ( .A(n3366), .ZN(n2336) );
  NAND2_X1 U2900 ( .A1(n2417), .A2(n2431), .ZN(n2460) );
  INV_X1 U2901 ( .A(n2401), .ZN(n2400) );
  NOR2_X1 U2902 ( .A1(n2404), .A2(n2402), .ZN(n2401) );
  AND2_X1 U2903 ( .A1(n2752), .A2(n2740), .ZN(n2238) );
  NOR2_X1 U2904 ( .A1(n4155), .A2(n3061), .ZN(n2239) );
  AND2_X1 U2905 ( .A1(n4118), .A2(n4106), .ZN(n2240) );
  OR2_X1 U2906 ( .A1(n3609), .A2(n3562), .ZN(n2241) );
  AND2_X1 U2907 ( .A1(n2345), .A2(n3061), .ZN(n2242) );
  AND2_X1 U2908 ( .A1(n2360), .A2(n4035), .ZN(n2243) );
  NAND4_X1 U2909 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .ZN(n3025)
         );
  NAND2_X1 U2910 ( .A1(n3577), .A2(n4393), .ZN(n2244) );
  AND3_X1 U2911 ( .A1(n2346), .A2(n2449), .A3(n2431), .ZN(n2462) );
  OR2_X1 U2912 ( .A1(n3987), .A2(n3432), .ZN(n2245) );
  NAND2_X1 U2913 ( .A1(n2676), .A2(n2322), .ZN(n2246) );
  OR2_X1 U2914 ( .A1(n3739), .A2(n2937), .ZN(n2247) );
  AND2_X1 U2915 ( .A1(n3359), .A2(n3073), .ZN(n2248) );
  NAND2_X1 U2916 ( .A1(n2449), .A2(n2429), .ZN(n2452) );
  NAND2_X1 U2917 ( .A1(n2568), .A2(n2569), .ZN(n2249) );
  NAND2_X1 U2918 ( .A1(n3512), .A2(n3048), .ZN(n2250) );
  AND2_X1 U2919 ( .A1(n4124), .A2(n4106), .ZN(n3116) );
  INV_X1 U2920 ( .A(n3355), .ZN(n2392) );
  NOR2_X1 U2921 ( .A1(n2571), .A2(IR_REG_21__SCAN_IN), .ZN(n2526) );
  INV_X1 U2922 ( .A(IR_REG_21__SCAN_IN), .ZN(n2569) );
  AND2_X1 U2923 ( .A1(n3921), .A2(n3068), .ZN(n2251) );
  NAND2_X1 U2924 ( .A1(n3478), .A2(n2757), .ZN(n3437) );
  OR2_X1 U2925 ( .A1(n4397), .A2(n4432), .ZN(n2252) );
  INV_X1 U2926 ( .A(IR_REG_25__SCAN_IN), .ZN(n2297) );
  AND4_X1 U2927 ( .A1(n2346), .A2(n2431), .A3(n2432), .A4(n2449), .ZN(n2466)
         );
  INV_X1 U2928 ( .A(n3991), .ZN(n3031) );
  NAND2_X1 U2929 ( .A1(n3705), .A2(n2341), .ZN(n4238) );
  NAND2_X1 U2930 ( .A1(n3666), .A2(n2382), .ZN(n2381) );
  NAND2_X1 U2931 ( .A1(n4415), .A2(n4417), .ZN(n3722) );
  NAND2_X1 U2932 ( .A1(n2328), .A2(n2333), .ZN(n3589) );
  INV_X1 U2933 ( .A(n3891), .ZN(n2294) );
  INV_X1 U2934 ( .A(n3292), .ZN(n2322) );
  NOR2_X1 U2935 ( .A1(n2486), .A2(IR_REG_13__SCAN_IN), .ZN(n2510) );
  AND2_X1 U2936 ( .A1(n4173), .A2(n4161), .ZN(n2253) );
  INV_X1 U2937 ( .A(n3322), .ZN(n3285) );
  OAI21_X1 U2938 ( .B1(n3144), .B2(n3191), .A(n2472), .ZN(n3322) );
  AND2_X1 U2939 ( .A1(n4227), .A2(n4214), .ZN(n2254) );
  AND2_X1 U2940 ( .A1(n4143), .A2(n3096), .ZN(n2255) );
  AND2_X1 U2941 ( .A1(n4257), .A2(n4226), .ZN(n2256) );
  AND2_X1 U2942 ( .A1(n2552), .A2(n2441), .ZN(n2257) );
  AND2_X1 U2943 ( .A1(n2938), .A2(n2327), .ZN(n2258) );
  INV_X1 U2944 ( .A(n2415), .ZN(n2414) );
  NAND2_X1 U2945 ( .A1(n2416), .A2(n3062), .ZN(n2415) );
  AND2_X1 U2946 ( .A1(n3978), .A2(n3098), .ZN(n2259) );
  AND2_X1 U2947 ( .A1(n2348), .A2(n2244), .ZN(n2260) );
  NOR2_X1 U2948 ( .A1(n4428), .A2(n4400), .ZN(n2261) );
  AND2_X1 U2949 ( .A1(n3218), .A2(n4210), .ZN(n2262) );
  NAND2_X1 U2950 ( .A1(n3717), .A2(n3981), .ZN(n2263) );
  INV_X1 U2951 ( .A(IR_REG_28__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U2952 ( .A1(n2999), .A2(n4441), .ZN(n2264) );
  INV_X1 U2953 ( .A(n4479), .ZN(n3183) );
  AND2_X1 U2954 ( .A1(n2464), .A2(n2463), .ZN(n4479) );
  INV_X1 U2955 ( .A(n2381), .ZN(n2380) );
  INV_X1 U2956 ( .A(IR_REG_29__SCAN_IN), .ZN(n2572) );
  OR2_X1 U2957 ( .A1(n2239), .A2(n2255), .ZN(n2265) );
  OR2_X1 U2958 ( .A1(n3985), .A2(n3567), .ZN(n2266) );
  AND2_X1 U2959 ( .A1(n2897), .A2(n3761), .ZN(n2267) );
  OR2_X1 U2960 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2268)
         );
  NAND2_X1 U2961 ( .A1(n3638), .A2(n3637), .ZN(n3636) );
  OAI21_X1 U2962 ( .B1(n3245), .B2(n2321), .A(n2319), .ZN(n3318) );
  INV_X1 U2963 ( .A(n4420), .ZN(n2342) );
  OAI21_X1 U2964 ( .B1(n3410), .B2(n3408), .A(n3916), .ZN(n3330) );
  XNOR2_X1 U2965 ( .A(n2524), .B(IR_REG_26__SCAN_IN), .ZN(n2551) );
  AND2_X1 U2966 ( .A1(n2806), .A2(n2805), .ZN(n2269) );
  INV_X1 U2967 ( .A(IR_REG_14__SCAN_IN), .ZN(n2507) );
  AND2_X1 U2968 ( .A1(n2888), .A2(n2887), .ZN(n3788) );
  INV_X1 U2969 ( .A(n3788), .ZN(n2309) );
  INV_X1 U2970 ( .A(n4192), .ZN(n4202) );
  AND2_X1 U2971 ( .A1(n3144), .A2(DATAI_22_), .ZN(n4192) );
  INV_X1 U2972 ( .A(n3055), .ZN(n2407) );
  INV_X1 U2973 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U2974 ( .A1(n2595), .A2(n4629), .ZN(n3251) );
  OR2_X1 U2975 ( .A1(n3396), .A2(n3261), .ZN(n3252) );
  INV_X1 U2976 ( .A(n3252), .ZN(n2337) );
  OAI21_X1 U2977 ( .B1(n2571), .B2(n2249), .A(IR_REG_31__SCAN_IN), .ZN(n2583)
         );
  NAND2_X1 U2978 ( .A1(n3222), .A2(n2636), .ZN(n3228) );
  AND2_X1 U2979 ( .A1(n2243), .A2(n2359), .ZN(n2270) );
  AND2_X1 U2980 ( .A1(n3144), .A2(DATAI_23_), .ZN(n3094) );
  INV_X1 U2981 ( .A(n3094), .ZN(n4179) );
  NAND2_X1 U2982 ( .A1(n2302), .A2(n3750), .ZN(n3222) );
  INV_X1 U2983 ( .A(IR_REG_16__SCAN_IN), .ZN(n2505) );
  INV_X1 U2984 ( .A(IR_REG_3__SCAN_IN), .ZN(n2454) );
  INV_X1 U2985 ( .A(n4393), .ZN(n2278) );
  INV_X1 U2986 ( .A(DATAI_0_), .ZN(n2343) );
  NAND2_X1 U2987 ( .A1(n3993), .A2(n3994), .ZN(n3992) );
  INV_X1 U2988 ( .A(n4037), .ZN(n2359) );
  INV_X1 U2989 ( .A(IR_REG_0__SCAN_IN), .ZN(n2344) );
  INV_X1 U2990 ( .A(n4044), .ZN(n2276) );
  INV_X1 U2991 ( .A(n4045), .ZN(n2277) );
  XNOR2_X1 U2992 ( .A(n3492), .B(n4522), .ZN(n4519) );
  OAI21_X1 U2993 ( .B1(n2279), .B2(n3674), .A(n4561), .ZN(n4566) );
  INV_X1 U2994 ( .A(n2281), .ZN(n4138) );
  OAI21_X1 U2995 ( .B1(n3063), .B2(n3897), .A(n3901), .ZN(n3447) );
  INV_X1 U2996 ( .A(n3878), .ZN(n3065) );
  NAND2_X1 U2997 ( .A1(n2292), .A2(n3902), .ZN(n3385) );
  NAND2_X1 U2998 ( .A1(n2295), .A2(n3894), .ZN(n3626) );
  OAI21_X2 U2999 ( .B1(n3357), .B2(n3354), .A(n3928), .ZN(n3463) );
  OR2_X1 U3000 ( .A1(n3101), .A2(n4262), .ZN(n3106) );
  AOI21_X2 U3001 ( .B1(n4115), .B2(n3837), .A(n3962), .ZN(n4097) );
  NAND2_X1 U3002 ( .A1(n3626), .A2(n3876), .ZN(n3652) );
  NAND2_X1 U3003 ( .A1(n3901), .A2(n3898), .ZN(n3063) );
  NAND2_X1 U3004 ( .A1(n4138), .A2(n3955), .ZN(n4115) );
  OAI21_X1 U3005 ( .B1(n3260), .B2(n3067), .A(n3911), .ZN(n3410) );
  NAND2_X2 U3006 ( .A1(n2440), .A2(n2439), .ZN(n2571) );
  NAND2_X1 U3007 ( .A1(n2576), .A2(n2575), .ZN(n2577) );
  OAI211_X1 U3008 ( .C1(n2301), .C2(n2264), .A(n2423), .B(n2300), .ZN(U3217)
         );
  NOR2_X1 U3009 ( .A1(n3221), .A2(n2303), .ZN(n2302) );
  XNOR2_X1 U3010 ( .A(n2632), .B(n2633), .ZN(n3221) );
  NAND2_X1 U3011 ( .A1(n3318), .A2(n2725), .ZN(n2736) );
  NAND2_X1 U3012 ( .A1(n2741), .A2(n2238), .ZN(n3478) );
  NAND3_X1 U3013 ( .A1(n2337), .A2(n2338), .A3(n2336), .ZN(n3369) );
  INV_X1 U3014 ( .A(n2609), .ZN(n4628) );
  MUX2_X1 U3015 ( .A(n2344), .B(n2343), .S(n2521), .Z(n2609) );
  NAND2_X1 U3016 ( .A1(n3578), .A2(REG1_REG_12__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U3017 ( .A1(n2236), .A2(n4459), .ZN(n2351) );
  INV_X1 U3018 ( .A(n3171), .ZN(n4474) );
  NAND2_X1 U3019 ( .A1(n4573), .A2(n4035), .ZN(n4585) );
  INV_X1 U3020 ( .A(n2364), .ZN(n4031) );
  NAND2_X1 U3021 ( .A1(n4485), .A2(n3173), .ZN(n3497) );
  NAND2_X1 U3022 ( .A1(n2368), .A2(n2365), .ZN(n3498) );
  NAND2_X1 U3023 ( .A1(n2366), .A2(n4485), .ZN(n2365) );
  NAND2_X1 U3024 ( .A1(n2370), .A2(n2367), .ZN(n2366) );
  NAND2_X1 U3025 ( .A1(n3173), .A2(n2371), .ZN(n2367) );
  INV_X1 U3026 ( .A(n2370), .ZN(n2369) );
  OAI21_X1 U3027 ( .B1(n3651), .B2(n2376), .A(n2373), .ZN(n2372) );
  OAI21_X1 U3028 ( .B1(n3651), .B2(n3052), .A(n2252), .ZN(n3667) );
  NAND2_X1 U3029 ( .A1(n2383), .A2(n2241), .ZN(n3603) );
  NAND3_X1 U3030 ( .A1(n2385), .A2(n2266), .A3(n2384), .ZN(n2383) );
  INV_X1 U3031 ( .A(n2390), .ZN(n2389) );
  NAND2_X1 U3032 ( .A1(n2391), .A2(n2390), .ZN(n3513) );
  NAND2_X1 U3033 ( .A1(n2392), .A2(n2245), .ZN(n2391) );
  NOR2_X1 U3034 ( .A1(n3376), .A2(n3071), .ZN(n2394) );
  NAND2_X1 U3035 ( .A1(n4132), .A2(n2411), .ZN(n2409) );
  AOI21_X1 U3036 ( .B1(n4132), .B2(n3062), .A(n2239), .ZN(n4113) );
  INV_X1 U3037 ( .A(n2571), .ZN(n2420) );
  NAND2_X1 U3038 ( .A1(n2421), .A2(n2419), .ZN(n3130) );
  NOR2_X1 U3039 ( .A1(n2571), .A2(n2570), .ZN(n2584) );
  OAI22_X1 U3040 ( .A1(n3386), .A2(n2971), .B1(n3457), .B2(n2627), .ZN(n2628)
         );
  NAND2_X1 U3041 ( .A1(n3130), .A2(n2577), .ZN(n2578) );
  NAND2_X1 U3042 ( .A1(n2583), .A2(n2443), .ZN(n2442) );
  NAND2_X1 U3043 ( .A1(n2521), .A2(DATAI_7_), .ZN(n2472) );
  NAND2_X1 U3044 ( .A1(n2521), .A2(DATAI_1_), .ZN(n2447) );
  OR2_X1 U3045 ( .A1(n4292), .A2(n3251), .ZN(n4294) );
  INV_X1 U3046 ( .A(n2579), .ZN(n4385) );
  AOI21_X2 U3047 ( .B1(n3805), .B2(n3807), .A(n3806), .ZN(n3733) );
  OR2_X1 U3048 ( .A1(n2609), .A2(n2627), .ZN(n2422) );
  AND2_X1 U3049 ( .A1(n2471), .A2(n2473), .ZN(n4395) );
  INV_X1 U3050 ( .A(IR_REG_31__SCAN_IN), .ZN(n2553) );
  AND2_X1 U3051 ( .A1(n3023), .A2(n3022), .ZN(n2423) );
  AND2_X1 U3052 ( .A1(n2694), .A2(n2693), .ZN(n2424) );
  NAND2_X1 U3053 ( .A1(n4615), .A2(REG1_REG_13__SCAN_IN), .ZN(n2425) );
  AND2_X1 U3054 ( .A1(n4613), .A2(REG1_REG_15__SCAN_IN), .ZN(n2426) );
  INV_X1 U3055 ( .A(n3978), .ZN(n4118) );
  AND3_X1 U3056 ( .A1(n2997), .A2(n2998), .A3(n4441), .ZN(n2427) );
  AND2_X1 U3057 ( .A1(n3144), .A2(DATAI_25_), .ZN(n4141) );
  INV_X1 U3058 ( .A(n4141), .ZN(n3061) );
  AND4_X1 U3059 ( .A1(n2916), .A2(n2915), .A3(n2914), .A4(n2913), .ZN(n4191)
         );
  AND4_X1 U3060 ( .A1(n2945), .A2(n2944), .A3(n2943), .A4(n2942), .ZN(n4155)
         );
  NOR2_X1 U3061 ( .A1(n3049), .A2(n3514), .ZN(n2428) );
  INV_X1 U3062 ( .A(IR_REG_4__SCAN_IN), .ZN(n2430) );
  AND2_X1 U3063 ( .A1(n3605), .A2(n3604), .ZN(n3936) );
  INV_X1 U3064 ( .A(n3941), .ZN(n3081) );
  AND2_X1 U3065 ( .A1(n3864), .A2(n4151), .ZN(n3949) );
  NAND2_X2 U3066 ( .A1(n2597), .A2(n3269), .ZN(n2627) );
  INV_X1 U3067 ( .A(n3481), .ZN(n2752) );
  INV_X1 U3068 ( .A(n4472), .ZN(n3182) );
  INV_X1 U3069 ( .A(n4609), .ZN(n4034) );
  NAND2_X1 U3070 ( .A1(n3031), .A2(n3261), .ZN(n3908) );
  INV_X1 U3071 ( .A(IR_REG_27__SCAN_IN), .ZN(n2443) );
  INV_X1 U3072 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2689) );
  AND2_X1 U3073 ( .A1(n3741), .A2(n3742), .ZN(n2938) );
  INV_X1 U3074 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2701) );
  AND2_X1 U3075 ( .A1(n2613), .A2(IR_REG_0__SCAN_IN), .ZN(n2614) );
  XNOR2_X1 U3076 ( .A(n3165), .B(n3163), .ZN(n3164) );
  NAND2_X1 U3077 ( .A1(n4175), .A2(n4192), .ZN(n3057) );
  NAND2_X1 U3078 ( .A1(n3715), .A2(n4420), .ZN(n3054) );
  NAND2_X1 U3079 ( .A1(n3652), .A2(n3078), .ZN(n3654) );
  OR2_X1 U3080 ( .A1(n3280), .A2(n3043), .ZN(n3045) );
  AND2_X1 U3081 ( .A1(n3907), .A2(n3904), .ZN(n3877) );
  INV_X1 U3082 ( .A(n4256), .ZN(n4142) );
  AND2_X1 U3083 ( .A1(n2553), .A2(n2297), .ZN(n2532) );
  NOR2_X1 U3084 ( .A1(n2690), .A2(n2689), .ZN(n2710) );
  OR2_X1 U3085 ( .A1(n2743), .A2(n4892), .ZN(n2758) );
  INV_X1 U3086 ( .A(n2896), .ZN(n3761) );
  OR3_X1 U3087 ( .A1(n2940), .A2(n3774), .A3(n3782), .ZN(n2951) );
  AND2_X1 U3088 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2838), .ZN(n2850) );
  NAND2_X1 U3089 ( .A1(n2521), .A2(DATAI_4_), .ZN(n2458) );
  NAND2_X1 U3090 ( .A1(n2878), .A2(REG3_REG_20__SCAN_IN), .ZN(n2901) );
  AND2_X1 U3091 ( .A1(n2850), .A2(REG3_REG_18__SCAN_IN), .ZN(n2865) );
  AND2_X1 U3092 ( .A1(n3009), .A2(n4268), .ZN(n4433) );
  INV_X1 U3093 ( .A(n4090), .ZN(n3021) );
  AND4_X1 U3094 ( .A1(n2907), .A2(n2906), .A3(n2905), .A4(n2904), .ZN(n4215)
         );
  AOI22_X1 U3095 ( .A1(n4079), .A2(n4078), .B1(n4077), .B2(n4076), .ZN(n4081)
         );
  NAND2_X1 U3096 ( .A1(n2678), .A2(REG3_REG_6__SCAN_IN), .ZN(n2690) );
  INV_X1 U3097 ( .A(n3134), .ZN(n3108) );
  INV_X1 U3098 ( .A(n4287), .ZN(n4255) );
  INV_X1 U3099 ( .A(n4226), .ZN(n4239) );
  INV_X1 U3100 ( .A(n3073), .ZN(n3477) );
  INV_X1 U3101 ( .A(n4388), .ZN(n2529) );
  INV_X1 U3102 ( .A(n3082), .ZN(n3717) );
  INV_X1 U3103 ( .A(n4433), .ZN(n3752) );
  NAND2_X1 U3104 ( .A1(n2808), .A2(REG3_REG_15__SCAN_IN), .ZN(n2817) );
  AND4_X1 U3105 ( .A1(n2930), .A2(n2929), .A3(n2928), .A4(n2927), .ZN(n4173)
         );
  AND4_X1 U3106 ( .A1(n2799), .A2(n2798), .A3(n2797), .A4(n2796), .ZN(n4431)
         );
  AND4_X1 U3107 ( .A1(n2763), .A2(n2762), .A3(n2761), .A4(n2760), .ZN(n3464)
         );
  INV_X1 U3108 ( .A(n4623), .ZN(n4489) );
  NAND2_X1 U3109 ( .A1(n4518), .A2(n3493), .ZN(n3496) );
  XNOR2_X1 U3110 ( .A(n4079), .B(n4078), .ZN(n4088) );
  INV_X1 U3111 ( .A(n3865), .ZN(n4189) );
  OR2_X1 U3112 ( .A1(n3942), .A2(n3825), .ZN(n3666) );
  AND2_X1 U3113 ( .A1(n4273), .A2(n3284), .ZN(n4237) );
  AOI21_X1 U3114 ( .B1(n3108), .B2(n3136), .A(n3135), .ZN(n3120) );
  AND2_X1 U3115 ( .A1(n4294), .A2(n4293), .ZN(n4295) );
  INV_X1 U3116 ( .A(n3140), .ZN(n3198) );
  AND2_X1 U3117 ( .A1(n2495), .A2(n2496), .ZN(n4613) );
  AND2_X1 U3118 ( .A1(n3160), .A2(n3159), .ZN(n4581) );
  INV_X1 U3119 ( .A(n4441), .ZN(n4418) );
  AND4_X1 U3120 ( .A1(n3018), .A2(n3017), .A3(n3016), .A4(n3015), .ZN(n3817)
         );
  INV_X1 U3121 ( .A(n4431), .ZN(n3983) );
  INV_X1 U3122 ( .A(n4396), .ZN(n3163) );
  INV_X1 U3123 ( .A(n4615), .ZN(n4534) );
  INV_X1 U3124 ( .A(n4556), .ZN(n4593) );
  INV_X1 U3125 ( .A(n4237), .ZN(n4275) );
  OR2_X1 U3126 ( .A1(n4089), .A2(n4333), .ZN(n3119) );
  INV_X1 U3127 ( .A(n4684), .ZN(n4682) );
  OR2_X1 U3128 ( .A1(n4089), .A2(n4379), .ZN(n3125) );
  INV_X1 U3129 ( .A(n4673), .ZN(n4672) );
  INV_X1 U3130 ( .A(n4685), .ZN(n4605) );
  AND2_X1 U3131 ( .A1(n2493), .A2(n2492), .ZN(n4543) );
  NOR2_X1 U3132 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2435)
         );
  NOR2_X1 U3133 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2434)
         );
  INV_X1 U3134 ( .A(n2486), .ZN(n2440) );
  NAND4_X1 U3135 ( .A1(n2518), .A2(n2506), .A3(n2515), .A4(n2559), .ZN(n2438)
         );
  NAND2_X1 U3136 ( .A1(n2443), .A2(IR_REG_28__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3137 ( .A1(n3144), .A2(DATAI_31_), .ZN(n3965) );
  INV_X1 U3138 ( .A(n2232), .ZN(n2448) );
  INV_X1 U3139 ( .A(n2230), .ZN(n3026) );
  NAND2_X1 U3140 ( .A1(n2452), .A2(IR_REG_31__SCAN_IN), .ZN(n2455) );
  XNOR2_X1 U3141 ( .A(n2455), .B(IR_REG_3__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U3142 ( .A1(n4636), .A2(n3394), .ZN(n3396) );
  NAND2_X1 U3143 ( .A1(n2455), .A2(n2454), .ZN(n2456) );
  NAND2_X1 U3144 ( .A1(n2456), .A2(IR_REG_31__SCAN_IN), .ZN(n2457) );
  XNOR2_X1 U3145 ( .A(n2457), .B(IR_REG_4__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U3146 ( .A1(n2460), .A2(IR_REG_31__SCAN_IN), .ZN(n2461) );
  MUX2_X1 U3147 ( .A(IR_REG_31__SCAN_IN), .B(n2461), .S(IR_REG_5__SCAN_IN), 
        .Z(n2464) );
  INV_X1 U31480 ( .A(n2462), .ZN(n2463) );
  MUX2_X1 U31490 ( .A(n4479), .B(DATAI_5_), .S(n2521), .Z(n3411) );
  NOR2_X1 U3150 ( .A1(n2462), .A2(n2553), .ZN(n2465) );
  MUX2_X1 U3151 ( .A(n2553), .B(n2465), .S(IR_REG_6__SCAN_IN), .Z(n2467) );
  OR2_X1 U3152 ( .A1(n2467), .A2(n2466), .ZN(n4623) );
  MUX2_X1 U3153 ( .A(n4489), .B(DATAI_6_), .S(n3144), .Z(n3331) );
  OR2_X1 U3154 ( .A1(n2466), .A2(n2553), .ZN(n2470) );
  INV_X1 U3155 ( .A(n2470), .ZN(n2468) );
  NAND2_X1 U3156 ( .A1(n2468), .A2(IR_REG_7__SCAN_IN), .ZN(n2471) );
  INV_X1 U3157 ( .A(IR_REG_7__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3158 ( .A1(n2470), .A2(n2469), .ZN(n2473) );
  NAND2_X1 U3159 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2474) );
  XNOR2_X1 U3160 ( .A(n2474), .B(IR_REG_8__SCAN_IN), .ZN(n4621) );
  MUX2_X1 U3161 ( .A(n4621), .B(DATAI_8_), .S(n3144), .Z(n3366) );
  NOR2_X1 U3162 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2475)
         );
  NAND2_X1 U3163 ( .A1(n2466), .A2(n2475), .ZN(n2477) );
  NAND2_X1 U3164 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  MUX2_X1 U3165 ( .A(IR_REG_31__SCAN_IN), .B(n2476), .S(IR_REG_9__SCAN_IN), 
        .Z(n2478) );
  MUX2_X1 U3166 ( .A(n3501), .B(DATAI_9_), .S(n3144), .Z(n3432) );
  NAND2_X1 U3167 ( .A1(n2480), .A2(IR_REG_31__SCAN_IN), .ZN(n2479) );
  XNOR2_X1 U3168 ( .A(n2479), .B(IR_REG_10__SCAN_IN), .ZN(n4617) );
  MUX2_X1 U3169 ( .A(n4617), .B(DATAI_10_), .S(n2521), .Z(n3073) );
  OAI21_X1 U3170 ( .B1(n2480), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2482) );
  OR2_X1 U3171 ( .A1(n2482), .A2(n2481), .ZN(n2483) );
  NAND2_X1 U3172 ( .A1(n2482), .A2(n2481), .ZN(n2484) );
  MUX2_X1 U3173 ( .A(n4394), .B(DATAI_11_), .S(n2521), .Z(n3517) );
  NAND2_X1 U3174 ( .A1(n2484), .A2(IR_REG_31__SCAN_IN), .ZN(n2485) );
  XNOR2_X1 U3175 ( .A(n2485), .B(IR_REG_12__SCAN_IN), .ZN(n4393) );
  MUX2_X1 U3176 ( .A(n4393), .B(DATAI_12_), .S(n3144), .Z(n3567) );
  NAND2_X1 U3177 ( .A1(n2486), .A2(IR_REG_31__SCAN_IN), .ZN(n2487) );
  MUX2_X1 U3178 ( .A(IR_REG_31__SCAN_IN), .B(n2487), .S(IR_REG_13__SCAN_IN), 
        .Z(n2488) );
  AND2_X1 U3179 ( .A1(n2488), .A2(n2490), .ZN(n4615) );
  INV_X1 U3180 ( .A(DATAI_13_), .ZN(n2489) );
  MUX2_X1 U3181 ( .A(n4534), .B(n2489), .S(n3144), .Z(n3076) );
  NAND2_X1 U3182 ( .A1(n2490), .A2(IR_REG_31__SCAN_IN), .ZN(n2491) );
  MUX2_X1 U3183 ( .A(n2491), .B(IR_REG_31__SCAN_IN), .S(n2507), .Z(n2493) );
  INV_X1 U3184 ( .A(n2494), .ZN(n2492) );
  MUX2_X1 U3185 ( .A(n4543), .B(DATAI_14_), .S(n2521), .Z(n3628) );
  OR2_X1 U3186 ( .A1(n2501), .A2(n2506), .ZN(n2495) );
  NAND2_X1 U3187 ( .A1(n2501), .A2(n2506), .ZN(n2496) );
  MUX2_X1 U3188 ( .A(n4613), .B(DATAI_15_), .S(n3144), .Z(n3077) );
  NAND2_X1 U3189 ( .A1(n2496), .A2(IR_REG_31__SCAN_IN), .ZN(n2497) );
  XNOR2_X1 U3190 ( .A(n2497), .B(n2505), .ZN(n4612) );
  INV_X1 U3191 ( .A(n4612), .ZN(n2498) );
  MUX2_X1 U3192 ( .A(n2498), .B(DATAI_16_), .S(n2521), .Z(n3672) );
  OR2_X1 U3193 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2499)
         );
  NAND2_X1 U3194 ( .A1(IR_REG_31__SCAN_IN), .A2(n2499), .ZN(n2500) );
  NAND2_X1 U3195 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  XNOR2_X1 U3196 ( .A(n2502), .B(n2504), .ZN(n4609) );
  INV_X1 U3197 ( .A(DATAI_17_), .ZN(n2503) );
  MUX2_X1 U3198 ( .A(n4034), .B(n2503), .S(n3144), .Z(n3082) );
  AND3_X1 U3199 ( .A1(n2506), .A2(n2505), .A3(n2504), .ZN(n2508) );
  AND2_X1 U3200 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  INV_X1 U3201 ( .A(n2516), .ZN(n2511) );
  NAND2_X1 U3202 ( .A1(n2511), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  XNOR2_X1 U3203 ( .A(n2512), .B(IR_REG_18__SCAN_IN), .ZN(n4052) );
  INV_X1 U3204 ( .A(DATAI_18_), .ZN(n2513) );
  MUX2_X1 U3205 ( .A(n4608), .B(n2513), .S(n3144), .Z(n4420) );
  AND2_X1 U3206 ( .A1(n2515), .A2(n2518), .ZN(n2514) );
  NAND2_X1 U3207 ( .A1(n2516), .A2(n2515), .ZN(n2517) );
  NAND2_X1 U3208 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2519) );
  INV_X1 U3209 ( .A(DATAI_19_), .ZN(n5039) );
  MUX2_X1 U32100 ( .A(n4058), .B(n5039), .S(n3144), .Z(n4264) );
  NAND2_X1 U32110 ( .A1(n2521), .A2(DATAI_20_), .ZN(n4226) );
  NAND2_X1 U32120 ( .A1(n2521), .A2(DATAI_26_), .ZN(n4126) );
  NAND2_X1 U32130 ( .A1(n2521), .A2(DATAI_27_), .ZN(n4106) );
  NAND2_X1 U32140 ( .A1(n3144), .A2(DATAI_28_), .ZN(n3118) );
  AND2_X1 U32150 ( .A1(n3144), .A2(DATAI_29_), .ZN(n4068) );
  INV_X1 U32160 ( .A(n4068), .ZN(n4082) );
  NAND2_X1 U32170 ( .A1(n3144), .A2(DATAI_30_), .ZN(n3820) );
  INV_X1 U32180 ( .A(n3820), .ZN(n4288) );
  INV_X1 U32190 ( .A(n2526), .ZN(n2560) );
  NAND2_X1 U32200 ( .A1(n2526), .A2(n2523), .ZN(n2535) );
  INV_X1 U32210 ( .A(IR_REG_23__SCAN_IN), .ZN(n2556) );
  AND2_X1 U32220 ( .A1(n2552), .A2(n2556), .ZN(n2525) );
  AND2_X1 U32230 ( .A1(n2526), .A2(n2525), .ZN(n2527) );
  NAND2_X1 U32240 ( .A1(n2569), .A2(n2257), .ZN(n2530) );
  NOR2_X1 U32250 ( .A1(n2571), .A2(n2530), .ZN(n2531) );
  NOR2_X1 U32260 ( .A1(n2531), .A2(n2553), .ZN(n2533) );
  NAND2_X1 U32270 ( .A1(n2535), .A2(n2534), .ZN(n2550) );
  NAND2_X1 U32280 ( .A1(n2550), .A2(n2529), .ZN(n2536) );
  MUX2_X1 U32290 ( .A(n2529), .B(n2536), .S(B_REG_SCAN_IN), .Z(n2537) );
  NOR2_X1 U32300 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_7__SCAN_IN), .ZN(n2541)
         );
  NOR4_X1 U32310 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2540) );
  NOR4_X1 U32320 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2539) );
  NOR4_X1 U32330 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2538) );
  AND4_X1 U32340 ( .A1(n2541), .A2(n2540), .A3(n2539), .A4(n2538), .ZN(n2547)
         );
  NOR4_X1 U32350 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2545) );
  NOR4_X1 U32360 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2544) );
  NOR4_X1 U32370 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2543) );
  NOR4_X1 U32380 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2542) );
  AND4_X1 U32390 ( .A1(n2545), .A2(n2544), .A3(n2543), .A4(n2542), .ZN(n2546)
         );
  NAND2_X1 U32400 ( .A1(n2547), .A2(n2546), .ZN(n3107) );
  INV_X1 U32410 ( .A(n3107), .ZN(n2548) );
  NAND2_X1 U32420 ( .A1(n2548), .A2(D_REG_1__SCAN_IN), .ZN(n2549) );
  INV_X1 U32430 ( .A(n2551), .ZN(n2563) );
  NAND2_X1 U32440 ( .A1(n2550), .A2(n2563), .ZN(n3109) );
  INV_X1 U32450 ( .A(n3109), .ZN(n3138) );
  AOI21_X1 U32460 ( .B1(n3108), .B2(n2549), .A(n3138), .ZN(n2989) );
  INV_X1 U32470 ( .A(n2550), .ZN(n4387) );
  INV_X1 U32480 ( .A(n2597), .ZN(n2613) );
  AND2_X1 U32490 ( .A1(n2526), .A2(n2552), .ZN(n2554) );
  NAND2_X1 U32500 ( .A1(n2557), .A2(n2556), .ZN(n2555) );
  NAND2_X1 U32510 ( .A1(n3142), .A2(STATE_REG_SCAN_IN), .ZN(n4606) );
  NAND2_X1 U32520 ( .A1(n2595), .A2(n4058), .ZN(n2990) );
  NAND2_X1 U32530 ( .A1(n2560), .A2(IR_REG_31__SCAN_IN), .ZN(n2561) );
  XNOR2_X1 U32540 ( .A(n2561), .B(n2552), .ZN(n2567) );
  AND2_X1 U32550 ( .A1(n2571), .A2(IR_REG_31__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32560 ( .A1(n2990), .A2(n3141), .ZN(n3110) );
  NAND3_X1 U32570 ( .A1(n2989), .A2(n3198), .A3(n3110), .ZN(n2564) );
  INV_X1 U32580 ( .A(D_REG_0__SCAN_IN), .ZN(n3136) );
  NOR2_X1 U32590 ( .A1(n4058), .A2(n4389), .ZN(n2565) );
  NAND2_X1 U32600 ( .A1(n2595), .A2(n2565), .ZN(n4668) );
  OR2_X1 U32610 ( .A1(n4668), .A2(n4390), .ZN(n3111) );
  AND2_X1 U32620 ( .A1(n4273), .A2(n4058), .ZN(n3286) );
  NAND2_X1 U32630 ( .A1(n4278), .A2(n4598), .ZN(n2590) );
  INV_X1 U32640 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4944) );
  OR2_X1 U32650 ( .A1(n4273), .A2(n4944), .ZN(n2588) );
  INV_X1 U32660 ( .A(n2595), .ZN(n4391) );
  OAI21_X1 U32670 ( .B1(n2574), .B2(n2553), .A(IR_REG_29__SCAN_IN), .ZN(n2576)
         );
  AND2_X2 U32680 ( .A1(n2579), .A2(n3131), .ZN(n2692) );
  NAND2_X1 U32690 ( .A1(n2692), .A2(REG1_REG_31__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U32700 ( .A1(n3206), .A2(REG2_REG_31__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U32710 ( .A1(n3207), .A2(REG0_REG_31__SCAN_IN), .ZN(n2580) );
  NAND3_X1 U32720 ( .A1(n2582), .A2(n2581), .A3(n2580), .ZN(n3839) );
  XNOR2_X1 U32730 ( .A(n2583), .B(IR_REG_27__SCAN_IN), .ZN(n4452) );
  OR2_X1 U32740 ( .A1(n2584), .A2(n2553), .ZN(n2586) );
  XNOR2_X1 U32750 ( .A(n2586), .B(n2585), .ZN(n3013) );
  NAND2_X1 U32760 ( .A1(n3013), .A2(n3141), .ZN(n4256) );
  AOI21_X1 U32770 ( .B1(n4452), .B2(B_REG_SCAN_IN), .A(n4256), .ZN(n4069) );
  NAND2_X1 U32780 ( .A1(n3839), .A2(n4069), .ZN(n4285) );
  OAI21_X1 U32790 ( .B1(n3965), .B2(n4255), .A(n4285), .ZN(n4279) );
  NAND2_X1 U32800 ( .A1(n4273), .A2(n4279), .ZN(n2587) );
  AND2_X1 U32810 ( .A1(n2588), .A2(n2587), .ZN(n2589) );
  NAND2_X1 U32820 ( .A1(n2590), .A2(n2589), .ZN(U3260) );
  NAND2_X1 U32830 ( .A1(n2603), .A2(REG2_REG_1__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U32840 ( .A1(n2651), .A2(REG0_REG_1__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U32850 ( .A1(n2692), .A2(REG1_REG_1__SCAN_IN), .ZN(n2591) );
  INV_X1 U32860 ( .A(n3025), .ZN(n3451) );
  INV_X1 U32870 ( .A(n3269), .ZN(n2596) );
  NAND2_X1 U32880 ( .A1(n4058), .A2(n4389), .ZN(n3005) );
  OR2_X2 U32890 ( .A1(n2627), .A2(n2598), .ZN(n2629) );
  NAND2_X1 U32900 ( .A1(n2231), .A2(n2600), .ZN(n2601) );
  XNOR2_X1 U32910 ( .A(n2621), .B(n2620), .ZN(n3748) );
  INV_X1 U32920 ( .A(n3748), .ZN(n2619) );
  NAND2_X1 U32930 ( .A1(n2650), .A2(REG3_REG_0__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U32940 ( .A1(n2692), .A2(REG1_REG_0__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U32950 ( .A1(n2603), .A2(REG2_REG_0__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U32960 ( .A1(n2651), .A2(REG0_REG_0__SCAN_IN), .ZN(n2604) );
  NAND4_X1 U32970 ( .A1(n2607), .A2(n2606), .A3(n2605), .A4(n2604), .ZN(n2608)
         );
  INV_X1 U32980 ( .A(n2608), .ZN(n3064) );
  OAI21_X1 U32990 ( .B1(n3064), .B2(n2972), .A(n2422), .ZN(n2610) );
  INV_X1 U33000 ( .A(n2610), .ZN(n2617) );
  INV_X1 U33010 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2611) );
  OR2_X1 U33020 ( .A1(n2597), .A2(n2611), .ZN(n2612) );
  NAND2_X1 U33030 ( .A1(n2617), .A2(n2612), .ZN(n3195) );
  NAND2_X1 U33040 ( .A1(n2608), .A2(n2658), .ZN(n2616) );
  AOI21_X1 U33050 ( .B1(n2600), .B2(n4628), .A(n2614), .ZN(n2615) );
  NAND2_X1 U33060 ( .A1(n2616), .A2(n2615), .ZN(n3194) );
  AOI22_X1 U33070 ( .A1(n3195), .A2(n3194), .B1(n2617), .B2(n2984), .ZN(n3749)
         );
  INV_X1 U33080 ( .A(n3749), .ZN(n2618) );
  NAND2_X1 U33090 ( .A1(n2619), .A2(n2618), .ZN(n3750) );
  NAND2_X1 U33100 ( .A1(n2621), .A2(n2620), .ZN(n2622) );
  NAND2_X1 U33110 ( .A1(n2977), .A2(REG3_REG_2__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U33120 ( .A1(n2234), .A2(REG1_REG_2__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U33130 ( .A1(n2603), .A2(REG2_REG_2__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U33140 ( .A1(n2651), .A2(REG0_REG_2__SCAN_IN), .ZN(n2623) );
  INV_X1 U33150 ( .A(n3448), .ZN(n3457) );
  XNOR2_X1 U33160 ( .A(n2628), .B(n2973), .ZN(n2632) );
  OR2_X1 U33170 ( .A1(n3386), .A2(n2629), .ZN(n2631) );
  NAND2_X1 U33180 ( .A1(n3448), .A2(n2600), .ZN(n2630) );
  NAND2_X1 U33190 ( .A1(n2631), .A2(n2630), .ZN(n2633) );
  INV_X1 U33200 ( .A(n2632), .ZN(n2635) );
  INV_X1 U33210 ( .A(n2633), .ZN(n2634) );
  NAND2_X1 U33220 ( .A1(n2635), .A2(n2634), .ZN(n2636) );
  INV_X1 U33230 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U33240 ( .A1(n2977), .A2(n2637), .ZN(n2641) );
  NAND2_X1 U33250 ( .A1(n2234), .A2(REG1_REG_3__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U33260 ( .A1(n2603), .A2(REG2_REG_3__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U33270 ( .A1(n2651), .A2(REG0_REG_3__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U33280 ( .A1(n3449), .A2(n2600), .ZN(n2643) );
  NAND2_X1 U33290 ( .A1(n3387), .A2(n2986), .ZN(n2642) );
  NAND2_X1 U33300 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  XNOR2_X1 U33310 ( .A(n2644), .B(n2973), .ZN(n2645) );
  AOI22_X1 U33320 ( .A1(n3449), .A2(n2658), .B1(n3387), .B2(n2600), .ZN(n2646)
         );
  XNOR2_X1 U33330 ( .A(n2645), .B(n2646), .ZN(n3229) );
  INV_X1 U33340 ( .A(n2645), .ZN(n2647) );
  AND2_X1 U33350 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  NAND2_X1 U33360 ( .A1(n2603), .A2(REG2_REG_4__SCAN_IN), .ZN(n2656) );
  INV_X1 U33370 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2649) );
  XNOR2_X1 U33380 ( .A(n2649), .B(REG3_REG_3__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U33390 ( .A1(n2650), .A2(n3236), .ZN(n2654) );
  NAND2_X1 U33400 ( .A1(n2692), .A2(REG1_REG_4__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U33410 ( .A1(n2651), .A2(REG0_REG_4__SCAN_IN), .ZN(n2652) );
  INV_X1 U33420 ( .A(n3261), .ZN(n3030) );
  OAI22_X1 U33430 ( .A1(n3031), .A2(n2971), .B1(n3030), .B2(n2627), .ZN(n2657)
         );
  XNOR2_X1 U33440 ( .A(n2657), .B(n2984), .ZN(n2661) );
  OR2_X1 U33450 ( .A1(n3031), .A2(n2629), .ZN(n2660) );
  NAND2_X1 U33460 ( .A1(n3261), .A2(n2600), .ZN(n2659) );
  NAND2_X1 U33470 ( .A1(n2660), .A2(n2659), .ZN(n2662) );
  XNOR2_X1 U33480 ( .A(n2661), .B(n2662), .ZN(n3238) );
  NAND2_X1 U33490 ( .A1(n3239), .A2(n3238), .ZN(n3237) );
  INV_X1 U33500 ( .A(n2661), .ZN(n2663) );
  NAND2_X1 U33510 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  NAND2_X1 U33520 ( .A1(n3237), .A2(n2664), .ZN(n3247) );
  NAND2_X1 U3353 ( .A1(n2651), .A2(REG0_REG_5__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U33540 ( .A1(n2235), .A2(REG1_REG_5__SCAN_IN), .ZN(n2668) );
  AOI21_X1 U3355 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2665) );
  NOR2_X1 U3356 ( .A1(n2665), .A2(n2678), .ZN(n3244) );
  NAND2_X1 U3357 ( .A1(n2977), .A2(n3244), .ZN(n2667) );
  NAND2_X1 U3358 ( .A1(n2603), .A2(REG2_REG_5__SCAN_IN), .ZN(n2666) );
  NAND4_X1 U3359 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .ZN(n3990)
         );
  NAND2_X1 U3360 ( .A1(n3990), .A2(n2600), .ZN(n2671) );
  NAND2_X1 U3361 ( .A1(n3411), .A2(n2986), .ZN(n2670) );
  NAND2_X1 U3362 ( .A1(n2671), .A2(n2670), .ZN(n2672) );
  XNOR2_X1 U3363 ( .A(n2672), .B(n2973), .ZN(n2675) );
  AOI22_X1 U3364 ( .A1(n3990), .A2(n2658), .B1(n3411), .B2(n2600), .ZN(n2673)
         );
  XNOR2_X1 U3365 ( .A(n2675), .B(n2673), .ZN(n3246) );
  NAND2_X1 U3366 ( .A1(n3247), .A2(n3246), .ZN(n3245) );
  INV_X1 U3367 ( .A(n2673), .ZN(n2674) );
  NAND2_X1 U3368 ( .A1(n2675), .A2(n2674), .ZN(n2676) );
  INV_X1 U3369 ( .A(n2678), .ZN(n2677) );
  INV_X1 U3370 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4868) );
  NAND2_X1 U3371 ( .A1(n2677), .A2(n4868), .ZN(n2679) );
  AND2_X1 U3372 ( .A1(n2679), .A2(n2690), .ZN(n4595) );
  NAND2_X1 U3373 ( .A1(n2977), .A2(n4595), .ZN(n2683) );
  NAND2_X1 U3374 ( .A1(n2235), .A2(REG1_REG_6__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3375 ( .A1(n2603), .A2(REG2_REG_6__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3376 ( .A1(n2651), .A2(REG0_REG_6__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3377 ( .A1(n3989), .A2(n2658), .ZN(n2685) );
  NAND2_X1 U3378 ( .A1(n3331), .A2(n2600), .ZN(n2684) );
  NAND2_X1 U3379 ( .A1(n2685), .A2(n2684), .ZN(n3292) );
  NAND2_X1 U3380 ( .A1(n3989), .A2(n2600), .ZN(n2687) );
  NAND2_X1 U3381 ( .A1(n3331), .A2(n2986), .ZN(n2686) );
  NAND2_X1 U3382 ( .A1(n2687), .A2(n2686), .ZN(n2688) );
  XNOR2_X1 U3383 ( .A(n2688), .B(n2973), .ZN(n3291) );
  AND2_X1 U3384 ( .A1(n2690), .A2(n2689), .ZN(n2691) );
  NOR2_X1 U3385 ( .A1(n2710), .A2(n2691), .ZN(n3323) );
  NAND2_X1 U3386 ( .A1(n2977), .A2(n3323), .ZN(n2695) );
  NAND2_X1 U3387 ( .A1(n2692), .A2(REG1_REG_7__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3388 ( .A1(n2651), .A2(REG0_REG_7__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3389 ( .A1(n2603), .A2(REG2_REG_7__SCAN_IN), .ZN(n2696) );
  OAI22_X1 U3390 ( .A1(n3349), .A2(n2972), .B1(n3285), .B2(n2627), .ZN(n2698)
         );
  XNOR2_X1 U3391 ( .A(n2698), .B(n2984), .ZN(n2727) );
  OR2_X1 U3392 ( .A1(n3349), .A2(n2629), .ZN(n2700) );
  NAND2_X1 U3393 ( .A1(n3322), .A2(n2600), .ZN(n2699) );
  NAND2_X1 U3394 ( .A1(n2700), .A2(n2699), .ZN(n2728) );
  XNOR2_X1 U3395 ( .A(n2727), .B(n2728), .ZN(n3343) );
  NAND2_X1 U3396 ( .A1(n2235), .A2(REG1_REG_9__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U3397 ( .A1(n2651), .A2(REG0_REG_9__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U3398 ( .A1(n2710), .A2(REG3_REG_8__SCAN_IN), .ZN(n2712) );
  NAND2_X1 U3399 ( .A1(n2712), .A2(n2701), .ZN(n2702) );
  AND2_X1 U3400 ( .A1(n2743), .A2(n2702), .ZN(n3433) );
  NAND2_X1 U3401 ( .A1(n2977), .A2(n3433), .ZN(n2704) );
  NAND2_X1 U3402 ( .A1(n3206), .A2(REG2_REG_9__SCAN_IN), .ZN(n2703) );
  NAND4_X1 U3403 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), .ZN(n3987)
         );
  NAND2_X1 U3404 ( .A1(n3987), .A2(n2600), .ZN(n2708) );
  NAND2_X1 U3405 ( .A1(n3432), .A2(n2986), .ZN(n2707) );
  NAND2_X1 U3406 ( .A1(n2708), .A2(n2707), .ZN(n2709) );
  XNOR2_X1 U3407 ( .A(n2709), .B(n2973), .ZN(n2737) );
  AOI22_X1 U3408 ( .A1(n3987), .A2(n2658), .B1(n3432), .B2(n2600), .ZN(n2738)
         );
  XNOR2_X1 U3409 ( .A(n2737), .B(n2738), .ZN(n3429) );
  INV_X1 U3410 ( .A(n3429), .ZN(n2724) );
  NAND2_X1 U3411 ( .A1(n2651), .A2(REG0_REG_8__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3412 ( .A1(n2235), .A2(REG1_REG_8__SCAN_IN), .ZN(n2715) );
  OR2_X1 U3413 ( .A1(n2710), .A2(REG3_REG_8__SCAN_IN), .ZN(n2711) );
  AND2_X1 U3414 ( .A1(n2712), .A2(n2711), .ZN(n3401) );
  NAND2_X1 U3415 ( .A1(n2977), .A2(n3401), .ZN(n2714) );
  NAND2_X1 U3416 ( .A1(n2603), .A2(REG2_REG_8__SCAN_IN), .ZN(n2713) );
  NAND4_X1 U3417 ( .A1(n2716), .A2(n2715), .A3(n2714), .A4(n2713), .ZN(n3274)
         );
  NAND2_X1 U3418 ( .A1(n3274), .A2(n2600), .ZN(n2718) );
  NAND2_X1 U3419 ( .A1(n3366), .A2(n2986), .ZN(n2717) );
  NAND2_X1 U3420 ( .A1(n2718), .A2(n2717), .ZN(n2719) );
  XNOR2_X1 U3421 ( .A(n2719), .B(n2973), .ZN(n2731) );
  INV_X1 U3422 ( .A(n2731), .ZN(n2723) );
  NAND2_X1 U3423 ( .A1(n3274), .A2(n2658), .ZN(n2721) );
  NAND2_X1 U3424 ( .A1(n3366), .A2(n2600), .ZN(n2720) );
  NAND2_X1 U3425 ( .A1(n2721), .A2(n2720), .ZN(n2730) );
  INV_X1 U3426 ( .A(n2730), .ZN(n2722) );
  NAND2_X1 U3427 ( .A1(n2723), .A2(n2722), .ZN(n3426) );
  AND2_X1 U3428 ( .A1(n3343), .A2(n2726), .ZN(n2725) );
  INV_X1 U3429 ( .A(n2726), .ZN(n2734) );
  INV_X1 U3430 ( .A(n2727), .ZN(n2729) );
  NAND2_X1 U3431 ( .A1(n2729), .A2(n2728), .ZN(n3344) );
  AND2_X1 U3432 ( .A1(n2731), .A2(n2730), .ZN(n3345) );
  INV_X1 U3433 ( .A(n3345), .ZN(n2732) );
  AND2_X1 U3434 ( .A1(n3344), .A2(n2732), .ZN(n3424) );
  AND2_X1 U3435 ( .A1(n3424), .A2(n3429), .ZN(n2733) );
  NAND2_X1 U3436 ( .A1(n2736), .A2(n2735), .ZN(n2741) );
  INV_X1 U3437 ( .A(n2737), .ZN(n2739) );
  NAND2_X1 U3438 ( .A1(n2739), .A2(n2738), .ZN(n2740) );
  NAND2_X1 U3439 ( .A1(n3207), .A2(REG0_REG_10__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U3440 ( .A1(n2235), .A2(REG1_REG_10__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U3441 ( .A1(n2743), .A2(n4892), .ZN(n2744) );
  AND2_X1 U3442 ( .A1(n2758), .A2(n2744), .ZN(n3484) );
  NAND2_X1 U3443 ( .A1(n2977), .A2(n3484), .ZN(n2746) );
  NAND2_X1 U3444 ( .A1(n3206), .A2(REG2_REG_10__SCAN_IN), .ZN(n2745) );
  NAND4_X1 U3445 ( .A1(n2748), .A2(n2747), .A3(n2746), .A4(n2745), .ZN(n3359)
         );
  NAND2_X1 U3446 ( .A1(n3359), .A2(n2600), .ZN(n2750) );
  NAND2_X1 U3447 ( .A1(n3073), .A2(n2986), .ZN(n2749) );
  NAND2_X1 U3448 ( .A1(n2750), .A2(n2749), .ZN(n2751) );
  XNOR2_X1 U3449 ( .A(n2751), .B(n2984), .ZN(n2753) );
  AOI22_X1 U3450 ( .A1(n3359), .A2(n2658), .B1(n3073), .B2(n2600), .ZN(n2754)
         );
  XNOR2_X1 U3451 ( .A(n2753), .B(n2754), .ZN(n3481) );
  INV_X1 U3452 ( .A(n2753), .ZN(n2756) );
  INV_X1 U3453 ( .A(n2754), .ZN(n2755) );
  NAND2_X1 U3454 ( .A1(n2756), .A2(n2755), .ZN(n2757) );
  NAND2_X1 U3455 ( .A1(n2651), .A2(REG0_REG_11__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U3456 ( .A1(n2235), .A2(REG1_REG_11__SCAN_IN), .ZN(n2762) );
  AND2_X1 U3457 ( .A1(n2758), .A2(n3439), .ZN(n2759) );
  NOR2_X1 U34580 ( .A1(n2767), .A2(n2759), .ZN(n3525) );
  NAND2_X1 U34590 ( .A1(n2977), .A2(n3525), .ZN(n2761) );
  NAND2_X1 U3460 ( .A1(n3206), .A2(REG2_REG_11__SCAN_IN), .ZN(n2760) );
  OAI22_X1 U3461 ( .A1(n3464), .A2(n2972), .B1(n3523), .B2(n2627), .ZN(n2764)
         );
  XNOR2_X1 U3462 ( .A(n2764), .B(n2984), .ZN(n3545) );
  OR2_X1 U3463 ( .A1(n3464), .A2(n2629), .ZN(n2766) );
  NAND2_X1 U3464 ( .A1(n3517), .A2(n2600), .ZN(n2765) );
  NAND2_X1 U3465 ( .A1(n3207), .A2(REG0_REG_12__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U3466 ( .A1(n2235), .A2(REG1_REG_12__SCAN_IN), .ZN(n2771) );
  NOR2_X1 U34670 ( .A1(n2767), .A2(REG3_REG_12__SCAN_IN), .ZN(n2768) );
  NOR2_X1 U3468 ( .A1(n2785), .A2(n2768), .ZN(n3570) );
  NAND2_X1 U34690 ( .A1(n2977), .A2(n3570), .ZN(n2770) );
  NAND2_X1 U3470 ( .A1(n3206), .A2(REG2_REG_12__SCAN_IN), .ZN(n2769) );
  NAND4_X1 U34710 ( .A1(n2772), .A2(n2771), .A3(n2770), .A4(n2769), .ZN(n3985)
         );
  NAND2_X1 U3472 ( .A1(n3985), .A2(n2600), .ZN(n2774) );
  NAND2_X1 U34730 ( .A1(n3567), .A2(n2986), .ZN(n2773) );
  NAND2_X1 U3474 ( .A1(n2774), .A2(n2773), .ZN(n2775) );
  XNOR2_X1 U34750 ( .A(n2775), .B(n2973), .ZN(n2778) );
  NAND2_X1 U3476 ( .A1(n3985), .A2(n2658), .ZN(n2777) );
  NAND2_X1 U34770 ( .A1(n3567), .A2(n2600), .ZN(n2776) );
  NAND2_X1 U3478 ( .A1(n2777), .A2(n2776), .ZN(n2779) );
  NAND2_X1 U34790 ( .A1(n2778), .A2(n2779), .ZN(n3541) );
  OAI21_X1 U3480 ( .B1(n3545), .B2(n3543), .A(n3541), .ZN(n2784) );
  NAND3_X1 U34810 ( .A1(n3545), .A2(n3543), .A3(n3541), .ZN(n2782) );
  INV_X1 U3482 ( .A(n2778), .ZN(n2781) );
  INV_X1 U34830 ( .A(n2779), .ZN(n2780) );
  NAND2_X1 U3484 ( .A1(n2781), .A2(n2780), .ZN(n3540) );
  AND2_X1 U34850 ( .A1(n2782), .A2(n3540), .ZN(n2783) );
  NAND2_X1 U3486 ( .A1(n3207), .A2(REG0_REG_13__SCAN_IN), .ZN(n2790) );
  NAND2_X1 U34870 ( .A1(n2235), .A2(REG1_REG_13__SCAN_IN), .ZN(n2789) );
  NOR2_X1 U3488 ( .A1(n2785), .A2(REG3_REG_13__SCAN_IN), .ZN(n2786) );
  NOR2_X1 U34890 ( .A1(n2794), .A2(n2786), .ZN(n3618) );
  NAND2_X1 U3490 ( .A1(n2977), .A2(n3618), .ZN(n2788) );
  NAND2_X1 U34910 ( .A1(n3206), .A2(REG2_REG_13__SCAN_IN), .ZN(n2787) );
  OAI22_X1 U3492 ( .A1(n3631), .A2(n2972), .B1(n3076), .B2(n2627), .ZN(n2791)
         );
  XNOR2_X1 U34930 ( .A(n2791), .B(n2984), .ZN(n3531) );
  OR2_X1 U3494 ( .A1(n3631), .A2(n2629), .ZN(n2793) );
  NAND2_X1 U34950 ( .A1(n3615), .A2(n2600), .ZN(n2792) );
  NAND2_X1 U3496 ( .A1(n2793), .A2(n2792), .ZN(n3532) );
  NAND2_X1 U34970 ( .A1(n3207), .A2(REG0_REG_14__SCAN_IN), .ZN(n2799) );
  NAND2_X1 U3498 ( .A1(n2235), .A2(REG1_REG_14__SCAN_IN), .ZN(n2798) );
  OR2_X1 U34990 ( .A1(n2794), .A2(REG3_REG_14__SCAN_IN), .ZN(n2795) );
  AND2_X1 U3500 ( .A1(n2795), .A2(n2807), .ZN(n3635) );
  NAND2_X1 U35010 ( .A1(n2977), .A2(n3635), .ZN(n2797) );
  NAND2_X1 U3502 ( .A1(n3206), .A2(REG2_REG_14__SCAN_IN), .ZN(n2796) );
  OAI22_X1 U35030 ( .A1(n4431), .A2(n2972), .B1(n3637), .B2(n2627), .ZN(n2800)
         );
  XNOR2_X1 U3504 ( .A(n2800), .B(n2973), .ZN(n2803) );
  OR2_X1 U35050 ( .A1(n4431), .A2(n2629), .ZN(n2802) );
  NAND2_X1 U35060 ( .A1(n3628), .A2(n2600), .ZN(n2801) );
  NAND2_X1 U35070 ( .A1(n2802), .A2(n2801), .ZN(n2804) );
  INV_X1 U35080 ( .A(n2803), .ZN(n2806) );
  INV_X1 U35090 ( .A(n2804), .ZN(n2805) );
  OAI21_X1 U35100 ( .B1(REG3_REG_15__SCAN_IN), .B2(n2808), .A(n2817), .ZN(
        n4445) );
  INV_X1 U35110 ( .A(n4445), .ZN(n2809) );
  NAND2_X1 U35120 ( .A1(n2977), .A2(n2809), .ZN(n2813) );
  NAND2_X1 U35130 ( .A1(n2235), .A2(REG1_REG_15__SCAN_IN), .ZN(n2812) );
  NAND2_X1 U35140 ( .A1(n2603), .A2(REG2_REG_15__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U35150 ( .A1(n3207), .A2(REG0_REG_15__SCAN_IN), .ZN(n2810) );
  NAND4_X1 U35160 ( .A1(n2813), .A2(n2812), .A3(n2811), .A4(n2810), .ZN(n3982)
         );
  NAND2_X1 U35170 ( .A1(n3982), .A2(n2600), .ZN(n2815) );
  NAND2_X1 U35180 ( .A1(n3077), .A2(n2986), .ZN(n2814) );
  NAND2_X1 U35190 ( .A1(n2815), .A2(n2814), .ZN(n2816) );
  XNOR2_X1 U35200 ( .A(n2816), .B(n2984), .ZN(n2830) );
  NOR2_X1 U35210 ( .A1(n2831), .A2(n2830), .ZN(n4403) );
  INV_X1 U35220 ( .A(n2817), .ZN(n2819) );
  INV_X1 U35230 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4398) );
  INV_X1 U35240 ( .A(n2838), .ZN(n2818) );
  OAI21_X1 U35250 ( .B1(REG3_REG_16__SCAN_IN), .B2(n2819), .A(n2818), .ZN(
        n4409) );
  INV_X1 U35260 ( .A(n4409), .ZN(n2820) );
  NAND2_X1 U35270 ( .A1(n2977), .A2(n2820), .ZN(n2824) );
  NAND2_X1 U35280 ( .A1(n2235), .A2(REG1_REG_16__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U35290 ( .A1(n2603), .A2(REG2_REG_16__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U35300 ( .A1(n3207), .A2(REG0_REG_16__SCAN_IN), .ZN(n2821) );
  INV_X1 U35310 ( .A(n3672), .ZN(n4400) );
  OAI22_X1 U35320 ( .A1(n4428), .A2(n2972), .B1(n4400), .B2(n2627), .ZN(n2825)
         );
  XNOR2_X1 U35330 ( .A(n2825), .B(n2984), .ZN(n2829) );
  OR2_X1 U35340 ( .A1(n4428), .A2(n2629), .ZN(n2827) );
  NAND2_X1 U35350 ( .A1(n3672), .A2(n2600), .ZN(n2826) );
  AND2_X1 U35360 ( .A1(n2827), .A2(n2826), .ZN(n2828) );
  NAND2_X1 U35370 ( .A1(n2829), .A2(n2828), .ZN(n2834) );
  OAI21_X1 U35380 ( .B1(n2829), .B2(n2828), .A(n2834), .ZN(n4405) );
  NOR2_X1 U35390 ( .A1(n4403), .A2(n4405), .ZN(n2837) );
  NAND2_X1 U35400 ( .A1(n2831), .A2(n2830), .ZN(n4436) );
  NAND2_X1 U35410 ( .A1(n3982), .A2(n2658), .ZN(n2833) );
  NAND2_X1 U35420 ( .A1(n3077), .A2(n2600), .ZN(n2832) );
  NAND2_X1 U35430 ( .A1(n2833), .A2(n2832), .ZN(n4437) );
  NAND2_X1 U35440 ( .A1(n4436), .A2(n4437), .ZN(n2836) );
  INV_X1 U35450 ( .A(n2834), .ZN(n2835) );
  AOI21_X1 U35460 ( .B1(n2837), .B2(n2836), .A(n2835), .ZN(n3710) );
  NOR2_X1 U35470 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2838), .ZN(n2839) );
  NOR2_X1 U35480 ( .A1(n2850), .A2(n2839), .ZN(n3718) );
  NAND2_X1 U35490 ( .A1(n2977), .A2(n3718), .ZN(n2843) );
  NAND2_X1 U35500 ( .A1(n2235), .A2(REG1_REG_17__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U35510 ( .A1(n2603), .A2(REG2_REG_17__SCAN_IN), .ZN(n2841) );
  NAND2_X1 U35520 ( .A1(n3207), .A2(REG0_REG_17__SCAN_IN), .ZN(n2840) );
  NAND4_X1 U35530 ( .A1(n2843), .A2(n2842), .A3(n2841), .A4(n2840), .ZN(n3981)
         );
  NAND2_X1 U35540 ( .A1(n3981), .A2(n2600), .ZN(n2845) );
  NAND2_X1 U35550 ( .A1(n3717), .A2(n2986), .ZN(n2844) );
  NAND2_X1 U35560 ( .A1(n2845), .A2(n2844), .ZN(n2846) );
  XNOR2_X1 U35570 ( .A(n2846), .B(n2984), .ZN(n2849) );
  NOR2_X1 U35580 ( .A1(n3082), .A2(n2971), .ZN(n2847) );
  AOI21_X1 U35590 ( .B1(n3981), .B2(n2658), .A(n2847), .ZN(n2848) );
  NOR2_X1 U35600 ( .A1(n2849), .A2(n2848), .ZN(n3713) );
  NAND2_X1 U35610 ( .A1(n2849), .A2(n2848), .ZN(n3711) );
  OAI21_X1 U35620 ( .B1(n3710), .B2(n3713), .A(n3711), .ZN(n4414) );
  NAND2_X1 U35630 ( .A1(n3207), .A2(REG0_REG_18__SCAN_IN), .ZN(n2857) );
  NAND2_X1 U35640 ( .A1(n2235), .A2(REG1_REG_18__SCAN_IN), .ZN(n2856) );
  INV_X1 U35650 ( .A(n2865), .ZN(n2853) );
  INV_X1 U35660 ( .A(n2850), .ZN(n2851) );
  INV_X1 U35670 ( .A(REG3_REG_18__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U35680 ( .A1(n2851), .A2(n5042), .ZN(n2852) );
  NAND2_X1 U35690 ( .A1(n2853), .A2(n2852), .ZN(n4427) );
  INV_X1 U35700 ( .A(n4427), .ZN(n3692) );
  NAND2_X1 U35710 ( .A1(n2977), .A2(n3692), .ZN(n2855) );
  NAND2_X1 U35720 ( .A1(n3206), .A2(REG2_REG_18__SCAN_IN), .ZN(n2854) );
  NAND4_X1 U35730 ( .A1(n2857), .A2(n2856), .A3(n2855), .A4(n2854), .ZN(n4259)
         );
  NAND2_X1 U35740 ( .A1(n4259), .A2(n2600), .ZN(n2859) );
  NAND2_X1 U35750 ( .A1(n2342), .A2(n2986), .ZN(n2858) );
  NAND2_X1 U35760 ( .A1(n2859), .A2(n2858), .ZN(n2860) );
  XNOR2_X1 U35770 ( .A(n2860), .B(n2984), .ZN(n4412) );
  NOR2_X1 U35780 ( .A1(n4420), .A2(n2972), .ZN(n2861) );
  AOI21_X1 U35790 ( .B1(n4259), .B2(n2658), .A(n2861), .ZN(n4413) );
  NAND2_X1 U35800 ( .A1(n4414), .A2(n2864), .ZN(n4415) );
  NAND2_X1 U35810 ( .A1(n4412), .A2(n4413), .ZN(n4417) );
  NAND2_X1 U3582 ( .A1(n2235), .A2(REG1_REG_19__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U3583 ( .A1(n3207), .A2(REG0_REG_19__SCAN_IN), .ZN(n2869) );
  NOR2_X1 U3584 ( .A1(n2865), .A2(REG3_REG_19__SCAN_IN), .ZN(n2866) );
  NOR2_X1 U3585 ( .A1(n2878), .A2(n2866), .ZN(n4267) );
  NAND2_X1 U3586 ( .A1(n2977), .A2(n4267), .ZN(n2868) );
  NAND2_X1 U3587 ( .A1(n3206), .A2(REG2_REG_19__SCAN_IN), .ZN(n2867) );
  NAND4_X1 U3588 ( .A1(n2870), .A2(n2869), .A3(n2868), .A4(n2867), .ZN(n4234)
         );
  NAND2_X1 U3589 ( .A1(n4234), .A2(n2600), .ZN(n2872) );
  INV_X1 U3590 ( .A(n4264), .ZN(n3860) );
  NAND2_X1 U3591 ( .A1(n3860), .A2(n2986), .ZN(n2871) );
  NAND2_X1 U3592 ( .A1(n2872), .A2(n2871), .ZN(n2873) );
  XNOR2_X1 U3593 ( .A(n2873), .B(n2973), .ZN(n2874) );
  OAI22_X1 U3594 ( .A1(n4410), .A2(n2629), .B1(n4264), .B2(n2972), .ZN(n2875)
         );
  XOR2_X1 U3595 ( .A(n2874), .B(n2875), .Z(n3723) );
  INV_X1 U3596 ( .A(n2874), .ZN(n2877) );
  INV_X1 U3597 ( .A(n2875), .ZN(n2876) );
  NAND2_X1 U3598 ( .A1(n3207), .A2(REG0_REG_20__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3599 ( .A1(n2235), .A2(REG1_REG_20__SCAN_IN), .ZN(n2881) );
  OAI21_X1 U3600 ( .B1(n2878), .B2(REG3_REG_20__SCAN_IN), .A(n2901), .ZN(n4242) );
  INV_X1 U3601 ( .A(n4242), .ZN(n3794) );
  NAND2_X1 U3602 ( .A1(n2977), .A2(n3794), .ZN(n2880) );
  NAND2_X1 U3603 ( .A1(n2603), .A2(REG2_REG_20__SCAN_IN), .ZN(n2879) );
  NAND4_X1 U3604 ( .A1(n2882), .A2(n2881), .A3(n2880), .A4(n2879), .ZN(n4222)
         );
  NAND2_X1 U3605 ( .A1(n4222), .A2(n2600), .ZN(n2884) );
  NAND2_X1 U3606 ( .A1(n4239), .A2(n2986), .ZN(n2883) );
  NAND2_X1 U3607 ( .A1(n2884), .A2(n2883), .ZN(n2885) );
  XNOR2_X1 U3608 ( .A(n2885), .B(n2984), .ZN(n2888) );
  NOR2_X1 U3609 ( .A1(n4226), .A2(n2971), .ZN(n2886) );
  AOI21_X1 U3610 ( .B1(n4222), .B2(n2658), .A(n2886), .ZN(n2887) );
  NOR2_X1 U3611 ( .A1(n2888), .A2(n2887), .ZN(n3789) );
  NAND2_X1 U3612 ( .A1(n3207), .A2(REG0_REG_21__SCAN_IN), .ZN(n2892) );
  NAND2_X1 U3613 ( .A1(n2235), .A2(REG1_REG_21__SCAN_IN), .ZN(n2891) );
  XNOR2_X1 U3614 ( .A(n2901), .B(REG3_REG_21__SCAN_IN), .ZN(n4211) );
  NAND2_X1 U3615 ( .A1(n2977), .A2(n4211), .ZN(n2890) );
  NAND2_X1 U3616 ( .A1(n2603), .A2(REG2_REG_21__SCAN_IN), .ZN(n2889) );
  OR2_X1 U3617 ( .A1(n4227), .A2(n2629), .ZN(n2894) );
  NAND2_X1 U3618 ( .A1(n4210), .A2(n2600), .ZN(n2893) );
  INV_X1 U3619 ( .A(n4210), .ZN(n4214) );
  OAI22_X1 U3620 ( .A1(n4227), .A2(n2972), .B1(n4214), .B2(n2627), .ZN(n2895)
         );
  XNOR2_X1 U3621 ( .A(n2895), .B(n2984), .ZN(n3762) );
  NAND2_X1 U3622 ( .A1(n2896), .A2(n3762), .ZN(n2898) );
  INV_X1 U3623 ( .A(n3762), .ZN(n2897) );
  AOI21_X1 U3624 ( .B1(n3760), .B2(n2898), .A(n2267), .ZN(n3798) );
  NAND2_X1 U3625 ( .A1(n3207), .A2(REG0_REG_22__SCAN_IN), .ZN(n2907) );
  NAND2_X1 U3626 ( .A1(n2235), .A2(REG1_REG_22__SCAN_IN), .ZN(n2906) );
  INV_X1 U3627 ( .A(n2901), .ZN(n2899) );
  AOI21_X1 U3628 ( .B1(n2899), .B2(REG3_REG_21__SCAN_IN), .A(
        REG3_REG_22__SCAN_IN), .ZN(n2902) );
  NAND2_X1 U3629 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2900) );
  OR2_X1 U3630 ( .A1(n2902), .A2(n2911), .ZN(n4199) );
  INV_X1 U3631 ( .A(n4199), .ZN(n2903) );
  NAND2_X1 U3632 ( .A1(n2977), .A2(n2903), .ZN(n2905) );
  NAND2_X1 U3633 ( .A1(n2603), .A2(REG2_REG_22__SCAN_IN), .ZN(n2904) );
  OR2_X1 U3634 ( .A1(n4215), .A2(n2629), .ZN(n2909) );
  NAND2_X1 U3635 ( .A1(n4192), .A2(n2600), .ZN(n2908) );
  NAND2_X1 U3636 ( .A1(n2909), .A2(n2908), .ZN(n2921) );
  OAI22_X1 U3637 ( .A1(n4215), .A2(n2972), .B1(n4202), .B2(n2627), .ZN(n2910)
         );
  XNOR2_X1 U3638 ( .A(n2910), .B(n2973), .ZN(n2920) );
  XOR2_X1 U3639 ( .A(n2921), .B(n2920), .Z(n3799) );
  NAND2_X1 U3640 ( .A1(n3207), .A2(REG0_REG_23__SCAN_IN), .ZN(n2916) );
  NAND2_X1 U3641 ( .A1(n2235), .A2(REG1_REG_23__SCAN_IN), .ZN(n2915) );
  OR2_X1 U3642 ( .A1(n2911), .A2(REG3_REG_23__SCAN_IN), .ZN(n2912) );
  AND2_X1 U3643 ( .A1(n2940), .A2(n2912), .ZN(n4180) );
  NAND2_X1 U3644 ( .A1(n2977), .A2(n4180), .ZN(n2914) );
  NAND2_X1 U3645 ( .A1(n3206), .A2(REG2_REG_23__SCAN_IN), .ZN(n2913) );
  OAI22_X1 U3646 ( .A1(n4191), .A2(n2972), .B1(n4179), .B2(n2627), .ZN(n2917)
         );
  XNOR2_X1 U3647 ( .A(n2917), .B(n2984), .ZN(n2926) );
  OR2_X1 U3648 ( .A1(n4191), .A2(n2629), .ZN(n2919) );
  NAND2_X1 U3649 ( .A1(n3094), .A2(n2600), .ZN(n2918) );
  NAND2_X1 U3650 ( .A1(n2919), .A2(n2918), .ZN(n2924) );
  XNOR2_X1 U3651 ( .A(n2926), .B(n2924), .ZN(n3741) );
  INV_X1 U3652 ( .A(n2920), .ZN(n2923) );
  INV_X1 U3653 ( .A(n2921), .ZN(n2922) );
  NAND2_X1 U3654 ( .A1(n2923), .A2(n2922), .ZN(n3742) );
  INV_X1 U3655 ( .A(n2924), .ZN(n2925) );
  NOR2_X1 U3656 ( .A1(n2926), .A2(n2925), .ZN(n2933) );
  NAND2_X1 U3657 ( .A1(n3207), .A2(REG0_REG_24__SCAN_IN), .ZN(n2930) );
  NAND2_X1 U3658 ( .A1(n2235), .A2(REG1_REG_24__SCAN_IN), .ZN(n2929) );
  XNOR2_X1 U3659 ( .A(n2940), .B(REG3_REG_24__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U3660 ( .A1(n2977), .A2(n4163), .ZN(n2928) );
  NAND2_X1 U3661 ( .A1(n2603), .A2(REG2_REG_24__SCAN_IN), .ZN(n2927) );
  OR2_X1 U3662 ( .A1(n4173), .A2(n2629), .ZN(n2932) );
  NAND2_X1 U3663 ( .A1(n3095), .A2(n2600), .ZN(n2931) );
  NAND2_X1 U3664 ( .A1(n2932), .A2(n2931), .ZN(n2934) );
  INV_X1 U3665 ( .A(n2933), .ZN(n2936) );
  INV_X1 U3666 ( .A(n2934), .ZN(n2935) );
  INV_X1 U3667 ( .A(n3095), .ZN(n4161) );
  OAI22_X1 U3668 ( .A1(n4173), .A2(n2972), .B1(n4161), .B2(n2627), .ZN(n2939)
         );
  XOR2_X1 U3669 ( .A(n2973), .B(n2939), .Z(n3780) );
  NAND2_X1 U3670 ( .A1(n2692), .A2(REG1_REG_25__SCAN_IN), .ZN(n2945) );
  NAND2_X1 U3671 ( .A1(n3207), .A2(REG0_REG_25__SCAN_IN), .ZN(n2944) );
  INV_X1 U3672 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3782) );
  INV_X1 U3673 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3774) );
  OAI21_X1 U3674 ( .B1(n2940), .B2(n3782), .A(n3774), .ZN(n2941) );
  AND2_X1 U3675 ( .A1(n2941), .A2(n2951), .ZN(n4134) );
  NAND2_X1 U3676 ( .A1(n2977), .A2(n4134), .ZN(n2943) );
  NAND2_X1 U3677 ( .A1(n2603), .A2(REG2_REG_25__SCAN_IN), .ZN(n2942) );
  OAI22_X1 U3678 ( .A1(n4155), .A2(n2972), .B1(n3061), .B2(n2627), .ZN(n2946)
         );
  XNOR2_X1 U3679 ( .A(n2946), .B(n2984), .ZN(n2950) );
  OR2_X1 U3680 ( .A1(n4155), .A2(n2629), .ZN(n2948) );
  NAND2_X1 U3681 ( .A1(n4141), .A2(n2600), .ZN(n2947) );
  AND2_X1 U3682 ( .A1(n2948), .A2(n2947), .ZN(n2949) );
  NAND2_X1 U3683 ( .A1(n2950), .A2(n2949), .ZN(n3770) );
  NOR2_X1 U3684 ( .A1(n2950), .A2(n2949), .ZN(n3772) );
  NAND2_X1 U3685 ( .A1(n2692), .A2(REG1_REG_26__SCAN_IN), .ZN(n2956) );
  NAND2_X1 U3686 ( .A1(n3207), .A2(REG0_REG_26__SCAN_IN), .ZN(n2955) );
  INV_X1 U3687 ( .A(REG3_REG_26__SCAN_IN), .ZN(n5043) );
  AND2_X1 U3688 ( .A1(n2951), .A2(n5043), .ZN(n2952) );
  NOR2_X1 U3689 ( .A1(n2965), .A2(n2952), .ZN(n4127) );
  NAND2_X1 U3690 ( .A1(n2977), .A2(n4127), .ZN(n2954) );
  NAND2_X1 U3691 ( .A1(n2603), .A2(REG2_REG_26__SCAN_IN), .ZN(n2953) );
  NAND4_X1 U3692 ( .A1(n2956), .A2(n2955), .A3(n2954), .A4(n2953), .ZN(n4143)
         );
  NAND2_X1 U3693 ( .A1(n4143), .A2(n2600), .ZN(n2958) );
  NAND2_X1 U3694 ( .A1(n3096), .A2(n2986), .ZN(n2957) );
  NAND2_X1 U3695 ( .A1(n2958), .A2(n2957), .ZN(n2959) );
  XNOR2_X1 U3696 ( .A(n2959), .B(n2984), .ZN(n2964) );
  INV_X1 U3697 ( .A(n2964), .ZN(n2962) );
  NOR2_X1 U3698 ( .A1(n4126), .A2(n2972), .ZN(n2960) );
  AOI21_X1 U3699 ( .B1(n4143), .B2(n2658), .A(n2960), .ZN(n2963) );
  INV_X1 U3700 ( .A(n2963), .ZN(n2961) );
  NAND2_X1 U3701 ( .A1(n2962), .A2(n2961), .ZN(n3807) );
  AND2_X1 U3702 ( .A1(n2964), .A2(n2963), .ZN(n3806) );
  NAND2_X1 U3703 ( .A1(n2692), .A2(REG1_REG_27__SCAN_IN), .ZN(n2970) );
  NAND2_X1 U3704 ( .A1(n3207), .A2(REG0_REG_27__SCAN_IN), .ZN(n2969) );
  NOR2_X1 U3705 ( .A1(n2965), .A2(REG3_REG_27__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3706 ( .A1(n2977), .A2(n3736), .ZN(n2968) );
  NAND2_X1 U3707 ( .A1(n3206), .A2(REG2_REG_27__SCAN_IN), .ZN(n2967) );
  NAND4_X1 U3708 ( .A1(n2970), .A2(n2969), .A3(n2968), .A4(n2967), .ZN(n3978)
         );
  OAI22_X1 U3709 ( .A1(n4118), .A2(n2629), .B1(n4106), .B2(n2971), .ZN(n2995)
         );
  OAI22_X1 U3710 ( .A1(n4118), .A2(n2972), .B1(n4106), .B2(n2627), .ZN(n2974)
         );
  XNOR2_X1 U3711 ( .A(n2974), .B(n2973), .ZN(n2996) );
  XOR2_X1 U3712 ( .A(n2995), .B(n2996), .Z(n3732) );
  NAND2_X1 U3713 ( .A1(n3207), .A2(REG0_REG_28__SCAN_IN), .ZN(n2981) );
  NAND2_X1 U3714 ( .A1(n2692), .A2(REG1_REG_28__SCAN_IN), .ZN(n2980) );
  NOR2_X1 U3715 ( .A1(n2975), .A2(REG3_REG_28__SCAN_IN), .ZN(n2976) );
  NAND2_X1 U3716 ( .A1(n2977), .A2(n3021), .ZN(n2979) );
  NAND2_X1 U3717 ( .A1(n3206), .A2(REG2_REG_28__SCAN_IN), .ZN(n2978) );
  NAND4_X1 U3718 ( .A1(n2981), .A2(n2980), .A3(n2979), .A4(n2978), .ZN(n4076)
         );
  NAND2_X1 U3719 ( .A1(n4076), .A2(n2658), .ZN(n2983) );
  INV_X1 U3720 ( .A(n3118), .ZN(n4077) );
  NAND2_X1 U3721 ( .A1(n4077), .A2(n2600), .ZN(n2982) );
  NAND2_X1 U3722 ( .A1(n2983), .A2(n2982), .ZN(n2985) );
  XNOR2_X1 U3723 ( .A(n2985), .B(n2984), .ZN(n2988) );
  AOI22_X1 U3724 ( .A1(n4076), .A2(n2600), .B1(n4077), .B2(n2986), .ZN(n2987)
         );
  XNOR2_X1 U3725 ( .A(n2988), .B(n2987), .ZN(n2999) );
  NAND2_X1 U3726 ( .A1(n3120), .A2(n2989), .ZN(n3012) );
  INV_X1 U3727 ( .A(n3012), .ZN(n2994) );
  NAND2_X1 U3728 ( .A1(n2990), .A2(n4629), .ZN(n2992) );
  INV_X1 U3729 ( .A(n3141), .ZN(n2991) );
  NAND2_X1 U3730 ( .A1(n2992), .A2(n2991), .ZN(n3001) );
  NOR2_X1 U3731 ( .A1(n3140), .A2(n3001), .ZN(n2993) );
  INV_X1 U3732 ( .A(n2999), .ZN(n2997) );
  NAND2_X1 U3733 ( .A1(n2996), .A2(n2995), .ZN(n2998) );
  INV_X1 U3734 ( .A(n2998), .ZN(n3000) );
  NAND3_X1 U3735 ( .A1(n3000), .A2(n4441), .A3(n2999), .ZN(n3023) );
  NAND2_X1 U3736 ( .A1(n3001), .A2(n4255), .ZN(n3002) );
  NAND2_X1 U3737 ( .A1(n3012), .A2(n3002), .ZN(n3003) );
  NAND2_X1 U3738 ( .A1(n3003), .A2(n3110), .ZN(n3196) );
  NAND2_X1 U3739 ( .A1(n2597), .A2(n3142), .ZN(n3004) );
  OAI21_X1 U3740 ( .B1(n3196), .B2(n3004), .A(STATE_REG_SCAN_IN), .ZN(n3007)
         );
  NOR2_X1 U3741 ( .A1(n4606), .A2(n3005), .ZN(n3006) );
  NAND2_X1 U3742 ( .A1(n3012), .A2(n3011), .ZN(n3197) );
  OR2_X1 U3743 ( .A1(n3140), .A2(n4255), .ZN(n3008) );
  OR2_X1 U3744 ( .A1(n3012), .A2(n3008), .ZN(n3009) );
  INV_X1 U3745 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3010) );
  OAI22_X1 U3746 ( .A1(n4433), .A2(n3118), .B1(STATE_REG_SCAN_IN), .B2(n3010), 
        .ZN(n3020) );
  INV_X1 U3747 ( .A(n3011), .ZN(n3973) );
  NOR2_X1 U3748 ( .A1(n3012), .A2(n3973), .ZN(n3014) );
  NAND2_X1 U3749 ( .A1(n3207), .A2(REG0_REG_29__SCAN_IN), .ZN(n3018) );
  NAND2_X1 U3750 ( .A1(n2692), .A2(REG1_REG_29__SCAN_IN), .ZN(n3017) );
  NAND2_X1 U3751 ( .A1(n2977), .A2(n4075), .ZN(n3016) );
  NAND2_X1 U3752 ( .A1(n3206), .A2(REG2_REG_29__SCAN_IN), .ZN(n3015) );
  OAI22_X1 U3753 ( .A1(n4118), .A2(n4430), .B1(n4429), .B2(n3817), .ZN(n3019)
         );
  AOI211_X1 U3754 ( .C1(n3021), .C2(n3812), .A(n3020), .B(n3019), .ZN(n3022)
         );
  XNOR2_X1 U3755 ( .A(n3269), .B(n4389), .ZN(n3024) );
  NAND2_X1 U3756 ( .A1(n3024), .A2(n4058), .ZN(n3613) );
  INV_X1 U3757 ( .A(n4106), .ZN(n3098) );
  AND2_X1 U3758 ( .A1(n2608), .A2(n4628), .ZN(n3305) );
  NAND2_X1 U3759 ( .A1(n3063), .A2(n3305), .ZN(n3307) );
  NAND2_X1 U3760 ( .A1(n3025), .A2(n2231), .ZN(n3027) );
  NAND2_X1 U3761 ( .A1(n3307), .A2(n3027), .ZN(n3444) );
  INV_X1 U3762 ( .A(n3444), .ZN(n3028) );
  NAND2_X1 U3763 ( .A1(n3386), .A2(n3448), .ZN(n3902) );
  NAND2_X1 U3764 ( .A1(n3753), .A2(n3457), .ZN(n3905) );
  NAND2_X1 U3765 ( .A1(n3028), .A2(n3065), .ZN(n3446) );
  NAND2_X1 U3766 ( .A1(n3386), .A2(n3457), .ZN(n3029) );
  NAND2_X1 U3767 ( .A1(n3446), .A2(n3029), .ZN(n3254) );
  NOR2_X1 U3768 ( .A1(n3449), .A2(n3387), .ZN(n3255) );
  NAND2_X1 U3769 ( .A1(n3991), .A2(n3030), .ZN(n3911) );
  NAND2_X1 U3770 ( .A1(n3991), .A2(n3261), .ZN(n3033) );
  INV_X1 U3771 ( .A(n3033), .ZN(n3032) );
  NOR2_X1 U3772 ( .A1(n3259), .A2(n3032), .ZN(n3035) );
  OR2_X1 U3773 ( .A1(n3255), .A2(n3035), .ZN(n3037) );
  NAND2_X1 U3774 ( .A1(n3449), .A2(n3387), .ZN(n3256) );
  AND2_X1 U3775 ( .A1(n3256), .A2(n3033), .ZN(n3034) );
  OR2_X1 U3776 ( .A1(n3035), .A2(n3034), .ZN(n3036) );
  OAI21_X1 U3777 ( .B1(n3254), .B2(n3037), .A(n3036), .ZN(n3415) );
  AND2_X1 U3778 ( .A1(n3990), .A2(n3411), .ZN(n3038) );
  OAI22_X1 U3779 ( .A1(n3415), .A2(n3038), .B1(n3411), .B2(n3990), .ZN(n3279)
         );
  NOR2_X1 U3780 ( .A1(n3989), .A2(n3331), .ZN(n3280) );
  AND2_X1 U3781 ( .A1(n3274), .A2(n3366), .ZN(n3040) );
  NAND2_X1 U3782 ( .A1(n3988), .A2(n3322), .ZN(n3039) );
  NAND2_X1 U3783 ( .A1(n2251), .A2(n3039), .ZN(n3372) );
  NAND2_X1 U3784 ( .A1(n3989), .A2(n3331), .ZN(n3281) );
  AND2_X1 U3785 ( .A1(n3281), .A2(n3039), .ZN(n3370) );
  INV_X1 U3786 ( .A(n3370), .ZN(n3041) );
  NOR2_X1 U3787 ( .A1(n3041), .A2(n3040), .ZN(n3042) );
  OR2_X1 U3788 ( .A1(n3043), .A2(n3042), .ZN(n3044) );
  OAI21_X1 U3789 ( .B1(n3279), .B2(n3045), .A(n3044), .ZN(n3047) );
  NAND2_X1 U3790 ( .A1(n3430), .A2(n2336), .ZN(n3046) );
  NAND2_X1 U3791 ( .A1(n3047), .A2(n3046), .ZN(n3355) );
  INV_X1 U3792 ( .A(n3987), .ZN(n3376) );
  INV_X1 U3793 ( .A(n3432), .ZN(n3071) );
  NAND2_X1 U3794 ( .A1(n3519), .A2(n3477), .ZN(n3512) );
  NAND2_X1 U3795 ( .A1(n3464), .A2(n3523), .ZN(n3048) );
  INV_X1 U3796 ( .A(n3048), .ZN(n3049) );
  NAND2_X1 U3797 ( .A1(n3464), .A2(n3517), .ZN(n3891) );
  INV_X1 U3798 ( .A(n3464), .ZN(n3986) );
  NAND2_X1 U3799 ( .A1(n3986), .A2(n3523), .ZN(n3935) );
  NAND2_X1 U3800 ( .A1(n3891), .A2(n3935), .ZN(n3514) );
  INV_X1 U3801 ( .A(n3985), .ZN(n3609) );
  INV_X1 U3802 ( .A(n3567), .ZN(n3562) );
  NOR2_X1 U3803 ( .A1(n3631), .A2(n3076), .ZN(n3050) );
  OAI22_X1 U3804 ( .A1(n3603), .A2(n3050), .B1(n3615), .B2(n3984), .ZN(n3625)
         );
  NAND2_X1 U3805 ( .A1(n4431), .A2(n3628), .ZN(n3895) );
  NAND2_X1 U3806 ( .A1(n3983), .A2(n3637), .ZN(n3823) );
  NAND2_X1 U3807 ( .A1(n3895), .A2(n3823), .ZN(n3624) );
  NAND2_X1 U3808 ( .A1(n3625), .A2(n3624), .ZN(n3623) );
  NAND2_X1 U3809 ( .A1(n3623), .A2(n3051), .ZN(n3651) );
  NOR2_X1 U3810 ( .A1(n3982), .A2(n3077), .ZN(n3052) );
  INV_X1 U3811 ( .A(n3982), .ZN(n4397) );
  INV_X1 U3812 ( .A(n3077), .ZN(n4432) );
  NOR2_X1 U3813 ( .A1(n4428), .A2(n3672), .ZN(n3942) );
  NAND2_X1 U3814 ( .A1(n4428), .A2(n3672), .ZN(n3944) );
  INV_X1 U3815 ( .A(n3981), .ZN(n4421) );
  NAND2_X1 U3816 ( .A1(n4421), .A2(n3082), .ZN(n3053) );
  NOR2_X1 U3817 ( .A1(n4259), .A2(n4420), .ZN(n4249) );
  AND2_X1 U3818 ( .A1(n4259), .A2(n4420), .ZN(n4250) );
  NOR2_X1 U3819 ( .A1(n4249), .A2(n4250), .ZN(n3862) );
  INV_X1 U3820 ( .A(n3862), .ZN(n3689) );
  NAND2_X1 U3821 ( .A1(n3690), .A2(n3689), .ZN(n3688) );
  NAND2_X1 U3822 ( .A1(n3688), .A2(n3054), .ZN(n4248) );
  NAND2_X1 U3823 ( .A1(n4234), .A2(n3860), .ZN(n3056) );
  INV_X1 U3824 ( .A(n4222), .ZN(n4257) );
  INV_X1 U3825 ( .A(n4227), .ZN(n3218) );
  NAND2_X1 U3826 ( .A1(n4215), .A2(n4192), .ZN(n4170) );
  INV_X1 U3827 ( .A(n4215), .ZN(n4175) );
  NAND2_X1 U3828 ( .A1(n4175), .A2(n4202), .ZN(n3089) );
  NAND2_X1 U3829 ( .A1(n4187), .A2(n3057), .ZN(n4168) );
  NAND2_X1 U3830 ( .A1(n4191), .A2(n4179), .ZN(n3059) );
  INV_X1 U3831 ( .A(n4191), .ZN(n3980) );
  INV_X1 U3832 ( .A(n4173), .ZN(n3979) );
  NAND2_X1 U3833 ( .A1(n3979), .A2(n3095), .ZN(n3060) );
  NAND2_X1 U3834 ( .A1(n4155), .A2(n3061), .ZN(n3062) );
  INV_X1 U3835 ( .A(n4155), .ZN(n4120) );
  NOR2_X1 U3836 ( .A1(n4143), .A2(n3096), .ZN(n3854) );
  INV_X1 U3837 ( .A(n4076), .ZN(n4099) );
  NAND2_X1 U3838 ( .A1(n4099), .A2(n4077), .ZN(n4063) );
  NAND2_X1 U3839 ( .A1(n4076), .A2(n3118), .ZN(n4065) );
  NAND2_X1 U3840 ( .A1(n4063), .A2(n4065), .ZN(n4078) );
  NAND2_X1 U3841 ( .A1(n3064), .A2(n4628), .ZN(n3897) );
  INV_X1 U3842 ( .A(n3449), .ZN(n3263) );
  NAND2_X1 U3843 ( .A1(n3263), .A2(n3387), .ZN(n3907) );
  NAND2_X1 U3844 ( .A1(n3449), .A2(n3394), .ZN(n3904) );
  NAND2_X1 U3845 ( .A1(n3385), .A2(n3877), .ZN(n3066) );
  NAND2_X1 U3846 ( .A1(n3066), .A2(n3907), .ZN(n3260) );
  INV_X1 U3847 ( .A(n3908), .ZN(n3067) );
  INV_X1 U3848 ( .A(n3411), .ZN(n3418) );
  AND2_X1 U3849 ( .A1(n3990), .A2(n3418), .ZN(n3408) );
  INV_X1 U3850 ( .A(n3990), .ZN(n3333) );
  NAND2_X1 U3851 ( .A1(n3333), .A2(n3411), .ZN(n3916) );
  NAND2_X1 U3852 ( .A1(n3989), .A2(n3329), .ZN(n3915) );
  INV_X1 U3853 ( .A(n3989), .ZN(n3319) );
  NAND2_X1 U3854 ( .A1(n3319), .A2(n3331), .ZN(n3913) );
  INV_X1 U3855 ( .A(n3068), .ZN(n3069) );
  NAND2_X1 U3856 ( .A1(n3430), .A2(n3366), .ZN(n3927) );
  NAND2_X1 U3857 ( .A1(n3375), .A2(n3927), .ZN(n3070) );
  NAND2_X1 U3858 ( .A1(n3274), .A2(n2336), .ZN(n3922) );
  AND2_X1 U3859 ( .A1(n3987), .A2(n3071), .ZN(n3354) );
  INV_X1 U3860 ( .A(n3354), .ZN(n3072) );
  NAND2_X1 U3861 ( .A1(n3376), .A2(n3432), .ZN(n3928) );
  NAND2_X1 U3862 ( .A1(n3359), .A2(n3477), .ZN(n3934) );
  NAND2_X1 U3863 ( .A1(n3463), .A2(n3934), .ZN(n3074) );
  NAND2_X1 U3864 ( .A1(n3519), .A2(n3073), .ZN(n3932) );
  NAND2_X1 U3865 ( .A1(n3074), .A2(n3932), .ZN(n3516) );
  NAND2_X1 U3866 ( .A1(n3516), .A2(n3935), .ZN(n3075) );
  NOR2_X1 U3867 ( .A1(n3985), .A2(n3562), .ZN(n3892) );
  NAND2_X1 U3868 ( .A1(n3985), .A2(n3562), .ZN(n3605) );
  NAND2_X1 U3869 ( .A1(n3984), .A2(n3076), .ZN(n3604) );
  NAND2_X1 U3870 ( .A1(n3631), .A2(n3615), .ZN(n3894) );
  INV_X1 U3871 ( .A(n3624), .ZN(n3876) );
  NAND2_X1 U3872 ( .A1(n4397), .A2(n3077), .ZN(n3893) );
  NAND2_X1 U3873 ( .A1(n3982), .A2(n4432), .ZN(n3824) );
  NAND2_X1 U3874 ( .A1(n3893), .A2(n3824), .ZN(n3873) );
  INV_X1 U3875 ( .A(n3895), .ZN(n3822) );
  NOR2_X1 U3876 ( .A1(n3873), .A2(n3822), .ZN(n3078) );
  NAND2_X1 U3877 ( .A1(n3654), .A2(n3824), .ZN(n3669) );
  INV_X1 U3878 ( .A(n3666), .ZN(n3851) );
  INV_X1 U3879 ( .A(n3942), .ZN(n3079) );
  AND2_X1 U3880 ( .A1(n4234), .A2(n4264), .ZN(n3080) );
  NOR2_X1 U3881 ( .A1(n4250), .A2(n3080), .ZN(n3085) );
  NAND2_X1 U3882 ( .A1(n3981), .A2(n3082), .ZN(n3697) );
  NAND2_X1 U3883 ( .A1(n3085), .A2(n3697), .ZN(n3941) );
  NOR2_X1 U3884 ( .A1(n3981), .A2(n3082), .ZN(n3698) );
  OR2_X1 U3885 ( .A1(n4249), .A2(n3698), .ZN(n3084) );
  NOR2_X1 U3886 ( .A1(n4234), .A2(n4264), .ZN(n3083) );
  AOI21_X1 U3887 ( .B1(n3085), .B2(n3084), .A(n3083), .ZN(n4228) );
  NAND2_X1 U3888 ( .A1(n4257), .A2(n4239), .ZN(n3086) );
  NAND2_X1 U3889 ( .A1(n4228), .A2(n3086), .ZN(n3947) );
  INV_X1 U3890 ( .A(n3947), .ZN(n3087) );
  NAND2_X1 U3891 ( .A1(n4229), .A2(n3087), .ZN(n3088) );
  NAND2_X1 U3892 ( .A1(n4222), .A2(n4226), .ZN(n3946) );
  NAND2_X1 U3893 ( .A1(n4227), .A2(n4210), .ZN(n4169) );
  AND2_X1 U3894 ( .A1(n4170), .A2(n4169), .ZN(n3951) );
  OR2_X1 U3895 ( .A1(n4191), .A2(n3094), .ZN(n3090) );
  NAND2_X1 U3896 ( .A1(n3090), .A2(n3089), .ZN(n3952) );
  INV_X1 U3897 ( .A(n3952), .ZN(n3093) );
  OR2_X1 U3898 ( .A1(n4227), .A2(n4210), .ZN(n3945) );
  INV_X1 U3899 ( .A(n3945), .ZN(n3091) );
  NAND2_X1 U3900 ( .A1(n3091), .A2(n4170), .ZN(n3092) );
  AND2_X1 U3901 ( .A1(n3093), .A2(n3092), .ZN(n3832) );
  NAND2_X1 U3902 ( .A1(n4173), .A2(n3095), .ZN(n3864) );
  NAND2_X1 U3903 ( .A1(n4191), .A2(n3094), .ZN(n4151) );
  NOR2_X1 U3904 ( .A1(n4173), .A2(n3095), .ZN(n3863) );
  NOR2_X1 U3905 ( .A1(n4155), .A2(n4141), .ZN(n3852) );
  NOR2_X1 U3906 ( .A1(n3863), .A2(n3852), .ZN(n3955) );
  NAND2_X1 U3907 ( .A1(n4155), .A2(n4141), .ZN(n4114) );
  INV_X1 U3908 ( .A(n4143), .ZN(n4098) );
  NAND2_X1 U3909 ( .A1(n4098), .A2(n3096), .ZN(n3097) );
  NAND2_X1 U3910 ( .A1(n4114), .A2(n3097), .ZN(n3953) );
  INV_X1 U3911 ( .A(n3953), .ZN(n3837) );
  AND2_X1 U3912 ( .A1(n4143), .A2(n4126), .ZN(n3962) );
  AND2_X1 U3913 ( .A1(n3978), .A2(n4106), .ZN(n3957) );
  INV_X1 U3914 ( .A(n3957), .ZN(n3099) );
  NAND2_X1 U3915 ( .A1(n4118), .A2(n3098), .ZN(n3815) );
  NAND2_X1 U3916 ( .A1(n4097), .A2(n4103), .ZN(n4096) );
  NAND2_X1 U3917 ( .A1(n4096), .A2(n3815), .ZN(n4066) );
  XNOR2_X1 U3918 ( .A(n4066), .B(n4078), .ZN(n3101) );
  NAND2_X1 U3919 ( .A1(n4391), .A2(n4390), .ZN(n3967) );
  INV_X1 U3920 ( .A(n4058), .ZN(n4392) );
  NAND2_X1 U3921 ( .A1(n4392), .A2(n4389), .ZN(n3100) );
  OAI22_X1 U3922 ( .A1(n3817), .A2(n4256), .B1(n4255), .B2(n3118), .ZN(n3102)
         );
  INV_X1 U3923 ( .A(n3102), .ZN(n3103) );
  INV_X1 U3924 ( .A(n3104), .ZN(n3105) );
  NAND2_X1 U3925 ( .A1(n3108), .A2(n3107), .ZN(n3115) );
  OAI21_X1 U3926 ( .B1(n3134), .B2(D_REG_1__SCAN_IN), .A(n3109), .ZN(n3114) );
  NAND2_X1 U3927 ( .A1(n3111), .A2(n3110), .ZN(n3112) );
  NOR2_X1 U3928 ( .A1(n3140), .A2(n3112), .ZN(n3113) );
  INV_X1 U3929 ( .A(n4083), .ZN(n3117) );
  OAI21_X1 U3930 ( .B1(n3116), .B2(n3118), .A(n3117), .ZN(n4089) );
  NAND2_X1 U3931 ( .A1(n4684), .A2(n2598), .ZN(n4333) );
  INV_X1 U3932 ( .A(n3120), .ZN(n3122) );
  INV_X1 U3933 ( .A(n3124), .ZN(n3126) );
  NAND2_X1 U3934 ( .A1(n4673), .A2(n2598), .ZN(n4379) );
  NAND2_X1 U3935 ( .A1(n3126), .A2(n3125), .ZN(U3514) );
  INV_X2 U3936 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND3_X1 U3937 ( .A1(n3127), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3129) );
  INV_X1 U3938 ( .A(DATAI_31_), .ZN(n3128) );
  OAI22_X1 U3939 ( .A1(n3130), .A2(n3129), .B1(STATE_REG_SCAN_IN), .B2(n3128), 
        .ZN(U3321) );
  INV_X1 U3940 ( .A(DATAI_29_), .ZN(n3133) );
  NAND2_X1 U3941 ( .A1(n3131), .A2(STATE_REG_SCAN_IN), .ZN(n3132) );
  OAI21_X1 U3942 ( .B1(STATE_REG_SCAN_IN), .B2(n3133), .A(n3132), .ZN(U3323)
         );
  AOI22_X1 U3943 ( .A1(n4685), .A2(n3136), .B1(n3135), .B2(n3137), .ZN(U3458)
         );
  INV_X1 U3944 ( .A(D_REG_1__SCAN_IN), .ZN(n4925) );
  AOI22_X1 U3945 ( .A1(n4685), .A2(n4925), .B1(n3138), .B2(n3137), .ZN(U3459)
         );
  INV_X1 U3946 ( .A(n3142), .ZN(n3139) );
  NAND2_X1 U3947 ( .A1(n3139), .A2(STATE_REG_SCAN_IN), .ZN(n3976) );
  NAND2_X1 U3948 ( .A1(n3140), .A2(n3976), .ZN(n3159) );
  NAND2_X1 U3949 ( .A1(n3142), .A2(n3141), .ZN(n3143) );
  AND2_X1 U3950 ( .A1(n3144), .A2(n3143), .ZN(n3158) );
  NAND2_X1 U3951 ( .A1(n3159), .A2(n3158), .ZN(n4455) );
  NOR2_X1 U3952 ( .A1(n4455), .A2(n4452), .ZN(n4577) );
  INV_X1 U3953 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3145) );
  MUX2_X1 U3954 ( .A(REG1_REG_1__SCAN_IN), .B(n3145), .S(n2232), .Z(n3993) );
  AND2_X1 U3955 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3994)
         );
  NAND2_X1 U3956 ( .A1(n2232), .A2(REG1_REG_1__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U3957 ( .A1(n3992), .A2(n4016), .ZN(n3148) );
  INV_X1 U3958 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3147) );
  MUX2_X1 U3959 ( .A(REG1_REG_2__SCAN_IN), .B(n3147), .S(n3146), .Z(n4015) );
  NAND2_X1 U3960 ( .A1(n3146), .A2(REG1_REG_2__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U3961 ( .A1(n4019), .A2(n3149), .ZN(n3165) );
  XOR2_X1 U3962 ( .A(n3164), .B(REG1_REG_3__SCAN_IN), .Z(n3157) );
  NAND2_X1 U3963 ( .A1(n4386), .A2(n4452), .ZN(n4008) );
  NOR2_X2 U3964 ( .A1(n4455), .A2(n4008), .ZN(n4588) );
  INV_X1 U3965 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3151) );
  MUX2_X1 U3966 ( .A(REG2_REG_1__SCAN_IN), .B(n3151), .S(n3150), .Z(n3995) );
  AND2_X1 U3967 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4000)
         );
  NAND2_X1 U3968 ( .A1(n3995), .A2(n4000), .ZN(n4010) );
  NAND2_X1 U3969 ( .A1(n2232), .A2(REG2_REG_1__SCAN_IN), .ZN(n4009) );
  NAND2_X1 U3970 ( .A1(n4010), .A2(n4009), .ZN(n3154) );
  INV_X1 U3971 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3152) );
  MUX2_X1 U3972 ( .A(REG2_REG_2__SCAN_IN), .B(n3152), .S(n3146), .Z(n3153) );
  NAND2_X1 U3973 ( .A1(n3154), .A2(n3153), .ZN(n4013) );
  NAND2_X1 U3974 ( .A1(n3146), .A2(REG2_REG_2__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U3975 ( .A1(n4013), .A2(n3155), .ZN(n3177) );
  XNOR2_X1 U3976 ( .A(n3177), .B(n3163), .ZN(n3176) );
  XOR2_X1 U3977 ( .A(n3176), .B(REG2_REG_3__SCAN_IN), .Z(n3156) );
  AOI22_X1 U3978 ( .A1(n4577), .A2(n3157), .B1(n4588), .B2(n3156), .ZN(n3162)
         );
  INV_X1 U3979 ( .A(n3158), .ZN(n3160) );
  NOR2_X1 U3980 ( .A1(STATE_REG_SCAN_IN), .A2(n2637), .ZN(n3232) );
  AOI21_X1 U3981 ( .B1(n4581), .B2(ADDR_REG_3__SCAN_IN), .A(n3232), .ZN(n3161)
         );
  OAI211_X1 U3982 ( .C1(n3163), .C2(n4593), .A(n3162), .B(n3161), .ZN(U3243)
         );
  MUX2_X1 U3983 ( .A(REG1_REG_7__SCAN_IN), .B(n2371), .S(n4395), .Z(n3175) );
  NAND2_X1 U3984 ( .A1(n3164), .A2(REG1_REG_3__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U3985 ( .A1(n3165), .A2(n4396), .ZN(n3166) );
  NAND2_X1 U3986 ( .A1(n3167), .A2(n3166), .ZN(n3169) );
  XNOR2_X1 U3987 ( .A(n3169), .B(n4461), .ZN(n4459) );
  INV_X1 U3988 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3168) );
  INV_X1 U3989 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4952) );
  MUX2_X1 U3990 ( .A(n4952), .B(REG1_REG_5__SCAN_IN), .S(n4479), .Z(n4475) );
  NAND2_X1 U3991 ( .A1(n3171), .A2(n3170), .ZN(n3172) );
  NAND2_X1 U3992 ( .A1(n4489), .A2(n3172), .ZN(n3173) );
  OAI21_X1 U3993 ( .B1(n3175), .B2(n3497), .A(n4577), .ZN(n3174) );
  AOI21_X1 U3994 ( .B1(n3175), .B2(n3497), .A(n3174), .ZN(n3193) );
  INV_X1 U3995 ( .A(n4395), .ZN(n3191) );
  INV_X1 U3996 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U3997 ( .A1(n3176), .A2(REG2_REG_3__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U3998 ( .A1(n3177), .A2(n4396), .ZN(n3178) );
  NAND2_X1 U3999 ( .A1(n3179), .A2(n3178), .ZN(n3180) );
  XNOR2_X1 U4000 ( .A(n3180), .B(n4461), .ZN(n4457) );
  NAND2_X1 U4001 ( .A1(n3180), .A2(n4461), .ZN(n3181) );
  MUX2_X1 U4002 ( .A(n3420), .B(REG2_REG_5__SCAN_IN), .S(n4479), .Z(n4472) );
  NAND2_X1 U4003 ( .A1(n4489), .A2(n3184), .ZN(n3185) );
  INV_X1 U4004 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3186) );
  MUX2_X1 U4005 ( .A(REG2_REG_7__SCAN_IN), .B(n3186), .S(n4395), .Z(n3187) );
  OAI211_X1 U4006 ( .C1(n3188), .C2(n3187), .A(n4588), .B(n3486), .ZN(n3190)
         );
  AND2_X1 U4007 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3321) );
  AOI21_X1 U4008 ( .B1(n4581), .B2(ADDR_REG_7__SCAN_IN), .A(n3321), .ZN(n3189)
         );
  OAI211_X1 U4009 ( .C1(n4593), .C2(n3191), .A(n3190), .B(n3189), .ZN(n3192)
         );
  OR2_X1 U4010 ( .A1(n3193), .A2(n3192), .ZN(U3247) );
  NOR2_X1 U4011 ( .A1(n4581), .A2(U4043), .ZN(U3148) );
  XNOR2_X1 U4012 ( .A(n3195), .B(n3194), .ZN(n4002) );
  INV_X1 U4013 ( .A(n3196), .ZN(n3199) );
  NAND3_X1 U4014 ( .A1(n3199), .A2(n3198), .A3(n3197), .ZN(n3756) );
  OAI22_X1 U4015 ( .A1(n4429), .A2(n3451), .B1(n4433), .B2(n2609), .ZN(n3200)
         );
  AOI21_X1 U4016 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3756), .A(n3200), .ZN(n3201)
         );
  OAI21_X1 U4017 ( .B1(n4002), .B2(n4418), .A(n3201), .ZN(U3229) );
  INV_X1 U4018 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4862) );
  INV_X1 U4019 ( .A(n4428), .ZN(n3202) );
  NAND2_X1 U4020 ( .A1(n3202), .A2(U4043), .ZN(n3203) );
  OAI21_X1 U4021 ( .B1(U4043), .B2(n4862), .A(n3203), .ZN(U3566) );
  INV_X1 U4022 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U4023 ( .A1(n4259), .A2(U4043), .ZN(n3204) );
  OAI21_X1 U4024 ( .B1(U4043), .B2(n4875), .A(n3204), .ZN(U3568) );
  INV_X1 U4025 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U4026 ( .A1(n3449), .A2(U4043), .ZN(n3205) );
  OAI21_X1 U4027 ( .B1(U4043), .B2(n4834), .A(n3205), .ZN(U3553) );
  INV_X1 U4028 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U4029 ( .A1(n2692), .A2(REG1_REG_30__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4030 ( .A1(n3206), .A2(REG2_REG_30__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4031 ( .A1(n3207), .A2(REG0_REG_30__SCAN_IN), .ZN(n3208) );
  NAND3_X1 U4032 ( .A1(n3210), .A2(n3209), .A3(n3208), .ZN(n4070) );
  NAND2_X1 U4033 ( .A1(n4070), .A2(U4043), .ZN(n3211) );
  OAI21_X1 U4034 ( .B1(U4043), .B2(n4898), .A(n3211), .ZN(U3580) );
  INV_X1 U4035 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4841) );
  NAND2_X1 U4036 ( .A1(n3359), .A2(U4043), .ZN(n3212) );
  OAI21_X1 U4037 ( .B1(U4043), .B2(n4841), .A(n3212), .ZN(U3560) );
  INV_X1 U4038 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U4039 ( .A1(n3839), .A2(U4043), .ZN(n3213) );
  OAI21_X1 U4040 ( .B1(U4043), .B2(n4955), .A(n3213), .ZN(U3581) );
  INV_X1 U4041 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4958) );
  NAND2_X1 U4042 ( .A1(n3753), .A2(U4043), .ZN(n3214) );
  OAI21_X1 U40430 ( .B1(U4043), .B2(n4958), .A(n3214), .ZN(U3552) );
  INV_X1 U4044 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U4045 ( .A1(n4234), .A2(U4043), .ZN(n3215) );
  OAI21_X1 U4046 ( .B1(U4043), .B2(n4840), .A(n3215), .ZN(U3569) );
  INV_X1 U4047 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U4048 ( .A1(n4175), .A2(U4043), .ZN(n3216) );
  OAI21_X1 U4049 ( .B1(U4043), .B2(n4968), .A(n3216), .ZN(U3572) );
  INV_X1 U4050 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U4051 ( .A1(n3274), .A2(U4043), .ZN(n3217) );
  OAI21_X1 U4052 ( .B1(U4043), .B2(n4833), .A(n3217), .ZN(U3558) );
  INV_X1 U4053 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U4054 ( .A1(n3218), .A2(U4043), .ZN(n3219) );
  OAI21_X1 U4055 ( .B1(U4043), .B2(n4843), .A(n3219), .ZN(U3571) );
  INV_X1 U4056 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U4057 ( .A1(n2608), .A2(U4043), .ZN(n3220) );
  OAI21_X1 U4058 ( .B1(U4043), .B2(n4931), .A(n3220), .ZN(U3550) );
  INV_X1 U4059 ( .A(n3222), .ZN(n3223) );
  AOI21_X1 U4060 ( .B1(n3221), .B2(n3224), .A(n3223), .ZN(n3227) );
  INV_X1 U4061 ( .A(n4429), .ZN(n3754) );
  AOI22_X1 U4062 ( .A1(n3754), .A2(n3449), .B1(n3752), .B2(n3448), .ZN(n3226)
         );
  INV_X1 U4063 ( .A(n4430), .ZN(n3755) );
  AOI22_X1 U4064 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3756), .B1(n3755), .B2(n3025), .ZN(n3225) );
  OAI211_X1 U4065 ( .C1(n3227), .C2(n4418), .A(n3226), .B(n3225), .ZN(U3234)
         );
  XNOR2_X1 U4066 ( .A(n3228), .B(n3229), .ZN(n3230) );
  NAND2_X1 U4067 ( .A1(n3230), .A2(n4441), .ZN(n3234) );
  OAI22_X1 U4068 ( .A1(n3031), .A2(n4429), .B1(n4430), .B2(n3386), .ZN(n3231)
         );
  AOI211_X1 U4069 ( .C1(n3387), .C2(n3752), .A(n3232), .B(n3231), .ZN(n3233)
         );
  OAI211_X1 U4070 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4446), .A(n3234), .B(n3233), 
        .ZN(U3215) );
  INV_X1 U4071 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U4072 ( .A1(n4120), .A2(U4043), .ZN(n3235) );
  OAI21_X1 U4073 ( .B1(U4043), .B2(n4904), .A(n3235), .ZN(U3575) );
  INV_X1 U4074 ( .A(n3236), .ZN(n3253) );
  OAI211_X1 U4075 ( .C1(n3239), .C2(n3238), .A(n3237), .B(n4441), .ZN(n3242)
         );
  AND2_X1 U4076 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4462) );
  OAI22_X1 U4077 ( .A1(n3263), .A2(n4430), .B1(n4429), .B2(n3333), .ZN(n3240)
         );
  AOI211_X1 U4078 ( .C1(n3261), .C2(n3752), .A(n4462), .B(n3240), .ZN(n3241)
         );
  OAI211_X1 U4079 ( .C1(n4446), .C2(n3253), .A(n3242), .B(n3241), .ZN(U3227)
         );
  NAND2_X1 U4080 ( .A1(n4004), .A2(DATAO_REG_29__SCAN_IN), .ZN(n3243) );
  OAI21_X1 U4081 ( .B1(n3817), .B2(n4004), .A(n3243), .ZN(U3579) );
  INV_X1 U4082 ( .A(n3244), .ZN(n3419) );
  OAI211_X1 U4083 ( .C1(n3247), .C2(n3246), .A(n3245), .B(n4441), .ZN(n3250)
         );
  AND2_X1 U4084 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4482) );
  OAI22_X1 U4085 ( .A1(n3031), .A2(n4430), .B1(n4429), .B2(n3319), .ZN(n3248)
         );
  AOI211_X1 U4086 ( .C1(n3411), .C2(n3752), .A(n4482), .B(n3248), .ZN(n3249)
         );
  OAI211_X1 U4087 ( .C1(n4446), .C2(n3419), .A(n3250), .B(n3249), .ZN(U3224)
         );
  AOI211_X1 U4088 ( .C1(n3261), .C2(n3396), .A(n3251), .B(n2337), .ZN(n4648)
         );
  NOR2_X1 U4089 ( .A1(n4268), .A2(n3253), .ZN(n3267) );
  OR2_X1 U4090 ( .A1(n3254), .A2(n3255), .ZN(n3257) );
  NAND2_X1 U4091 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  XNOR2_X1 U4092 ( .A(n3259), .B(n3258), .ZN(n3268) );
  INV_X1 U4093 ( .A(n3259), .ZN(n3879) );
  XNOR2_X1 U4094 ( .A(n3260), .B(n3879), .ZN(n3265) );
  AOI22_X1 U4095 ( .A1(n3990), .A2(n4142), .B1(n4287), .B2(n3261), .ZN(n3262)
         );
  OAI21_X1 U4096 ( .B1(n3263), .B2(n4195), .A(n3262), .ZN(n3264) );
  AOI21_X1 U4097 ( .B1(n3265), .B2(n4197), .A(n3264), .ZN(n3266) );
  OAI21_X1 U4098 ( .B1(n3268), .B2(n3613), .A(n3266), .ZN(n4647) );
  AOI211_X1 U4099 ( .C1(n4648), .C2(n4058), .A(n3267), .B(n4647), .ZN(n3272)
         );
  INV_X2 U4100 ( .A(n4273), .ZN(n4604) );
  INV_X1 U4101 ( .A(n3268), .ZN(n4650) );
  OR2_X1 U4102 ( .A1(n3269), .A2(n4058), .ZN(n3283) );
  INV_X1 U4103 ( .A(n3283), .ZN(n3270) );
  NAND2_X1 U4104 ( .A1(n4273), .A2(n3270), .ZN(n3641) );
  INV_X1 U4105 ( .A(n3641), .ZN(n4599) );
  AOI22_X1 U4106 ( .A1(n4650), .A2(n4599), .B1(REG2_REG_4__SCAN_IN), .B2(n4604), .ZN(n3271) );
  OAI21_X1 U4107 ( .B1(n3272), .B2(n4604), .A(n3271), .ZN(U3286) );
  XNOR2_X1 U4108 ( .A(n3273), .B(n2251), .ZN(n3278) );
  NAND2_X1 U4109 ( .A1(n3989), .A2(n4260), .ZN(n3276) );
  NAND2_X1 U4110 ( .A1(n3274), .A2(n4142), .ZN(n3275) );
  OAI211_X1 U4111 ( .C1(n4255), .C2(n3285), .A(n3276), .B(n3275), .ZN(n3277)
         );
  AOI21_X1 U4112 ( .B1(n3278), .B2(n4197), .A(n3277), .ZN(n4660) );
  OR2_X1 U4113 ( .A1(n3279), .A2(n3280), .ZN(n3371) );
  NAND2_X1 U4114 ( .A1(n3371), .A2(n3281), .ZN(n3282) );
  XNOR2_X1 U4115 ( .A(n3282), .B(n2251), .ZN(n4657) );
  NAND2_X1 U4116 ( .A1(n3613), .A2(n3283), .ZN(n3284) );
  OAI211_X1 U4117 ( .C1(n3327), .C2(n3285), .A(n2598), .B(n3367), .ZN(n4658)
         );
  INV_X1 U4118 ( .A(n3286), .ZN(n3694) );
  NOR2_X1 U4119 ( .A1(n4658), .A2(n3694), .ZN(n3289) );
  INV_X1 U4120 ( .A(n3323), .ZN(n3287) );
  OAI22_X1 U4121 ( .A1(n4273), .A2(n3186), .B1(n3287), .B2(n4268), .ZN(n3288)
         );
  AOI211_X1 U4122 ( .C1(n4657), .C2(n4237), .A(n3289), .B(n3288), .ZN(n3290)
         );
  OAI21_X1 U4123 ( .B1(n4604), .B2(n4660), .A(n3290), .ZN(U3283) );
  XOR2_X1 U4124 ( .A(n3292), .B(n3291), .Z(n3293) );
  XNOR2_X1 U4125 ( .A(n3294), .B(n3293), .ZN(n3298) );
  NOR2_X1 U4126 ( .A1(STATE_REG_SCAN_IN), .A2(n4868), .ZN(n4484) );
  OAI22_X1 U4127 ( .A1(n3333), .A2(n4430), .B1(n4429), .B2(n3349), .ZN(n3295)
         );
  AOI211_X1 U4128 ( .C1(n3331), .C2(n3752), .A(n4484), .B(n3295), .ZN(n3297)
         );
  NAND2_X1 U4129 ( .A1(n3812), .A2(n4595), .ZN(n3296) );
  OAI211_X1 U4130 ( .C1(n3298), .C2(n4418), .A(n3297), .B(n3296), .ZN(U3236)
         );
  NAND2_X1 U4131 ( .A1(n2608), .A2(n2609), .ZN(n3899) );
  AND2_X1 U4132 ( .A1(n3897), .A2(n3899), .ZN(n4624) );
  AOI21_X1 U4133 ( .B1(n4262), .B2(n3613), .A(n4624), .ZN(n3299) );
  AOI21_X1 U4134 ( .B1(n4142), .B2(n3025), .A(n3299), .ZN(n4625) );
  AND2_X1 U4135 ( .A1(n4058), .A2(n4629), .ZN(n3300) );
  OAI21_X1 U4136 ( .B1(n4287), .B2(n3300), .A(n4628), .ZN(n3301) );
  AOI21_X1 U4137 ( .B1(n4625), .B2(n3301), .A(n4604), .ZN(n3302) );
  INV_X1 U4138 ( .A(n3302), .ZN(n3304) );
  AOI22_X1 U4139 ( .A1(n4604), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4594), .ZN(n3303) );
  OAI211_X1 U4140 ( .C1(n4624), .C2(n3641), .A(n3304), .B(n3303), .ZN(U3290)
         );
  OR2_X1 U4141 ( .A1(n3063), .A2(n3305), .ZN(n3306) );
  NAND2_X1 U4142 ( .A1(n3307), .A2(n3306), .ZN(n4631) );
  NAND2_X1 U4143 ( .A1(n2231), .A2(n4287), .ZN(n3309) );
  NAND2_X1 U4144 ( .A1(n2608), .A2(n4260), .ZN(n3308) );
  OAI211_X1 U4145 ( .C1(n3386), .C2(n4256), .A(n3309), .B(n3308), .ZN(n3310)
         );
  INV_X1 U4146 ( .A(n3310), .ZN(n3313) );
  XNOR2_X1 U4147 ( .A(n3063), .B(n3897), .ZN(n3311) );
  NAND2_X1 U4148 ( .A1(n3311), .A2(n4197), .ZN(n3312) );
  OAI211_X1 U4149 ( .C1(n4631), .C2(n3613), .A(n3313), .B(n3312), .ZN(n4632)
         );
  MUX2_X1 U4150 ( .A(n4632), .B(REG2_REG_1__SCAN_IN), .S(n4604), .Z(n3314) );
  INV_X1 U4151 ( .A(n3314), .ZN(n3317) );
  INV_X1 U4152 ( .A(n3315), .ZN(n3458) );
  AOI21_X1 U4153 ( .B1(n4628), .B2(n2231), .A(n3458), .ZN(n4634) );
  AOI22_X1 U4154 ( .A1(n4598), .A2(n4634), .B1(REG3_REG_1__SCAN_IN), .B2(n4594), .ZN(n3316) );
  OAI211_X1 U4155 ( .C1(n4631), .C2(n3641), .A(n3317), .B(n3316), .ZN(U3289)
         );
  XNOR2_X1 U4156 ( .A(n3318), .B(n3343), .ZN(n3326) );
  OAI22_X1 U4157 ( .A1(n3319), .A2(n4430), .B1(n4429), .B2(n3430), .ZN(n3320)
         );
  AOI211_X1 U4158 ( .C1(n3322), .C2(n3752), .A(n3321), .B(n3320), .ZN(n3325)
         );
  NAND2_X1 U4159 ( .A1(n3812), .A2(n3323), .ZN(n3324) );
  OAI211_X1 U4160 ( .C1(n3326), .C2(n4418), .A(n3325), .B(n3324), .ZN(U3210)
         );
  INV_X1 U4161 ( .A(n3327), .ZN(n3328) );
  OAI21_X1 U4162 ( .B1(n3416), .B2(n3329), .A(n3328), .ZN(n4596) );
  INV_X1 U4163 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4906) );
  INV_X1 U4164 ( .A(n4668), .ZN(n4649) );
  AND2_X1 U4165 ( .A1(n3913), .A2(n3915), .ZN(n3855) );
  XNOR2_X1 U4166 ( .A(n3279), .B(n3855), .ZN(n3334) );
  INV_X1 U4167 ( .A(n3334), .ZN(n4600) );
  XNOR2_X1 U4168 ( .A(n3330), .B(n3855), .ZN(n3337) );
  AOI22_X1 U4169 ( .A1(n3988), .A2(n4142), .B1(n4287), .B2(n3331), .ZN(n3332)
         );
  OAI21_X1 U4170 ( .B1(n3333), .B2(n4195), .A(n3332), .ZN(n3336) );
  NOR2_X1 U4171 ( .A1(n3334), .A2(n3613), .ZN(n3335) );
  AOI211_X1 U4172 ( .C1(n3337), .C2(n4197), .A(n3336), .B(n3335), .ZN(n4603)
         );
  INV_X1 U4173 ( .A(n4603), .ZN(n3338) );
  AOI21_X1 U4174 ( .B1(n4649), .B2(n4600), .A(n3338), .ZN(n3340) );
  MUX2_X1 U4175 ( .A(n4906), .B(n3340), .S(n4673), .Z(n3339) );
  OAI21_X1 U4176 ( .B1(n4596), .B2(n4379), .A(n3339), .ZN(U3479) );
  INV_X1 U4177 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3341) );
  MUX2_X1 U4178 ( .A(n3341), .B(n3340), .S(n4684), .Z(n3342) );
  OAI21_X1 U4179 ( .B1(n4596), .B2(n4333), .A(n3342), .ZN(U3524) );
  NAND2_X1 U4180 ( .A1(n3318), .A2(n3343), .ZN(n3425) );
  NAND2_X1 U4181 ( .A1(n3425), .A2(n3344), .ZN(n3348) );
  INV_X1 U4182 ( .A(n3426), .ZN(n3346) );
  NOR2_X1 U4183 ( .A1(n3346), .A2(n3345), .ZN(n3347) );
  XNOR2_X1 U4184 ( .A(n3348), .B(n3347), .ZN(n3353) );
  INV_X1 U4185 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4976) );
  NOR2_X1 U4186 ( .A1(STATE_REG_SCAN_IN), .A2(n4976), .ZN(n4496) );
  OAI22_X1 U4187 ( .A1(n3349), .A2(n4430), .B1(n4429), .B2(n3376), .ZN(n3350)
         );
  AOI211_X1 U4188 ( .C1(n3366), .C2(n3752), .A(n4496), .B(n3350), .ZN(n3352)
         );
  NAND2_X1 U4189 ( .A1(n3812), .A2(n3401), .ZN(n3351) );
  OAI211_X1 U4190 ( .C1(n3353), .C2(n4418), .A(n3352), .B(n3351), .ZN(U3218)
         );
  AND2_X1 U4191 ( .A1(n3072), .A2(n3928), .ZN(n3857) );
  XNOR2_X1 U4192 ( .A(n3355), .B(n3857), .ZN(n4662) );
  INV_X1 U4193 ( .A(n3857), .ZN(n3356) );
  XNOR2_X1 U4194 ( .A(n3357), .B(n3356), .ZN(n3358) );
  NAND2_X1 U4195 ( .A1(n3358), .A2(n4197), .ZN(n3361) );
  AOI22_X1 U4196 ( .A1(n3359), .A2(n4142), .B1(n4287), .B2(n3432), .ZN(n3360)
         );
  OAI211_X1 U4197 ( .C1(n3430), .C2(n4195), .A(n3361), .B(n3360), .ZN(n4664)
         );
  NAND2_X1 U4198 ( .A1(n4664), .A2(n4273), .ZN(n3365) );
  AOI21_X1 U4199 ( .B1(n3432), .B2(n3369), .A(n3469), .ZN(n4665) );
  INV_X1 U4200 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3490) );
  INV_X1 U4201 ( .A(n3433), .ZN(n3362) );
  OAI22_X1 U4202 ( .A1(n4273), .A2(n3490), .B1(n3362), .B2(n4268), .ZN(n3363)
         );
  AOI21_X1 U4203 ( .B1(n4665), .B2(n4598), .A(n3363), .ZN(n3364) );
  OAI211_X1 U4204 ( .C1(n4662), .C2(n4275), .A(n3365), .B(n3364), .ZN(U3281)
         );
  NAND2_X1 U4205 ( .A1(n3367), .A2(n3366), .ZN(n3368) );
  NAND2_X1 U4206 ( .A1(n3369), .A2(n3368), .ZN(n3403) );
  INV_X1 U4207 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4208 ( .A1(n3371), .A2(n3370), .ZN(n3373) );
  AND2_X1 U4209 ( .A1(n3373), .A2(n3372), .ZN(n3374) );
  AND2_X1 U4210 ( .A1(n3927), .A2(n3922), .ZN(n3856) );
  XNOR2_X1 U4211 ( .A(n3374), .B(n3856), .ZN(n3405) );
  XNOR2_X1 U4212 ( .A(n3375), .B(n3856), .ZN(n3379) );
  OAI22_X1 U4213 ( .A1(n3376), .A2(n4256), .B1(n4255), .B2(n2336), .ZN(n3377)
         );
  AOI21_X1 U4214 ( .B1(n4260), .B2(n3988), .A(n3377), .ZN(n3378) );
  OAI21_X1 U4215 ( .B1(n3379), .B2(n4262), .A(n3378), .ZN(n3400) );
  AOI21_X1 U4216 ( .B1(n3405), .B2(n4656), .A(n3400), .ZN(n3382) );
  MUX2_X1 U4217 ( .A(n3380), .B(n3382), .S(n4673), .Z(n3381) );
  OAI21_X1 U4218 ( .B1(n3403), .B2(n4379), .A(n3381), .ZN(U3483) );
  INV_X1 U4219 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4812) );
  MUX2_X1 U4220 ( .A(n4812), .B(n3382), .S(n4684), .Z(n3383) );
  OAI21_X1 U4221 ( .B1(n3403), .B2(n4333), .A(n3383), .ZN(U3526) );
  INV_X1 U4222 ( .A(n3877), .ZN(n3384) );
  XNOR2_X1 U4223 ( .A(n3254), .B(n3384), .ZN(n4643) );
  INV_X1 U4224 ( .A(n3613), .ZN(n3633) );
  NAND2_X1 U4225 ( .A1(n4643), .A2(n3633), .ZN(n3393) );
  XNOR2_X1 U4226 ( .A(n3385), .B(n3877), .ZN(n3391) );
  OR2_X1 U4227 ( .A1(n3386), .A2(n4195), .ZN(n3389) );
  NAND2_X1 U4228 ( .A1(n3387), .A2(n4287), .ZN(n3388) );
  OAI211_X1 U4229 ( .C1(n3031), .C2(n4256), .A(n3389), .B(n3388), .ZN(n3390)
         );
  AOI21_X1 U4230 ( .B1(n3391), .B2(n4197), .A(n3390), .ZN(n3392) );
  AND2_X1 U4231 ( .A1(n3393), .A2(n3392), .ZN(n4645) );
  OR2_X1 U4232 ( .A1(n4636), .A2(n3394), .ZN(n3395) );
  NAND2_X1 U4233 ( .A1(n3396), .A2(n3395), .ZN(n4641) );
  AOI22_X1 U4234 ( .A1(n4604), .A2(REG2_REG_3__SCAN_IN), .B1(n4594), .B2(n2637), .ZN(n3397) );
  OAI21_X1 U4235 ( .B1(n4266), .B2(n4641), .A(n3397), .ZN(n3398) );
  AOI21_X1 U4236 ( .B1(n4643), .B2(n4599), .A(n3398), .ZN(n3399) );
  OAI21_X1 U4237 ( .B1(n4645), .B2(n4604), .A(n3399), .ZN(U3287) );
  INV_X1 U4238 ( .A(n3400), .ZN(n3407) );
  AOI22_X1 U4239 ( .A1(n4604), .A2(REG2_REG_8__SCAN_IN), .B1(n3401), .B2(n4594), .ZN(n3402) );
  OAI21_X1 U4240 ( .B1(n3403), .B2(n4266), .A(n3402), .ZN(n3404) );
  AOI21_X1 U4241 ( .B1(n3405), .B2(n4237), .A(n3404), .ZN(n3406) );
  OAI21_X1 U4242 ( .B1(n3407), .B2(n4604), .A(n3406), .ZN(U3282) );
  INV_X1 U4243 ( .A(n3408), .ZN(n3910) );
  AND2_X1 U4244 ( .A1(n3910), .A2(n3916), .ZN(n3884) );
  INV_X1 U4245 ( .A(n3884), .ZN(n3409) );
  XNOR2_X1 U4246 ( .A(n3410), .B(n3409), .ZN(n3414) );
  AOI22_X1 U4247 ( .A1(n3989), .A2(n4142), .B1(n4287), .B2(n3411), .ZN(n3412)
         );
  OAI21_X1 U4248 ( .B1(n3031), .B2(n4195), .A(n3412), .ZN(n3413) );
  AOI21_X1 U4249 ( .B1(n3414), .B2(n4197), .A(n3413), .ZN(n4652) );
  XNOR2_X1 U4250 ( .A(n3415), .B(n3884), .ZN(n4655) );
  INV_X1 U4251 ( .A(n3416), .ZN(n3417) );
  OAI21_X1 U4252 ( .B1(n2337), .B2(n3418), .A(n3417), .ZN(n4653) );
  NOR2_X1 U4253 ( .A1(n4653), .A2(n4266), .ZN(n3422) );
  OAI22_X1 U4254 ( .A1(n4273), .A2(n3420), .B1(n3419), .B2(n4268), .ZN(n3421)
         );
  AOI211_X1 U4255 ( .C1(n4655), .C2(n4237), .A(n3422), .B(n3421), .ZN(n3423)
         );
  OAI21_X1 U4256 ( .B1(n4604), .B2(n4652), .A(n3423), .ZN(U3285) );
  NAND2_X1 U4257 ( .A1(n3425), .A2(n3424), .ZN(n3427) );
  NAND2_X1 U4258 ( .A1(n3427), .A2(n3426), .ZN(n3428) );
  XOR2_X1 U4259 ( .A(n3429), .B(n3428), .Z(n3436) );
  AND2_X1 U4260 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4506) );
  OAI22_X1 U4261 ( .A1(n3430), .A2(n4430), .B1(n4429), .B2(n3519), .ZN(n3431)
         );
  AOI211_X1 U4262 ( .C1(n3432), .C2(n3752), .A(n4506), .B(n3431), .ZN(n3435)
         );
  NAND2_X1 U4263 ( .A1(n3812), .A2(n3433), .ZN(n3434) );
  OAI211_X1 U4264 ( .C1(n3436), .C2(n4418), .A(n3435), .B(n3434), .ZN(U3228)
         );
  INV_X1 U4265 ( .A(n3543), .ZN(n3542) );
  XNOR2_X1 U4266 ( .A(n3545), .B(n3542), .ZN(n3438) );
  XNOR2_X1 U4267 ( .A(n3437), .B(n3438), .ZN(n3443) );
  NOR2_X1 U4268 ( .A1(STATE_REG_SCAN_IN), .A2(n3439), .ZN(n3509) );
  OAI22_X1 U4269 ( .A1(n3519), .A2(n4430), .B1(n4429), .B2(n3609), .ZN(n3440)
         );
  AOI211_X1 U4270 ( .C1(n3517), .C2(n3752), .A(n3509), .B(n3440), .ZN(n3442)
         );
  NAND2_X1 U4271 ( .A1(n3812), .A2(n3525), .ZN(n3441) );
  OAI211_X1 U4272 ( .C1(n3443), .C2(n4418), .A(n3442), .B(n3441), .ZN(U3233)
         );
  NAND2_X1 U4273 ( .A1(n3444), .A2(n3878), .ZN(n3445) );
  NAND2_X1 U4274 ( .A1(n3446), .A2(n3445), .ZN(n4640) );
  INV_X1 U4275 ( .A(n4640), .ZN(n3462) );
  XNOR2_X1 U4276 ( .A(n3447), .B(n3065), .ZN(n3455) );
  NAND2_X1 U4277 ( .A1(n4640), .A2(n3633), .ZN(n3454) );
  AOI22_X1 U4278 ( .A1(n3449), .A2(n4142), .B1(n4287), .B2(n3448), .ZN(n3450)
         );
  OAI21_X1 U4279 ( .B1(n3451), .B2(n4195), .A(n3450), .ZN(n3452) );
  INV_X1 U4280 ( .A(n3452), .ZN(n3453) );
  OAI211_X1 U4281 ( .C1(n3455), .C2(n4262), .A(n3454), .B(n3453), .ZN(n4638)
         );
  MUX2_X1 U4282 ( .A(n4638), .B(REG2_REG_2__SCAN_IN), .S(n4604), .Z(n3456) );
  INV_X1 U4283 ( .A(n3456), .ZN(n3461) );
  NOR2_X1 U4284 ( .A1(n3458), .A2(n3457), .ZN(n4637) );
  NOR3_X1 U4285 ( .A1(n4266), .A2(n4636), .A3(n4637), .ZN(n3459) );
  AOI21_X1 U4286 ( .B1(n4594), .B2(REG3_REG_2__SCAN_IN), .A(n3459), .ZN(n3460)
         );
  OAI211_X1 U4287 ( .C1(n3462), .C2(n3641), .A(n3461), .B(n3460), .ZN(U3288)
         );
  AND2_X1 U4288 ( .A1(n3932), .A2(n3934), .ZN(n3858) );
  XOR2_X1 U4289 ( .A(n3858), .B(n3463), .Z(n3467) );
  OAI22_X1 U4290 ( .A1(n3464), .A2(n4256), .B1(n4255), .B2(n3477), .ZN(n3465)
         );
  AOI21_X1 U4291 ( .B1(n4260), .B2(n3987), .A(n3465), .ZN(n3466) );
  OAI21_X1 U4292 ( .B1(n3467), .B2(n4262), .A(n3466), .ZN(n3553) );
  INV_X1 U4293 ( .A(n3553), .ZN(n3474) );
  XNOR2_X1 U4294 ( .A(n3468), .B(n3858), .ZN(n3554) );
  NOR2_X1 U4295 ( .A1(n3469), .A2(n3477), .ZN(n3470) );
  OR2_X1 U4296 ( .A1(n3524), .A2(n3470), .ZN(n3559) );
  AOI22_X1 U4297 ( .A1(n4604), .A2(REG2_REG_10__SCAN_IN), .B1(n3484), .B2(
        n4594), .ZN(n3471) );
  OAI21_X1 U4298 ( .B1(n3559), .B2(n4266), .A(n3471), .ZN(n3472) );
  AOI21_X1 U4299 ( .B1(n3554), .B2(n4237), .A(n3472), .ZN(n3473) );
  OAI21_X1 U4300 ( .B1(n3474), .B2(n4604), .A(n3473), .ZN(U3280) );
  AOI22_X1 U4301 ( .A1(n3755), .A2(n3987), .B1(n3754), .B2(n3986), .ZN(n3476)
         );
  NOR2_X1 U4302 ( .A1(n4892), .A2(STATE_REG_SCAN_IN), .ZN(n4516) );
  INV_X1 U4303 ( .A(n4516), .ZN(n3475) );
  OAI211_X1 U4304 ( .C1(n4433), .C2(n3477), .A(n3476), .B(n3475), .ZN(n3483)
         );
  INV_X1 U4305 ( .A(n3478), .ZN(n3479) );
  AOI211_X1 U4306 ( .C1(n3481), .C2(n3480), .A(n4418), .B(n3479), .ZN(n3482)
         );
  AOI211_X1 U4307 ( .C1(n3484), .C2(n3812), .A(n3483), .B(n3482), .ZN(n3485)
         );
  INV_X1 U4308 ( .A(n3485), .ZN(U3214) );
  INV_X1 U4309 ( .A(n4394), .ZN(n3581) );
  NAND2_X1 U4310 ( .A1(n4395), .A2(REG2_REG_7__SCAN_IN), .ZN(n3487) );
  NAND2_X1 U4311 ( .A1(n4621), .A2(n3488), .ZN(n3489) );
  INV_X1 U4312 ( .A(n4621), .ZN(n4502) );
  XNOR2_X1 U4313 ( .A(n3488), .B(n4502), .ZN(n4499) );
  NAND2_X1 U4314 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4499), .ZN(n4498) );
  INV_X1 U4315 ( .A(n3501), .ZN(n4620) );
  AOI22_X1 U4316 ( .A1(n3501), .A2(REG2_REG_9__SCAN_IN), .B1(n3490), .B2(n4620), .ZN(n4510) );
  NAND2_X1 U4317 ( .A1(n3501), .A2(REG2_REG_9__SCAN_IN), .ZN(n3491) );
  INV_X1 U4318 ( .A(n4617), .ZN(n4522) );
  NAND2_X1 U4319 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4519), .ZN(n4518) );
  NAND2_X1 U4320 ( .A1(n4617), .A2(n3492), .ZN(n3493) );
  INV_X1 U4321 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3494) );
  MUX2_X1 U4322 ( .A(REG2_REG_11__SCAN_IN), .B(n3494), .S(n4394), .Z(n3495) );
  NAND2_X1 U4323 ( .A1(n3496), .A2(n3495), .ZN(n3580) );
  OAI211_X1 U4324 ( .C1(n3496), .C2(n3495), .A(n3580), .B(n4588), .ZN(n3511)
         );
  INV_X1 U4325 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4515) );
  NOR2_X1 U4326 ( .A1(n4502), .A2(n3498), .ZN(n3499) );
  XOR2_X1 U4327 ( .A(n4621), .B(n3498), .Z(n4495) );
  NOR2_X1 U4328 ( .A1(n4812), .A2(n4495), .ZN(n4494) );
  NOR2_X1 U4329 ( .A1(n3499), .A2(n4494), .ZN(n4505) );
  NAND2_X1 U4330 ( .A1(n3501), .A2(REG1_REG_9__SCAN_IN), .ZN(n3500) );
  OAI21_X1 U4331 ( .B1(n3501), .B2(REG1_REG_9__SCAN_IN), .A(n3500), .ZN(n4504)
         );
  NOR2_X1 U4332 ( .A1(n4505), .A2(n4504), .ZN(n4503) );
  NOR2_X1 U4333 ( .A1(n3502), .A2(n4522), .ZN(n3503) );
  INV_X1 U4334 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3504) );
  MUX2_X1 U4335 ( .A(n3504), .B(REG1_REG_11__SCAN_IN), .S(n4394), .Z(n3506) );
  INV_X1 U4336 ( .A(n3576), .ZN(n3505) );
  AOI211_X1 U4337 ( .C1(n3507), .C2(n3506), .A(n3505), .B(n4583), .ZN(n3508)
         );
  AOI211_X1 U4338 ( .C1(n4581), .C2(ADDR_REG_11__SCAN_IN), .A(n3509), .B(n3508), .ZN(n3510) );
  OAI211_X1 U4339 ( .C1(n4593), .C2(n3581), .A(n3511), .B(n3510), .ZN(U3251)
         );
  NAND2_X1 U4340 ( .A1(n3513), .A2(n3512), .ZN(n3515) );
  INV_X1 U4341 ( .A(n3514), .ZN(n3885) );
  XNOR2_X1 U4342 ( .A(n3515), .B(n3885), .ZN(n4669) );
  XNOR2_X1 U4343 ( .A(n3516), .B(n3885), .ZN(n3521) );
  AOI22_X1 U4344 ( .A1(n3985), .A2(n4142), .B1(n4287), .B2(n3517), .ZN(n3518)
         );
  OAI21_X1 U4345 ( .B1(n3519), .B2(n4195), .A(n3518), .ZN(n3520) );
  AOI21_X1 U4346 ( .B1(n3521), .B2(n4197), .A(n3520), .ZN(n3522) );
  OAI21_X1 U4347 ( .B1(n4669), .B2(n3613), .A(n3522), .ZN(n4671) );
  INV_X1 U4348 ( .A(n4671), .ZN(n3530) );
  INV_X1 U4349 ( .A(n4669), .ZN(n3528) );
  OAI21_X1 U4350 ( .B1(n3524), .B2(n3523), .A(n3568), .ZN(n4667) );
  AOI22_X1 U4351 ( .A1(n4604), .A2(REG2_REG_11__SCAN_IN), .B1(n3525), .B2(
        n4594), .ZN(n3526) );
  OAI21_X1 U4352 ( .B1(n4667), .B2(n4266), .A(n3526), .ZN(n3527) );
  AOI21_X1 U4353 ( .B1(n3528), .B2(n4599), .A(n3527), .ZN(n3529) );
  OAI21_X1 U4354 ( .B1(n3530), .B2(n4604), .A(n3529), .ZN(U3279) );
  XOR2_X1 U4355 ( .A(n3532), .B(n3531), .Z(n3533) );
  XNOR2_X1 U4356 ( .A(n3534), .B(n3533), .ZN(n3539) );
  INV_X1 U4357 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3535) );
  NOR2_X1 U4358 ( .A1(STATE_REG_SCAN_IN), .A2(n3535), .ZN(n4526) );
  OAI22_X1 U4359 ( .A1(n3609), .A2(n4430), .B1(n4429), .B2(n4431), .ZN(n3536)
         );
  AOI211_X1 U4360 ( .C1(n3615), .C2(n3752), .A(n4526), .B(n3536), .ZN(n3538)
         );
  NAND2_X1 U4361 ( .A1(n3812), .A2(n3618), .ZN(n3537) );
  OAI211_X1 U4362 ( .C1(n3539), .C2(n4418), .A(n3538), .B(n3537), .ZN(U3231)
         );
  NAND2_X1 U4363 ( .A1(n3541), .A2(n3540), .ZN(n3548) );
  NOR2_X1 U4364 ( .A1(n3437), .A2(n3542), .ZN(n3546) );
  INV_X1 U4365 ( .A(n3437), .ZN(n3544) );
  OAI22_X1 U4366 ( .A1(n3546), .A2(n3545), .B1(n3544), .B2(n3543), .ZN(n3547)
         );
  XOR2_X1 U4367 ( .A(n3548), .B(n3547), .Z(n3552) );
  AOI22_X1 U4368 ( .A1(n3755), .A2(n3986), .B1(n3754), .B2(n3984), .ZN(n3549)
         );
  NAND2_X1 U4369 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n3583) );
  OAI211_X1 U4370 ( .C1(n4433), .C2(n3562), .A(n3549), .B(n3583), .ZN(n3550)
         );
  AOI21_X1 U4371 ( .B1(n3570), .B2(n3812), .A(n3550), .ZN(n3551) );
  OAI21_X1 U4372 ( .B1(n3552), .B2(n4418), .A(n3551), .ZN(U3221) );
  INV_X1 U4373 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3555) );
  AOI21_X1 U4374 ( .B1(n3554), .B2(n4656), .A(n3553), .ZN(n3557) );
  MUX2_X1 U4375 ( .A(n3555), .B(n3557), .S(n4673), .Z(n3556) );
  OAI21_X1 U4376 ( .B1(n3559), .B2(n4379), .A(n3556), .ZN(U3487) );
  MUX2_X1 U4377 ( .A(n4515), .B(n3557), .S(n4684), .Z(n3558) );
  OAI21_X1 U4378 ( .B1(n3559), .B2(n4333), .A(n3558), .ZN(U3528) );
  INV_X1 U4379 ( .A(n3605), .ZN(n3560) );
  OR2_X1 U4380 ( .A1(n3560), .A2(n3892), .ZN(n3883) );
  XNOR2_X1 U4381 ( .A(n3561), .B(n3883), .ZN(n3565) );
  OAI22_X1 U4382 ( .A1(n3631), .A2(n4256), .B1(n4255), .B2(n3562), .ZN(n3563)
         );
  AOI21_X1 U4383 ( .B1(n4260), .B2(n3986), .A(n3563), .ZN(n3564) );
  OAI21_X1 U4384 ( .B1(n3565), .B2(n4262), .A(n3564), .ZN(n3596) );
  INV_X1 U4385 ( .A(n3596), .ZN(n3574) );
  XNOR2_X1 U4386 ( .A(n3566), .B(n3883), .ZN(n3597) );
  NAND2_X1 U4387 ( .A1(n3568), .A2(n3567), .ZN(n3569) );
  NAND2_X1 U4388 ( .A1(n3616), .A2(n3569), .ZN(n3602) );
  AOI22_X1 U4389 ( .A1(n4604), .A2(REG2_REG_12__SCAN_IN), .B1(n3570), .B2(
        n4594), .ZN(n3571) );
  OAI21_X1 U4390 ( .B1(n3602), .B2(n4266), .A(n3571), .ZN(n3572) );
  AOI21_X1 U4391 ( .B1(n3597), .B2(n4237), .A(n3572), .ZN(n3573) );
  OAI21_X1 U4392 ( .B1(n3574), .B2(n4604), .A(n3573), .ZN(U3278) );
  INV_X1 U4393 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U4394 ( .A1(n4394), .A2(REG1_REG_11__SCAN_IN), .ZN(n3575) );
  OR2_X1 U4395 ( .A1(n3577), .A2(n4393), .ZN(n3578) );
  AOI211_X1 U4396 ( .C1(n4879), .C2(n3579), .A(n2260), .B(n4583), .ZN(n3588)
         );
  OAI211_X1 U4397 ( .C1(n3582), .C2(REG2_REG_12__SCAN_IN), .A(n4588), .B(n4041), .ZN(n3586) );
  INV_X1 U4398 ( .A(n3583), .ZN(n3584) );
  AOI21_X1 U4399 ( .B1(n4581), .B2(ADDR_REG_12__SCAN_IN), .A(n3584), .ZN(n3585) );
  OAI211_X1 U4400 ( .C1(n4593), .C2(n2278), .A(n3586), .B(n3585), .ZN(n3587)
         );
  OR2_X1 U4401 ( .A1(n3588), .A2(n3587), .ZN(U3252) );
  NOR2_X1 U4402 ( .A1(n2269), .A2(n3590), .ZN(n3591) );
  XNOR2_X1 U4403 ( .A(n3589), .B(n3591), .ZN(n3595) );
  AOI22_X1 U4404 ( .A1(n3755), .A2(n3984), .B1(n3754), .B2(n3982), .ZN(n3592)
         );
  NAND2_X1 U4405 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4544) );
  OAI211_X1 U4406 ( .C1(n4433), .C2(n3637), .A(n3592), .B(n4544), .ZN(n3593)
         );
  AOI21_X1 U4407 ( .B1(n3635), .B2(n3812), .A(n3593), .ZN(n3594) );
  OAI21_X1 U4408 ( .B1(n3595), .B2(n4418), .A(n3594), .ZN(U3212) );
  AOI21_X1 U4409 ( .B1(n4656), .B2(n3597), .A(n3596), .ZN(n3599) );
  MUX2_X1 U4410 ( .A(n4879), .B(n3599), .S(n4684), .Z(n3598) );
  OAI21_X1 U4411 ( .B1(n3602), .B2(n4333), .A(n3598), .ZN(U3530) );
  INV_X1 U4412 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3600) );
  MUX2_X1 U4413 ( .A(n3600), .B(n3599), .S(n4673), .Z(n3601) );
  OAI21_X1 U4414 ( .B1(n3602), .B2(n4379), .A(n3601), .ZN(U3491) );
  NAND2_X1 U4415 ( .A1(n3894), .A2(n3604), .ZN(n3871) );
  XNOR2_X1 U4416 ( .A(n3603), .B(n3871), .ZN(n3614) );
  NAND2_X1 U4417 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  XNOR2_X1 U4418 ( .A(n3607), .B(n3871), .ZN(n3611) );
  AOI22_X1 U4419 ( .A1(n3983), .A2(n4142), .B1(n4287), .B2(n3615), .ZN(n3608)
         );
  OAI21_X1 U4420 ( .B1(n3609), .B2(n4195), .A(n3608), .ZN(n3610) );
  AOI21_X1 U4421 ( .B1(n3611), .B2(n4197), .A(n3610), .ZN(n3612) );
  OAI21_X1 U4422 ( .B1(n3614), .B2(n3613), .A(n3612), .ZN(n3644) );
  INV_X1 U4423 ( .A(n3644), .ZN(n3622) );
  INV_X1 U4424 ( .A(n3614), .ZN(n3645) );
  AND2_X1 U4425 ( .A1(n3616), .A2(n3615), .ZN(n3617) );
  OR2_X1 U4426 ( .A1(n3638), .A2(n3617), .ZN(n3650) );
  AOI22_X1 U4427 ( .A1(n4604), .A2(REG2_REG_13__SCAN_IN), .B1(n3618), .B2(
        n4594), .ZN(n3619) );
  OAI21_X1 U4428 ( .B1(n3650), .B2(n4266), .A(n3619), .ZN(n3620) );
  AOI21_X1 U4429 ( .B1(n3645), .B2(n4599), .A(n3620), .ZN(n3621) );
  OAI21_X1 U4430 ( .B1(n3622), .B2(n4604), .A(n3621), .ZN(U3277) );
  OAI21_X1 U4431 ( .B1(n3625), .B2(n3624), .A(n3623), .ZN(n3634) );
  OAI21_X1 U4432 ( .B1(n3876), .B2(n3626), .A(n3652), .ZN(n3627) );
  NAND2_X1 U4433 ( .A1(n3627), .A2(n4197), .ZN(n3630) );
  AOI22_X1 U4434 ( .A1(n3982), .A2(n4142), .B1(n4287), .B2(n3628), .ZN(n3629)
         );
  OAI211_X1 U4435 ( .C1(n3631), .C2(n4195), .A(n3630), .B(n3629), .ZN(n3632)
         );
  AOI21_X1 U4436 ( .B1(n3634), .B2(n3633), .A(n3632), .ZN(n4351) );
  INV_X1 U4437 ( .A(n3634), .ZN(n4352) );
  AOI22_X1 U4438 ( .A1(n4604), .A2(REG2_REG_14__SCAN_IN), .B1(n3635), .B2(
        n4594), .ZN(n3640) );
  OR2_X1 U4439 ( .A1(n3638), .A2(n3637), .ZN(n4349) );
  NAND3_X1 U4440 ( .A1(n3636), .A2(n4349), .A3(n4598), .ZN(n3639) );
  OAI211_X1 U4441 ( .C1(n4352), .C2(n3641), .A(n3640), .B(n3639), .ZN(n3642)
         );
  INV_X1 U4442 ( .A(n3642), .ZN(n3643) );
  OAI21_X1 U4443 ( .B1(n4604), .B2(n4351), .A(n3643), .ZN(U3276) );
  INV_X1 U4444 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3646) );
  AOI21_X1 U4445 ( .B1(n4649), .B2(n3645), .A(n3644), .ZN(n3648) );
  MUX2_X1 U4446 ( .A(n3646), .B(n3648), .S(n4673), .Z(n3647) );
  OAI21_X1 U4447 ( .B1(n3650), .B2(n4379), .A(n3647), .ZN(U3493) );
  INV_X1 U4448 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4023) );
  MUX2_X1 U4449 ( .A(n4023), .B(n3648), .S(n4684), .Z(n3649) );
  OAI21_X1 U4450 ( .B1(n4333), .B2(n3650), .A(n3649), .ZN(U3531) );
  XNOR2_X1 U4451 ( .A(n3651), .B(n3873), .ZN(n3679) );
  INV_X1 U4452 ( .A(n3679), .ZN(n3664) );
  INV_X1 U4453 ( .A(n3652), .ZN(n3653) );
  OAI21_X1 U4454 ( .B1(n3653), .B2(n3822), .A(n3873), .ZN(n3655) );
  NAND3_X1 U4455 ( .A1(n3655), .A2(n4197), .A3(n3654), .ZN(n3658) );
  OAI22_X1 U4456 ( .A1(n4428), .A2(n4256), .B1(n4255), .B2(n4432), .ZN(n3656)
         );
  INV_X1 U4457 ( .A(n3656), .ZN(n3657) );
  OAI211_X1 U4458 ( .C1(n4431), .C2(n4195), .A(n3658), .B(n3657), .ZN(n3678)
         );
  INV_X1 U4459 ( .A(n3636), .ZN(n3659) );
  OAI21_X1 U4460 ( .B1(n3659), .B2(n4432), .A(n3673), .ZN(n3683) );
  NOR2_X1 U4461 ( .A1(n3683), .A2(n4266), .ZN(n3662) );
  INV_X1 U4462 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3660) );
  OAI22_X1 U4463 ( .A1(n4273), .A2(n3660), .B1(n4445), .B2(n4268), .ZN(n3661)
         );
  AOI211_X1 U4464 ( .C1(n3678), .C2(n4273), .A(n3662), .B(n3661), .ZN(n3663)
         );
  OAI21_X1 U4465 ( .B1(n3664), .B2(n4275), .A(n3663), .ZN(U3275) );
  OAI21_X1 U4466 ( .B1(n3667), .B2(n3666), .A(n3665), .ZN(n4348) );
  OAI211_X1 U4467 ( .C1(n3669), .C2(n3851), .A(n3668), .B(n4197), .ZN(n3671)
         );
  AOI22_X1 U4468 ( .A1(n3981), .A2(n4142), .B1(n3672), .B2(n4287), .ZN(n3670)
         );
  OAI211_X1 U4469 ( .C1(n4397), .C2(n4195), .A(n3671), .B(n3670), .ZN(n4343)
         );
  NAND2_X1 U4470 ( .A1(n3673), .A2(n3672), .ZN(n4344) );
  AND3_X1 U4471 ( .A1(n4345), .A2(n4598), .A3(n4344), .ZN(n3676) );
  INV_X1 U4472 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3674) );
  OAI22_X1 U4473 ( .A1(n4273), .A2(n3674), .B1(n4409), .B2(n4268), .ZN(n3675)
         );
  AOI211_X1 U4474 ( .C1(n4343), .C2(n4273), .A(n3676), .B(n3675), .ZN(n3677)
         );
  OAI21_X1 U4475 ( .B1(n4348), .B2(n4275), .A(n3677), .ZN(U3274) );
  INV_X1 U4476 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4977) );
  AOI21_X1 U4477 ( .B1(n3679), .B2(n4656), .A(n3678), .ZN(n3681) );
  MUX2_X1 U4478 ( .A(n4977), .B(n3681), .S(n4673), .Z(n3680) );
  OAI21_X1 U4479 ( .B1(n3683), .B2(n4379), .A(n3680), .ZN(U3497) );
  INV_X1 U4480 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4029) );
  MUX2_X1 U4481 ( .A(n4029), .B(n3681), .S(n4684), .Z(n3682) );
  OAI21_X1 U4482 ( .B1(n4333), .B2(n3683), .A(n3682), .ZN(U3533) );
  AOI21_X1 U4483 ( .B1(n3684), .B2(n3697), .A(n3698), .ZN(n4252) );
  XNOR2_X1 U4484 ( .A(n4252), .B(n3689), .ZN(n3687) );
  AOI22_X1 U4485 ( .A1(n4234), .A2(n4142), .B1(n2342), .B2(n4287), .ZN(n3685)
         );
  OAI21_X1 U4486 ( .B1(n4421), .B2(n4195), .A(n3685), .ZN(n3686) );
  AOI21_X1 U4487 ( .B1(n3687), .B2(n4197), .A(n3686), .ZN(n4336) );
  OAI21_X1 U4488 ( .B1(n3690), .B2(n3689), .A(n3688), .ZN(n4334) );
  XNOR2_X1 U4489 ( .A(n3705), .B(n2342), .ZN(n3691) );
  NAND2_X1 U4490 ( .A1(n3691), .A2(n2598), .ZN(n4335) );
  AOI22_X1 U4491 ( .A1(n4604), .A2(REG2_REG_18__SCAN_IN), .B1(n3692), .B2(
        n4594), .ZN(n3693) );
  OAI21_X1 U4492 ( .B1(n4335), .B2(n3694), .A(n3693), .ZN(n3695) );
  AOI21_X1 U4493 ( .B1(n4334), .B2(n4237), .A(n3695), .ZN(n3696) );
  OAI21_X1 U4494 ( .B1(n4604), .B2(n4336), .A(n3696), .ZN(U3272) );
  INV_X1 U4495 ( .A(n3697), .ZN(n3699) );
  OR2_X1 U4496 ( .A1(n3699), .A2(n3698), .ZN(n3859) );
  XNOR2_X1 U4497 ( .A(n3700), .B(n3859), .ZN(n4342) );
  XNOR2_X1 U4498 ( .A(n3701), .B(n3859), .ZN(n3704) );
  AOI22_X1 U4499 ( .A1(n4259), .A2(n4142), .B1(n4287), .B2(n3717), .ZN(n3702)
         );
  OAI21_X1 U4500 ( .B1(n4428), .B2(n4195), .A(n3702), .ZN(n3703) );
  AOI21_X1 U4501 ( .B1(n3704), .B2(n4197), .A(n3703), .ZN(n4341) );
  AOI22_X1 U4502 ( .A1(n4604), .A2(REG2_REG_17__SCAN_IN), .B1(n3718), .B2(
        n4594), .ZN(n3707) );
  INV_X1 U4503 ( .A(n3705), .ZN(n4339) );
  NAND2_X1 U4504 ( .A1(n4345), .A2(n3717), .ZN(n4338) );
  NAND3_X1 U4505 ( .A1(n4339), .A2(n4598), .A3(n4338), .ZN(n3706) );
  OAI211_X1 U4506 ( .C1(n4341), .C2(n4604), .A(n3707), .B(n3706), .ZN(n3708)
         );
  INV_X1 U4507 ( .A(n3708), .ZN(n3709) );
  OAI21_X1 U4508 ( .B1(n4342), .B2(n4275), .A(n3709), .ZN(U3273) );
  INV_X1 U4509 ( .A(n3711), .ZN(n3712) );
  NOR2_X1 U4510 ( .A1(n3713), .A2(n3712), .ZN(n3714) );
  XNOR2_X1 U4511 ( .A(n3710), .B(n3714), .ZN(n3721) );
  AND2_X1 U4512 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4569) );
  INV_X1 U4513 ( .A(n4259), .ZN(n3715) );
  OAI22_X1 U4514 ( .A1(n4428), .A2(n4430), .B1(n4429), .B2(n3715), .ZN(n3716)
         );
  AOI211_X1 U4515 ( .C1(n3717), .C2(n3752), .A(n4569), .B(n3716), .ZN(n3720)
         );
  NAND2_X1 U4516 ( .A1(n3812), .A2(n3718), .ZN(n3719) );
  OAI211_X1 U4517 ( .C1(n3721), .C2(n4418), .A(n3720), .B(n3719), .ZN(U3225)
         );
  XOR2_X1 U4518 ( .A(n3723), .B(n3722), .Z(n3727) );
  AOI22_X1 U4519 ( .A1(n3755), .A2(n4259), .B1(n3754), .B2(n4222), .ZN(n3724)
         );
  NAND2_X1 U4520 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4057) );
  OAI211_X1 U4521 ( .C1(n4433), .C2(n4264), .A(n3724), .B(n4057), .ZN(n3725)
         );
  AOI21_X1 U4522 ( .B1(n4267), .B2(n3812), .A(n3725), .ZN(n3726) );
  OAI21_X1 U4523 ( .B1(n3727), .B2(n4418), .A(n3726), .ZN(U3216) );
  INV_X1 U4524 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3731) );
  INV_X1 U4525 ( .A(n4379), .ZN(n3728) );
  NAND2_X1 U4526 ( .A1(n4278), .A2(n3728), .ZN(n3730) );
  NAND2_X1 U4527 ( .A1(n4279), .A2(n4673), .ZN(n3729) );
  OAI211_X1 U4528 ( .C1(n4673), .C2(n3731), .A(n3730), .B(n3729), .ZN(U3517)
         );
  XNOR2_X1 U4529 ( .A(n3733), .B(n3732), .ZN(n3738) );
  INV_X1 U4530 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4967) );
  OAI22_X1 U4531 ( .A1(n4433), .A2(n4106), .B1(STATE_REG_SCAN_IN), .B2(n4967), 
        .ZN(n3735) );
  OAI22_X1 U4532 ( .A1(n4098), .A2(n4430), .B1(n4429), .B2(n4099), .ZN(n3734)
         );
  AOI211_X1 U4533 ( .C1(n3736), .C2(n3812), .A(n3735), .B(n3734), .ZN(n3737)
         );
  OAI21_X1 U4534 ( .B1(n3738), .B2(n4418), .A(n3737), .ZN(U3211) );
  INV_X1 U4535 ( .A(n3739), .ZN(n3740) );
  NAND2_X1 U4536 ( .A1(n3740), .A2(n4441), .ZN(n3747) );
  AOI21_X1 U4537 ( .B1(n3797), .B2(n3742), .A(n3741), .ZN(n3746) );
  INV_X1 U4538 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4946) );
  OAI22_X1 U4539 ( .A1(n4433), .A2(n4179), .B1(STATE_REG_SCAN_IN), .B2(n4946), 
        .ZN(n3744) );
  OAI22_X1 U4540 ( .A1(n4215), .A2(n4430), .B1(n4429), .B2(n4173), .ZN(n3743)
         );
  AOI211_X1 U4541 ( .C1(n4180), .C2(n3812), .A(n3744), .B(n3743), .ZN(n3745)
         );
  OAI21_X1 U4542 ( .B1(n3747), .B2(n3746), .A(n3745), .ZN(U3213) );
  AOI21_X1 U4543 ( .B1(n3749), .B2(n3748), .A(n4418), .ZN(n3751) );
  NAND2_X1 U4544 ( .A1(n3751), .A2(n3750), .ZN(n3759) );
  AOI22_X1 U4545 ( .A1(n3754), .A2(n3753), .B1(n3752), .B2(n2231), .ZN(n3758)
         );
  AOI22_X1 U4546 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3756), .B1(n3755), .B2(n2608), .ZN(n3757) );
  NAND3_X1 U4547 ( .A1(n3759), .A2(n3758), .A3(n3757), .ZN(U3219) );
  XNOR2_X1 U4548 ( .A(n3762), .B(n3761), .ZN(n3763) );
  XNOR2_X1 U4549 ( .A(n3760), .B(n3763), .ZN(n3768) );
  INV_X1 U4550 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3764) );
  OAI22_X1 U4551 ( .A1(n4433), .A2(n4214), .B1(STATE_REG_SCAN_IN), .B2(n3764), 
        .ZN(n3766) );
  OAI22_X1 U4552 ( .A1(n4257), .A2(n4430), .B1(n4429), .B2(n4215), .ZN(n3765)
         );
  AOI211_X1 U4553 ( .C1(n4211), .C2(n3812), .A(n3766), .B(n3765), .ZN(n3767)
         );
  OAI21_X1 U4554 ( .B1(n3768), .B2(n4418), .A(n3767), .ZN(U3220) );
  INV_X1 U4555 ( .A(n3770), .ZN(n3771) );
  NOR2_X1 U4556 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  XNOR2_X1 U4557 ( .A(n3769), .B(n3773), .ZN(n3778) );
  OAI22_X1 U4558 ( .A1(n4433), .A2(n3061), .B1(STATE_REG_SCAN_IN), .B2(n3774), 
        .ZN(n3776) );
  OAI22_X1 U4559 ( .A1(n4173), .A2(n4430), .B1(n4429), .B2(n4098), .ZN(n3775)
         );
  AOI211_X1 U4560 ( .C1(n4134), .C2(n3812), .A(n3776), .B(n3775), .ZN(n3777)
         );
  OAI21_X1 U4561 ( .B1(n3778), .B2(n4418), .A(n3777), .ZN(U3222) );
  NAND2_X1 U4562 ( .A1(n3779), .A2(n2247), .ZN(n3781) );
  XNOR2_X1 U4563 ( .A(n3781), .B(n3780), .ZN(n3786) );
  OAI22_X1 U4564 ( .A1(n4433), .A2(n4161), .B1(STATE_REG_SCAN_IN), .B2(n3782), 
        .ZN(n3784) );
  OAI22_X1 U4565 ( .A1(n4191), .A2(n4430), .B1(n4429), .B2(n4155), .ZN(n3783)
         );
  AOI211_X1 U4566 ( .C1(n4163), .C2(n3812), .A(n3784), .B(n3783), .ZN(n3785)
         );
  OAI21_X1 U4567 ( .B1(n3786), .B2(n4418), .A(n3785), .ZN(U3226) );
  OR2_X1 U4568 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  AOI22_X1 U4569 ( .A1(n3787), .A2(n2309), .B1(n3791), .B2(n3790), .ZN(n3796)
         );
  INV_X1 U4570 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4932) );
  OAI22_X1 U4571 ( .A1(n4433), .A2(n4226), .B1(STATE_REG_SCAN_IN), .B2(n4932), 
        .ZN(n3793) );
  OAI22_X1 U4572 ( .A1(n4410), .A2(n4430), .B1(n4429), .B2(n4227), .ZN(n3792)
         );
  AOI211_X1 U4573 ( .C1(n3794), .C2(n3812), .A(n3793), .B(n3792), .ZN(n3795)
         );
  OAI21_X1 U4574 ( .B1(n3796), .B2(n4418), .A(n3795), .ZN(U3230) );
  OAI21_X1 U4575 ( .B1(n3799), .B2(n3798), .A(n3797), .ZN(n3800) );
  NAND2_X1 U4576 ( .A1(n3800), .A2(n4441), .ZN(n3804) );
  NOR2_X1 U4577 ( .A1(n4433), .A2(n4202), .ZN(n3802) );
  OAI22_X1 U4578 ( .A1(n4191), .A2(n4429), .B1(n4430), .B2(n4227), .ZN(n3801)
         );
  AOI211_X1 U4579 ( .C1(REG3_REG_22__SCAN_IN), .C2(U3149), .A(n3802), .B(n3801), .ZN(n3803) );
  OAI211_X1 U4580 ( .C1(n4446), .C2(n4199), .A(n3804), .B(n3803), .ZN(U3232)
         );
  INV_X1 U4581 ( .A(n3806), .ZN(n3808) );
  NAND2_X1 U4582 ( .A1(n3808), .A2(n3807), .ZN(n3809) );
  XNOR2_X1 U4583 ( .A(n3805), .B(n3809), .ZN(n3814) );
  OAI22_X1 U4584 ( .A1(n4433), .A2(n4126), .B1(STATE_REG_SCAN_IN), .B2(n5043), 
        .ZN(n3811) );
  OAI22_X1 U4585 ( .A1(n4155), .A2(n4430), .B1(n4429), .B2(n4118), .ZN(n3810)
         );
  AOI211_X1 U4586 ( .C1(n4127), .C2(n3812), .A(n3811), .B(n3810), .ZN(n3813)
         );
  OAI21_X1 U4587 ( .B1(n3814), .B2(n4418), .A(n3813), .ZN(U3237) );
  NAND2_X1 U4588 ( .A1(n4063), .A2(n3815), .ZN(n3835) );
  INV_X1 U4589 ( .A(n3835), .ZN(n3818) );
  OR2_X1 U4590 ( .A1(n3817), .A2(n4068), .ZN(n3848) );
  NAND2_X1 U4591 ( .A1(n3848), .A2(n4065), .ZN(n3961) );
  OR2_X1 U4592 ( .A1(n4070), .A2(n3820), .ZN(n3816) );
  NAND2_X1 U4593 ( .A1(n3839), .A2(n3965), .ZN(n3843) );
  AND2_X1 U4594 ( .A1(n3816), .A2(n3843), .ZN(n3874) );
  NAND2_X1 U4595 ( .A1(n3817), .A2(n4068), .ZN(n3847) );
  OAI211_X1 U4596 ( .C1(n3818), .C2(n3961), .A(n3874), .B(n3847), .ZN(n3819)
         );
  INV_X1 U4597 ( .A(n3819), .ZN(n3971) );
  NAND2_X1 U4598 ( .A1(n4070), .A2(n3820), .ZN(n3841) );
  INV_X1 U4599 ( .A(n3949), .ZN(n3833) );
  INV_X1 U4600 ( .A(n3946), .ZN(n3830) );
  INV_X1 U4601 ( .A(n3893), .ZN(n3821) );
  NOR4_X1 U4602 ( .A1(n3626), .A2(n3825), .A3(n3822), .A4(n3821), .ZN(n3827)
         );
  NAND2_X1 U4603 ( .A1(n3824), .A2(n3823), .ZN(n3926) );
  NAND2_X1 U4604 ( .A1(n3926), .A2(n3893), .ZN(n3940) );
  NOR2_X1 U4605 ( .A1(n3940), .A2(n3825), .ZN(n3826) );
  NOR4_X1 U4606 ( .A1(n3827), .A2(n3942), .A3(n3826), .A4(n3941), .ZN(n3828)
         );
  NOR2_X1 U4607 ( .A1(n3828), .A2(n3947), .ZN(n3829) );
  OAI21_X1 U4608 ( .B1(n3830), .B2(n3829), .A(n3951), .ZN(n3831) );
  OAI221_X1 U4609 ( .B1(n3833), .B2(n3832), .C1(n3833), .C2(n3831), .A(n3955), 
        .ZN(n3838) );
  INV_X1 U4610 ( .A(n3847), .ZN(n3834) );
  NOR2_X1 U4611 ( .A1(n3835), .A2(n3834), .ZN(n3836) );
  NAND4_X1 U4612 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3874), .ZN(n3840)
         );
  OR2_X1 U4613 ( .A1(n3839), .A2(n3965), .ZN(n3842) );
  OAI211_X1 U4614 ( .C1(n3965), .C2(n3841), .A(n3840), .B(n3842), .ZN(n3963)
         );
  INV_X1 U4615 ( .A(n3963), .ZN(n3846) );
  INV_X1 U4616 ( .A(n3967), .ZN(n3845) );
  NAND2_X1 U4617 ( .A1(n3842), .A2(n3841), .ZN(n3969) );
  AOI21_X1 U4618 ( .B1(n3969), .B2(n3843), .A(n4391), .ZN(n3844) );
  AOI21_X1 U4619 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(n3970) );
  NAND2_X1 U4620 ( .A1(n3848), .A2(n3847), .ZN(n4080) );
  INV_X1 U4621 ( .A(n4080), .ZN(n3850) );
  INV_X1 U4622 ( .A(n4078), .ZN(n3849) );
  AND4_X1 U4623 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n4103), .ZN(n3890)
         );
  INV_X1 U4624 ( .A(n4114), .ZN(n3853) );
  OR2_X1 U4625 ( .A1(n3853), .A2(n3852), .ZN(n4139) );
  OR2_X1 U4626 ( .A1(n2255), .A2(n3854), .ZN(n4117) );
  NAND4_X1 U4627 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3868)
         );
  INV_X1 U4628 ( .A(n3859), .ZN(n3861) );
  XNOR2_X1 U4629 ( .A(n4234), .B(n3860), .ZN(n4254) );
  XNOR2_X1 U4630 ( .A(n4222), .B(n4239), .ZN(n4235) );
  NAND4_X1 U4631 ( .A1(n3862), .A2(n3861), .A3(n4254), .A4(n4235), .ZN(n3867)
         );
  INV_X1 U4632 ( .A(n3863), .ZN(n4137) );
  AND2_X1 U4633 ( .A1(n4137), .A2(n3864), .ZN(n4153) );
  AND2_X1 U4634 ( .A1(n3945), .A2(n4169), .ZN(n4207) );
  XNOR2_X1 U4635 ( .A(n4191), .B(n4179), .ZN(n4172) );
  NAND4_X1 U4636 ( .A1(n4153), .A2(n3865), .A3(n4207), .A4(n4172), .ZN(n3866)
         );
  NOR3_X1 U4637 ( .A1(n3868), .A2(n3867), .A3(n3866), .ZN(n3870) );
  NAND3_X1 U4638 ( .A1(n4117), .A2(n3870), .A3(n3869), .ZN(n3872) );
  NOR3_X1 U4639 ( .A1(n4139), .A2(n3872), .A3(n3871), .ZN(n3889) );
  INV_X1 U4640 ( .A(n3873), .ZN(n3875) );
  NAND4_X1 U4641 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n4624), .ZN(n3882)
         );
  INV_X1 U4642 ( .A(n3063), .ZN(n3880) );
  NAND4_X1 U4643 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  NOR2_X1 U4644 ( .A1(n3882), .A2(n3881), .ZN(n3888) );
  INV_X1 U4645 ( .A(n3883), .ZN(n3886) );
  AND4_X1 U4646 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n2251), .ZN(n3887)
         );
  NAND4_X1 U4647 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3959)
         );
  OAI21_X1 U4648 ( .B1(n2294), .B2(n3892), .A(n3936), .ZN(n3896) );
  NAND4_X1 U4649 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3939)
         );
  INV_X1 U4650 ( .A(n3940), .ZN(n3933) );
  INV_X1 U4651 ( .A(n3897), .ZN(n3900) );
  OAI211_X1 U4652 ( .C1(n3900), .C2(n4390), .A(n3899), .B(n3898), .ZN(n3903)
         );
  NAND3_X1 U4653 ( .A1(n3903), .A2(n3902), .A3(n3901), .ZN(n3906) );
  NAND3_X1 U4654 ( .A1(n3906), .A2(n3905), .A3(n3904), .ZN(n3909) );
  NAND3_X1 U4655 ( .A1(n3909), .A2(n3908), .A3(n3907), .ZN(n3912) );
  NAND4_X1 U4656 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3915), .ZN(n3914)
         );
  NAND3_X1 U4657 ( .A1(n3914), .A2(n2251), .A3(n3913), .ZN(n3920) );
  INV_X1 U4658 ( .A(n3926), .ZN(n3919) );
  INV_X1 U4659 ( .A(n3915), .ZN(n3917) );
  NOR2_X1 U4660 ( .A1(n3917), .A2(n3916), .ZN(n3918) );
  AOI22_X1 U4661 ( .A1(n3920), .A2(n3919), .B1(n3918), .B2(n3940), .ZN(n3925)
         );
  INV_X1 U4662 ( .A(n3921), .ZN(n3924) );
  INV_X1 U4663 ( .A(n3922), .ZN(n3923) );
  NOR3_X1 U4664 ( .A1(n3925), .A2(n3924), .A3(n3923), .ZN(n3930) );
  AOI21_X1 U4665 ( .B1(n3928), .B2(n3927), .A(n3926), .ZN(n3929) );
  OAI21_X1 U4666 ( .B1(n3930), .B2(n3929), .A(n3072), .ZN(n3931) );
  OAI21_X1 U4667 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(n3937) );
  AND4_X1 U4668 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3938)
         );
  AOI21_X1 U4669 ( .B1(n3940), .B2(n3939), .A(n3938), .ZN(n3943) );
  AOI211_X1 U4670 ( .C1(n3944), .C2(n3943), .A(n3942), .B(n3941), .ZN(n3948)
         );
  OAI211_X1 U4671 ( .C1(n3948), .C2(n3947), .A(n3946), .B(n3945), .ZN(n3950)
         );
  OAI221_X1 U4672 ( .B1(n3952), .B2(n3951), .C1(n3952), .C2(n3950), .A(n3949), 
        .ZN(n3954) );
  AOI21_X1 U4673 ( .B1(n3955), .B2(n3954), .A(n3953), .ZN(n3956) );
  OR4_X1 U4674 ( .A1(n3957), .A2(n3962), .A3(n3956), .A4(n3961), .ZN(n3958) );
  MUX2_X1 U4675 ( .A(n3959), .B(n3958), .S(n2595), .Z(n3968) );
  INV_X1 U4676 ( .A(n4103), .ZN(n3960) );
  NOR4_X1 U4677 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  AOI21_X1 U4678 ( .B1(n4288), .B2(n3965), .A(n3964), .ZN(n3966) );
  OAI222_X1 U4679 ( .A1(n3971), .A2(n3970), .B1(n3969), .B2(n3968), .C1(n3967), 
        .C2(n3966), .ZN(n3972) );
  XNOR2_X1 U4680 ( .A(n3972), .B(n4392), .ZN(n3977) );
  NOR2_X1 U4681 ( .A1(n3973), .A2(n4008), .ZN(n3975) );
  OAI21_X1 U4682 ( .B1(n3976), .B2(n4389), .A(B_REG_SCAN_IN), .ZN(n3974) );
  OAI22_X1 U4683 ( .A1(n3977), .A2(n3976), .B1(n3975), .B2(n3974), .ZN(U3239)
         );
  MUX2_X1 U4684 ( .A(n4076), .B(DATAO_REG_28__SCAN_IN), .S(n4004), .Z(U3578)
         );
  MUX2_X1 U4685 ( .A(n3978), .B(DATAO_REG_27__SCAN_IN), .S(n4004), .Z(U3577)
         );
  MUX2_X1 U4686 ( .A(n4143), .B(DATAO_REG_26__SCAN_IN), .S(n4004), .Z(U3576)
         );
  MUX2_X1 U4687 ( .A(DATAO_REG_24__SCAN_IN), .B(n3979), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4688 ( .A(DATAO_REG_23__SCAN_IN), .B(n3980), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4689 ( .A(n4222), .B(DATAO_REG_20__SCAN_IN), .S(n4004), .Z(U3570)
         );
  MUX2_X1 U4690 ( .A(n3981), .B(DATAO_REG_17__SCAN_IN), .S(n4004), .Z(U3567)
         );
  MUX2_X1 U4691 ( .A(n3982), .B(DATAO_REG_15__SCAN_IN), .S(n4004), .Z(U3565)
         );
  MUX2_X1 U4692 ( .A(DATAO_REG_14__SCAN_IN), .B(n3983), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4693 ( .A(DATAO_REG_13__SCAN_IN), .B(n3984), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4694 ( .A(n3985), .B(DATAO_REG_12__SCAN_IN), .S(n4004), .Z(U3562)
         );
  MUX2_X1 U4695 ( .A(DATAO_REG_11__SCAN_IN), .B(n3986), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4696 ( .A(n3987), .B(DATAO_REG_9__SCAN_IN), .S(n4004), .Z(U3559) );
  MUX2_X1 U4697 ( .A(DATAO_REG_7__SCAN_IN), .B(n3988), .S(U4043), .Z(U3557) );
  MUX2_X1 U4698 ( .A(n3989), .B(DATAO_REG_6__SCAN_IN), .S(n4004), .Z(U3556) );
  MUX2_X1 U4699 ( .A(n3990), .B(DATAO_REG_5__SCAN_IN), .S(n4004), .Z(U3555) );
  MUX2_X1 U4700 ( .A(DATAO_REG_4__SCAN_IN), .B(n3991), .S(U4043), .Z(U3554) );
  MUX2_X1 U4701 ( .A(DATAO_REG_1__SCAN_IN), .B(n3025), .S(U4043), .Z(U3551) );
  OAI211_X1 U4702 ( .C1(n3994), .C2(n3993), .A(n4577), .B(n3992), .ZN(n3999)
         );
  OAI211_X1 U4703 ( .C1(n4000), .C2(n3995), .A(n4588), .B(n4010), .ZN(n3998)
         );
  AOI22_X1 U4704 ( .A1(n4581), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3997) );
  NAND2_X1 U4705 ( .A1(n4556), .A2(n2232), .ZN(n3996) );
  NAND4_X1 U4706 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(U3241)
         );
  INV_X1 U4707 ( .A(n4000), .ZN(n4007) );
  INV_X1 U4708 ( .A(n4452), .ZN(n4001) );
  NAND3_X1 U4709 ( .A1(n4002), .A2(n4386), .A3(n4001), .ZN(n4006) );
  INV_X1 U4710 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U4711 ( .A1(n4452), .A2(n4894), .ZN(n4003) );
  NAND2_X1 U4712 ( .A1(n4386), .A2(n4003), .ZN(n4450) );
  AOI21_X1 U4713 ( .B1(n4450), .B2(n2344), .A(n4004), .ZN(n4005) );
  OAI211_X1 U4714 ( .C1(n4008), .C2(n4007), .A(n4006), .B(n4005), .ZN(n4467)
         );
  AOI22_X1 U4715 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4581), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4022) );
  MUX2_X1 U4716 ( .A(n3152), .B(REG2_REG_2__SCAN_IN), .S(n3146), .Z(n4011) );
  NAND3_X1 U4717 ( .A1(n4011), .A2(n4010), .A3(n4009), .ZN(n4012) );
  AND3_X1 U4718 ( .A1(n4013), .A2(n4012), .A3(n4588), .ZN(n4014) );
  AOI21_X1 U4719 ( .B1(n4556), .B2(n3146), .A(n4014), .ZN(n4021) );
  INV_X1 U4720 ( .A(n4015), .ZN(n4017) );
  NAND3_X1 U4721 ( .A1(n4017), .A2(n3992), .A3(n4016), .ZN(n4018) );
  NAND3_X1 U4722 ( .A1(n4577), .A2(n4019), .A3(n4018), .ZN(n4020) );
  NAND4_X1 U4723 ( .A1(n4467), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(U3242)
         );
  AOI22_X1 U4724 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4534), .B1(n4615), .B2(
        n4023), .ZN(n4524) );
  INV_X1 U4725 ( .A(n4523), .ZN(n4024) );
  NAND2_X1 U4726 ( .A1(n4024), .A2(n2425), .ZN(n4025) );
  NAND2_X1 U4727 ( .A1(n4025), .A2(n4543), .ZN(n4027) );
  NAND2_X1 U4728 ( .A1(n4027), .A2(n4026), .ZN(n4540) );
  INV_X1 U4729 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4539) );
  INV_X1 U4730 ( .A(n4027), .ZN(n4028) );
  INV_X1 U4731 ( .A(n4613), .ZN(n4030) );
  AOI22_X1 U4732 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4030), .B1(n4613), .B2(
        n4029), .ZN(n4548) );
  INV_X1 U4733 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U4734 ( .A1(n4031), .A2(n4612), .ZN(n4032) );
  INV_X1 U4735 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4736 ( .A1(n4034), .A2(n4033), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4609), .ZN(n4575) );
  NAND2_X1 U4737 ( .A1(n4034), .A2(n4033), .ZN(n4035) );
  INV_X1 U4738 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4818) );
  AOI22_X1 U4739 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4608), .B1(n4052), .B2(
        n4818), .ZN(n4584) );
  NAND2_X1 U4740 ( .A1(n4052), .A2(REG1_REG_18__SCAN_IN), .ZN(n4036) );
  XNOR2_X1 U4741 ( .A(n4392), .B(REG1_REG_19__SCAN_IN), .ZN(n4037) );
  NAND2_X1 U4742 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4052), .ZN(n4038) );
  OAI21_X1 U4743 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4052), .A(n4038), .ZN(n4587) );
  NAND2_X1 U4744 ( .A1(n4393), .A2(n4039), .ZN(n4040) );
  NAND2_X1 U4745 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4530), .ZN(n4043) );
  INV_X1 U4746 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4537) );
  NOR2_X1 U4747 ( .A1(n4045), .A2(n4535), .ZN(n4553) );
  NAND2_X1 U4748 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4613), .ZN(n4046) );
  OAI21_X1 U4749 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4613), .A(n4046), .ZN(n4552) );
  NOR2_X1 U4750 ( .A1(n4553), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U4751 ( .A1(n4048), .A2(n4612), .ZN(n4049) );
  NAND2_X1 U4752 ( .A1(n4049), .A2(n4561), .ZN(n4571) );
  NOR2_X1 U4753 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4609), .ZN(n4050) );
  AOI21_X1 U4754 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4609), .A(n4050), .ZN(n4572) );
  NAND2_X1 U4755 ( .A1(n4571), .A2(n4572), .ZN(n4570) );
  INV_X1 U4756 ( .A(n4050), .ZN(n4051) );
  AND2_X1 U4757 ( .A1(n4052), .A2(REG2_REG_18__SCAN_IN), .ZN(n4053) );
  NOR2_X1 U4758 ( .A1(n4586), .A2(n4053), .ZN(n4055) );
  XNOR2_X1 U4759 ( .A(n4058), .B(REG2_REG_19__SCAN_IN), .ZN(n4054) );
  XNOR2_X1 U4760 ( .A(n4055), .B(n4054), .ZN(n4060) );
  NAND2_X1 U4761 ( .A1(n4581), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4056) );
  OAI211_X1 U4762 ( .C1(n4593), .C2(n4058), .A(n4057), .B(n4056), .ZN(n4059)
         );
  AOI21_X1 U4763 ( .B1(n4060), .B2(n4588), .A(n4059), .ZN(n4061) );
  OAI21_X1 U4764 ( .B1(n4062), .B2(n4583), .A(n4061), .ZN(U3259) );
  INV_X1 U4765 ( .A(n4063), .ZN(n4064) );
  AOI21_X1 U4766 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4067) );
  XNOR2_X1 U4767 ( .A(n4067), .B(n4080), .ZN(n4073) );
  AOI22_X1 U4768 ( .A1(n4070), .A2(n4069), .B1(n4068), .B2(n4287), .ZN(n4071)
         );
  OAI21_X1 U4769 ( .B1(n4099), .B2(n4195), .A(n4071), .ZN(n4072) );
  INV_X1 U4770 ( .A(n4293), .ZN(n4074) );
  AOI21_X1 U4771 ( .B1(n4075), .B2(n4594), .A(n4074), .ZN(n4087) );
  XNOR2_X1 U4772 ( .A(n4081), .B(n4080), .ZN(n4291) );
  NAND2_X1 U4773 ( .A1(n4291), .A2(n4237), .ZN(n4086) );
  OAI21_X1 U4774 ( .B1(n4083), .B2(n4082), .A(n4284), .ZN(n4292) );
  INV_X1 U4775 ( .A(n4292), .ZN(n4084) );
  AOI22_X1 U4776 ( .A1(n4084), .A2(n4598), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4604), .ZN(n4085) );
  OAI211_X1 U4777 ( .C1(n4604), .C2(n4087), .A(n4086), .B(n4085), .ZN(U3354)
         );
  INV_X1 U4778 ( .A(n4089), .ZN(n4094) );
  INV_X1 U4779 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4091) );
  OAI22_X1 U4780 ( .A1(n4273), .A2(n4091), .B1(n4090), .B2(n4268), .ZN(n4093)
         );
  NOR2_X1 U4781 ( .A1(n2228), .A2(n4604), .ZN(n4092) );
  AOI211_X2 U4782 ( .C1(n4598), .C2(n4094), .A(n4093), .B(n4092), .ZN(n4095)
         );
  OAI21_X1 U4783 ( .B1(n4088), .B2(n4275), .A(n4095), .ZN(U3262) );
  OAI21_X1 U4784 ( .B1(n4097), .B2(n4103), .A(n4096), .ZN(n4102) );
  NOR2_X1 U4785 ( .A1(n4098), .A2(n4195), .ZN(n4101) );
  OAI22_X1 U4786 ( .A1(n4099), .A2(n4256), .B1(n4255), .B2(n4106), .ZN(n4100)
         );
  AOI211_X1 U4787 ( .C1(n4102), .C2(n4197), .A(n4101), .B(n4100), .ZN(n4298)
         );
  XNOR2_X1 U4788 ( .A(n4104), .B(n4103), .ZN(n4297) );
  NAND2_X1 U4789 ( .A1(n4297), .A2(n4237), .ZN(n4112) );
  INV_X1 U4790 ( .A(n3116), .ZN(n4105) );
  OAI21_X1 U4791 ( .B1(n4124), .B2(n4106), .A(n4105), .ZN(n4300) );
  INV_X1 U4792 ( .A(n4300), .ZN(n4110) );
  INV_X1 U4793 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4108) );
  OAI22_X1 U4794 ( .A1(n4273), .A2(n4108), .B1(n4107), .B2(n4268), .ZN(n4109)
         );
  AOI21_X1 U4795 ( .B1(n4110), .B2(n4598), .A(n4109), .ZN(n4111) );
  OAI211_X1 U4796 ( .C1(n4298), .C2(n4604), .A(n4112), .B(n4111), .ZN(U3263)
         );
  XOR2_X1 U4797 ( .A(n4117), .B(n4113), .Z(n4302) );
  INV_X1 U4798 ( .A(n4302), .ZN(n4131) );
  NAND2_X1 U4799 ( .A1(n4115), .A2(n4114), .ZN(n4116) );
  XOR2_X1 U4800 ( .A(n4117), .B(n4116), .Z(n4122) );
  OAI22_X1 U4801 ( .A1(n4118), .A2(n4256), .B1(n4255), .B2(n4126), .ZN(n4119)
         );
  AOI21_X1 U4802 ( .B1(n4260), .B2(n4120), .A(n4119), .ZN(n4121) );
  OAI21_X1 U4803 ( .B1(n4122), .B2(n4262), .A(n4121), .ZN(n4301) );
  INV_X1 U4804 ( .A(n4123), .ZN(n4133) );
  INV_X1 U4805 ( .A(n4124), .ZN(n4125) );
  OAI21_X1 U4806 ( .B1(n4133), .B2(n4126), .A(n4125), .ZN(n4361) );
  AOI22_X1 U4807 ( .A1(n4604), .A2(REG2_REG_26__SCAN_IN), .B1(n4127), .B2(
        n4594), .ZN(n4128) );
  OAI21_X1 U4808 ( .B1(n4361), .B2(n4266), .A(n4128), .ZN(n4129) );
  AOI21_X1 U4809 ( .B1(n4301), .B2(n4273), .A(n4129), .ZN(n4130) );
  OAI21_X1 U4810 ( .B1(n4131), .B2(n4275), .A(n4130), .ZN(U3264) );
  XNOR2_X1 U4811 ( .A(n4132), .B(n4139), .ZN(n4308) );
  AOI21_X1 U4812 ( .B1(n4141), .B2(n4160), .A(n4133), .ZN(n4305) );
  INV_X1 U4813 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4136) );
  INV_X1 U4814 ( .A(n4134), .ZN(n4135) );
  OAI22_X1 U4815 ( .A1(n4273), .A2(n4136), .B1(n4135), .B2(n4268), .ZN(n4148)
         );
  NAND2_X1 U4816 ( .A1(n4138), .A2(n4137), .ZN(n4140) );
  XNOR2_X1 U4817 ( .A(n4140), .B(n4139), .ZN(n4146) );
  AOI22_X1 U4818 ( .A1(n4143), .A2(n4142), .B1(n4287), .B2(n4141), .ZN(n4144)
         );
  OAI21_X1 U4819 ( .B1(n4173), .B2(n4195), .A(n4144), .ZN(n4145) );
  AOI21_X1 U4820 ( .B1(n4146), .B2(n4197), .A(n4145), .ZN(n4307) );
  NOR2_X1 U4821 ( .A1(n4307), .A2(n4604), .ZN(n4147) );
  AOI211_X1 U4822 ( .C1(n4305), .C2(n4598), .A(n4148), .B(n4147), .ZN(n4149)
         );
  OAI21_X1 U4823 ( .B1(n4308), .B2(n4275), .A(n4149), .ZN(U3265) );
  XOR2_X1 U4824 ( .A(n4153), .B(n4150), .Z(n4310) );
  INV_X1 U4825 ( .A(n4310), .ZN(n4167) );
  NAND2_X1 U4826 ( .A1(n4152), .A2(n4151), .ZN(n4154) );
  XNOR2_X1 U4827 ( .A(n4154), .B(n4153), .ZN(n4158) );
  NOR2_X1 U4828 ( .A1(n4191), .A2(n4195), .ZN(n4157) );
  OAI22_X1 U4829 ( .A1(n4155), .A2(n4256), .B1(n4255), .B2(n4161), .ZN(n4156)
         );
  AOI211_X1 U4830 ( .C1(n4158), .C2(n4197), .A(n4157), .B(n4156), .ZN(n4159)
         );
  INV_X1 U4831 ( .A(n4159), .ZN(n4309) );
  INV_X1 U4832 ( .A(n4178), .ZN(n4162) );
  OAI21_X1 U4833 ( .B1(n4162), .B2(n4161), .A(n4160), .ZN(n4366) );
  AOI22_X1 U4834 ( .A1(n4604), .A2(REG2_REG_24__SCAN_IN), .B1(n4163), .B2(
        n4594), .ZN(n4164) );
  OAI21_X1 U4835 ( .B1(n4366), .B2(n4266), .A(n4164), .ZN(n4165) );
  AOI21_X1 U4836 ( .B1(n4309), .B2(n4273), .A(n4165), .ZN(n4166) );
  OAI21_X1 U4837 ( .B1(n4167), .B2(n4275), .A(n4166), .ZN(U3266) );
  XNOR2_X1 U4838 ( .A(n4168), .B(n4172), .ZN(n4314) );
  INV_X1 U4839 ( .A(n4314), .ZN(n4186) );
  INV_X1 U4840 ( .A(n4207), .ZN(n4216) );
  OR2_X1 U4841 ( .A1(n4217), .A2(n4216), .ZN(n4219) );
  OAI21_X1 U4842 ( .B1(n4190), .B2(n4189), .A(n4170), .ZN(n4171) );
  XOR2_X1 U4843 ( .A(n4172), .B(n4171), .Z(n4177) );
  OAI22_X1 U4844 ( .A1(n4173), .A2(n4256), .B1(n4255), .B2(n4179), .ZN(n4174)
         );
  AOI21_X1 U4845 ( .B1(n4260), .B2(n4175), .A(n4174), .ZN(n4176) );
  OAI21_X1 U4846 ( .B1(n4177), .B2(n4262), .A(n4176), .ZN(n4313) );
  OAI21_X1 U4847 ( .B1(n4318), .B2(n4179), .A(n4178), .ZN(n4370) );
  NOR2_X1 U4848 ( .A1(n4370), .A2(n4266), .ZN(n4184) );
  INV_X1 U4849 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4182) );
  INV_X1 U4850 ( .A(n4180), .ZN(n4181) );
  OAI22_X1 U4851 ( .A1(n4273), .A2(n4182), .B1(n4181), .B2(n4268), .ZN(n4183)
         );
  AOI211_X1 U4852 ( .C1(n4313), .C2(n4273), .A(n4184), .B(n4183), .ZN(n4185)
         );
  OAI21_X1 U4853 ( .B1(n4186), .B2(n4275), .A(n4185), .ZN(U3267) );
  OAI21_X1 U4854 ( .B1(n4188), .B2(n4189), .A(n4187), .ZN(n4321) );
  XNOR2_X1 U4855 ( .A(n4190), .B(n4189), .ZN(n4198) );
  OR2_X1 U4856 ( .A1(n4191), .A2(n4256), .ZN(n4194) );
  NAND2_X1 U4857 ( .A1(n4192), .A2(n4287), .ZN(n4193) );
  OAI211_X1 U4858 ( .C1(n4227), .C2(n4195), .A(n4194), .B(n4193), .ZN(n4196)
         );
  AOI21_X1 U4859 ( .B1(n4198), .B2(n4197), .A(n4196), .ZN(n4320) );
  INV_X1 U4860 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4200) );
  OAI22_X1 U4861 ( .A1(n4273), .A2(n4200), .B1(n4199), .B2(n4268), .ZN(n4201)
         );
  INV_X1 U4862 ( .A(n4201), .ZN(n4204) );
  NOR2_X1 U4863 ( .A1(n4209), .A2(n4202), .ZN(n4317) );
  OR3_X1 U4864 ( .A1(n4318), .A2(n4317), .A3(n4266), .ZN(n4203) );
  OAI211_X1 U4865 ( .C1(n4320), .C2(n4604), .A(n4204), .B(n4203), .ZN(n4205)
         );
  INV_X1 U4866 ( .A(n4205), .ZN(n4206) );
  OAI21_X1 U4867 ( .B1(n4321), .B2(n4275), .A(n4206), .ZN(U3268) );
  XNOR2_X1 U4868 ( .A(n4208), .B(n4207), .ZN(n4325) );
  AOI21_X1 U4869 ( .B1(n4210), .B2(n4241), .A(n4209), .ZN(n4322) );
  INV_X1 U4870 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4213) );
  INV_X1 U4871 ( .A(n4211), .ZN(n4212) );
  OAI22_X1 U4872 ( .A1(n4273), .A2(n4213), .B1(n4212), .B2(n4268), .ZN(n4224)
         );
  OAI22_X1 U4873 ( .A1(n4215), .A2(n4256), .B1(n4255), .B2(n4214), .ZN(n4221)
         );
  NAND2_X1 U4874 ( .A1(n4217), .A2(n4216), .ZN(n4218) );
  AOI21_X1 U4875 ( .B1(n4219), .B2(n4218), .A(n4262), .ZN(n4220) );
  AOI211_X1 U4876 ( .C1(n4260), .C2(n4222), .A(n4221), .B(n4220), .ZN(n4324)
         );
  NOR2_X1 U4877 ( .A1(n4324), .A2(n4604), .ZN(n4223) );
  AOI211_X1 U4878 ( .C1(n4322), .C2(n4598), .A(n4224), .B(n4223), .ZN(n4225)
         );
  OAI21_X1 U4879 ( .B1(n4325), .B2(n4275), .A(n4225), .ZN(U3269) );
  OAI22_X1 U4880 ( .A1(n4227), .A2(n4256), .B1(n4255), .B2(n4226), .ZN(n4233)
         );
  NAND2_X1 U4881 ( .A1(n4229), .A2(n4228), .ZN(n4230) );
  XOR2_X1 U4882 ( .A(n4235), .B(n4230), .Z(n4231) );
  NOR2_X1 U4883 ( .A1(n4231), .A2(n4262), .ZN(n4232) );
  AOI211_X1 U4884 ( .C1(n4260), .C2(n4234), .A(n4233), .B(n4232), .ZN(n4326)
         );
  XNOR2_X1 U4885 ( .A(n4236), .B(n4235), .ZN(n4328) );
  NAND2_X1 U4886 ( .A1(n4328), .A2(n4237), .ZN(n4247) );
  NAND2_X1 U4887 ( .A1(n4238), .A2(n4239), .ZN(n4240) );
  NAND2_X1 U4888 ( .A1(n4241), .A2(n4240), .ZN(n4375) );
  INV_X1 U4889 ( .A(n4375), .ZN(n4245) );
  INV_X1 U4890 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4243) );
  OAI22_X1 U4891 ( .A1(n4273), .A2(n4243), .B1(n4242), .B2(n4268), .ZN(n4244)
         );
  AOI21_X1 U4892 ( .B1(n4245), .B2(n4598), .A(n4244), .ZN(n4246) );
  OAI211_X1 U4893 ( .C1(n4604), .C2(n4326), .A(n4247), .B(n4246), .ZN(U3270)
         );
  XOR2_X1 U4894 ( .A(n4254), .B(n4248), .Z(n4331) );
  INV_X1 U4895 ( .A(n4331), .ZN(n4276) );
  INV_X1 U4896 ( .A(n4249), .ZN(n4251) );
  AOI21_X1 U4897 ( .B1(n4252), .B2(n4251), .A(n4250), .ZN(n4253) );
  XOR2_X1 U4898 ( .A(n4254), .B(n4253), .Z(n4263) );
  OAI22_X1 U4899 ( .A1(n4257), .A2(n4256), .B1(n4255), .B2(n4264), .ZN(n4258)
         );
  AOI21_X1 U4900 ( .B1(n4260), .B2(n4259), .A(n4258), .ZN(n4261) );
  OAI21_X1 U4901 ( .B1(n4263), .B2(n4262), .A(n4261), .ZN(n4330) );
  OAI21_X1 U4902 ( .B1(n4265), .B2(n4264), .A(n4238), .ZN(n4380) );
  NOR2_X1 U4903 ( .A1(n4380), .A2(n4266), .ZN(n4272) );
  INV_X1 U4904 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4270) );
  INV_X1 U4905 ( .A(n4267), .ZN(n4269) );
  OAI22_X1 U4906 ( .A1(n4273), .A2(n4270), .B1(n4269), .B2(n4268), .ZN(n4271)
         );
  AOI211_X1 U4907 ( .C1(n4330), .C2(n4273), .A(n4272), .B(n4271), .ZN(n4274)
         );
  OAI21_X1 U4908 ( .B1(n4276), .B2(n4275), .A(n4274), .ZN(U3271) );
  INV_X1 U4909 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4282) );
  INV_X1 U4910 ( .A(n4333), .ZN(n4277) );
  NAND2_X1 U4911 ( .A1(n4278), .A2(n4277), .ZN(n4281) );
  NAND2_X1 U4912 ( .A1(n4279), .A2(n4684), .ZN(n4280) );
  OAI211_X1 U4913 ( .C1(n4684), .C2(n4282), .A(n4281), .B(n4280), .ZN(U3549)
         );
  AOI21_X1 U4914 ( .B1(n4288), .B2(n4284), .A(n4283), .ZN(n4447) );
  INV_X1 U4915 ( .A(n4447), .ZN(n4355) );
  INV_X1 U4916 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4289) );
  INV_X1 U4917 ( .A(n4285), .ZN(n4286) );
  AOI21_X1 U4918 ( .B1(n4288), .B2(n4287), .A(n4286), .ZN(n4449) );
  MUX2_X1 U4919 ( .A(n4289), .B(n4449), .S(n4684), .Z(n4290) );
  OAI21_X1 U4920 ( .B1(n4355), .B2(n4333), .A(n4290), .ZN(U3548) );
  NAND2_X1 U4921 ( .A1(n4291), .A2(n4656), .ZN(n4296) );
  NAND2_X1 U4922 ( .A1(n4296), .A2(n4295), .ZN(n4356) );
  MUX2_X1 U4923 ( .A(REG1_REG_29__SCAN_IN), .B(n4356), .S(n4684), .Z(U3547) );
  NAND2_X1 U4924 ( .A1(n4297), .A2(n4656), .ZN(n4299) );
  OAI211_X1 U4925 ( .C1(n3251), .C2(n4300), .A(n4299), .B(n4298), .ZN(n4357)
         );
  MUX2_X1 U4926 ( .A(REG1_REG_27__SCAN_IN), .B(n4357), .S(n4684), .Z(U3545) );
  INV_X1 U4927 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4303) );
  AOI21_X1 U4928 ( .B1(n4302), .B2(n4656), .A(n4301), .ZN(n4358) );
  MUX2_X1 U4929 ( .A(n4303), .B(n4358), .S(n4684), .Z(n4304) );
  OAI21_X1 U4930 ( .B1(n4333), .B2(n4361), .A(n4304), .ZN(U3544) );
  NAND2_X1 U4931 ( .A1(n4305), .A2(n2598), .ZN(n4306) );
  OAI211_X1 U4932 ( .C1(n4308), .C2(n4661), .A(n4307), .B(n4306), .ZN(n4362)
         );
  MUX2_X1 U4933 ( .A(REG1_REG_25__SCAN_IN), .B(n4362), .S(n4684), .Z(U3543) );
  INV_X1 U4934 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4311) );
  AOI21_X1 U4935 ( .B1(n4310), .B2(n4656), .A(n4309), .ZN(n4363) );
  MUX2_X1 U4936 ( .A(n4311), .B(n4363), .S(n4684), .Z(n4312) );
  OAI21_X1 U4937 ( .B1(n4333), .B2(n4366), .A(n4312), .ZN(U3542) );
  INV_X1 U4938 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4315) );
  AOI21_X1 U4939 ( .B1(n4314), .B2(n4656), .A(n4313), .ZN(n4367) );
  MUX2_X1 U4940 ( .A(n4315), .B(n4367), .S(n4684), .Z(n4316) );
  OAI21_X1 U4941 ( .B1(n4333), .B2(n4370), .A(n4316), .ZN(U3541) );
  OR3_X1 U4942 ( .A1(n4318), .A2(n4317), .A3(n3251), .ZN(n4319) );
  OAI211_X1 U4943 ( .C1(n4321), .C2(n4661), .A(n4320), .B(n4319), .ZN(n4371)
         );
  MUX2_X1 U4944 ( .A(REG1_REG_22__SCAN_IN), .B(n4371), .S(n4684), .Z(U3540) );
  NAND2_X1 U4945 ( .A1(n4322), .A2(n2598), .ZN(n4323) );
  OAI211_X1 U4946 ( .C1(n4325), .C2(n4661), .A(n4324), .B(n4323), .ZN(n4372)
         );
  MUX2_X1 U4947 ( .A(REG1_REG_21__SCAN_IN), .B(n4372), .S(n4684), .Z(U3539) );
  INV_X1 U4948 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4909) );
  INV_X1 U4949 ( .A(n4326), .ZN(n4327) );
  AOI21_X1 U4950 ( .B1(n4328), .B2(n4656), .A(n4327), .ZN(n4373) );
  MUX2_X1 U4951 ( .A(n4909), .B(n4373), .S(n4684), .Z(n4329) );
  OAI21_X1 U4952 ( .B1(n4333), .B2(n4375), .A(n4329), .ZN(U3538) );
  INV_X1 U4953 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4953) );
  AOI21_X1 U4954 ( .B1(n4331), .B2(n4656), .A(n4330), .ZN(n4376) );
  MUX2_X1 U4955 ( .A(n4953), .B(n4376), .S(n4684), .Z(n4332) );
  OAI21_X1 U4956 ( .B1(n4333), .B2(n4380), .A(n4332), .ZN(U3537) );
  INV_X1 U4957 ( .A(n4334), .ZN(n4337) );
  OAI211_X1 U4958 ( .C1(n4337), .C2(n4661), .A(n4336), .B(n4335), .ZN(n4381)
         );
  MUX2_X1 U4959 ( .A(REG1_REG_18__SCAN_IN), .B(n4381), .S(n4684), .Z(U3536) );
  NAND3_X1 U4960 ( .A1(n4339), .A2(n2598), .A3(n4338), .ZN(n4340) );
  OAI211_X1 U4961 ( .C1(n4342), .C2(n4661), .A(n4341), .B(n4340), .ZN(n4382)
         );
  MUX2_X1 U4962 ( .A(REG1_REG_17__SCAN_IN), .B(n4382), .S(n4684), .Z(U3535) );
  INV_X1 U4963 ( .A(n4343), .ZN(n4347) );
  NAND3_X1 U4964 ( .A1(n4345), .A2(n2598), .A3(n4344), .ZN(n4346) );
  OAI211_X1 U4965 ( .C1(n4348), .C2(n4661), .A(n4347), .B(n4346), .ZN(n4383)
         );
  MUX2_X1 U4966 ( .A(REG1_REG_16__SCAN_IN), .B(n4383), .S(n4684), .Z(U3534) );
  NAND3_X1 U4967 ( .A1(n3636), .A2(n4349), .A3(n2598), .ZN(n4350) );
  OAI211_X1 U4968 ( .C1(n4352), .C2(n4668), .A(n4351), .B(n4350), .ZN(n4384)
         );
  MUX2_X1 U4969 ( .A(REG1_REG_14__SCAN_IN), .B(n4384), .S(n4684), .Z(U3532) );
  INV_X1 U4970 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4353) );
  MUX2_X1 U4971 ( .A(n4353), .B(n4449), .S(n4673), .Z(n4354) );
  OAI21_X1 U4972 ( .B1(n4355), .B2(n4379), .A(n4354), .ZN(U3516) );
  MUX2_X1 U4973 ( .A(REG0_REG_29__SCAN_IN), .B(n4356), .S(n4673), .Z(U3515) );
  MUX2_X1 U4974 ( .A(REG0_REG_27__SCAN_IN), .B(n4357), .S(n4673), .Z(U3513) );
  INV_X1 U4975 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4359) );
  MUX2_X1 U4976 ( .A(n4359), .B(n4358), .S(n4673), .Z(n4360) );
  OAI21_X1 U4977 ( .B1(n4361), .B2(n4379), .A(n4360), .ZN(U3512) );
  MUX2_X1 U4978 ( .A(REG0_REG_25__SCAN_IN), .B(n4362), .S(n4673), .Z(U3511) );
  INV_X1 U4979 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4364) );
  MUX2_X1 U4980 ( .A(n4364), .B(n4363), .S(n4673), .Z(n4365) );
  OAI21_X1 U4981 ( .B1(n4366), .B2(n4379), .A(n4365), .ZN(U3510) );
  INV_X1 U4982 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4368) );
  MUX2_X1 U4983 ( .A(n4368), .B(n4367), .S(n4673), .Z(n4369) );
  OAI21_X1 U4984 ( .B1(n4370), .B2(n4379), .A(n4369), .ZN(U3509) );
  MUX2_X1 U4985 ( .A(REG0_REG_22__SCAN_IN), .B(n4371), .S(n4673), .Z(U3508) );
  MUX2_X1 U4986 ( .A(REG0_REG_21__SCAN_IN), .B(n4372), .S(n4673), .Z(U3507) );
  INV_X1 U4987 ( .A(REG0_REG_20__SCAN_IN), .ZN(n5053) );
  MUX2_X1 U4988 ( .A(n5053), .B(n4373), .S(n4673), .Z(n4374) );
  OAI21_X1 U4989 ( .B1(n4375), .B2(n4379), .A(n4374), .ZN(U3506) );
  INV_X1 U4990 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4377) );
  MUX2_X1 U4991 ( .A(n4377), .B(n4376), .S(n4673), .Z(n4378) );
  OAI21_X1 U4992 ( .B1(n4380), .B2(n4379), .A(n4378), .ZN(U3505) );
  MUX2_X1 U4993 ( .A(REG0_REG_18__SCAN_IN), .B(n4381), .S(n4673), .Z(U3503) );
  MUX2_X1 U4994 ( .A(REG0_REG_17__SCAN_IN), .B(n4382), .S(n4673), .Z(U3501) );
  MUX2_X1 U4995 ( .A(REG0_REG_16__SCAN_IN), .B(n4383), .S(n4673), .Z(U3499) );
  MUX2_X1 U4996 ( .A(REG0_REG_14__SCAN_IN), .B(n4384), .S(n4673), .Z(U3495) );
  MUX2_X1 U4997 ( .A(DATAI_30_), .B(n4385), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4998 ( .A(n4386), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U4999 ( .A(n4452), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5000 ( .A(n2551), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5001 ( .A(DATAI_25_), .B(n4387), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5002 ( .A(n4388), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5003 ( .A(n4389), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5004 ( .A(n4390), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5005 ( .A(DATAI_20_), .B(n4391), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5006 ( .A(n4392), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5007 ( .A(n4543), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5008 ( .A(n4393), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5009 ( .A(n4394), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5010 ( .A(n4395), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5011 ( .A(n4479), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5012 ( .A(DATAI_4_), .B(n4461), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5013 ( .A(DATAI_3_), .B(n4396), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5014 ( .A(n3146), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5015 ( .A(n2232), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI22_X1 U5016 ( .A1(n4421), .A2(n4429), .B1(n4430), .B2(n4397), .ZN(n4402)
         );
  NOR2_X1 U5017 ( .A1(STATE_REG_SCAN_IN), .A2(n4398), .ZN(n4560) );
  INV_X1 U5018 ( .A(n4560), .ZN(n4399) );
  OAI21_X1 U5019 ( .B1(n4433), .B2(n4400), .A(n4399), .ZN(n4401) );
  NOR2_X1 U5020 ( .A1(n4402), .A2(n4401), .ZN(n4408) );
  OR2_X1 U5021 ( .A1(n4403), .A2(n4437), .ZN(n4440) );
  NAND2_X1 U5022 ( .A1(n4440), .A2(n4436), .ZN(n4404) );
  XOR2_X1 U5023 ( .A(n4405), .B(n4404), .Z(n4406) );
  NAND2_X1 U5024 ( .A1(n4406), .A2(n4441), .ZN(n4407) );
  OAI211_X1 U5025 ( .C1(n4446), .C2(n4409), .A(n4408), .B(n4407), .ZN(U3223)
         );
  OAI22_X1 U5026 ( .A1(n4429), .A2(n4410), .B1(STATE_REG_SCAN_IN), .B2(n5042), 
        .ZN(n4411) );
  INV_X1 U5027 ( .A(n4411), .ZN(n4426) );
  XOR2_X1 U5028 ( .A(n4413), .B(n4412), .Z(n4416) );
  OAI21_X1 U5029 ( .B1(n4416), .B2(n4414), .A(n4415), .ZN(n4424) );
  INV_X1 U5030 ( .A(n4417), .ZN(n4419) );
  AOI21_X1 U5031 ( .B1(n4414), .B2(n4419), .A(n4418), .ZN(n4423) );
  OAI22_X1 U5032 ( .A1(n4430), .A2(n4421), .B1(n4433), .B2(n4420), .ZN(n4422)
         );
  AOI21_X1 U5033 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(n4425) );
  OAI211_X1 U5034 ( .C1(n4446), .C2(n4427), .A(n4426), .B(n4425), .ZN(U3235)
         );
  OAI22_X1 U5035 ( .A1(n4431), .A2(n4430), .B1(n4429), .B2(n4428), .ZN(n4435)
         );
  NAND2_X1 U5036 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4557) );
  OAI21_X1 U5037 ( .B1(n4433), .B2(n4432), .A(n4557), .ZN(n4434) );
  NOR2_X1 U5038 ( .A1(n4435), .A2(n4434), .ZN(n4444) );
  INV_X1 U5039 ( .A(n4436), .ZN(n4439) );
  OAI21_X1 U5040 ( .B1(n4403), .B2(n4439), .A(n4437), .ZN(n4438) );
  OAI21_X1 U5041 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n4442) );
  NAND2_X1 U5042 ( .A1(n4442), .A2(n4441), .ZN(n4443) );
  OAI211_X1 U5043 ( .C1(n4446), .C2(n4445), .A(n4444), .B(n4443), .ZN(U3238)
         );
  AOI22_X1 U5044 ( .A1(n4447), .A2(n4598), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4604), .ZN(n4448) );
  OAI21_X1 U5045 ( .B1(n4604), .B2(n4449), .A(n4448), .ZN(U3261) );
  INV_X1 U5046 ( .A(n4450), .ZN(n4451) );
  OAI21_X1 U5047 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4452), .A(n4451), .ZN(n4453)
         );
  XNOR2_X1 U5048 ( .A(n4453), .B(n2344), .ZN(n4456) );
  AOI22_X1 U5049 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4581), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4454) );
  OAI21_X1 U5050 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(U3240) );
  XNOR2_X1 U5051 ( .A(n4457), .B(REG2_REG_4__SCAN_IN), .ZN(n4458) );
  NAND2_X1 U5052 ( .A1(n4588), .A2(n4458), .ZN(n4466) );
  XNOR2_X1 U5053 ( .A(n4459), .B(REG1_REG_4__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U5054 ( .A1(n4577), .A2(n4460), .ZN(n4465) );
  NAND2_X1 U5055 ( .A1(n4556), .A2(n4461), .ZN(n4464) );
  AOI21_X1 U5056 ( .B1(n4581), .B2(ADDR_REG_4__SCAN_IN), .A(n4462), .ZN(n4463)
         );
  AND4_X1 U5057 ( .A1(n4466), .A2(n4465), .A3(n4464), .A4(n4463), .ZN(n4468)
         );
  NAND2_X1 U5058 ( .A1(n4468), .A2(n4467), .ZN(U3244) );
  INV_X1 U5059 ( .A(n4469), .ZN(n4473) );
  INV_X1 U5060 ( .A(n4470), .ZN(n4471) );
  INV_X1 U5061 ( .A(n4588), .ZN(n4550) );
  AOI211_X1 U5062 ( .C1(n4473), .C2(n4472), .A(n4471), .B(n4550), .ZN(n4478)
         );
  AOI211_X1 U5063 ( .C1(n4476), .C2(n4475), .A(n4474), .B(n4583), .ZN(n4477)
         );
  AOI211_X1 U5064 ( .C1(n4556), .C2(n4479), .A(n4478), .B(n4477), .ZN(n4480)
         );
  INV_X1 U5065 ( .A(n4480), .ZN(n4481) );
  AOI211_X1 U5066 ( .C1(n4581), .C2(ADDR_REG_5__SCAN_IN), .A(n4482), .B(n4481), 
        .ZN(n4483) );
  INV_X1 U5067 ( .A(n4483), .ZN(U3245) );
  AOI21_X1 U5068 ( .B1(n4581), .B2(ADDR_REG_6__SCAN_IN), .A(n4484), .ZN(n4493)
         );
  OAI211_X1 U5069 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4486), .A(n4577), .B(n4485), 
        .ZN(n4492) );
  OAI211_X1 U5070 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4488), .A(n4588), .B(n4487), 
        .ZN(n4491) );
  NAND2_X1 U5071 ( .A1(n4489), .A2(n4556), .ZN(n4490) );
  NAND4_X1 U5072 ( .A1(n4493), .A2(n4492), .A3(n4491), .A4(n4490), .ZN(U3246)
         );
  AOI211_X1 U5073 ( .C1(n4812), .C2(n4495), .A(n4494), .B(n4583), .ZN(n4497)
         );
  AOI211_X1 U5074 ( .C1(n4581), .C2(ADDR_REG_8__SCAN_IN), .A(n4497), .B(n4496), 
        .ZN(n4501) );
  OAI211_X1 U5075 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4499), .A(n4588), .B(n4498), 
        .ZN(n4500) );
  OAI211_X1 U5076 ( .C1(n4593), .C2(n4502), .A(n4501), .B(n4500), .ZN(U3248)
         );
  AOI211_X1 U5077 ( .C1(n4505), .C2(n4504), .A(n4503), .B(n4583), .ZN(n4507)
         );
  AOI211_X1 U5078 ( .C1(n4581), .C2(ADDR_REG_9__SCAN_IN), .A(n4507), .B(n4506), 
        .ZN(n4512) );
  OAI211_X1 U5079 ( .C1(n4510), .C2(n4509), .A(n4588), .B(n4508), .ZN(n4511)
         );
  OAI211_X1 U5080 ( .C1(n4593), .C2(n4620), .A(n4512), .B(n4511), .ZN(U3249)
         );
  AOI211_X1 U5081 ( .C1(n4515), .C2(n4514), .A(n4513), .B(n4583), .ZN(n4517)
         );
  AOI211_X1 U5082 ( .C1(n4581), .C2(ADDR_REG_10__SCAN_IN), .A(n4517), .B(n4516), .ZN(n4521) );
  OAI211_X1 U5083 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4519), .A(n4588), .B(n4518), .ZN(n4520) );
  OAI211_X1 U5084 ( .C1(n4593), .C2(n4522), .A(n4521), .B(n4520), .ZN(U3250)
         );
  AOI211_X1 U5085 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4583), .ZN(n4527)
         );
  AOI211_X1 U5086 ( .C1(n4581), .C2(ADDR_REG_13__SCAN_IN), .A(n4527), .B(n4526), .ZN(n4533) );
  INV_X1 U5087 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5088 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4615), .B1(n4534), .B2(
        n4528), .ZN(n4531) );
  AOI21_X1 U5089 ( .B1(n4531), .B2(n4530), .A(n4550), .ZN(n4529) );
  OAI21_X1 U5090 ( .B1(n4531), .B2(n4530), .A(n4529), .ZN(n4532) );
  OAI211_X1 U5091 ( .C1(n4593), .C2(n4534), .A(n4533), .B(n4532), .ZN(U3253)
         );
  NAND2_X1 U5092 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4581), .ZN(n4546) );
  AOI211_X1 U5093 ( .C1(n4537), .C2(n4536), .A(n4535), .B(n4550), .ZN(n4542)
         );
  AOI211_X1 U5094 ( .C1(n4540), .C2(n4539), .A(n4538), .B(n4583), .ZN(n4541)
         );
  AOI211_X1 U5095 ( .C1(n4556), .C2(n4543), .A(n4542), .B(n4541), .ZN(n4545)
         );
  NAND3_X1 U5096 ( .A1(n4546), .A2(n4545), .A3(n4544), .ZN(U3254) );
  INV_X1 U5097 ( .A(n4581), .ZN(n4559) );
  INV_X1 U5098 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n5036) );
  AOI211_X1 U5099 ( .C1(n4549), .C2(n4548), .A(n4547), .B(n4583), .ZN(n4555)
         );
  AOI211_X1 U5100 ( .C1(n4553), .C2(n4552), .A(n4551), .B(n4550), .ZN(n4554)
         );
  AOI211_X1 U5101 ( .C1(n4556), .C2(n4613), .A(n4555), .B(n4554), .ZN(n4558)
         );
  OAI211_X1 U5102 ( .C1(n4559), .C2(n5036), .A(n4558), .B(n4557), .ZN(U3255)
         );
  AOI21_X1 U5103 ( .B1(n4581), .B2(ADDR_REG_16__SCAN_IN), .A(n4560), .ZN(n4568) );
  OAI21_X1 U5104 ( .B1(n4564), .B2(n4563), .A(n4562), .ZN(n4565) );
  AOI22_X1 U5105 ( .A1(n4588), .A2(n4566), .B1(n4577), .B2(n4565), .ZN(n4567)
         );
  OAI211_X1 U5106 ( .C1(n4612), .C2(n4593), .A(n4568), .B(n4567), .ZN(U3256)
         );
  AOI21_X1 U5107 ( .B1(n4581), .B2(ADDR_REG_17__SCAN_IN), .A(n4569), .ZN(n4580) );
  OAI21_X1 U5108 ( .B1(n4572), .B2(n4571), .A(n4570), .ZN(n4578) );
  OAI21_X1 U5109 ( .B1(n4575), .B2(n4574), .A(n4573), .ZN(n4576) );
  AOI22_X1 U5110 ( .A1(n4588), .A2(n4578), .B1(n4577), .B2(n4576), .ZN(n4579)
         );
  OAI211_X1 U5111 ( .C1(n4034), .C2(n4593), .A(n4580), .B(n4579), .ZN(U3257)
         );
  AOI22_X1 U5112 ( .A1(ADDR_REG_18__SCAN_IN), .A2(n4581), .B1(
        REG3_REG_18__SCAN_IN), .B2(U3149), .ZN(n4592) );
  OAI211_X1 U5113 ( .C1(n4608), .C2(n4593), .A(n4592), .B(n4591), .ZN(U3258)
         );
  AOI22_X1 U5114 ( .A1(n4595), .A2(n4594), .B1(REG2_REG_6__SCAN_IN), .B2(n4604), .ZN(n4602) );
  INV_X1 U5115 ( .A(n4596), .ZN(n4597) );
  AOI22_X1 U5116 ( .A1(n4600), .A2(n4599), .B1(n4598), .B2(n4597), .ZN(n4601)
         );
  OAI211_X1 U5117 ( .C1(n4604), .C2(n4603), .A(n4602), .B(n4601), .ZN(U3284)
         );
  INV_X1 U5118 ( .A(D_REG_31__SCAN_IN), .ZN(n4865) );
  NOR2_X1 U5119 ( .A1(n4605), .A2(n4865), .ZN(U3291) );
  AND2_X1 U5120 ( .A1(D_REG_30__SCAN_IN), .A2(n4685), .ZN(U3292) );
  AND2_X1 U5121 ( .A1(D_REG_29__SCAN_IN), .A2(n4685), .ZN(U3293) );
  AND2_X1 U5122 ( .A1(n4685), .A2(D_REG_28__SCAN_IN), .ZN(U3294) );
  INV_X1 U5123 ( .A(D_REG_27__SCAN_IN), .ZN(n4794) );
  NOR2_X1 U5124 ( .A1(n4605), .A2(n4794), .ZN(U3295) );
  AND2_X1 U5125 ( .A1(D_REG_26__SCAN_IN), .A2(n4685), .ZN(U3296) );
  AND2_X1 U5126 ( .A1(D_REG_25__SCAN_IN), .A2(n4685), .ZN(U3297) );
  AND2_X1 U5127 ( .A1(D_REG_24__SCAN_IN), .A2(n4685), .ZN(U3298) );
  AND2_X1 U5128 ( .A1(D_REG_23__SCAN_IN), .A2(n4685), .ZN(U3299) );
  INV_X1 U5129 ( .A(D_REG_22__SCAN_IN), .ZN(n4922) );
  NOR2_X1 U5130 ( .A1(n4605), .A2(n4922), .ZN(U3300) );
  AND2_X1 U5131 ( .A1(D_REG_21__SCAN_IN), .A2(n4685), .ZN(U3301) );
  AND2_X1 U5132 ( .A1(D_REG_20__SCAN_IN), .A2(n4685), .ZN(U3302) );
  AND2_X1 U5133 ( .A1(n4685), .A2(D_REG_19__SCAN_IN), .ZN(U3303) );
  AND2_X1 U5134 ( .A1(D_REG_18__SCAN_IN), .A2(n4685), .ZN(U3304) );
  AND2_X1 U5135 ( .A1(D_REG_17__SCAN_IN), .A2(n4685), .ZN(U3305) );
  AND2_X1 U5136 ( .A1(D_REG_16__SCAN_IN), .A2(n4685), .ZN(U3306) );
  INV_X1 U5137 ( .A(D_REG_15__SCAN_IN), .ZN(n4791) );
  NOR2_X1 U5138 ( .A1(n4605), .A2(n4791), .ZN(U3307) );
  INV_X1 U5139 ( .A(D_REG_14__SCAN_IN), .ZN(n4942) );
  NOR2_X1 U5140 ( .A1(n4605), .A2(n4942), .ZN(U3308) );
  AND2_X1 U5141 ( .A1(n4685), .A2(D_REG_13__SCAN_IN), .ZN(U3309) );
  AND2_X1 U5142 ( .A1(D_REG_12__SCAN_IN), .A2(n4685), .ZN(U3310) );
  INV_X1 U5143 ( .A(D_REG_10__SCAN_IN), .ZN(n4792) );
  NOR2_X1 U5144 ( .A1(n4605), .A2(n4792), .ZN(U3312) );
  AND2_X1 U5145 ( .A1(n4685), .A2(D_REG_9__SCAN_IN), .ZN(U3313) );
  AND2_X1 U5146 ( .A1(D_REG_8__SCAN_IN), .A2(n4685), .ZN(U3314) );
  AND2_X1 U5147 ( .A1(n4685), .A2(D_REG_7__SCAN_IN), .ZN(U3315) );
  AND2_X1 U5148 ( .A1(D_REG_6__SCAN_IN), .A2(n4685), .ZN(U3316) );
  AND2_X1 U5149 ( .A1(D_REG_5__SCAN_IN), .A2(n4685), .ZN(U3317) );
  INV_X1 U5150 ( .A(D_REG_4__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5151 ( .A1(n4605), .A2(n4779), .ZN(U3318) );
  AND2_X1 U5152 ( .A1(D_REG_3__SCAN_IN), .A2(n4685), .ZN(U3319) );
  INV_X1 U5153 ( .A(D_REG_2__SCAN_IN), .ZN(n4783) );
  NOR2_X1 U5154 ( .A1(n4605), .A2(n4783), .ZN(U3320) );
  OAI21_X1 U5155 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4606), .ZN(
        n4607) );
  INV_X1 U5156 ( .A(n4607), .ZN(U3329) );
  AOI22_X1 U5157 ( .A1(STATE_REG_SCAN_IN), .A2(n4608), .B1(n2513), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5158 ( .A1(U3149), .A2(n4609), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4610) );
  INV_X1 U5159 ( .A(n4610), .ZN(U3335) );
  INV_X1 U5160 ( .A(DATAI_16_), .ZN(n4611) );
  AOI22_X1 U5161 ( .A1(STATE_REG_SCAN_IN), .A2(n4612), .B1(n4611), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5162 ( .A1(U3149), .A2(n4613), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4614) );
  INV_X1 U5163 ( .A(n4614), .ZN(U3337) );
  OAI22_X1 U5164 ( .A1(U3149), .A2(n4615), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4616) );
  INV_X1 U5165 ( .A(n4616), .ZN(U3339) );
  OAI22_X1 U5166 ( .A1(U3149), .A2(n4617), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4618) );
  INV_X1 U5167 ( .A(n4618), .ZN(U3342) );
  INV_X1 U5168 ( .A(DATAI_9_), .ZN(n4619) );
  AOI22_X1 U5169 ( .A1(STATE_REG_SCAN_IN), .A2(n4620), .B1(n4619), .B2(U3149), 
        .ZN(U3343) );
  OAI22_X1 U5170 ( .A1(U3149), .A2(n4621), .B1(DATAI_8_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4622) );
  INV_X1 U5171 ( .A(n4622), .ZN(U3344) );
  INV_X1 U5172 ( .A(DATAI_6_), .ZN(n4866) );
  AOI22_X1 U5173 ( .A1(STATE_REG_SCAN_IN), .A2(n4623), .B1(n4866), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5174 ( .A1(STATE_REG_SCAN_IN), .A2(n2344), .B1(n2343), .B2(U3149), 
        .ZN(U3352) );
  NOR2_X1 U5175 ( .A1(n4624), .A2(n4668), .ZN(n4627) );
  INV_X1 U5176 ( .A(n4625), .ZN(n4626) );
  AOI211_X1 U5177 ( .C1(n4629), .C2(n4628), .A(n4627), .B(n4626), .ZN(n4674)
         );
  INV_X1 U5178 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U5179 ( .A1(n4673), .A2(n4674), .B1(n4630), .B2(n4672), .ZN(U3467)
         );
  NOR2_X1 U5180 ( .A1(n4631), .A2(n4668), .ZN(n4633) );
  AOI211_X1 U5181 ( .C1(n2598), .C2(n4634), .A(n4633), .B(n4632), .ZN(n4675)
         );
  INV_X1 U5182 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5183 ( .A1(n4673), .A2(n4675), .B1(n4635), .B2(n4672), .ZN(U3469)
         );
  NOR3_X1 U5184 ( .A1(n4637), .A2(n4636), .A3(n3251), .ZN(n4639) );
  AOI211_X1 U5185 ( .C1(n4649), .C2(n4640), .A(n4639), .B(n4638), .ZN(n4676)
         );
  INV_X1 U5186 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4880) );
  AOI22_X1 U5187 ( .A1(n4673), .A2(n4676), .B1(n4880), .B2(n4672), .ZN(U3471)
         );
  NOR2_X1 U5188 ( .A1(n4641), .A2(n3251), .ZN(n4642) );
  AOI21_X1 U5189 ( .B1(n4643), .B2(n4649), .A(n4642), .ZN(n4644) );
  AND2_X1 U5190 ( .A1(n4645), .A2(n4644), .ZN(n4677) );
  INV_X1 U5191 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U5192 ( .A1(n4673), .A2(n4677), .B1(n4646), .B2(n4672), .ZN(U3473)
         );
  AOI211_X1 U5193 ( .C1(n4650), .C2(n4649), .A(n4648), .B(n4647), .ZN(n4678)
         );
  INV_X1 U5194 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4651) );
  AOI22_X1 U5195 ( .A1(n4673), .A2(n4678), .B1(n4651), .B2(n4672), .ZN(U3475)
         );
  OAI21_X1 U5196 ( .B1(n3251), .B2(n4653), .A(n4652), .ZN(n4654) );
  AOI21_X1 U5197 ( .B1(n4655), .B2(n4656), .A(n4654), .ZN(n4679) );
  INV_X1 U5198 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U5199 ( .A1(n4673), .A2(n4679), .B1(n4973), .B2(n4672), .ZN(U3477)
         );
  NAND2_X1 U5200 ( .A1(n4657), .A2(n4656), .ZN(n4659) );
  AND3_X1 U5201 ( .A1(n4660), .A2(n4659), .A3(n4658), .ZN(n4680) );
  INV_X1 U5202 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U5203 ( .A1(n4673), .A2(n4680), .B1(n4863), .B2(n4672), .ZN(U3481)
         );
  NOR2_X1 U5204 ( .A1(n4662), .A2(n4661), .ZN(n4663) );
  AOI211_X1 U5205 ( .C1(n2598), .C2(n4665), .A(n4664), .B(n4663), .ZN(n4681)
         );
  INV_X1 U5206 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5207 ( .A1(n4673), .A2(n4681), .B1(n4666), .B2(n4672), .ZN(U3485)
         );
  OAI22_X1 U5208 ( .A1(n4669), .A2(n4668), .B1(n3251), .B2(n4667), .ZN(n4670)
         );
  NOR2_X1 U5209 ( .A1(n4671), .A2(n4670), .ZN(n4683) );
  INV_X1 U5210 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U5211 ( .A1(n4673), .A2(n4683), .B1(n4797), .B2(n4672), .ZN(U3489)
         );
  AOI22_X1 U5212 ( .A1(n4684), .A2(n4674), .B1(n2611), .B2(n4682), .ZN(U3518)
         );
  AOI22_X1 U5213 ( .A1(n4684), .A2(n4675), .B1(n3145), .B2(n4682), .ZN(U3519)
         );
  AOI22_X1 U5214 ( .A1(n4684), .A2(n4676), .B1(n3147), .B2(n4682), .ZN(U3520)
         );
  INV_X1 U5215 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U5216 ( .A1(n4684), .A2(n4677), .B1(n4860), .B2(n4682), .ZN(U3521)
         );
  AOI22_X1 U5217 ( .A1(n4684), .A2(n4678), .B1(n3168), .B2(n4682), .ZN(U3522)
         );
  AOI22_X1 U5218 ( .A1(n4684), .A2(n4679), .B1(n4952), .B2(n4682), .ZN(U3523)
         );
  AOI22_X1 U5219 ( .A1(n4684), .A2(n4680), .B1(n2371), .B2(n4682), .ZN(U3525)
         );
  INV_X1 U5220 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4890) );
  AOI22_X1 U5221 ( .A1(n4684), .A2(n4681), .B1(n4890), .B2(n4682), .ZN(U3527)
         );
  AOI22_X1 U5222 ( .A1(n4684), .A2(n4683), .B1(n3504), .B2(n4682), .ZN(U3529)
         );
  NAND2_X1 U5223 ( .A1(n4685), .A2(D_REG_11__SCAN_IN), .ZN(n5075) );
  AOI22_X1 U5224 ( .A1(DATAI_19_), .A2(keyinput244), .B1(DATAI_22_), .B2(
        keyinput154), .ZN(n4686) );
  OAI221_X1 U5225 ( .B1(DATAI_19_), .B2(keyinput244), .C1(DATAI_22_), .C2(
        keyinput154), .A(n4686), .ZN(n4693) );
  AOI22_X1 U5226 ( .A1(DATAI_18_), .A2(keyinput176), .B1(DATAI_14_), .B2(
        keyinput246), .ZN(n4687) );
  OAI221_X1 U5227 ( .B1(DATAI_18_), .B2(keyinput176), .C1(DATAI_14_), .C2(
        keyinput246), .A(n4687), .ZN(n4692) );
  AOI22_X1 U5228 ( .A1(DATAI_12_), .A2(keyinput129), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput234), .ZN(n4688) );
  OAI221_X1 U5229 ( .B1(DATAI_12_), .B2(keyinput129), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput234), .A(n4688), .ZN(n4691) );
  AOI22_X1 U5230 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput187), .B1(
        REG3_REG_23__SCAN_IN), .B2(keyinput133), .ZN(n4689) );
  OAI221_X1 U5231 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput187), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput133), .A(n4689), .ZN(n4690) );
  NOR4_X1 U5232 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4721)
         );
  AOI22_X1 U5233 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput245), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput232), .ZN(n4694) );
  OAI221_X1 U5234 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput245), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput232), .A(n4694), .ZN(n4701) );
  AOI22_X1 U5235 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput134), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput145), .ZN(n4695) );
  OAI221_X1 U5236 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput134), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput145), .A(n4695), .ZN(n4700) );
  AOI22_X1 U5237 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput144), .B1(
        REG3_REG_13__SCAN_IN), .B2(keyinput236), .ZN(n4696) );
  OAI221_X1 U5238 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput144), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput236), .A(n4696), .ZN(n4699) );
  AOI22_X1 U5239 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput132), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput166), .ZN(n4697) );
  OAI221_X1 U5240 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput132), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput166), .A(n4697), .ZN(n4698) );
  NOR4_X1 U5241 ( .A1(n4701), .A2(n4700), .A3(n4699), .A4(n4698), .ZN(n4720)
         );
  AOI22_X1 U5242 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput170), .B1(
        IR_REG_11__SCAN_IN), .B2(keyinput182), .ZN(n4702) );
  OAI221_X1 U5243 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput170), .C1(
        IR_REG_11__SCAN_IN), .C2(keyinput182), .A(n4702), .ZN(n4709) );
  AOI22_X1 U5244 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput214), .B1(
        IR_REG_19__SCAN_IN), .B2(keyinput137), .ZN(n4703) );
  OAI221_X1 U5245 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput214), .C1(
        IR_REG_19__SCAN_IN), .C2(keyinput137), .A(n4703), .ZN(n4708) );
  AOI22_X1 U5246 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput146), .B1(
        IR_REG_24__SCAN_IN), .B2(keyinput228), .ZN(n4704) );
  OAI221_X1 U5247 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput146), .C1(
        IR_REG_24__SCAN_IN), .C2(keyinput228), .A(n4704), .ZN(n4707) );
  AOI22_X1 U5248 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput223), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput230), .ZN(n4705) );
  OAI221_X1 U5249 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput223), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput230), .A(n4705), .ZN(n4706) );
  NOR4_X1 U5250 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(n4719)
         );
  AOI22_X1 U5251 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput222), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput253), .ZN(n4710) );
  OAI221_X1 U5252 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput222), .C1(
        D_REG_13__SCAN_IN), .C2(keyinput253), .A(n4710), .ZN(n4717) );
  AOI22_X1 U5253 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput209), .B1(
        D_REG_19__SCAN_IN), .B2(keyinput212), .ZN(n4711) );
  OAI221_X1 U5254 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput209), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput212), .A(n4711), .ZN(n4716) );
  AOI22_X1 U5255 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput243), .B1(
        D_REG_28__SCAN_IN), .B2(keyinput250), .ZN(n4712) );
  OAI221_X1 U5256 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput243), .C1(
        D_REG_28__SCAN_IN), .C2(keyinput250), .A(n4712), .ZN(n4715) );
  AOI22_X1 U5257 ( .A1(REG0_REG_2__SCAN_IN), .A2(keyinput198), .B1(
        REG0_REG_5__SCAN_IN), .B2(keyinput148), .ZN(n4713) );
  OAI221_X1 U5258 ( .B1(REG0_REG_2__SCAN_IN), .B2(keyinput198), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput148), .A(n4713), .ZN(n4714) );
  NOR4_X1 U5259 ( .A1(n4717), .A2(n4716), .A3(n4715), .A4(n4714), .ZN(n4718)
         );
  NAND4_X1 U5260 ( .A1(n4721), .A2(n4720), .A3(n4719), .A4(n4718), .ZN(n4857)
         );
  AOI22_X1 U5261 ( .A1(REG0_REG_19__SCAN_IN), .A2(keyinput217), .B1(
        REG0_REG_20__SCAN_IN), .B2(keyinput204), .ZN(n4722) );
  OAI221_X1 U5262 ( .B1(REG0_REG_19__SCAN_IN), .B2(keyinput217), .C1(
        REG0_REG_20__SCAN_IN), .C2(keyinput204), .A(n4722), .ZN(n4729) );
  AOI22_X1 U5263 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput174), .B1(
        REG0_REG_28__SCAN_IN), .B2(keyinput162), .ZN(n4723) );
  OAI221_X1 U5264 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput174), .C1(
        REG0_REG_28__SCAN_IN), .C2(keyinput162), .A(n4723), .ZN(n4728) );
  AOI22_X1 U5265 ( .A1(REG1_REG_5__SCAN_IN), .A2(keyinput164), .B1(
        REG1_REG_9__SCAN_IN), .B2(keyinput179), .ZN(n4724) );
  OAI221_X1 U5266 ( .B1(REG1_REG_5__SCAN_IN), .B2(keyinput164), .C1(
        REG1_REG_9__SCAN_IN), .C2(keyinput179), .A(n4724), .ZN(n4727) );
  AOI22_X1 U5267 ( .A1(REG1_REG_12__SCAN_IN), .A2(keyinput199), .B1(
        REG1_REG_19__SCAN_IN), .B2(keyinput172), .ZN(n4725) );
  OAI221_X1 U5268 ( .B1(REG1_REG_12__SCAN_IN), .B2(keyinput199), .C1(
        REG1_REG_19__SCAN_IN), .C2(keyinput172), .A(n4725), .ZN(n4726) );
  NOR4_X1 U5269 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4757)
         );
  AOI22_X1 U5270 ( .A1(REG1_REG_30__SCAN_IN), .A2(keyinput165), .B1(
        REG1_REG_25__SCAN_IN), .B2(keyinput221), .ZN(n4730) );
  OAI221_X1 U5271 ( .B1(REG1_REG_30__SCAN_IN), .B2(keyinput165), .C1(
        REG1_REG_25__SCAN_IN), .C2(keyinput221), .A(n4730), .ZN(n4737) );
  AOI22_X1 U5272 ( .A1(REG2_REG_0__SCAN_IN), .A2(keyinput171), .B1(
        REG2_REG_2__SCAN_IN), .B2(keyinput169), .ZN(n4731) );
  OAI221_X1 U5273 ( .B1(REG2_REG_0__SCAN_IN), .B2(keyinput171), .C1(
        REG2_REG_2__SCAN_IN), .C2(keyinput169), .A(n4731), .ZN(n4736) );
  AOI22_X1 U5274 ( .A1(REG2_REG_11__SCAN_IN), .A2(keyinput143), .B1(
        REG2_REG_10__SCAN_IN), .B2(keyinput140), .ZN(n4732) );
  OAI221_X1 U5275 ( .B1(REG2_REG_11__SCAN_IN), .B2(keyinput143), .C1(
        REG2_REG_10__SCAN_IN), .C2(keyinput140), .A(n4732), .ZN(n4735) );
  AOI22_X1 U5276 ( .A1(REG2_REG_12__SCAN_IN), .A2(keyinput160), .B1(
        REG2_REG_17__SCAN_IN), .B2(keyinput197), .ZN(n4733) );
  OAI221_X1 U5277 ( .B1(REG2_REG_12__SCAN_IN), .B2(keyinput160), .C1(
        REG2_REG_17__SCAN_IN), .C2(keyinput197), .A(n4733), .ZN(n4734) );
  NOR4_X1 U5278 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4756)
         );
  AOI22_X1 U5279 ( .A1(REG2_REG_18__SCAN_IN), .A2(keyinput157), .B1(
        REG2_REG_22__SCAN_IN), .B2(keyinput219), .ZN(n4738) );
  OAI221_X1 U5280 ( .B1(REG2_REG_18__SCAN_IN), .B2(keyinput157), .C1(
        REG2_REG_22__SCAN_IN), .C2(keyinput219), .A(n4738), .ZN(n4745) );
  AOI22_X1 U5281 ( .A1(REG2_REG_31__SCAN_IN), .A2(keyinput185), .B1(
        REG2_REG_20__SCAN_IN), .B2(keyinput150), .ZN(n4739) );
  OAI221_X1 U5282 ( .B1(REG2_REG_31__SCAN_IN), .B2(keyinput185), .C1(
        REG2_REG_20__SCAN_IN), .C2(keyinput150), .A(n4739), .ZN(n4744) );
  AOI22_X1 U5283 ( .A1(ADDR_REG_12__SCAN_IN), .A2(keyinput194), .B1(
        ADDR_REG_13__SCAN_IN), .B2(keyinput130), .ZN(n4740) );
  OAI221_X1 U5284 ( .B1(ADDR_REG_12__SCAN_IN), .B2(keyinput194), .C1(
        ADDR_REG_13__SCAN_IN), .C2(keyinput130), .A(n4740), .ZN(n4743) );
  AOI22_X1 U5285 ( .A1(ADDR_REG_7__SCAN_IN), .A2(keyinput163), .B1(
        ADDR_REG_9__SCAN_IN), .B2(keyinput192), .ZN(n4741) );
  OAI221_X1 U5286 ( .B1(ADDR_REG_7__SCAN_IN), .B2(keyinput163), .C1(
        ADDR_REG_9__SCAN_IN), .C2(keyinput192), .A(n4741), .ZN(n4742) );
  NOR4_X1 U5287 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4755)
         );
  AOI22_X1 U5288 ( .A1(ADDR_REG_0__SCAN_IN), .A2(keyinput195), .B1(
        ADDR_REG_1__SCAN_IN), .B2(keyinput252), .ZN(n4746) );
  OAI221_X1 U5289 ( .B1(ADDR_REG_0__SCAN_IN), .B2(keyinput195), .C1(
        ADDR_REG_1__SCAN_IN), .C2(keyinput252), .A(n4746), .ZN(n4753) );
  AOI22_X1 U5290 ( .A1(DATAO_REG_13__SCAN_IN), .A2(keyinput211), .B1(
        DATAO_REG_2__SCAN_IN), .B2(keyinput184), .ZN(n4747) );
  OAI221_X1 U5291 ( .B1(DATAO_REG_13__SCAN_IN), .B2(keyinput211), .C1(
        DATAO_REG_2__SCAN_IN), .C2(keyinput184), .A(n4747), .ZN(n4752) );
  AOI22_X1 U5292 ( .A1(DATAO_REG_16__SCAN_IN), .A2(keyinput251), .B1(
        DATAO_REG_28__SCAN_IN), .B2(keyinput191), .ZN(n4748) );
  OAI221_X1 U5293 ( .B1(DATAO_REG_16__SCAN_IN), .B2(keyinput251), .C1(
        DATAO_REG_28__SCAN_IN), .C2(keyinput191), .A(n4748), .ZN(n4751) );
  AOI22_X1 U5294 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput152), .B1(
        DATAO_REG_25__SCAN_IN), .B2(keyinput151), .ZN(n4749) );
  OAI221_X1 U5295 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput152), .C1(
        DATAO_REG_25__SCAN_IN), .C2(keyinput151), .A(n4749), .ZN(n4750) );
  NOR4_X1 U5296 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(n4754)
         );
  NAND4_X1 U5297 ( .A1(n4757), .A2(n4756), .A3(n4755), .A4(n4754), .ZN(n4856)
         );
  AOI22_X1 U5298 ( .A1(DATAO_REG_30__SCAN_IN), .A2(keyinput183), .B1(
        REG3_REG_6__SCAN_IN), .B2(keyinput226), .ZN(n4758) );
  OAI221_X1 U5299 ( .B1(DATAO_REG_30__SCAN_IN), .B2(keyinput183), .C1(
        REG3_REG_6__SCAN_IN), .C2(keyinput226), .A(n4758), .ZN(n4766) );
  AOI22_X1 U5300 ( .A1(ADDR_REG_11__SCAN_IN), .A2(keyinput240), .B1(
        ADDR_REG_19__SCAN_IN), .B2(keyinput229), .ZN(n4759) );
  OAI221_X1 U5301 ( .B1(ADDR_REG_11__SCAN_IN), .B2(keyinput240), .C1(
        ADDR_REG_19__SCAN_IN), .C2(keyinput229), .A(n4759), .ZN(n4765) );
  AOI22_X1 U5302 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput136), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput147), .ZN(n4760) );
  OAI221_X1 U5303 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput136), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput147), .A(n4760), .ZN(n4764) );
  INV_X1 U5304 ( .A(DATAI_30_), .ZN(n5040) );
  INV_X1 U5305 ( .A(DATAI_26_), .ZN(n4762) );
  AOI22_X1 U5306 ( .A1(n5040), .A2(keyinput248), .B1(n4762), .B2(keyinput238), 
        .ZN(n4761) );
  OAI221_X1 U5307 ( .B1(n5040), .B2(keyinput248), .C1(n4762), .C2(keyinput238), 
        .A(n4761), .ZN(n4763) );
  NOR4_X1 U5308 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n4805)
         );
  AOI22_X1 U5309 ( .A1(n4866), .A2(keyinput247), .B1(keyinput135), .B2(n2343), 
        .ZN(n4767) );
  OAI221_X1 U5310 ( .B1(n4866), .B2(keyinput247), .C1(n2343), .C2(keyinput135), 
        .A(n4767), .ZN(n4777) );
  INV_X1 U5311 ( .A(DATAI_11_), .ZN(n4770) );
  INV_X1 U5312 ( .A(DATAI_5_), .ZN(n4769) );
  AOI22_X1 U5313 ( .A1(n4770), .A2(keyinput235), .B1(n4769), .B2(keyinput201), 
        .ZN(n4768) );
  OAI221_X1 U5314 ( .B1(n4770), .B2(keyinput235), .C1(n4769), .C2(keyinput201), 
        .A(n4768), .ZN(n4776) );
  INV_X1 U5315 ( .A(DATAI_4_), .ZN(n4972) );
  AOI22_X1 U5316 ( .A1(n4972), .A2(keyinput156), .B1(n4892), .B2(keyinput186), 
        .ZN(n4771) );
  OAI221_X1 U5317 ( .B1(n4972), .B2(keyinput156), .C1(n4892), .C2(keyinput186), 
        .A(n4771), .ZN(n4775) );
  XNOR2_X1 U5318 ( .A(IR_REG_1__SCAN_IN), .B(keyinput167), .ZN(n4773) );
  XNOR2_X1 U5319 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput189), .ZN(n4772) );
  NAND2_X1 U5320 ( .A1(n4773), .A2(n4772), .ZN(n4774) );
  NOR4_X1 U5321 ( .A1(n4777), .A2(n4776), .A3(n4775), .A4(n4774), .ZN(n4804)
         );
  AOI22_X1 U5322 ( .A1(n4925), .A2(keyinput131), .B1(keyinput208), .B2(n4779), 
        .ZN(n4778) );
  OAI221_X1 U5323 ( .B1(n4925), .B2(keyinput131), .C1(n4779), .C2(keyinput208), 
        .A(n4778), .ZN(n4789) );
  AOI22_X1 U5324 ( .A1(n4781), .A2(keyinput142), .B1(keyinput177), .B2(n2505), 
        .ZN(n4780) );
  OAI221_X1 U5325 ( .B1(n4781), .B2(keyinput142), .C1(n2505), .C2(keyinput177), 
        .A(n4780), .ZN(n4788) );
  AOI22_X1 U5326 ( .A1(n2297), .A2(keyinput141), .B1(keyinput216), .B2(n4783), 
        .ZN(n4782) );
  OAI221_X1 U5327 ( .B1(n2297), .B2(keyinput141), .C1(n4783), .C2(keyinput216), 
        .A(n4782), .ZN(n4787) );
  XOR2_X1 U5328 ( .A(n2454), .B(keyinput149), .Z(n4785) );
  XNOR2_X1 U5329 ( .A(IR_REG_12__SCAN_IN), .B(keyinput239), .ZN(n4784) );
  NAND2_X1 U5330 ( .A1(n4785), .A2(n4784), .ZN(n4786) );
  NOR4_X1 U5331 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(n4803)
         );
  AOI22_X1 U5332 ( .A1(n4792), .A2(keyinput128), .B1(keyinput213), .B2(n4791), 
        .ZN(n4790) );
  OAI221_X1 U5333 ( .B1(n4792), .B2(keyinput128), .C1(n4791), .C2(keyinput213), 
        .A(n4790), .ZN(n4801) );
  AOI22_X1 U5334 ( .A1(n4794), .A2(keyinput241), .B1(keyinput139), .B2(n4922), 
        .ZN(n4793) );
  OAI221_X1 U5335 ( .B1(n4794), .B2(keyinput241), .C1(n4922), .C2(keyinput139), 
        .A(n4793), .ZN(n4800) );
  AOI22_X1 U5336 ( .A1(n4906), .A2(keyinput158), .B1(keyinput255), .B2(n4863), 
        .ZN(n4795) );
  OAI221_X1 U5337 ( .B1(n4906), .B2(keyinput158), .C1(n4863), .C2(keyinput255), 
        .A(n4795), .ZN(n4799) );
  AOI22_X1 U5338 ( .A1(n4977), .A2(keyinput237), .B1(keyinput173), .B2(n4797), 
        .ZN(n4796) );
  OAI221_X1 U5339 ( .B1(n4977), .B2(keyinput237), .C1(n4797), .C2(keyinput173), 
        .A(n4796), .ZN(n4798) );
  NOR4_X1 U5340 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n4802)
         );
  NAND4_X1 U5341 ( .A1(n4805), .A2(n4804), .A3(n4803), .A4(n4802), .ZN(n4855)
         );
  INV_X1 U5342 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4923) );
  INV_X1 U5343 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4910) );
  AOI22_X1 U5344 ( .A1(n4923), .A2(keyinput138), .B1(keyinput159), .B2(n4910), 
        .ZN(n4806) );
  OAI221_X1 U5345 ( .B1(n4923), .B2(keyinput138), .C1(n4910), .C2(keyinput159), 
        .A(n4806), .ZN(n4816) );
  INV_X1 U5346 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4938) );
  INV_X1 U5347 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4808) );
  AOI22_X1 U5348 ( .A1(n4938), .A2(keyinput233), .B1(n4808), .B2(keyinput218), 
        .ZN(n4807) );
  OAI221_X1 U5349 ( .B1(n4938), .B2(keyinput233), .C1(n4808), .C2(keyinput218), 
        .A(n4807), .ZN(n4815) );
  INV_X1 U5350 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5351 ( .A1(n3147), .A2(keyinput207), .B1(n4810), .B2(keyinput225), 
        .ZN(n4809) );
  OAI221_X1 U5352 ( .B1(n3147), .B2(keyinput207), .C1(n4810), .C2(keyinput225), 
        .A(n4809), .ZN(n4814) );
  AOI22_X1 U5353 ( .A1(n4860), .A2(keyinput254), .B1(n4812), .B2(keyinput196), 
        .ZN(n4811) );
  OAI221_X1 U5354 ( .B1(n4860), .B2(keyinput254), .C1(n4812), .C2(keyinput196), 
        .A(n4811), .ZN(n4813) );
  NOR4_X1 U5355 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4853)
         );
  AOI22_X1 U5356 ( .A1(n4818), .A2(keyinput202), .B1(n4909), .B2(keyinput155), 
        .ZN(n4817) );
  OAI221_X1 U5357 ( .B1(n4818), .B2(keyinput202), .C1(n4909), .C2(keyinput155), 
        .A(n4817), .ZN(n4825) );
  INV_X1 U5358 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4876) );
  INV_X1 U5359 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4928) );
  AOI22_X1 U5360 ( .A1(n4876), .A2(keyinput206), .B1(keyinput205), .B2(n4928), 
        .ZN(n4819) );
  OAI221_X1 U5361 ( .B1(n4876), .B2(keyinput206), .C1(n4928), .C2(keyinput205), 
        .A(n4819), .ZN(n4824) );
  AOI22_X1 U5362 ( .A1(n3674), .A2(keyinput188), .B1(n4182), .B2(keyinput161), 
        .ZN(n4820) );
  OAI221_X1 U5363 ( .B1(n3674), .B2(keyinput188), .C1(n4182), .C2(keyinput161), 
        .A(n4820), .ZN(n4823) );
  INV_X1 U5364 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4869) );
  AOI22_X1 U5365 ( .A1(n4869), .A2(keyinput227), .B1(n4091), .B2(keyinput231), 
        .ZN(n4821) );
  OAI221_X1 U5366 ( .B1(n4869), .B2(keyinput227), .C1(n4091), .C2(keyinput231), 
        .A(n4821), .ZN(n4822) );
  NOR4_X1 U5367 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n4852)
         );
  INV_X1 U5368 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4827) );
  AOI22_X1 U5369 ( .A1(n4827), .A2(keyinput210), .B1(keyinput224), .B2(n5036), 
        .ZN(n4826) );
  OAI221_X1 U5370 ( .B1(n4827), .B2(keyinput210), .C1(n5036), .C2(keyinput224), 
        .A(n4826), .ZN(n4838) );
  INV_X1 U5371 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4830) );
  INV_X1 U5372 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5373 ( .A1(n4830), .A2(keyinput168), .B1(keyinput153), .B2(n4829), 
        .ZN(n4828) );
  OAI221_X1 U5374 ( .B1(n4830), .B2(keyinput168), .C1(n4829), .C2(keyinput153), 
        .A(n4828), .ZN(n4837) );
  INV_X1 U5375 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4960) );
  AOI22_X1 U5376 ( .A1(n4960), .A2(keyinput180), .B1(keyinput193), .B2(n4931), 
        .ZN(n4831) );
  OAI221_X1 U5377 ( .B1(n4960), .B2(keyinput180), .C1(n4931), .C2(keyinput193), 
        .A(n4831), .ZN(n4836) );
  AOI22_X1 U5378 ( .A1(n4834), .A2(keyinput178), .B1(n4833), .B2(keyinput215), 
        .ZN(n4832) );
  OAI221_X1 U5379 ( .B1(n4834), .B2(keyinput178), .C1(n4833), .C2(keyinput215), 
        .A(n4832), .ZN(n4835) );
  NOR4_X1 U5380 ( .A1(n4838), .A2(n4837), .A3(n4836), .A4(n4835), .ZN(n4851)
         );
  AOI22_X1 U5381 ( .A1(n4841), .A2(keyinput242), .B1(keyinput175), .B2(n4840), 
        .ZN(n4839) );
  OAI221_X1 U5382 ( .B1(n4841), .B2(keyinput242), .C1(n4840), .C2(keyinput175), 
        .A(n4839), .ZN(n4849) );
  AOI22_X1 U5383 ( .A1(n4875), .A2(keyinput203), .B1(keyinput181), .B2(n4843), 
        .ZN(n4842) );
  OAI221_X1 U5384 ( .B1(n4875), .B2(keyinput203), .C1(n4843), .C2(keyinput181), 
        .A(n4842), .ZN(n4848) );
  AOI22_X1 U5385 ( .A1(n4968), .A2(keyinput249), .B1(n5043), .B2(keyinput220), 
        .ZN(n4844) );
  OAI221_X1 U5386 ( .B1(n4968), .B2(keyinput249), .C1(n5043), .C2(keyinput220), 
        .A(n4844), .ZN(n4847) );
  AOI22_X1 U5387 ( .A1(n3774), .A2(keyinput190), .B1(keyinput200), .B2(n5042), 
        .ZN(n4845) );
  OAI221_X1 U5388 ( .B1(n3774), .B2(keyinput190), .C1(n5042), .C2(keyinput200), 
        .A(n4845), .ZN(n4846) );
  NOR4_X1 U5389 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n4850)
         );
  NAND4_X1 U5390 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4854)
         );
  NOR4_X1 U5391 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n5073)
         );
  INV_X1 U5392 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4859) );
  AOI22_X1 U5393 ( .A1(n4860), .A2(keyinput126), .B1(keyinput64), .B2(n4859), 
        .ZN(n4858) );
  OAI221_X1 U5394 ( .B1(n4860), .B2(keyinput126), .C1(n4859), .C2(keyinput64), 
        .A(n4858), .ZN(n4873) );
  AOI22_X1 U5395 ( .A1(n4863), .A2(keyinput127), .B1(keyinput123), .B2(n4862), 
        .ZN(n4861) );
  OAI221_X1 U5396 ( .B1(n4863), .B2(keyinput127), .C1(n4862), .C2(keyinput123), 
        .A(n4861), .ZN(n4872) );
  AOI22_X1 U5397 ( .A1(n4866), .A2(keyinput119), .B1(n4865), .B2(keyinput115), 
        .ZN(n4864) );
  OAI221_X1 U5398 ( .B1(n4866), .B2(keyinput119), .C1(n4865), .C2(keyinput115), 
        .A(n4864), .ZN(n4871) );
  AOI22_X1 U5399 ( .A1(n4869), .A2(keyinput99), .B1(n4868), .B2(keyinput98), 
        .ZN(n4867) );
  OAI221_X1 U5400 ( .B1(n4869), .B2(keyinput99), .C1(n4868), .C2(keyinput98), 
        .A(n4867), .ZN(n4870) );
  NOR4_X1 U5401 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), .ZN(n4920)
         );
  AOI22_X1 U5402 ( .A1(n4876), .A2(keyinput78), .B1(keyinput75), .B2(n4875), 
        .ZN(n4874) );
  OAI221_X1 U5403 ( .B1(n4876), .B2(keyinput78), .C1(n4875), .C2(keyinput75), 
        .A(n4874), .ZN(n4887) );
  AOI22_X1 U5404 ( .A1(n4200), .A2(keyinput91), .B1(keyinput79), .B2(n3147), 
        .ZN(n4877) );
  OAI221_X1 U5405 ( .B1(n4200), .B2(keyinput91), .C1(n3147), .C2(keyinput79), 
        .A(n4877), .ZN(n4886) );
  AOI22_X1 U5406 ( .A1(n4880), .A2(keyinput70), .B1(n4879), .B2(keyinput71), 
        .ZN(n4878) );
  OAI221_X1 U5407 ( .B1(n4880), .B2(keyinput70), .C1(n4879), .C2(keyinput71), 
        .A(n4878), .ZN(n4885) );
  INV_X1 U5408 ( .A(D_REG_11__SCAN_IN), .ZN(n4881) );
  XOR2_X1 U5409 ( .A(keyinput94), .B(n4881), .Z(n4883) );
  XNOR2_X1 U5410 ( .A(IR_REG_27__SCAN_IN), .B(keyinput95), .ZN(n4882) );
  NAND2_X1 U5411 ( .A1(n4883), .A2(n4882), .ZN(n4884) );
  NOR4_X1 U5412 ( .A1(n4887), .A2(n4886), .A3(n4885), .A4(n4884), .ZN(n4919)
         );
  INV_X1 U5413 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4889) );
  AOI22_X1 U5414 ( .A1(n4890), .A2(keyinput51), .B1(n4889), .B2(keyinput46), 
        .ZN(n4888) );
  OAI221_X1 U5415 ( .B1(n4890), .B2(keyinput51), .C1(n4889), .C2(keyinput46), 
        .A(n4888), .ZN(n4902) );
  INV_X1 U5416 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U5417 ( .A1(n4893), .A2(keyinput67), .B1(n4892), .B2(keyinput58), 
        .ZN(n4891) );
  OAI221_X1 U5418 ( .B1(n4893), .B2(keyinput67), .C1(n4892), .C2(keyinput58), 
        .A(n4891), .ZN(n4901) );
  XOR2_X1 U5419 ( .A(n4894), .B(keyinput43), .Z(n4897) );
  XNOR2_X1 U5420 ( .A(IR_REG_11__SCAN_IN), .B(keyinput54), .ZN(n4896) );
  XNOR2_X1 U5421 ( .A(IR_REG_7__SCAN_IN), .B(keyinput38), .ZN(n4895) );
  NAND3_X1 U5422 ( .A1(n4897), .A2(n4896), .A3(n4895), .ZN(n4900) );
  XNOR2_X1 U5423 ( .A(n4898), .B(keyinput55), .ZN(n4899) );
  NOR4_X1 U5424 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), .ZN(n4918)
         );
  AOI22_X1 U5425 ( .A1(n4243), .A2(keyinput22), .B1(keyinput23), .B2(n4904), 
        .ZN(n4903) );
  OAI221_X1 U5426 ( .B1(n4243), .B2(keyinput22), .C1(n4904), .C2(keyinput23), 
        .A(n4903), .ZN(n4916) );
  INV_X1 U5427 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4907) );
  AOI22_X1 U5428 ( .A1(n4907), .A2(keyinput35), .B1(n4906), .B2(keyinput30), 
        .ZN(n4905) );
  OAI221_X1 U5429 ( .B1(n4907), .B2(keyinput35), .C1(n4906), .C2(keyinput30), 
        .A(n4905), .ZN(n4915) );
  AOI22_X1 U5430 ( .A1(n4910), .A2(keyinput31), .B1(n4909), .B2(keyinput27), 
        .ZN(n4908) );
  OAI221_X1 U5431 ( .B1(n4910), .B2(keyinput31), .C1(n4909), .C2(keyinput27), 
        .A(n4908), .ZN(n4914) );
  XNOR2_X1 U5432 ( .A(IR_REG_23__SCAN_IN), .B(keyinput18), .ZN(n4912) );
  XNOR2_X1 U5433 ( .A(keyinput15), .B(REG2_REG_11__SCAN_IN), .ZN(n4911) );
  NAND2_X1 U5434 ( .A1(n4912), .A2(n4911), .ZN(n4913) );
  NOR4_X1 U5435 ( .A1(n4916), .A2(n4915), .A3(n4914), .A4(n4913), .ZN(n4917)
         );
  NAND4_X1 U5436 ( .A1(n4920), .A2(n4919), .A3(n4918), .A4(n4917), .ZN(n5072)
         );
  AOI22_X1 U5437 ( .A1(n4923), .A2(keyinput10), .B1(n4922), .B2(keyinput11), 
        .ZN(n4921) );
  OAI221_X1 U5438 ( .B1(n4923), .B2(keyinput10), .C1(n4922), .C2(keyinput11), 
        .A(n4921), .ZN(n4936) );
  INV_X1 U5439 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U5440 ( .A1(n4926), .A2(keyinput2), .B1(n4925), .B2(keyinput3), 
        .ZN(n4924) );
  OAI221_X1 U5441 ( .B1(n4926), .B2(keyinput2), .C1(n4925), .C2(keyinput3), 
        .A(n4924), .ZN(n4935) );
  INV_X1 U5442 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4929) );
  AOI22_X1 U5443 ( .A1(n4929), .A2(keyinput69), .B1(keyinput77), .B2(n4928), 
        .ZN(n4927) );
  OAI221_X1 U5444 ( .B1(n4929), .B2(keyinput69), .C1(n4928), .C2(keyinput77), 
        .A(n4927), .ZN(n4934) );
  AOI22_X1 U5445 ( .A1(n4932), .A2(keyinput61), .B1(keyinput65), .B2(n4931), 
        .ZN(n4930) );
  OAI221_X1 U5446 ( .B1(n4932), .B2(keyinput61), .C1(n4931), .C2(keyinput65), 
        .A(n4930), .ZN(n4933) );
  NOR4_X1 U5447 ( .A1(n4936), .A2(n4935), .A3(n4934), .A4(n4933), .ZN(n4986)
         );
  INV_X1 U5448 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4939) );
  AOI22_X1 U5449 ( .A1(n4939), .A2(keyinput101), .B1(n4938), .B2(keyinput105), 
        .ZN(n4937) );
  OAI221_X1 U5450 ( .B1(n4939), .B2(keyinput101), .C1(n4938), .C2(keyinput105), 
        .A(n4937), .ZN(n4950) );
  INV_X1 U5451 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U5452 ( .A1(n4942), .A2(keyinput81), .B1(keyinput93), .B2(n4941), 
        .ZN(n4940) );
  OAI221_X1 U5453 ( .B1(n4942), .B2(keyinput81), .C1(n4941), .C2(keyinput93), 
        .A(n4940), .ZN(n4949) );
  AOI22_X1 U5454 ( .A1(n4944), .A2(keyinput57), .B1(n2505), .B2(keyinput49), 
        .ZN(n4943) );
  OAI221_X1 U5455 ( .B1(n4944), .B2(keyinput57), .C1(n2505), .C2(keyinput49), 
        .A(n4943), .ZN(n4948) );
  AOI22_X1 U5456 ( .A1(n2454), .A2(keyinput21), .B1(keyinput5), .B2(n4946), 
        .ZN(n4945) );
  OAI221_X1 U5457 ( .B1(n2454), .B2(keyinput21), .C1(n4946), .C2(keyinput5), 
        .A(n4945), .ZN(n4947) );
  NOR4_X1 U5458 ( .A1(n4950), .A2(n4949), .A3(n4948), .A4(n4947), .ZN(n4985)
         );
  AOI22_X1 U5459 ( .A1(n4953), .A2(keyinput44), .B1(keyinput36), .B2(n4952), 
        .ZN(n4951) );
  OAI221_X1 U5460 ( .B1(n4953), .B2(keyinput44), .C1(n4952), .C2(keyinput36), 
        .A(n4951), .ZN(n4964) );
  INV_X1 U5461 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4956) );
  AOI22_X1 U5462 ( .A1(n4956), .A2(keyinput16), .B1(keyinput24), .B2(n4955), 
        .ZN(n4954) );
  OAI221_X1 U5463 ( .B1(n4956), .B2(keyinput16), .C1(n4955), .C2(keyinput24), 
        .A(n4954), .ZN(n4963) );
  AOI22_X1 U5464 ( .A1(n2513), .A2(keyinput48), .B1(keyinput56), .B2(n4958), 
        .ZN(n4957) );
  OAI221_X1 U5465 ( .B1(n2513), .B2(keyinput48), .C1(n4958), .C2(keyinput56), 
        .A(n4957), .ZN(n4962) );
  AOI22_X1 U5466 ( .A1(n3674), .A2(keyinput60), .B1(keyinput52), .B2(n4960), 
        .ZN(n4959) );
  OAI221_X1 U5467 ( .B1(n3674), .B2(keyinput60), .C1(n4960), .C2(keyinput52), 
        .A(n4959), .ZN(n4961) );
  NOR4_X1 U5468 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n4984)
         );
  INV_X1 U5469 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4966) );
  AOI22_X1 U5470 ( .A1(n4967), .A2(keyinput8), .B1(keyinput12), .B2(n4966), 
        .ZN(n4965) );
  OAI221_X1 U5471 ( .B1(n4967), .B2(keyinput8), .C1(n4966), .C2(keyinput12), 
        .A(n4965), .ZN(n4970) );
  XNOR2_X1 U5472 ( .A(n4968), .B(keyinput121), .ZN(n4969) );
  NOR2_X1 U5473 ( .A1(n4970), .A2(n4969), .ZN(n4982) );
  AOI22_X1 U5474 ( .A1(n4973), .A2(keyinput20), .B1(keyinput28), .B2(n4972), 
        .ZN(n4971) );
  OAI221_X1 U5475 ( .B1(n4973), .B2(keyinput20), .C1(n4972), .C2(keyinput28), 
        .A(n4971), .ZN(n4974) );
  INV_X1 U5476 ( .A(n4974), .ZN(n4981) );
  AOI22_X1 U5477 ( .A1(n4977), .A2(keyinput109), .B1(n4976), .B2(keyinput117), 
        .ZN(n4975) );
  OAI221_X1 U5478 ( .B1(n4977), .B2(keyinput109), .C1(n4976), .C2(keyinput117), 
        .A(n4975), .ZN(n4978) );
  INV_X1 U5479 ( .A(n4978), .ZN(n4980) );
  XNOR2_X1 U5480 ( .A(IR_REG_5__SCAN_IN), .B(keyinput4), .ZN(n4979) );
  AND4_X1 U5481 ( .A1(n4982), .A2(n4981), .A3(n4980), .A4(n4979), .ZN(n4983)
         );
  NAND4_X1 U5482 ( .A1(n4986), .A2(n4985), .A3(n4984), .A4(n4983), .ZN(n5071)
         );
  AOI22_X1 U5483 ( .A1(ADDR_REG_12__SCAN_IN), .A2(keyinput66), .B1(
        REG3_REG_25__SCAN_IN), .B2(keyinput62), .ZN(n4987) );
  OAI221_X1 U5484 ( .B1(ADDR_REG_12__SCAN_IN), .B2(keyinput66), .C1(
        REG3_REG_25__SCAN_IN), .C2(keyinput62), .A(n4987), .ZN(n4994) );
  AOI22_X1 U5485 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput74), .B1(
        IR_REG_15__SCAN_IN), .B2(keyinput86), .ZN(n4988) );
  OAI221_X1 U5486 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput74), .C1(
        IR_REG_15__SCAN_IN), .C2(keyinput86), .A(n4988), .ZN(n4993) );
  AOI22_X1 U5487 ( .A1(DATAI_22_), .A2(keyinput26), .B1(REG0_REG_28__SCAN_IN), 
        .B2(keyinput34), .ZN(n4989) );
  OAI221_X1 U5488 ( .B1(DATAI_22_), .B2(keyinput26), .C1(REG0_REG_28__SCAN_IN), 
        .C2(keyinput34), .A(n4989), .ZN(n4992) );
  AOI22_X1 U5489 ( .A1(DATAO_REG_3__SCAN_IN), .A2(keyinput50), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput42), .ZN(n4990) );
  OAI221_X1 U5490 ( .B1(DATAO_REG_3__SCAN_IN), .B2(keyinput50), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput42), .A(n4990), .ZN(n4991) );
  NOR4_X1 U5491 ( .A1(n4994), .A2(n4993), .A3(n4992), .A4(n4991), .ZN(n5069)
         );
  AOI22_X1 U5492 ( .A1(DATAI_14_), .A2(keyinput118), .B1(D_REG_28__SCAN_IN), 
        .B2(keyinput122), .ZN(n4995) );
  OAI221_X1 U5493 ( .B1(DATAI_14_), .B2(keyinput118), .C1(D_REG_28__SCAN_IN), 
        .C2(keyinput122), .A(n4995), .ZN(n5002) );
  AOI22_X1 U5494 ( .A1(DATAO_REG_10__SCAN_IN), .A2(keyinput114), .B1(DATAI_26_), .B2(keyinput110), .ZN(n4996) );
  OAI221_X1 U5495 ( .B1(DATAO_REG_10__SCAN_IN), .B2(keyinput114), .C1(
        DATAI_26_), .C2(keyinput110), .A(n4996), .ZN(n5001) );
  AOI22_X1 U5496 ( .A1(ADDR_REG_16__SCAN_IN), .A2(keyinput82), .B1(
        REG0_REG_25__SCAN_IN), .B2(keyinput90), .ZN(n4997) );
  OAI221_X1 U5497 ( .B1(ADDR_REG_16__SCAN_IN), .B2(keyinput82), .C1(
        REG0_REG_25__SCAN_IN), .C2(keyinput90), .A(n4997), .ZN(n5000) );
  AOI22_X1 U5498 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput102), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput106), .ZN(n4998) );
  OAI221_X1 U5499 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput102), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput106), .A(n4998), .ZN(n4999) );
  NOR4_X1 U5500 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5068)
         );
  OAI22_X1 U5501 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput9), .B1(keyinput111), 
        .B2(IR_REG_12__SCAN_IN), .ZN(n5003) );
  AOI221_X1 U5502 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput9), .C1(
        IR_REG_12__SCAN_IN), .C2(keyinput111), .A(n5003), .ZN(n5010) );
  OAI22_X1 U5503 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput59), .B1(DATAI_11_), 
        .B2(keyinput107), .ZN(n5004) );
  AOI221_X1 U5504 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput59), .C1(keyinput107), .C2(DATAI_11_), .A(n5004), .ZN(n5009) );
  OAI22_X1 U5505 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput104), .B1(keyinput40), .B2(ADDR_REG_3__SCAN_IN), .ZN(n5005) );
  AOI221_X1 U5506 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput104), .C1(
        ADDR_REG_3__SCAN_IN), .C2(keyinput40), .A(n5005), .ZN(n5008) );
  OAI22_X1 U5507 ( .A1(DATAO_REG_28__SCAN_IN), .A2(keyinput63), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput87), .ZN(n5006) );
  AOI221_X1 U5508 ( .B1(DATAO_REG_28__SCAN_IN), .B2(keyinput63), .C1(
        keyinput87), .C2(DATAO_REG_8__SCAN_IN), .A(n5006), .ZN(n5007) );
  NAND4_X1 U5509 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n5066)
         );
  OAI22_X1 U5510 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput19), .B1(DATAI_0_), .B2(
        keyinput7), .ZN(n5011) );
  AOI221_X1 U5511 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput19), .C1(keyinput7), 
        .C2(DATAI_0_), .A(n5011), .ZN(n5018) );
  OAI22_X1 U5512 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput14), .B1(
        REG3_REG_5__SCAN_IN), .B2(keyinput6), .ZN(n5012) );
  AOI221_X1 U5513 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput14), .C1(keyinput6), 
        .C2(REG3_REG_5__SCAN_IN), .A(n5012), .ZN(n5017) );
  OAI22_X1 U5514 ( .A1(REG2_REG_28__SCAN_IN), .A2(keyinput103), .B1(
        DATAO_REG_13__SCAN_IN), .B2(keyinput83), .ZN(n5013) );
  AOI221_X1 U5515 ( .B1(REG2_REG_28__SCAN_IN), .B2(keyinput103), .C1(
        keyinput83), .C2(DATAO_REG_13__SCAN_IN), .A(n5013), .ZN(n5016) );
  OAI22_X1 U5516 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput39), .B1(
        DATAO_REG_19__SCAN_IN), .B2(keyinput47), .ZN(n5014) );
  AOI221_X1 U5517 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput39), .C1(keyinput47), 
        .C2(DATAO_REG_19__SCAN_IN), .A(n5014), .ZN(n5015) );
  NAND4_X1 U5518 ( .A1(n5018), .A2(n5017), .A3(n5016), .A4(n5015), .ZN(n5065)
         );
  AOI22_X1 U5519 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput113), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput125), .ZN(n5019) );
  OAI221_X1 U5520 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput113), .C1(
        D_REG_13__SCAN_IN), .C2(keyinput125), .A(n5019), .ZN(n5026) );
  AOI22_X1 U5521 ( .A1(DATAO_REG_21__SCAN_IN), .A2(keyinput53), .B1(
        REG0_REG_11__SCAN_IN), .B2(keyinput45), .ZN(n5020) );
  OAI221_X1 U5522 ( .B1(DATAO_REG_21__SCAN_IN), .B2(keyinput53), .C1(
        REG0_REG_11__SCAN_IN), .C2(keyinput45), .A(n5020), .ZN(n5025) );
  AOI22_X1 U5523 ( .A1(ADDR_REG_5__SCAN_IN), .A2(keyinput25), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput17), .ZN(n5021) );
  OAI221_X1 U5524 ( .B1(ADDR_REG_5__SCAN_IN), .B2(keyinput25), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput17), .A(n5021), .ZN(n5024) );
  AOI22_X1 U5525 ( .A1(REG0_REG_19__SCAN_IN), .A2(keyinput89), .B1(
        REG0_REG_29__SCAN_IN), .B2(keyinput97), .ZN(n5022) );
  OAI221_X1 U5526 ( .B1(REG0_REG_19__SCAN_IN), .B2(keyinput89), .C1(
        REG0_REG_29__SCAN_IN), .C2(keyinput97), .A(n5022), .ZN(n5023) );
  NOR4_X1 U5527 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n5063)
         );
  AOI22_X1 U5528 ( .A1(REG1_REG_8__SCAN_IN), .A2(keyinput68), .B1(
        D_REG_10__SCAN_IN), .B2(keyinput0), .ZN(n5027) );
  OAI221_X1 U5529 ( .B1(REG1_REG_8__SCAN_IN), .B2(keyinput68), .C1(
        D_REG_10__SCAN_IN), .C2(keyinput0), .A(n5027), .ZN(n5034) );
  AOI22_X1 U5530 ( .A1(ADDR_REG_1__SCAN_IN), .A2(keyinput124), .B1(
        D_REG_19__SCAN_IN), .B2(keyinput84), .ZN(n5028) );
  OAI221_X1 U5531 ( .B1(ADDR_REG_1__SCAN_IN), .B2(keyinput124), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput84), .A(n5028), .ZN(n5033) );
  AOI22_X1 U5532 ( .A1(DATAI_5_), .A2(keyinput73), .B1(D_REG_15__SCAN_IN), 
        .B2(keyinput85), .ZN(n5029) );
  OAI221_X1 U5533 ( .B1(DATAI_5_), .B2(keyinput73), .C1(D_REG_15__SCAN_IN), 
        .C2(keyinput85), .A(n5029), .ZN(n5032) );
  AOI22_X1 U5534 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput88), .B1(
        D_REG_4__SCAN_IN), .B2(keyinput80), .ZN(n5030) );
  OAI221_X1 U5535 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput88), .C1(
        D_REG_4__SCAN_IN), .C2(keyinput80), .A(n5030), .ZN(n5031) );
  NOR4_X1 U5536 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n5062)
         );
  INV_X1 U5537 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n5037) );
  AOI22_X1 U5538 ( .A1(n5037), .A2(keyinput112), .B1(n5036), .B2(keyinput96), 
        .ZN(n5035) );
  OAI221_X1 U5539 ( .B1(n5037), .B2(keyinput112), .C1(n5036), .C2(keyinput96), 
        .A(n5035), .ZN(n5049) );
  AOI22_X1 U5540 ( .A1(n5040), .A2(keyinput120), .B1(n5039), .B2(keyinput116), 
        .ZN(n5038) );
  OAI221_X1 U5541 ( .B1(n5040), .B2(keyinput120), .C1(n5039), .C2(keyinput116), 
        .A(n5038), .ZN(n5048) );
  AOI22_X1 U5542 ( .A1(n5043), .A2(keyinput92), .B1(keyinput72), .B2(n5042), 
        .ZN(n5041) );
  OAI221_X1 U5543 ( .B1(n5043), .B2(keyinput92), .C1(n5042), .C2(keyinput72), 
        .A(n5041), .ZN(n5047) );
  XNOR2_X1 U5544 ( .A(IR_REG_24__SCAN_IN), .B(keyinput100), .ZN(n5045) );
  XNOR2_X1 U5545 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput108), .ZN(n5044) );
  NAND2_X1 U5546 ( .A1(n5045), .A2(n5044), .ZN(n5046) );
  NOR4_X1 U5547 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .ZN(n5061)
         );
  AOI22_X1 U5548 ( .A1(REG1_REG_30__SCAN_IN), .A2(keyinput37), .B1(
        REG2_REG_2__SCAN_IN), .B2(keyinput41), .ZN(n5050) );
  OAI221_X1 U5549 ( .B1(REG1_REG_30__SCAN_IN), .B2(keyinput37), .C1(
        REG2_REG_2__SCAN_IN), .C2(keyinput41), .A(n5050), .ZN(n5059) );
  AOI22_X1 U5550 ( .A1(DATAI_12_), .A2(keyinput1), .B1(IR_REG_25__SCAN_IN), 
        .B2(keyinput13), .ZN(n5051) );
  OAI221_X1 U5551 ( .B1(DATAI_12_), .B2(keyinput1), .C1(IR_REG_25__SCAN_IN), 
        .C2(keyinput13), .A(n5051), .ZN(n5058) );
  INV_X1 U5552 ( .A(REG2_REG_12__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U5553 ( .A1(n5054), .A2(keyinput32), .B1(n5053), .B2(keyinput76), 
        .ZN(n5052) );
  OAI221_X1 U5554 ( .B1(n5054), .B2(keyinput32), .C1(n5053), .C2(keyinput76), 
        .A(n5052), .ZN(n5057) );
  AOI22_X1 U5555 ( .A1(REG2_REG_18__SCAN_IN), .A2(keyinput29), .B1(
        REG2_REG_23__SCAN_IN), .B2(keyinput33), .ZN(n5055) );
  OAI221_X1 U5556 ( .B1(REG2_REG_18__SCAN_IN), .B2(keyinput29), .C1(
        REG2_REG_23__SCAN_IN), .C2(keyinput33), .A(n5055), .ZN(n5056) );
  NOR4_X1 U5557 ( .A1(n5059), .A2(n5058), .A3(n5057), .A4(n5056), .ZN(n5060)
         );
  NAND4_X1 U5558 ( .A1(n5063), .A2(n5062), .A3(n5061), .A4(n5060), .ZN(n5064)
         );
  NOR3_X1 U5559 ( .A1(n5066), .A2(n5065), .A3(n5064), .ZN(n5067) );
  NAND3_X1 U5560 ( .A1(n5069), .A2(n5068), .A3(n5067), .ZN(n5070) );
  NOR4_X1 U5561 ( .A1(n5073), .A2(n5072), .A3(n5071), .A4(n5070), .ZN(n5074)
         );
  XNOR2_X1 U5562 ( .A(n5075), .B(n5074), .ZN(U3311) );
  CLKBUF_X1 U2473 ( .A(n2692), .Z(n2742) );
  CLKBUF_X1 U2483 ( .A(n2651), .Z(n3207) );
  NAND3_X1 U2598 ( .A1(n2551), .A2(n4388), .A3(n4387), .ZN(n2597) );
endmodule

