

module b22_C_SARLock_k_128_5 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525;

  INV_X4 U7314 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X2 U7315 ( .A1(n9472), .A2(n9471), .ZN(n12837) );
  INV_X1 U7316 ( .A(n14997), .ZN(n13202) );
  XNOR2_X1 U7317 ( .A(n14465), .B(n14466), .ZN(n14467) );
  XNOR2_X1 U7318 ( .A(n14425), .B(n7059), .ZN(n14465) );
  NAND2_X1 U7319 ( .A1(n7060), .A2(n14424), .ZN(n14425) );
  INV_X1 U7320 ( .A(n12423), .ZN(n12456) );
  NAND2_X1 U7321 ( .A1(n10802), .A2(n12764), .ZN(n12229) );
  INV_X2 U7322 ( .A(n6570), .ZN(n6571) );
  INV_X2 U7323 ( .A(n6572), .ZN(n6575) );
  CLKBUF_X2 U7325 ( .A(n9138), .Z(n12056) );
  INV_X1 U7326 ( .A(n9003), .ZN(n7135) );
  OAI211_X1 U7327 ( .C1(n10749), .C2(n6567), .A(n9098), .B(n9097), .ZN(n11015)
         );
  CLKBUF_X2 U7328 ( .A(n8339), .Z(n8654) );
  NAND2_X2 U7329 ( .A1(n9064), .A2(n13186), .ZN(n9121) );
  CLKBUF_X2 U7330 ( .A(n8928), .Z(n6582) );
  INV_X1 U7331 ( .A(n8016), .ZN(n9999) );
  AND2_X1 U7332 ( .A1(n8246), .A2(n13730), .ZN(n8299) );
  CLKBUF_X1 U7333 ( .A(n8745), .Z(n6577) );
  AND2_X1 U7334 ( .A1(n7564), .A2(n7563), .ZN(n7746) );
  INV_X2 U7335 ( .A(n9945), .ZN(n9957) );
  NAND2_X1 U7337 ( .A1(n6566), .A2(n9957), .ZN(n9138) );
  INV_X1 U7338 ( .A(n12059), .ZN(n6572) );
  XNOR2_X1 U7339 ( .A(n12837), .B(n12847), .ZN(n12829) );
  OR2_X1 U7340 ( .A1(n12966), .A2(n9620), .ZN(n9622) );
  INV_X1 U7341 ( .A(n12213), .ZN(n12211) );
  NAND2_X1 U7342 ( .A1(n8653), .A2(n8659), .ZN(n8277) );
  INV_X1 U7343 ( .A(n13915), .ZN(n10610) );
  AND4_X2 U7344 ( .A1(n7686), .A2(n7279), .A3(n7278), .A4(n7277), .ZN(n7795)
         );
  OAI21_X1 U7345 ( .B1(n7552), .B2(n9947), .A(n6787), .ZN(n7549) );
  INV_X1 U7346 ( .A(n15116), .ZN(n7159) );
  INV_X1 U7347 ( .A(n12634), .ZN(n11492) );
  INV_X1 U7348 ( .A(n6572), .ZN(n6574) );
  INV_X1 U7349 ( .A(n9677), .ZN(n7968) );
  INV_X1 U7350 ( .A(n13914), .ZN(n10896) );
  INV_X1 U7351 ( .A(n8009), .ZN(n7699) );
  OAI211_X1 U7352 ( .C1(n8064), .C2(n6956), .A(n6955), .B(n6599), .ZN(n10892)
         );
  OR2_X1 U7353 ( .A1(n14392), .A2(n7918), .ZN(n7647) );
  AOI21_X1 U7355 ( .B1(n12577), .B2(n12862), .A(n12312), .ZN(n12314) );
  INV_X1 U7356 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9056) );
  OR2_X1 U7357 ( .A1(n8634), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U7358 ( .A1(n6788), .A2(n14464), .ZN(n14468) );
  INV_X1 U7359 ( .A(n10803), .ZN(n10777) );
  XNOR2_X1 U7360 ( .A(n9543), .B(n9544), .ZN(n10802) );
  NAND2_X1 U7361 ( .A1(n8647), .A2(n8648), .ZN(n11557) );
  XNOR2_X1 U7362 ( .A(n14467), .B(n14468), .ZN(n15515) );
  OR2_X1 U7363 ( .A1(n9601), .A2(n15122), .ZN(n6565) );
  INV_X1 U7364 ( .A(n9141), .ZN(n6570) );
  XNOR2_X1 U7365 ( .A(n7643), .B(n7642), .ZN(n14653) );
  NAND2_X1 U7366 ( .A1(n7651), .A2(n14400), .ZN(n8009) );
  NOR3_X1 U7367 ( .A1(n14266), .A2(n14265), .A3(n7544), .ZN(n14363) );
  AND2_X1 U7368 ( .A1(n14264), .A2(n14626), .ZN(n7544) );
  OAI21_X2 U7369 ( .B1(n9363), .B2(n9362), .A(n9364), .ZN(n9380) );
  AND2_X1 U7370 ( .A1(n7003), .A2(n7964), .ZN(n8091) );
  INV_X1 U7371 ( .A(n7066), .ZN(n14081) );
  NAND2_X1 U7372 ( .A1(n12431), .A2(n12733), .ZN(n6566) );
  NAND2_X1 U7373 ( .A1(n12431), .A2(n12733), .ZN(n6567) );
  NAND2_X1 U7374 ( .A1(n12431), .A2(n12733), .ZN(n10662) );
  OAI21_X2 U7375 ( .B1(n9829), .B2(n9830), .A(n9828), .ZN(n9834) );
  OAI22_X1 U7376 ( .A1(n12084), .A2(n12083), .B1(n12211), .B2(n12082), .ZN(
        n12085) );
  OR2_X1 U7377 ( .A1(n9060), .A2(n9056), .ZN(n9057) );
  BUF_X4 U7378 ( .A(n7699), .Z(n7757) );
  AND3_X4 U7379 ( .A1(n8373), .A2(n8224), .A3(n8306), .ZN(n8252) );
  AND2_X2 U7380 ( .A1(n8219), .A2(n8218), .ZN(n8373) );
  AND4_X2 U7381 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n8224)
         );
  NOR2_X2 U7382 ( .A1(n14469), .A2(n14470), .ZN(n14471) );
  OAI21_X2 U7383 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9700) );
  NAND4_X2 U7384 ( .A1(n7722), .A2(n7721), .A3(n7720), .A4(n7719), .ZN(n13914)
         );
  NAND2_X1 U7385 ( .A1(n8653), .A2(n8659), .ZN(n6568) );
  NAND2_X1 U7386 ( .A1(n8653), .A2(n8659), .ZN(n6569) );
  BUF_X2 U7387 ( .A(n8277), .Z(n10017) );
  INV_X4 U7388 ( .A(n10017), .ZN(n8529) );
  OAI21_X2 U7389 ( .B1(n12995), .B2(n9617), .A(n12142), .ZN(n12977) );
  NAND2_X2 U7390 ( .A1(n9276), .A2(n12137), .ZN(n12995) );
  NAND2_X2 U7391 ( .A1(n8349), .A2(n8348), .ZN(n14983) );
  NAND2_X4 U7392 ( .A1(n10806), .A2(n10805), .ZN(n10809) );
  NOR2_X2 U7393 ( .A1(n13918), .A2(n10771), .ZN(n9686) );
  NAND2_X2 U7394 ( .A1(n8446), .A2(n8445), .ZN(n14598) );
  NAND2_X4 U7395 ( .A1(n8256), .A2(n8255), .ZN(n13674) );
  XNOR2_X2 U7396 ( .A(n8279), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8246) );
  NAND2_X4 U7397 ( .A1(n9668), .A2(n9667), .ZN(n9835) );
  NAND2_X2 U7398 ( .A1(n9670), .A2(n11532), .ZN(n9668) );
  NOR2_X2 U7399 ( .A1(n10900), .A2(n10899), .ZN(n12443) );
  NOR2_X2 U7400 ( .A1(n10377), .A2(n10376), .ZN(n10900) );
  NAND2_X2 U7401 ( .A1(n7970), .A2(n7969), .ZN(n14325) );
  XNOR2_X2 U7402 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14453) );
  NAND2_X2 U7403 ( .A1(n6624), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9075) );
  OR2_X1 U7404 ( .A1(n8044), .A2(n7112), .ZN(n7675) );
  NAND2_X2 U7405 ( .A1(n7928), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7674) );
  XNOR2_X2 U7406 ( .A(n8092), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8143) );
  NAND2_X2 U7407 ( .A1(n8532), .A2(n8531), .ZN(n13583) );
  INV_X1 U7408 ( .A(n6572), .ZN(n6573) );
  NAND2_X4 U7409 ( .A1(n8275), .A2(n6747), .ZN(n10337) );
  OR2_X2 U7410 ( .A1(n8274), .A2(n9948), .ZN(n8275) );
  NAND2_X2 U7411 ( .A1(n8380), .A2(n8379), .ZN(n15003) );
  XNOR2_X2 U7412 ( .A(n7960), .B(n7946), .ZN(n11461) );
  NAND2_X2 U7413 ( .A1(n7958), .A2(n7945), .ZN(n7960) );
  NOR2_X2 U7415 ( .A1(n14507), .A2(n14506), .ZN(n14649) );
  AND2_X2 U7416 ( .A1(n6742), .A2(n6741), .ZN(n14507) );
  NAND2_X4 U7417 ( .A1(n9902), .A2(n9901), .ZN(n13217) );
  NAND2_X2 U7418 ( .A1(n6569), .A2(n9945), .ZN(n8273) );
  NAND2_X2 U7419 ( .A1(n8358), .A2(n8357), .ZN(n14991) );
  NAND2_X2 U7420 ( .A1(n8430), .A2(n8429), .ZN(n11237) );
  NAND2_X2 U7421 ( .A1(n8474), .A2(n8473), .ZN(n11676) );
  NAND2_X2 U7422 ( .A1(n7137), .A2(n7138), .ZN(n13456) );
  NOR2_X2 U7423 ( .A1(n6743), .A2(n14649), .ZN(n14543) );
  AND2_X2 U7424 ( .A1(n6746), .A2(n6745), .ZN(n6743) );
  NAND2_X1 U7425 ( .A1(n13284), .A2(n13219), .ZN(n13351) );
  OR2_X1 U7426 ( .A1(n12929), .A2(n6633), .ZN(n7182) );
  NOR2_X1 U7427 ( .A1(n12036), .A2(n12035), .ZN(n13191) );
  NAND2_X1 U7428 ( .A1(n11599), .A2(n11598), .ZN(n11731) );
  NAND2_X2 U7429 ( .A1(n9764), .A2(n9749), .ZN(n11830) );
  NAND2_X1 U7430 ( .A1(n7849), .A2(n7848), .ZN(n7034) );
  INV_X2 U7431 ( .A(n15129), .ZN(n6576) );
  INV_X1 U7432 ( .A(n10809), .ZN(n7398) );
  INV_X2 U7433 ( .A(n12635), .ZN(n11266) );
  INV_X1 U7434 ( .A(n15142), .ZN(n10999) );
  INV_X1 U7435 ( .A(n12636), .ZN(n13015) );
  INV_X1 U7436 ( .A(n9835), .ZN(n9827) );
  INV_X2 U7437 ( .A(n8993), .ZN(n8848) );
  NAND2_X2 U7438 ( .A1(n14317), .A2(n12417), .ZN(n10375) );
  CLKBUF_X1 U7439 ( .A(n8745), .Z(n6585) );
  CLKBUF_X2 U7440 ( .A(n12733), .Z(n12725) );
  NOR2_X2 U7441 ( .A1(n11557), .A2(n9024), .ZN(n9035) );
  BUF_X2 U7442 ( .A(n8299), .Z(n6579) );
  INV_X1 U7443 ( .A(n14040), .ZN(n10460) );
  NOR2_X1 U7444 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8227) );
  NAND2_X1 U7445 ( .A1(n9834), .A2(n9833), .ZN(n9836) );
  OR2_X1 U7446 ( .A1(n9042), .A2(n9041), .ZN(n6779) );
  AOI21_X1 U7447 ( .B1(n14060), .B2(n14626), .A(n7044), .ZN(n7043) );
  OR2_X1 U7448 ( .A1(n13103), .A2(n13011), .ZN(n9594) );
  AOI21_X1 U7449 ( .B1(n12314), .B2(n6608), .A(n6718), .ZN(n12316) );
  MUX2_X1 U7450 ( .A(n13109), .B(n13108), .S(n15177), .Z(n13110) );
  MUX2_X1 U7451 ( .A(n13038), .B(n13108), .S(n15192), .Z(n13039) );
  NOR2_X1 U7452 ( .A1(n13459), .A2(n7201), .ZN(n13424) );
  NAND2_X1 U7453 ( .A1(n8633), .A2(n8632), .ZN(n8937) );
  OR2_X1 U7454 ( .A1(n13617), .A2(n8652), .ZN(n8631) );
  NAND2_X1 U7455 ( .A1(n8621), .A2(n8620), .ZN(n13617) );
  NAND2_X1 U7456 ( .A1(n7671), .A2(n7670), .ZN(n7066) );
  NAND2_X1 U7457 ( .A1(n8066), .A2(n8065), .ZN(n14270) );
  OAI211_X1 U7458 ( .C1(n6978), .C2(n8013), .A(n6671), .B(n6772), .ZN(n14126)
         );
  XNOR2_X1 U7459 ( .A(n7668), .B(n7669), .ZN(n13733) );
  NAND2_X1 U7460 ( .A1(n13827), .A2(n13826), .ZN(n13825) );
  NAND2_X1 U7461 ( .A1(n7182), .A2(n7181), .ZN(n12887) );
  AOI21_X1 U7462 ( .B1(n6590), .B2(n6628), .A(n7151), .ZN(n7150) );
  NAND2_X1 U7463 ( .A1(n8052), .A2(n8051), .ZN(n14135) );
  NAND2_X1 U7464 ( .A1(n13755), .A2(n12368), .ZN(n13827) );
  NAND2_X1 U7465 ( .A1(n7162), .A2(n7160), .ZN(n12929) );
  NAND2_X1 U7466 ( .A1(n12197), .A2(n12200), .ZN(n12845) );
  CLKBUF_X1 U7467 ( .A(n14172), .Z(n6770) );
  OAI21_X1 U7468 ( .B1(n7508), .B2(n13191), .A(n7509), .ZN(n7507) );
  AOI21_X1 U7469 ( .B1(n14233), .B2(n14246), .A(n8123), .ZN(n14217) );
  NAND2_X1 U7470 ( .A1(n8569), .A2(n8568), .ZN(n13537) );
  NAND2_X2 U7471 ( .A1(n8003), .A2(n8002), .ZN(n14384) );
  NAND2_X1 U7472 ( .A1(n7999), .A2(n7984), .ZN(n11530) );
  NAND2_X1 U7473 ( .A1(n12005), .A2(n6980), .ZN(n12326) );
  XNOR2_X1 U7474 ( .A(n7610), .B(n15431), .ZN(n8014) );
  NAND3_X1 U7475 ( .A1(n7299), .A2(n7298), .A3(n7300), .ZN(n12005) );
  NAND2_X1 U7476 ( .A1(n11818), .A2(n7415), .ZN(n12281) );
  OAI21_X1 U7477 ( .B1(n11237), .B2(n8441), .A(n8442), .ZN(n11400) );
  AND2_X1 U7478 ( .A1(n6886), .A2(n6885), .ZN(n14634) );
  NAND2_X1 U7479 ( .A1(n8496), .A2(n8495), .ZN(n13687) );
  OR2_X1 U7480 ( .A1(n14617), .A2(n13885), .ZN(n9764) );
  NAND2_X1 U7481 ( .A1(n6755), .A2(n6754), .ZN(n6885) );
  OR2_X1 U7482 ( .A1(n7944), .A2(n10511), .ZN(n7958) );
  NAND2_X1 U7483 ( .A1(n11713), .A2(n7536), .ZN(n11848) );
  NAND2_X1 U7484 ( .A1(n7903), .A2(n7902), .ZN(n14351) );
  NAND2_X1 U7485 ( .A1(n8464), .A2(n8463), .ZN(n14589) );
  NAND2_X1 U7486 ( .A1(n7883), .A2(n7882), .ZN(n14617) );
  NAND2_X1 U7487 ( .A1(n7914), .A2(n7913), .ZN(n7598) );
  NAND2_X1 U7488 ( .A1(n6888), .A2(n14531), .ZN(n14630) );
  NAND2_X1 U7489 ( .A1(n8422), .A2(n8421), .ZN(n14938) );
  NAND2_X1 U7490 ( .A1(n7028), .A2(n7024), .ZN(n7588) );
  NAND2_X1 U7491 ( .A1(n8436), .A2(n8435), .ZN(n11431) );
  NAND2_X1 U7492 ( .A1(n7814), .A2(n7813), .ZN(n11716) );
  NAND2_X1 U7493 ( .A1(n8395), .A2(n8394), .ZN(n10951) );
  AND2_X2 U7494 ( .A1(n6604), .A2(n10599), .ZN(n7209) );
  NAND2_X1 U7495 ( .A1(n7808), .A2(n7807), .ZN(n7810) );
  NAND2_X1 U7496 ( .A1(n6893), .A2(n14474), .ZN(n14476) );
  NOR2_X2 U7497 ( .A1(n10680), .A2(n12754), .ZN(n15080) );
  AND2_X1 U7498 ( .A1(n12091), .A2(n12092), .ZN(n9605) );
  AND2_X1 U7499 ( .A1(n12081), .A2(n12086), .ZN(n13018) );
  MUX2_X1 U7500 ( .A(n9688), .B(n9689), .S(n9835), .Z(n9694) );
  OR2_X2 U7501 ( .A1(n10936), .A2(n10777), .ZN(n12213) );
  NAND4_X1 U7502 ( .A1(n9125), .A2(n9124), .A3(n9123), .A4(n9122), .ZN(n12635)
         );
  BUF_X2 U7503 ( .A(n9835), .Z(n6809) );
  CLKBUF_X3 U7504 ( .A(n9119), .Z(n12061) );
  OR2_X2 U7505 ( .A1(n10021), .A2(P2_U3088), .ZN(n13379) );
  CLKBUF_X1 U7506 ( .A(n9100), .Z(n9244) );
  INV_X4 U7507 ( .A(n10913), .ZN(n12423) );
  INV_X1 U7508 ( .A(n12417), .ZN(n12458) );
  NAND4_X2 U7509 ( .A1(n7693), .A2(n7695), .A3(n7694), .A4(n7696), .ZN(n13918)
         );
  CLKBUF_X2 U7510 ( .A(n7672), .Z(n6584) );
  NAND2_X1 U7511 ( .A1(n7757), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7700) );
  CLKBUF_X1 U7512 ( .A(n10260), .Z(n14254) );
  AND2_X1 U7513 ( .A1(n9061), .A2(n13181), .ZN(n9063) );
  INV_X2 U7514 ( .A(n8274), .ZN(n8958) );
  NAND2_X1 U7515 ( .A1(n8297), .A2(n8296), .ZN(n8750) );
  AND2_X1 U7516 ( .A1(n9383), .A2(n9054), .ZN(n9542) );
  BUF_X2 U7517 ( .A(n7928), .Z(n7741) );
  OR2_X1 U7518 ( .A1(n8149), .A2(n14652), .ZN(n7693) );
  NAND2_X1 U7519 ( .A1(n10262), .A2(n10261), .ZN(n10913) );
  XNOR2_X1 U7520 ( .A(n7487), .B(n8644), .ZN(n8745) );
  MUX2_X1 U7521 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9059), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9061) );
  AND2_X1 U7522 ( .A1(n7649), .A2(n14400), .ZN(n7928) );
  BUF_X2 U7523 ( .A(n8299), .Z(n6580) );
  NAND2_X1 U7524 ( .A1(n8190), .A2(n8183), .ZN(n10262) );
  INV_X1 U7525 ( .A(n7651), .ZN(n7649) );
  NAND2_X2 U7526 ( .A1(n7651), .A2(n7650), .ZN(n8044) );
  OR2_X1 U7527 ( .A1(n9076), .A2(n6861), .ZN(n9058) );
  OR2_X1 U7528 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  INV_X1 U7529 ( .A(n8294), .ZN(n13730) );
  XNOR2_X1 U7530 ( .A(n8096), .B(n8095), .ZN(n11532) );
  XNOR2_X1 U7531 ( .A(n8094), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8150) );
  MUX2_X1 U7532 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8232), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8234) );
  NAND2_X1 U7533 ( .A1(n8152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U7534 ( .A1(n7967), .A2(n8156), .ZN(n14040) );
  XNOR2_X1 U7535 ( .A(n8239), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U7536 ( .A1(n7189), .A2(n7188), .ZN(n9076) );
  XNOR2_X1 U7537 ( .A(n8167), .B(n8166), .ZN(n14414) );
  INV_X1 U7538 ( .A(n14392), .ZN(n14393) );
  XNOR2_X1 U7539 ( .A(n7132), .B(n7648), .ZN(n14400) );
  AND2_X1 U7540 ( .A1(n9218), .A2(n7191), .ZN(n7188) );
  OR2_X1 U7541 ( .A1(n8237), .A2(n13724), .ZN(n8231) );
  NAND2_X1 U7542 ( .A1(n8238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8239) );
  XNOR2_X1 U7543 ( .A(n8528), .B(P2_IR_REG_19__SCAN_IN), .ZN(n11409) );
  NAND2_X2 U7544 ( .A1(n9957), .A2(P3_U3151), .ZN(n14525) );
  NOR2_X1 U7545 ( .A1(n8163), .A2(n7431), .ZN(n14392) );
  AND2_X1 U7546 ( .A1(n8707), .A2(n7483), .ZN(n8237) );
  OAI21_X1 U7547 ( .B1(n8163), .B2(n7433), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7132) );
  NAND2_X1 U7548 ( .A1(n7280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U7549 ( .A1(n14419), .A2(n7054), .ZN(n14452) );
  AND3_X1 U7550 ( .A1(n7638), .A2(n7637), .A3(n7636), .ZN(n8154) );
  AND3_X1 U7551 ( .A1(n7149), .A2(n7148), .A3(n7147), .ZN(n8230) );
  NAND4_X1 U7552 ( .A1(n8227), .A2(n8417), .A3(n8226), .A4(n8225), .ZN(n8526)
         );
  AND2_X1 U7553 ( .A1(n6884), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14454) );
  NOR2_X1 U7554 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8218) );
  NOR2_X1 U7555 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n8219) );
  NOR3_X1 U7556 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n7632) );
  NOR2_X1 U7557 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7277) );
  NOR2_X1 U7558 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7278) );
  NOR2_X1 U7559 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7279) );
  INV_X1 U7560 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8644) );
  INV_X1 U7561 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8726) );
  NOR2_X1 U7562 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n8215) );
  INV_X1 U7563 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8417) );
  INV_X1 U7564 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8523) );
  INV_X1 U7565 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8225) );
  INV_X1 U7566 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8226) );
  XNOR2_X1 U7567 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14451) );
  NOR2_X1 U7568 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n8216) );
  NOR2_X2 U7569 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10681) );
  INV_X4 U7570 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X4 U7571 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7572 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8223) );
  INV_X1 U7573 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9186) );
  OR2_X1 U7574 ( .A1(n14529), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6895) );
  NAND4_X2 U7576 ( .A1(n8331), .A2(n8330), .A3(n8329), .A4(n8328), .ZN(n13378)
         );
  NOR2_X1 U7577 ( .A1(n8882), .A2(n8881), .ZN(n8889) );
  NOR2_X2 U7578 ( .A1(n12800), .A2(n12799), .ZN(n12798) );
  OR2_X1 U7579 ( .A1(n8832), .A2(n8831), .ZN(n6648) );
  INV_X1 U7580 ( .A(n6748), .ZN(n6747) );
  BUF_X8 U7581 ( .A(n9827), .Z(n6578) );
  NAND2_X1 U7582 ( .A1(n9902), .A2(n9901), .ZN(n6581) );
  AOI21_X2 U7583 ( .B1(n12228), .B2(n12227), .A(n12257), .ZN(n12262) );
  XNOR2_X2 U7584 ( .A(n8231), .B(n8236), .ZN(n8653) );
  XNOR2_X1 U7585 ( .A(n10315), .B(n9907), .ZN(n10328) );
  BUF_X4 U7586 ( .A(n8928), .Z(n6583) );
  INV_X1 U7588 ( .A(n8149), .ZN(n7672) );
  NOR2_X2 U7589 ( .A1(n13630), .A2(n13484), .ZN(n13472) );
  NAND2_X1 U7590 ( .A1(n8609), .A2(n8608), .ZN(n13630) );
  NOR2_X2 U7591 ( .A1(n14240), .A2(n14332), .ZN(n7068) );
  XNOR2_X2 U7592 ( .A(n14420), .B(n7050), .ZN(n14460) );
  NAND2_X2 U7593 ( .A1(n7053), .A2(n7051), .ZN(n14420) );
  XNOR2_X1 U7594 ( .A(n14449), .B(n14423), .ZN(n14450) );
  CLKBUF_X2 U7595 ( .A(n14653), .Z(n6586) );
  XNOR2_X2 U7596 ( .A(n14422), .B(n7061), .ZN(n14449) );
  XNOR2_X2 U7597 ( .A(n7641), .B(n7646), .ZN(n14401) );
  NOR2_X2 U7598 ( .A1(n14637), .A2(n6890), .ZN(n14642) );
  NOR2_X1 U7599 ( .A1(n14270), .A2(n14101), .ZN(n7065) );
  NAND2_X1 U7600 ( .A1(n10994), .A2(n6646), .ZN(n11137) );
  OAI21_X1 U7601 ( .B1(n12779), .B2(n12780), .A(n12068), .ZN(n12256) );
  NAND2_X1 U7602 ( .A1(n12447), .A2(n13186), .ZN(n9119) );
  OR2_X1 U7603 ( .A1(n12711), .A2(n12710), .ZN(n12712) );
  AOI21_X1 U7604 ( .B1(n6597), .B2(n12898), .A(n6662), .ZN(n7181) );
  NAND2_X1 U7605 ( .A1(n9151), .A2(n9150), .ZN(n9156) );
  AOI21_X1 U7606 ( .B1(n7284), .B2(n7286), .A(n6639), .ZN(n7281) );
  NAND2_X1 U7607 ( .A1(n12326), .A2(n7284), .ZN(n7282) );
  NAND2_X1 U7608 ( .A1(n11719), .A2(n7301), .ZN(n7300) );
  NOR2_X1 U7609 ( .A1(n7302), .A2(n7303), .ZN(n7301) );
  INV_X1 U7610 ( .A(n11718), .ZN(n7303) );
  NAND2_X1 U7611 ( .A1(n14533), .A2(n14532), .ZN(n14531) );
  NAND2_X1 U7612 ( .A1(n8748), .A2(n14969), .ZN(n8751) );
  INV_X1 U7613 ( .A(n8780), .ZN(n6781) );
  NOR2_X1 U7614 ( .A1(n7932), .A2(n10451), .ZN(n7339) );
  INV_X1 U7615 ( .A(n7822), .ZN(n7578) );
  OAI21_X1 U7616 ( .B1(n7552), .B2(n6928), .A(n6927), .ZN(n7557) );
  NAND2_X1 U7617 ( .A1(n7552), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6927) );
  INV_X1 U7618 ( .A(n12308), .ZN(n7412) );
  INV_X1 U7619 ( .A(n12568), .ZN(n6818) );
  INV_X1 U7620 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9051) );
  NAND2_X1 U7621 ( .A1(n12075), .A2(n12077), .ZN(n10810) );
  OR2_X1 U7622 ( .A1(n13101), .A2(n12792), .ZN(n12224) );
  OR2_X1 U7623 ( .A1(n12816), .A2(n12805), .ZN(n12205) );
  AND2_X1 U7624 ( .A1(n12928), .A2(n9624), .ZN(n7226) );
  NOR2_X1 U7625 ( .A1(n7225), .A2(n6851), .ZN(n6848) );
  INV_X1 U7626 ( .A(n7226), .ZN(n7225) );
  OR2_X1 U7627 ( .A1(n9625), .A2(n12162), .ZN(n12231) );
  NAND2_X1 U7628 ( .A1(n9547), .A2(n6632), .ZN(n7528) );
  INV_X1 U7629 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9054) );
  AND2_X1 U7630 ( .A1(n7526), .A2(n7405), .ZN(n9383) );
  AND2_X1 U7631 ( .A1(n7407), .A2(n7406), .ZN(n7405) );
  AND2_X1 U7632 ( .A1(n9128), .A2(n6840), .ZN(n6839) );
  INV_X1 U7633 ( .A(n7418), .ZN(n7417) );
  INV_X1 U7634 ( .A(n9250), .ZN(n7092) );
  AND2_X1 U7635 ( .A1(n9241), .A2(n9238), .ZN(n7093) );
  INV_X1 U7636 ( .A(n7110), .ZN(n7103) );
  INV_X1 U7637 ( .A(n8680), .ZN(n7460) );
  INV_X1 U7638 ( .A(n13370), .ZN(n11191) );
  AOI21_X1 U7639 ( .B1(n6944), .B2(n6946), .A(n6940), .ZN(n6939) );
  INV_X1 U7640 ( .A(n8135), .ZN(n6940) );
  OR2_X1 U7641 ( .A1(n13815), .A2(n14235), .ZN(n9773) );
  NAND2_X1 U7642 ( .A1(n7266), .A2(n6638), .ZN(n11338) );
  NAND2_X1 U7643 ( .A1(n7627), .A2(n7626), .ZN(n7668) );
  NAND2_X1 U7644 ( .A1(n8076), .A2(n7625), .ZN(n7627) );
  NAND2_X1 U7645 ( .A1(n7013), .A2(n7015), .ZN(n7622) );
  AND2_X1 U7646 ( .A1(n7016), .A2(n15326), .ZN(n7015) );
  NAND2_X1 U7647 ( .A1(n8038), .A2(n6610), .ZN(n7013) );
  OR2_X1 U7648 ( .A1(n7018), .A2(n7017), .ZN(n7016) );
  XNOR2_X1 U7649 ( .A(n7581), .B(SI_11_), .ZN(n7835) );
  OAI21_X1 U7650 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n15296), .A(n14434), .ZN(
        n14480) );
  NAND2_X1 U7651 ( .A1(n6682), .A2(n7398), .ZN(n7397) );
  OR2_X1 U7652 ( .A1(n12263), .A2(n10801), .ZN(n10806) );
  NAND2_X1 U7653 ( .A1(n6587), .A2(n6601), .ZN(n6825) );
  NAND2_X1 U7654 ( .A1(n6830), .A2(n7408), .ZN(n6829) );
  XNOR2_X1 U7655 ( .A(n7398), .B(n10999), .ZN(n11134) );
  NAND2_X1 U7656 ( .A1(n11731), .A2(n6650), .ZN(n11818) );
  INV_X1 U7657 ( .A(n11734), .ZN(n7416) );
  INV_X1 U7658 ( .A(n6814), .ZN(n6812) );
  NAND2_X1 U7659 ( .A1(n10778), .A2(n10777), .ZN(n12263) );
  AND2_X1 U7660 ( .A1(n12788), .A2(n15114), .ZN(n6859) );
  OR2_X1 U7661 ( .A1(n12816), .A2(n12825), .ZN(n7240) );
  NAND2_X1 U7662 ( .A1(n12828), .A2(n7234), .ZN(n7241) );
  INV_X1 U7663 ( .A(n12825), .ZN(n12805) );
  NAND2_X1 U7664 ( .A1(n12938), .A2(n12937), .ZN(n7227) );
  AND4_X1 U7665 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12780) );
  NAND2_X1 U7666 ( .A1(n12058), .A2(n12057), .ZN(n12779) );
  AOI21_X1 U7667 ( .B1(n12625), .B2(n12985), .A(n9643), .ZN(n9644) );
  AOI21_X1 U7668 ( .B1(n7185), .B2(n12928), .A(n9625), .ZN(n7184) );
  NAND2_X1 U7669 ( .A1(n9355), .A2(n9354), .ZN(n13076) );
  INV_X1 U7670 ( .A(n12056), .ZN(n9457) );
  INV_X1 U7671 ( .A(n10662), .ZN(n9387) );
  INV_X1 U7672 ( .A(n9244), .ZN(n12055) );
  NAND2_X1 U7673 ( .A1(n9557), .A2(n9573), .ZN(n10010) );
  NAND2_X1 U7674 ( .A1(n9316), .A2(n9315), .ZN(n9332) );
  NAND2_X1 U7675 ( .A1(n9168), .A2(n7110), .ZN(n7107) );
  NOR2_X1 U7676 ( .A1(n7097), .A2(n9131), .ZN(n7096) );
  AND2_X1 U7677 ( .A1(n9949), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9131) );
  INV_X1 U7678 ( .A(n9104), .ZN(n7097) );
  NAND2_X1 U7679 ( .A1(n13472), .A2(n7199), .ZN(n7198) );
  AND2_X1 U7680 ( .A1(n7200), .A2(n6701), .ZN(n7199) );
  NOR2_X1 U7681 ( .A1(n8937), .A2(n13228), .ZN(n7200) );
  NAND2_X1 U7682 ( .A1(n13478), .A2(n6641), .ZN(n7009) );
  AOI21_X1 U7683 ( .B1(n7139), .B2(n7142), .A(n6637), .ZN(n7138) );
  INV_X1 U7684 ( .A(n8607), .ZN(n7142) );
  AOI21_X1 U7685 ( .B1(n6613), .B2(n8539), .A(n7156), .ZN(n7155) );
  INV_X1 U7686 ( .A(n8553), .ZN(n7156) );
  OR2_X1 U7687 ( .A1(n13577), .A2(n8539), .ZN(n7158) );
  OAI21_X1 U7688 ( .B1(n11590), .B2(n6669), .A(n7476), .ZN(n11811) );
  OR2_X1 U7689 ( .A1(n7478), .A2(n7477), .ZN(n7476) );
  INV_X1 U7690 ( .A(n8687), .ZN(n7477) );
  NAND2_X1 U7691 ( .A1(n7211), .A2(n7210), .ZN(n11803) );
  INV_X1 U7692 ( .A(n10231), .ZN(n7195) );
  OR2_X1 U7693 ( .A1(n13424), .A2(n6917), .ZN(n7146) );
  NAND2_X1 U7694 ( .A1(n6920), .A2(n6918), .ZN(n6917) );
  AOI21_X1 U7695 ( .B1(n6919), .B2(n8937), .A(n13202), .ZN(n6918) );
  INV_X2 U7696 ( .A(n8273), .ZN(n8530) );
  INV_X1 U7697 ( .A(n14400), .ZN(n7650) );
  INV_X1 U7698 ( .A(n9879), .ZN(n8203) );
  AOI21_X1 U7699 ( .B1(n14109), .B2(n14108), .A(n7539), .ZN(n14100) );
  NAND2_X1 U7700 ( .A1(n14100), .A2(n14099), .ZN(n14098) );
  NAND2_X1 U7701 ( .A1(n14113), .A2(n8142), .ZN(n14114) );
  NAND2_X1 U7702 ( .A1(n14144), .A2(n6947), .ZN(n6943) );
  OR2_X1 U7703 ( .A1(n14144), .A2(n6946), .ZN(n6942) );
  NAND2_X1 U7704 ( .A1(n6961), .A2(n6959), .ZN(n7113) );
  AND2_X1 U7705 ( .A1(n7956), .A2(n6960), .ZN(n6959) );
  NAND2_X1 U7706 ( .A1(n11655), .A2(n14536), .ZN(n11654) );
  NAND2_X1 U7707 ( .A1(n8080), .A2(n8079), .ZN(n14101) );
  NAND2_X1 U7708 ( .A1(n7343), .A2(n7623), .ZN(n8076) );
  OAI21_X1 U7709 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n15476), .A(n14437), .ZN(
        n14444) );
  OAI22_X1 U7710 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14492), .B1(n14491), 
        .B2(n14490), .ZN(n14497) );
  NAND2_X1 U7711 ( .A1(n10823), .A2(n10822), .ZN(n10994) );
  INV_X1 U7712 ( .A(n10821), .ZN(n10822) );
  INV_X1 U7713 ( .A(n12712), .ZN(n6872) );
  NOR2_X1 U7714 ( .A1(n12736), .A2(n12737), .ZN(n12755) );
  NAND2_X1 U7715 ( .A1(n7495), .A2(n12031), .ZN(n7494) );
  NOR2_X1 U7716 ( .A1(n7498), .A2(n12032), .ZN(n7492) );
  AND2_X1 U7717 ( .A1(n11995), .A2(n11994), .ZN(n6980) );
  OAI21_X1 U7718 ( .B1(n14533), .B2(n14532), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n6888) );
  NOR2_X1 U7719 ( .A1(n14638), .A2(n14639), .ZN(n14637) );
  AOI21_X1 U7720 ( .B1(n9903), .B2(n8992), .A(n8746), .ZN(n8760) );
  AND2_X1 U7721 ( .A1(n10337), .A2(n8968), .ZN(n8746) );
  INV_X1 U7722 ( .A(n6689), .ZN(n7375) );
  INV_X1 U7723 ( .A(n8773), .ZN(n6793) );
  INV_X1 U7724 ( .A(n8800), .ZN(n7364) );
  NAND2_X1 U7725 ( .A1(n8792), .A2(n6643), .ZN(n7363) );
  NAND2_X1 U7726 ( .A1(n8796), .A2(n6642), .ZN(n7362) );
  INV_X1 U7727 ( .A(n9765), .ZN(n6767) );
  NAND2_X1 U7728 ( .A1(n8836), .A2(n6712), .ZN(n7382) );
  NOR2_X1 U7729 ( .A1(n8836), .A2(n6712), .ZN(n7383) );
  OR2_X1 U7730 ( .A1(n9785), .A2(n9787), .ZN(n6801) );
  AND2_X1 U7731 ( .A1(n8863), .A2(n8864), .ZN(n7372) );
  NAND2_X1 U7732 ( .A1(n7371), .A2(n7370), .ZN(n7369) );
  INV_X1 U7733 ( .A(n8864), .ZN(n7371) );
  INV_X1 U7734 ( .A(n8863), .ZN(n7370) );
  NOR2_X1 U7735 ( .A1(n7392), .A2(n6618), .ZN(n7387) );
  AOI21_X1 U7736 ( .B1(n8887), .B2(n8888), .A(n8892), .ZN(n7392) );
  NAND2_X1 U7737 ( .A1(n7391), .A2(n8890), .ZN(n7390) );
  NAND2_X1 U7738 ( .A1(n8887), .A2(n8888), .ZN(n7391) );
  NOR2_X1 U7739 ( .A1(n8887), .A2(n8888), .ZN(n7389) );
  OR4_X1 U7740 ( .A1(n12829), .A2(n13127), .A3(n12627), .A4(n12845), .ZN(
        n12193) );
  AOI21_X1 U7741 ( .B1(n6676), .B2(n7932), .A(n7338), .ZN(n7337) );
  NOR2_X1 U7742 ( .A1(n7597), .A2(SI_17_), .ZN(n7338) );
  OR2_X1 U7743 ( .A1(n6686), .A2(n9493), .ZN(n7175) );
  INV_X1 U7744 ( .A(n12192), .ZN(n7176) );
  AND2_X1 U7745 ( .A1(n6614), .A2(n9219), .ZN(n6840) );
  NAND2_X1 U7746 ( .A1(n7352), .A2(n8907), .ZN(n7351) );
  INV_X1 U7747 ( .A(n7355), .ZN(n7352) );
  INV_X1 U7748 ( .A(n8026), .ZN(n7123) );
  NAND2_X1 U7749 ( .A1(n8110), .A2(n8109), .ZN(n7271) );
  INV_X1 U7750 ( .A(n7579), .ZN(n7333) );
  OR2_X1 U7751 ( .A1(n12804), .A2(n13033), .ZN(n12218) );
  NOR2_X1 U7752 ( .A1(n7411), .A2(n6832), .ZN(n6831) );
  INV_X1 U7753 ( .A(n12305), .ZN(n6832) );
  INV_X1 U7754 ( .A(n12561), .ZN(n7409) );
  OAI21_X1 U7755 ( .B1(n11127), .B2(n11103), .A(n11118), .ZN(n11162) );
  INV_X1 U7756 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U7757 ( .A1(n12808), .A2(n12815), .ZN(n7239) );
  NOR2_X1 U7758 ( .A1(n12813), .A2(n7235), .ZN(n7234) );
  INV_X1 U7759 ( .A(n7530), .ZN(n7235) );
  OR2_X1 U7760 ( .A1(n9447), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9462) );
  AND2_X1 U7761 ( .A1(n12100), .A2(n12104), .ZN(n12237) );
  INV_X1 U7762 ( .A(n7240), .ZN(n7233) );
  NOR2_X1 U7763 ( .A1(n12801), .A2(n7230), .ZN(n7229) );
  INV_X1 U7764 ( .A(n7234), .ZN(n7230) );
  AND2_X1 U7765 ( .A1(n12789), .A2(n7239), .ZN(n7238) );
  NOR2_X1 U7766 ( .A1(n7175), .A2(n7174), .ZN(n7173) );
  INV_X1 U7767 ( .A(n12200), .ZN(n7174) );
  INV_X1 U7768 ( .A(n7175), .ZN(n7172) );
  OR2_X1 U7769 ( .A1(n13037), .A2(n12815), .ZN(n12214) );
  INV_X1 U7770 ( .A(n12829), .ZN(n12823) );
  NAND2_X1 U7771 ( .A1(n12841), .A2(n12200), .ZN(n12824) );
  INV_X1 U7772 ( .A(n12845), .ZN(n12842) );
  OR2_X1 U7773 ( .A1(n13130), .A2(n12862), .ZN(n12187) );
  OR2_X1 U7774 ( .A1(n13136), .A2(n12880), .ZN(n12182) );
  AOI21_X1 U7775 ( .B1(n7083), .B2(n9453), .A(n6731), .ZN(n7082) );
  INV_X1 U7776 ( .A(n9443), .ZN(n7083) );
  NAND2_X1 U7777 ( .A1(n7081), .A2(n7079), .ZN(n9469) );
  NOR2_X1 U7778 ( .A1(n7080), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7079) );
  INV_X1 U7779 ( .A(n7082), .ZN(n7080) );
  INV_X1 U7780 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9576) );
  AND3_X1 U7781 ( .A1(n6602), .A2(n9052), .A3(n6681), .ZN(n9547) );
  INV_X1 U7782 ( .A(n7088), .ZN(n7087) );
  OAI21_X1 U7783 ( .B1(n9331), .B2(n7089), .A(n9346), .ZN(n7088) );
  INV_X1 U7784 ( .A(n9333), .ZN(n7089) );
  NOR2_X1 U7785 ( .A1(n9179), .A2(n7111), .ZN(n7110) );
  INV_X1 U7786 ( .A(n9167), .ZN(n7111) );
  AND2_X1 U7787 ( .A1(n8982), .A2(n8967), .ZN(n8974) );
  CLKBUF_X1 U7788 ( .A(n8279), .Z(n8291) );
  OR2_X1 U7789 ( .A1(n8937), .A2(n13617), .ZN(n7201) );
  NOR2_X1 U7790 ( .A1(n13647), .A2(n13537), .ZN(n6929) );
  NAND2_X1 U7791 ( .A1(n13547), .A2(n6929), .ZN(n6930) );
  AND2_X1 U7792 ( .A1(n13532), .A2(n7475), .ZN(n7474) );
  NAND2_X1 U7793 ( .A1(n8696), .A2(n8697), .ZN(n7475) );
  NAND2_X1 U7794 ( .A1(n15000), .A2(n14999), .ZN(n7453) );
  OAI21_X1 U7795 ( .B1(n7135), .B2(n7452), .A(n8669), .ZN(n7451) );
  INV_X1 U7796 ( .A(n8668), .ZN(n7452) );
  XNOR2_X1 U7797 ( .A(n10386), .B(n13378), .ZN(n9003) );
  XNOR2_X1 U7798 ( .A(n9903), .B(n10337), .ZN(n10191) );
  NAND2_X1 U7799 ( .A1(n7212), .A2(n7213), .ZN(n11585) );
  INV_X1 U7800 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7484) );
  INV_X1 U7801 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8236) );
  INV_X1 U7802 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7149) );
  INV_X1 U7803 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7147) );
  INV_X1 U7804 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8222) );
  INV_X1 U7805 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8220) );
  AND2_X1 U7806 ( .A1(n13870), .A2(n6988), .ZN(n6987) );
  OR2_X1 U7807 ( .A1(n13785), .A2(n6989), .ZN(n6988) );
  INV_X1 U7808 ( .A(n12410), .ZN(n6989) );
  AND2_X1 U7809 ( .A1(n8150), .A2(n11532), .ZN(n10261) );
  INV_X1 U7810 ( .A(n10369), .ZN(n8097) );
  NAND2_X1 U7811 ( .A1(n7002), .A2(n7001), .ZN(n10367) );
  NAND2_X1 U7812 ( .A1(n12423), .A2(n13770), .ZN(n7001) );
  OR2_X1 U7813 ( .A1(n10375), .A2(n10496), .ZN(n7002) );
  NOR2_X1 U7814 ( .A1(n14125), .A2(n6948), .ZN(n6947) );
  INV_X1 U7815 ( .A(n8133), .ZN(n6948) );
  INV_X1 U7816 ( .A(n8134), .ZN(n6946) );
  NAND2_X1 U7817 ( .A1(n7122), .A2(n8012), .ZN(n6977) );
  INV_X1 U7818 ( .A(n6977), .ZN(n6979) );
  OR2_X1 U7819 ( .A1(n14192), .A2(n14191), .ZN(n8013) );
  OR2_X1 U7820 ( .A1(n7273), .A2(n7272), .ZN(n7049) );
  INV_X1 U7821 ( .A(n8127), .ZN(n7272) );
  AND2_X1 U7822 ( .A1(n14208), .A2(n8124), .ZN(n7273) );
  NOR2_X1 U7823 ( .A1(n7943), .A2(n6965), .ZN(n6964) );
  INV_X1 U7824 ( .A(n7931), .ZN(n6965) );
  OR2_X1 U7825 ( .A1(n14351), .A2(n13799), .ZN(n9766) );
  OR2_X1 U7826 ( .A1(n14716), .A2(n13915), .ZN(n8099) );
  INV_X1 U7827 ( .A(n10261), .ZN(n10259) );
  NAND2_X1 U7828 ( .A1(n7320), .A2(n7325), .ZN(n8948) );
  OAI21_X1 U7829 ( .B1(n7538), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8153) );
  INV_X1 U7830 ( .A(n8161), .ZN(n8158) );
  NAND2_X1 U7831 ( .A1(n7540), .A2(n7006), .ZN(n7005) );
  INV_X1 U7832 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U7833 ( .A1(n8000), .A2(n7609), .ZN(n7610) );
  INV_X1 U7834 ( .A(n7982), .ZN(n7605) );
  NAND2_X1 U7835 ( .A1(n7007), .A2(n7602), .ZN(n7980) );
  NAND2_X1 U7836 ( .A1(n7594), .A2(n15328), .ZN(n7597) );
  INV_X1 U7837 ( .A(n7030), .ZN(n7029) );
  OAI21_X1 U7838 ( .B1(n7032), .B2(n7031), .A(SI_14_), .ZN(n7030) );
  AND2_X1 U7839 ( .A1(n7584), .A2(n10216), .ZN(n7024) );
  INV_X1 U7840 ( .A(n7341), .ZN(n7340) );
  INV_X1 U7841 ( .A(n7556), .ZN(n6934) );
  AND2_X2 U7842 ( .A1(n7037), .A2(n7039), .ZN(n7552) );
  INV_X1 U7843 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7038) );
  INV_X1 U7844 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7059) );
  AOI22_X1 U7845 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14429), .B1(n14473), .B2(
        n14428), .ZN(n14431) );
  XNOR2_X1 U7846 ( .A(n11134), .B(n11266), .ZN(n10996) );
  NAND2_X1 U7847 ( .A1(n12281), .A2(n12280), .ZN(n12282) );
  NAND2_X1 U7848 ( .A1(n7394), .A2(n7397), .ZN(n7396) );
  INV_X1 U7849 ( .A(n6620), .ZN(n6822) );
  INV_X1 U7850 ( .A(n12540), .ZN(n6824) );
  AND2_X1 U7851 ( .A1(n10662), .A2(n10679), .ZN(n10796) );
  NAND2_X1 U7852 ( .A1(n6815), .A2(n6719), .ZN(n6814) );
  OR2_X1 U7853 ( .A1(n6817), .A2(n6816), .ZN(n6815) );
  INV_X1 U7854 ( .A(n12489), .ZN(n6816) );
  NAND2_X1 U7855 ( .A1(n12223), .A2(n12779), .ZN(n7178) );
  NOR2_X1 U7856 ( .A1(n11099), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7253) );
  OR2_X1 U7857 ( .A1(n10752), .A2(n7257), .ZN(n7252) );
  OR2_X1 U7858 ( .A1(n7254), .A2(n9111), .ZN(n7250) );
  INV_X1 U7859 ( .A(n9099), .ZN(n7414) );
  NOR2_X1 U7860 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n6912) );
  NAND2_X1 U7861 ( .A1(n6734), .A2(n6600), .ZN(n7263) );
  AND2_X1 U7862 ( .A1(n7263), .A2(n7262), .ZN(n15049) );
  INV_X1 U7863 ( .A(n15050), .ZN(n7262) );
  AOI21_X1 U7864 ( .B1(n15059), .B2(n15058), .A(n6905), .ZN(n6904) );
  INV_X1 U7865 ( .A(n11156), .ZN(n6905) );
  AND2_X1 U7866 ( .A1(n6898), .A2(n6897), .ZN(n15096) );
  INV_X1 U7867 ( .A(n11469), .ZN(n6897) );
  NAND2_X1 U7868 ( .A1(n6881), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U7869 ( .A1(n11466), .A2(n6881), .ZN(n6879) );
  INV_X1 U7870 ( .A(n15102), .ZN(n6881) );
  NAND2_X1 U7871 ( .A1(n6870), .A2(n6869), .ZN(n7249) );
  INV_X1 U7872 ( .A(n11535), .ZN(n6869) );
  OAI22_X1 U7873 ( .A1(n15096), .A2(n15095), .B1(n11470), .B2(n11471), .ZN(
        n11541) );
  AND2_X1 U7874 ( .A1(n7249), .A2(n7248), .ZN(n12638) );
  NAND2_X1 U7875 ( .A1(n11887), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U7876 ( .A1(n6882), .A2(n12651), .ZN(n7260) );
  NAND2_X1 U7877 ( .A1(n7260), .A2(n12676), .ZN(n7259) );
  AND2_X1 U7878 ( .A1(n12748), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U7879 ( .A1(n12824), .A2(n12823), .ZN(n12822) );
  AND2_X1 U7880 ( .A1(n12205), .A2(n12206), .ZN(n12813) );
  NAND2_X1 U7881 ( .A1(n12844), .A2(n9630), .ZN(n12828) );
  NAND2_X1 U7882 ( .A1(n12846), .A2(n12845), .ZN(n12844) );
  INV_X1 U7883 ( .A(n12890), .ZN(n12862) );
  OR2_X1 U7884 ( .A1(n9419), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9434) );
  AOI21_X1 U7885 ( .B1(n7163), .B2(n7165), .A(n7161), .ZN(n7160) );
  INV_X1 U7886 ( .A(n12169), .ZN(n7161) );
  NAND2_X1 U7887 ( .A1(n7227), .A2(n7226), .ZN(n12921) );
  NAND2_X1 U7888 ( .A1(n6849), .A2(n6850), .ZN(n12938) );
  NAND2_X1 U7889 ( .A1(n9622), .A2(n6852), .ZN(n6849) );
  NAND2_X1 U7890 ( .A1(n6868), .A2(n7216), .ZN(n12996) );
  NAND2_X1 U7891 ( .A1(n7217), .A2(n9616), .ZN(n7216) );
  INV_X1 U7892 ( .A(n7220), .ZN(n7217) );
  NAND2_X1 U7893 ( .A1(n6867), .A2(n9613), .ZN(n11664) );
  AND2_X1 U7894 ( .A1(n12112), .A2(n12111), .ZN(n12235) );
  AND2_X1 U7895 ( .A1(n12110), .A2(n12105), .ZN(n12233) );
  OR2_X1 U7896 ( .A1(n11263), .A2(n12237), .ZN(n11362) );
  NOR2_X1 U7897 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9142) );
  NAND2_X1 U7898 ( .A1(n15113), .A2(n15112), .ZN(n15111) );
  AOI22_X1 U7899 ( .A1(n12889), .A2(n9628), .B1(n12880), .B2(n9627), .ZN(
        n12878) );
  INV_X1 U7900 ( .A(n15117), .ZN(n13016) );
  NAND2_X1 U7901 ( .A1(n12211), .A2(n10796), .ZN(n15120) );
  INV_X1 U7902 ( .A(n12166), .ZN(n7187) );
  AND2_X1 U7903 ( .A1(n6700), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U7904 ( .A1(n6848), .A2(n6846), .ZN(n6845) );
  NAND2_X1 U7905 ( .A1(n7226), .A2(n12160), .ZN(n7224) );
  INV_X1 U7906 ( .A(n6848), .ZN(n6847) );
  OR2_X1 U7907 ( .A1(n12596), .A2(n12941), .ZN(n12166) );
  INV_X1 U7908 ( .A(n12231), .ZN(n12909) );
  NAND2_X1 U7909 ( .A1(n9337), .A2(n9336), .ZN(n13079) );
  AND2_X1 U7910 ( .A1(n11906), .A2(n9614), .ZN(n7220) );
  OR2_X1 U7911 ( .A1(n11664), .A2(n9615), .ZN(n7221) );
  AND2_X1 U7912 ( .A1(n7221), .A2(n9614), .ZN(n11907) );
  AND2_X1 U7913 ( .A1(n12132), .A2(n12137), .ZN(n12244) );
  INV_X1 U7914 ( .A(n15155), .ZN(n15172) );
  AND2_X1 U7915 ( .A1(n10782), .A2(n10016), .ZN(n11073) );
  NAND2_X1 U7916 ( .A1(n9559), .A2(n9558), .ZN(n10780) );
  OAI21_X1 U7917 ( .B1(n10010), .B2(P3_D_REG_0__SCAN_IN), .A(n9561), .ZN(
        n10801) );
  NAND2_X1 U7918 ( .A1(n9532), .A2(n9531), .ZN(n12044) );
  NAND2_X1 U7919 ( .A1(n7074), .A2(n9497), .ZN(n9521) );
  INV_X1 U7920 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9553) );
  AND2_X1 U7921 ( .A1(n9547), .A2(n9576), .ZN(n6838) );
  NAND2_X1 U7922 ( .A1(n9442), .A2(n9441), .ZN(n9444) );
  AND2_X1 U7923 ( .A1(n9541), .A2(n9544), .ZN(n7423) );
  INV_X1 U7924 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9544) );
  INV_X1 U7925 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U7926 ( .A1(n9296), .A2(n9295), .ZN(n9314) );
  NOR2_X1 U7927 ( .A1(n9245), .A2(n7420), .ZN(n9272) );
  OAI21_X1 U7928 ( .B1(n9239), .B2(n7092), .A(n7090), .ZN(n9271) );
  INV_X1 U7929 ( .A(n7091), .ZN(n7090) );
  NAND2_X1 U7930 ( .A1(n9239), .A2(n7093), .ZN(n9251) );
  OR2_X1 U7931 ( .A1(n9237), .A2(n9236), .ZN(n9239) );
  AND2_X1 U7932 ( .A1(n7106), .A2(n7108), .ZN(n7105) );
  INV_X1 U7933 ( .A(n9182), .ZN(n7106) );
  NAND2_X1 U7934 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n7109), .ZN(n7108) );
  INV_X1 U7935 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7109) );
  XNOR2_X1 U7936 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n9178) );
  NAND2_X1 U7937 ( .A1(n9156), .A2(n9155), .ZN(n9168) );
  NAND2_X1 U7938 ( .A1(n7095), .A2(n7094), .ZN(n9151) );
  AND2_X1 U7939 ( .A1(n7098), .A2(n9133), .ZN(n7094) );
  INV_X1 U7940 ( .A(n9135), .ZN(n7098) );
  NAND2_X1 U7941 ( .A1(n10681), .A2(n9045), .ZN(n9099) );
  NAND2_X1 U7942 ( .A1(n9103), .A2(n9102), .ZN(n9105) );
  AND2_X1 U7943 ( .A1(n13313), .A2(n13205), .ZN(n13208) );
  OR2_X1 U7944 ( .A1(n7502), .A2(n11232), .ZN(n7501) );
  INV_X1 U7945 ( .A(n11183), .ZN(n7502) );
  INV_X1 U7946 ( .A(n11419), .ZN(n7500) );
  AND2_X1 U7947 ( .A1(n11940), .A2(n11941), .ZN(n7498) );
  INV_X1 U7948 ( .A(n11939), .ZN(n7493) );
  NAND2_X1 U7949 ( .A1(n7497), .A2(n7496), .ZN(n7495) );
  OR2_X1 U7950 ( .A1(n7498), .A2(n7499), .ZN(n7497) );
  INV_X1 U7951 ( .A(n11944), .ZN(n7496) );
  NAND2_X1 U7952 ( .A1(n7523), .A2(n7522), .ZN(n11448) );
  INV_X1 U7953 ( .A(n11424), .ZN(n7523) );
  XNOR2_X1 U7954 ( .A(n6581), .B(n10337), .ZN(n10315) );
  NAND2_X1 U7955 ( .A1(n14571), .A2(n11877), .ZN(n11939) );
  NOR2_X1 U7956 ( .A1(n9022), .A2(n6751), .ZN(n6750) );
  INV_X1 U7957 ( .A(n13466), .ZN(n6751) );
  AND4_X1 U7958 ( .A1(n8251), .A2(n8250), .A3(n8249), .A4(n8248), .ZN(n13343)
         );
  NAND2_X1 U7959 ( .A1(n14406), .A2(n8958), .ZN(n7025) );
  NAND2_X1 U7960 ( .A1(n7470), .A2(n6619), .ZN(n7469) );
  NAND2_X1 U7961 ( .A1(n13503), .A2(n8598), .ZN(n13490) );
  NAND2_X1 U7962 ( .A1(n13490), .A2(n13489), .ZN(n13488) );
  NOR2_X1 U7963 ( .A1(n6930), .A2(n8905), .ZN(n13506) );
  XNOR2_X1 U7964 ( .A(n13635), .B(n13357), .ZN(n13489) );
  AND2_X1 U7965 ( .A1(n13500), .A2(n8585), .ZN(n13516) );
  NAND2_X1 U7966 ( .A1(n8564), .A2(n8998), .ZN(n13528) );
  NOR2_X1 U7967 ( .A1(n13557), .A2(n13657), .ZN(n13547) );
  NAND2_X1 U7968 ( .A1(n7158), .A2(n8540), .ZN(n13565) );
  INV_X1 U7969 ( .A(n13564), .ZN(n7157) );
  NAND2_X1 U7970 ( .A1(n6914), .A2(n6913), .ZN(n13557) );
  INV_X1 U7971 ( .A(n13713), .ZN(n6913) );
  NAND2_X1 U7972 ( .A1(n6756), .A2(n8521), .ZN(n13577) );
  NAND2_X1 U7973 ( .A1(n11954), .A2(n6621), .ZN(n13600) );
  XNOR2_X1 U7974 ( .A(n13674), .B(n13364), .ZN(n13603) );
  NAND2_X1 U7975 ( .A1(n11956), .A2(n11955), .ZN(n11954) );
  INV_X1 U7976 ( .A(n14589), .ZN(n6915) );
  NOR2_X1 U7977 ( .A1(n8686), .A2(n7479), .ZN(n7478) );
  INV_X1 U7978 ( .A(n8685), .ZN(n7479) );
  NAND2_X1 U7979 ( .A1(n7459), .A2(n8679), .ZN(n7458) );
  INV_X1 U7980 ( .A(n14940), .ZN(n7463) );
  NAND2_X1 U7981 ( .A1(n10383), .A2(n7135), .ZN(n10382) );
  NAND2_X1 U7982 ( .A1(n10188), .A2(n8665), .ZN(n10229) );
  INV_X1 U7983 ( .A(n13530), .ZN(n14992) );
  OR2_X1 U7984 ( .A1(n13202), .A2(n13581), .ZN(n9930) );
  AND2_X1 U7985 ( .A1(n13430), .A2(n15024), .ZN(n6926) );
  INV_X1 U7986 ( .A(n13487), .ZN(n13635) );
  INV_X1 U7987 ( .A(n15018), .ZN(n14597) );
  MUX2_X1 U7988 ( .A(n8278), .B(n13743), .S(n8277), .Z(n14969) );
  NOR2_X1 U7989 ( .A1(n8719), .A2(n13742), .ZN(n14958) );
  INV_X1 U7990 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8645) );
  INV_X1 U7991 ( .A(n13904), .ZN(n12328) );
  AND2_X1 U7992 ( .A1(n13793), .A2(n6994), .ZN(n6993) );
  NAND2_X1 U7993 ( .A1(n12340), .A2(n13880), .ZN(n6994) );
  NOR2_X1 U7994 ( .A1(n12340), .A2(n13880), .ZN(n6995) );
  INV_X1 U7995 ( .A(n12387), .ZN(n7000) );
  AND2_X1 U7996 ( .A1(n13746), .A2(n6999), .ZN(n6998) );
  OR2_X1 U7997 ( .A1(n13848), .A2(n7000), .ZN(n6999) );
  NAND2_X1 U7998 ( .A1(n13774), .A2(n12380), .ZN(n13847) );
  OR2_X1 U7999 ( .A1(n7885), .A2(n7884), .ZN(n7905) );
  NAND2_X1 U8001 ( .A1(n12338), .A2(n12339), .ZN(n13877) );
  NAND2_X1 U8002 ( .A1(n6992), .A2(n12340), .ZN(n13878) );
  INV_X1 U8003 ( .A(n12338), .ZN(n6992) );
  AND2_X1 U8004 ( .A1(n9845), .A2(n7541), .ZN(n6763) );
  INV_X1 U8005 ( .A(n8044), .ZN(n8020) );
  INV_X1 U8006 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7642) );
  INV_X1 U8007 ( .A(n8089), .ZN(n7131) );
  NOR2_X1 U8008 ( .A1(n14108), .A2(n6945), .ZN(n6944) );
  NOR2_X1 U8009 ( .A1(n6947), .A2(n6946), .ZN(n6945) );
  OAI22_X1 U8010 ( .A1(n14126), .A2(n14123), .B1(n14371), .B2(n14143), .ZN(
        n14109) );
  INV_X1 U8011 ( .A(n13894), .ZN(n14143) );
  INV_X1 U8012 ( .A(n13896), .ZN(n14141) );
  INV_X1 U8013 ( .A(n14147), .ZN(n7035) );
  INV_X1 U8014 ( .A(n14146), .ZN(n7036) );
  OAI21_X1 U8015 ( .B1(n14177), .B2(n14179), .A(n8130), .ZN(n14162) );
  NAND2_X1 U8016 ( .A1(n8030), .A2(n8029), .ZN(n14172) );
  NAND2_X1 U8017 ( .A1(n8013), .A2(n8012), .ZN(n14180) );
  NAND2_X1 U8018 ( .A1(n14180), .A2(n14179), .ZN(n14178) );
  AND2_X1 U8019 ( .A1(n7978), .A2(n7994), .ZN(n6957) );
  XNOR2_X1 U8020 ( .A(n14315), .B(n13899), .ZN(n14208) );
  NAND2_X1 U8021 ( .A1(n8125), .A2(n7273), .ZN(n14204) );
  XNOR2_X1 U8022 ( .A(n14325), .B(n14237), .ZN(n14227) );
  INV_X1 U8023 ( .A(n6964), .ZN(n6963) );
  AOI21_X1 U8024 ( .B1(n6964), .B2(n9873), .A(n9772), .ZN(n6962) );
  NAND2_X1 U8025 ( .A1(n8120), .A2(n6644), .ZN(n12019) );
  NAND2_X1 U8026 ( .A1(n11966), .A2(n9873), .ZN(n8120) );
  NAND2_X1 U8027 ( .A1(n7114), .A2(n7115), .ZN(n11970) );
  AOI21_X1 U8028 ( .B1(n7116), .B2(n11840), .A(n6659), .ZN(n7115) );
  NAND2_X1 U8029 ( .A1(n11970), .A2(n11969), .ZN(n11968) );
  NAND2_X1 U8030 ( .A1(n7118), .A2(n11830), .ZN(n11837) );
  INV_X1 U8031 ( .A(n11839), .ZN(n7118) );
  AOI21_X1 U8032 ( .B1(n7276), .B2(n7275), .A(n6658), .ZN(n7274) );
  INV_X1 U8033 ( .A(n8112), .ZN(n7275) );
  AND4_X1 U8034 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n13840)
         );
  AOI21_X1 U8035 ( .B1(n11289), .B2(n6969), .A(n6656), .ZN(n6968) );
  OR2_X1 U8036 ( .A1(n11277), .A2(n11289), .ZN(n11278) );
  NAND2_X1 U8037 ( .A1(n11337), .A2(n11341), .ZN(n11336) );
  AND2_X1 U8038 ( .A1(n9864), .A2(n9860), .ZN(n7124) );
  OR2_X1 U8039 ( .A1(n9677), .A2(n9949), .ZN(n6955) );
  OAI22_X1 U8040 ( .A1(n10497), .A2(n7698), .B1(n13917), .B2(n13770), .ZN(
        n10453) );
  OR2_X1 U8041 ( .A1(n9998), .A2(n13934), .ZN(n14142) );
  NAND2_X1 U8042 ( .A1(n10493), .A2(n6759), .ZN(n9859) );
  NAND2_X1 U8043 ( .A1(n10771), .A2(n6760), .ZN(n6759) );
  INV_X1 U8044 ( .A(n13918), .ZN(n6760) );
  NAND2_X1 U8045 ( .A1(n9679), .A2(n9678), .ZN(n14047) );
  AND2_X1 U8046 ( .A1(n7937), .A2(n7936), .ZN(n14338) );
  AND2_X1 U8047 ( .A1(n7851), .A2(n7850), .ZN(n14536) );
  NAND2_X1 U8048 ( .A1(n10459), .A2(n8192), .ZN(n14744) );
  OR2_X1 U8049 ( .A1(n8143), .A2(n8150), .ZN(n10401) );
  OAI211_X1 U8050 ( .C1(n7668), .C2(n7319), .A(n7315), .B(n7313), .ZN(n12276)
         );
  NAND2_X1 U8051 ( .A1(n7325), .A2(n8924), .ZN(n7319) );
  OAI21_X1 U8052 ( .B1(n7321), .B2(n8924), .A(n7316), .ZN(n7315) );
  INV_X1 U8053 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7646) );
  NAND2_X1 U8054 ( .A1(n7622), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U8055 ( .A1(n7014), .A2(n6609), .ZN(n7623) );
  CLKBUF_X1 U8056 ( .A(n8163), .Z(n8164) );
  AND2_X1 U8057 ( .A1(n8160), .A2(n8159), .ZN(n8190) );
  NOR2_X1 U8058 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  OR2_X1 U8059 ( .A1(n8153), .A2(n7636), .ZN(n8160) );
  NOR2_X1 U8060 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n8157) );
  NOR2_X1 U8061 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7307) );
  OR2_X1 U8062 ( .A1(n7983), .A2(n7982), .ZN(n7999) );
  OAI21_X1 U8063 ( .B1(n7960), .B2(n7959), .A(n7958), .ZN(n7962) );
  NAND2_X1 U8064 ( .A1(n7330), .A2(n7579), .ZN(n7836) );
  NAND2_X1 U8065 ( .A1(n7810), .A2(n7334), .ZN(n7330) );
  XNOR2_X1 U8066 ( .A(n6949), .B(n7823), .ZN(n10149) );
  NAND2_X1 U8067 ( .A1(n7810), .A2(n7577), .ZN(n6949) );
  INV_X1 U8068 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U8069 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7055), .ZN(n7054) );
  INV_X1 U8070 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7055) );
  OAI21_X1 U8071 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14439), .A(n14438), .ZN(
        n14486) );
  INV_X1 U8072 ( .A(n14646), .ZN(n6741) );
  OR2_X1 U8073 ( .A1(n14645), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U8074 ( .A1(n12604), .A2(n12605), .B1(n12805), .B2(n12482), .ZN(
        n12510) );
  XNOR2_X1 U8075 ( .A(n12313), .B(n12881), .ZN(n7413) );
  INV_X1 U8076 ( .A(n12914), .ZN(n12941) );
  NAND2_X1 U8077 ( .A1(n11137), .A2(n11136), .ZN(n11490) );
  INV_X1 U8078 ( .A(n12627), .ZN(n12881) );
  INV_X1 U8079 ( .A(n12629), .ZN(n12583) );
  INV_X1 U8080 ( .A(n15038), .ZN(n12609) );
  NAND2_X1 U8081 ( .A1(n9485), .A2(n9484), .ZN(n12816) );
  OR2_X1 U8082 ( .A1(n12056), .A2(n15326), .ZN(n9484) );
  AND2_X1 U8083 ( .A1(n11064), .A2(n11073), .ZN(n12270) );
  AND3_X1 U8084 ( .A1(n7100), .A2(n7099), .A3(n6606), .ZN(n12260) );
  NOR2_X1 U8085 ( .A1(n12256), .A2(n12258), .ZN(n7100) );
  NAND4_X1 U8086 ( .A1(n9492), .A2(n9491), .A3(n9490), .A4(n9489), .ZN(n12825)
         );
  NAND4_X1 U8087 ( .A1(n9148), .A2(n9147), .A3(n9146), .A4(n9145), .ZN(n12634)
         );
  OR2_X1 U8088 ( .A1(n11468), .A2(n11670), .ZN(n6871) );
  XNOR2_X1 U8089 ( .A(n11533), .B(n11539), .ZN(n11468) );
  XNOR2_X1 U8090 ( .A(n7259), .B(n14528), .ZN(n12669) );
  NAND2_X1 U8091 ( .A1(n12712), .A2(n12739), .ZN(n12748) );
  NAND2_X1 U8092 ( .A1(n7526), .A2(n7407), .ZN(n9351) );
  NOR2_X1 U8093 ( .A1(n12755), .A2(n6627), .ZN(n12756) );
  NOR2_X1 U8094 ( .A1(n12771), .A2(n12770), .ZN(n12773) );
  NAND2_X1 U8095 ( .A1(n6858), .A2(n6716), .ZN(n13032) );
  NAND2_X1 U8096 ( .A1(n6860), .A2(n6859), .ZN(n6858) );
  NAND2_X1 U8097 ( .A1(n9446), .A2(n9445), .ZN(n12872) );
  AND3_X1 U8098 ( .A1(n9190), .A2(n9189), .A3(n9188), .ZN(n15154) );
  OAI21_X1 U8099 ( .B1(n13103), .B2(n13095), .A(n9654), .ZN(n9655) );
  XNOR2_X1 U8100 ( .A(n9632), .B(n9631), .ZN(n9645) );
  NOR2_X1 U8101 ( .A1(n7246), .A2(n7244), .ZN(n7243) );
  NOR2_X1 U8102 ( .A1(n9644), .A2(n15176), .ZN(n7244) );
  NAND2_X1 U8103 ( .A1(n7247), .A2(n13100), .ZN(n7246) );
  NOR2_X1 U8104 ( .A1(n13032), .A2(n6857), .ZN(n13104) );
  AND2_X1 U8105 ( .A1(n13033), .A2(n15155), .ZN(n6857) );
  OAI21_X1 U8106 ( .B1(n11424), .B2(n7519), .A(n7518), .ZN(n14572) );
  NAND2_X1 U8107 ( .A1(n6630), .A2(n7522), .ZN(n7519) );
  NAND2_X1 U8108 ( .A1(n10322), .A2(n9913), .ZN(n9925) );
  AND2_X1 U8109 ( .A1(n13197), .A2(n13196), .ZN(n6769) );
  NAND2_X1 U8110 ( .A1(n8508), .A2(n8507), .ZN(n13679) );
  AND2_X1 U8111 ( .A1(n13244), .A2(n6679), .ZN(n7506) );
  AND2_X1 U8112 ( .A1(n13337), .A2(n13218), .ZN(n13219) );
  NAND2_X1 U8113 ( .A1(n10244), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14581) );
  OR2_X1 U8114 ( .A1(n14412), .A2(n8274), .ZN(n8609) );
  NAND2_X1 U8115 ( .A1(n9932), .A2(n15200), .ZN(n14578) );
  NOR4_X1 U8116 ( .A1(n9030), .A2(n11409), .A3(n9029), .A4(n11694), .ZN(n9031)
         );
  INV_X1 U8117 ( .A(n13341), .ZN(n13357) );
  OAI21_X1 U8118 ( .B1(n13438), .B2(n13604), .A(n13437), .ZN(n6797) );
  OR2_X1 U8119 ( .A1(n15035), .A2(n13530), .ZN(n7143) );
  NAND2_X1 U8120 ( .A1(n7146), .A2(n8662), .ZN(n7020) );
  NAND2_X1 U8121 ( .A1(n7288), .A2(n6622), .ZN(n7287) );
  INV_X1 U8122 ( .A(n13836), .ZN(n7288) );
  NAND2_X1 U8123 ( .A1(n12326), .A2(n7289), .ZN(n7283) );
  NAND2_X1 U8124 ( .A1(n13856), .A2(n12360), .ZN(n13754) );
  AND2_X1 U8125 ( .A1(n12007), .A2(n6636), .ZN(n7298) );
  NAND2_X1 U8126 ( .A1(n12402), .A2(n12401), .ZN(n13784) );
  AND2_X1 U8127 ( .A1(n7925), .A2(n7924), .ZN(n14344) );
  INV_X1 U8128 ( .A(n13889), .ZN(n14613) );
  OR2_X1 U8129 ( .A1(n14412), .A2(n8064), .ZN(n8066) );
  NAND2_X1 U8130 ( .A1(n10918), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14622) );
  NAND2_X1 U8131 ( .A1(n6806), .A2(n6805), .ZN(n6804) );
  NAND2_X1 U8132 ( .A1(n9842), .A2(n9843), .ZN(n6805) );
  INV_X1 U8133 ( .A(n9857), .ZN(n6806) );
  INV_X1 U8134 ( .A(n13840), .ZN(n13905) );
  NAND2_X1 U8135 ( .A1(n14098), .A2(n8089), .ZN(n6976) );
  AOI21_X1 U8136 ( .B1(n14097), .B2(n14741), .A(n14096), .ZN(n14263) );
  INV_X1 U8137 ( .A(n14703), .ZN(n14244) );
  NOR2_X1 U8138 ( .A1(n14712), .A2(n14329), .ZN(n14121) );
  AND2_X1 U8139 ( .A1(n14064), .A2(n14062), .ZN(n7045) );
  OR2_X1 U8140 ( .A1(n7064), .A2(n14381), .ZN(n7535) );
  XNOR2_X1 U8141 ( .A(n8139), .B(n9880), .ZN(n14073) );
  NAND2_X1 U8142 ( .A1(n15524), .A2(n15525), .ZN(n14457) );
  INV_X1 U8143 ( .A(n14483), .ZN(n6894) );
  INV_X1 U8144 ( .A(n14631), .ZN(n6754) );
  NAND2_X1 U8145 ( .A1(n6739), .A2(n6738), .ZN(n6889) );
  INV_X1 U8146 ( .A(n14643), .ZN(n6738) );
  NAND2_X1 U8147 ( .A1(n8749), .A2(n8750), .ZN(n6780) );
  OR2_X1 U8148 ( .A1(n7439), .A2(n9714), .ZN(n7438) );
  INV_X1 U8149 ( .A(n9713), .ZN(n7439) );
  OAI21_X1 U8150 ( .B1(n8779), .B2(n7373), .A(n7374), .ZN(n8793) );
  NAND2_X1 U8151 ( .A1(n8787), .A2(n6689), .ZN(n7374) );
  OR2_X1 U8152 ( .A1(n7445), .A2(n9723), .ZN(n7444) );
  INV_X1 U8153 ( .A(n9722), .ZN(n7445) );
  INV_X1 U8154 ( .A(n8799), .ZN(n7365) );
  OR2_X1 U8155 ( .A1(n7442), .A2(n9732), .ZN(n7441) );
  INV_X1 U8156 ( .A(n9731), .ZN(n7442) );
  NOR2_X1 U8157 ( .A1(n8824), .A2(n8827), .ZN(n7385) );
  INV_X1 U8158 ( .A(n8824), .ZN(n7384) );
  AOI21_X1 U8159 ( .B1(n6766), .B2(n7436), .A(n7435), .ZN(n9774) );
  NOR2_X1 U8160 ( .A1(n9769), .A2(n9770), .ZN(n7435) );
  AOI21_X1 U8161 ( .B1(n9769), .B2(n9770), .A(n6661), .ZN(n7436) );
  NAND2_X1 U8162 ( .A1(n6799), .A2(n7430), .ZN(n9790) );
  AND2_X1 U8163 ( .A1(n8845), .A2(n8846), .ZN(n7393) );
  NAND2_X1 U8164 ( .A1(n7368), .A2(n8871), .ZN(n7367) );
  NAND2_X1 U8165 ( .A1(n7372), .A2(n7369), .ZN(n7368) );
  AND2_X1 U8166 ( .A1(n6791), .A2(n7369), .ZN(n6790) );
  INV_X1 U8167 ( .A(n8871), .ZN(n6791) );
  NAND2_X1 U8168 ( .A1(n7379), .A2(n8875), .ZN(n7378) );
  INV_X1 U8169 ( .A(n6675), .ZN(n7379) );
  NAND2_X1 U8170 ( .A1(n7447), .A2(n9805), .ZN(n7446) );
  NAND2_X1 U8171 ( .A1(n9815), .A2(n7429), .ZN(n7428) );
  AOI21_X1 U8172 ( .B1(n8889), .B2(n7388), .A(n7386), .ZN(n8897) );
  NOR2_X1 U8173 ( .A1(n6618), .A2(n7389), .ZN(n7388) );
  AND2_X1 U8174 ( .A1(n7390), .A2(n7387), .ZN(n7386) );
  AND2_X1 U8175 ( .A1(n12210), .A2(n12209), .ZN(n12212) );
  NAND2_X1 U8176 ( .A1(n8903), .A2(n7356), .ZN(n7355) );
  INV_X1 U8177 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8221) );
  NOR2_X2 U8178 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8524) );
  AND2_X1 U8179 ( .A1(n9826), .A2(n7426), .ZN(n7425) );
  INV_X1 U8180 ( .A(n9824), .ZN(n7426) );
  INV_X1 U8181 ( .A(n8924), .ZN(n7318) );
  NAND2_X1 U8182 ( .A1(n7669), .A2(n7630), .ZN(n7327) );
  AOI21_X1 U8183 ( .B1(n6592), .B2(n7339), .A(n6720), .ZN(n7336) );
  OAI21_X1 U8184 ( .B1(n7598), .B2(n7339), .A(n7337), .ZN(n7944) );
  NOR2_X1 U8185 ( .A1(n7585), .A2(n7033), .ZN(n7032) );
  INV_X1 U8186 ( .A(n7583), .ZN(n7033) );
  INV_X1 U8187 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7042) );
  INV_X1 U8188 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7041) );
  INV_X1 U8189 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7040) );
  INV_X1 U8190 ( .A(n6831), .ZN(n6830) );
  NAND2_X1 U8191 ( .A1(n10753), .A2(n7254), .ZN(n7256) );
  NAND2_X1 U8192 ( .A1(n10759), .A2(n10758), .ZN(n11100) );
  AND2_X1 U8193 ( .A1(n7257), .A2(n10752), .ZN(n7254) );
  NAND2_X1 U8194 ( .A1(n15052), .A2(n6774), .ZN(n11214) );
  OR2_X1 U8195 ( .A1(n15065), .A2(n11145), .ZN(n6774) );
  NOR2_X1 U8196 ( .A1(n15049), .A2(n7261), .ZN(n11197) );
  NOR2_X1 U8197 ( .A1(n15065), .A2(n11146), .ZN(n7261) );
  OAI21_X1 U8198 ( .B1(n11897), .B2(n11914), .A(n11889), .ZN(n12654) );
  OR2_X1 U8199 ( .A1(n9473), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U8200 ( .A1(n12855), .A2(n12863), .ZN(n12200) );
  AND2_X1 U8201 ( .A1(n12160), .A2(n7164), .ZN(n7163) );
  OR2_X1 U8202 ( .A1(n12956), .A2(n7165), .ZN(n7164) );
  INV_X1 U8203 ( .A(n12152), .ZN(n7165) );
  NOR2_X1 U8204 ( .A1(n6853), .A2(n9623), .ZN(n6852) );
  INV_X1 U8205 ( .A(n9621), .ZN(n6853) );
  NOR2_X1 U8206 ( .A1(n7218), .A2(n6866), .ZN(n6865) );
  INV_X1 U8207 ( .A(n9613), .ZN(n6866) );
  NAND2_X1 U8208 ( .A1(n7219), .A2(n9616), .ZN(n7218) );
  INV_X1 U8209 ( .A(n9615), .ZN(n7219) );
  NAND2_X1 U8210 ( .A1(n11919), .A2(n12239), .ZN(n6867) );
  INV_X1 U8211 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U8212 ( .A1(n11302), .A2(n13015), .ZN(n12094) );
  INV_X1 U8213 ( .A(n7184), .ZN(n7183) );
  INV_X1 U8214 ( .A(n6852), .ZN(n6846) );
  NAND2_X1 U8215 ( .A1(n6566), .A2(n9945), .ZN(n9100) );
  NAND2_X1 U8216 ( .A1(n9074), .A2(n6864), .ZN(n6861) );
  NAND2_X1 U8217 ( .A1(n9219), .A2(n9055), .ZN(n7190) );
  INV_X1 U8218 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U8219 ( .A1(n7419), .A2(n9050), .ZN(n7418) );
  INV_X1 U8220 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U8221 ( .A1(n9282), .A2(n9281), .ZN(n9294) );
  NAND2_X1 U8222 ( .A1(n9279), .A2(n9278), .ZN(n9282) );
  NAND2_X1 U8223 ( .A1(n9049), .A2(n7421), .ZN(n7420) );
  INV_X1 U8224 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9049) );
  INV_X1 U8225 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9280) );
  OAI21_X1 U8226 ( .B1(n7093), .B2(n7092), .A(n9268), .ZN(n7091) );
  INV_X1 U8227 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9048) );
  INV_X1 U8228 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9047) );
  NOR2_X1 U8229 ( .A1(n8510), .A2(n8509), .ZN(n8258) );
  AND3_X1 U8230 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8335) );
  AND2_X1 U8231 ( .A1(n7353), .A2(n7351), .ZN(n7350) );
  INV_X1 U8232 ( .A(n8906), .ZN(n7353) );
  NOR2_X1 U8233 ( .A1(n8976), .A2(n8975), .ZN(n7346) );
  AND2_X1 U8234 ( .A1(n8619), .A2(n7140), .ZN(n7139) );
  NAND2_X1 U8235 ( .A1(n7141), .A2(n8607), .ZN(n7140) );
  INV_X1 U8236 ( .A(n13489), .ZN(n7141) );
  INV_X1 U8237 ( .A(n13500), .ZN(n7151) );
  INV_X1 U8238 ( .A(n14598), .ZN(n7212) );
  NOR2_X1 U8239 ( .A1(n8449), .A2(n8242), .ZN(n8450) );
  AND2_X1 U8240 ( .A1(n8363), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8381) );
  OAI21_X1 U8241 ( .B1(n14991), .B2(n8371), .A(n8372), .ZN(n10733) );
  INV_X1 U8242 ( .A(n6922), .ZN(n6919) );
  NOR2_X1 U8243 ( .A1(n13617), .A2(n13228), .ZN(n6922) );
  NAND2_X1 U8244 ( .A1(n13472), .A2(n13623), .ZN(n13459) );
  AND2_X1 U8245 ( .A1(n8230), .A2(n7484), .ZN(n7483) );
  INV_X1 U8246 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8522) );
  AND2_X1 U8247 ( .A1(n8475), .A2(n8523), .ZN(n8724) );
  AND2_X1 U8248 ( .A1(n14611), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U8249 ( .A1(n7287), .A2(n7290), .ZN(n7285) );
  INV_X1 U8250 ( .A(n7287), .ZN(n7286) );
  OR4_X1 U8251 ( .A1(n14099), .A2(n14125), .A3(n14108), .A4(n9877), .ZN(n9878)
         );
  OR4_X1 U8252 ( .A1(n14147), .A2(n14173), .A3(n14179), .A4(n9876), .ZN(n9877)
         );
  OR2_X1 U8253 ( .A1(n9681), .A2(n9680), .ZN(n9849) );
  NAND2_X1 U8254 ( .A1(n6962), .A2(n6963), .ZN(n6960) );
  AND2_X1 U8255 ( .A1(n7926), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7938) );
  INV_X1 U8256 ( .A(n7892), .ZN(n7117) );
  NOR2_X1 U8257 ( .A1(n11279), .A2(n7265), .ZN(n6967) );
  INV_X1 U8258 ( .A(n7821), .ZN(n6969) );
  AOI21_X1 U8259 ( .B1(n7269), .B2(n7268), .A(n6660), .ZN(n7267) );
  INV_X1 U8260 ( .A(n8109), .ZN(n7268) );
  OR2_X1 U8261 ( .A1(n11052), .A2(n7270), .ZN(n7266) );
  AND2_X1 U8262 ( .A1(n7321), .A2(n7318), .ZN(n7314) );
  AOI21_X1 U8263 ( .B1(n7325), .B2(n7323), .A(n7322), .ZN(n7321) );
  INV_X1 U8264 ( .A(n8944), .ZN(n7322) );
  INV_X1 U8265 ( .A(n7630), .ZN(n7323) );
  NAND2_X1 U8266 ( .A1(n7321), .A2(n7317), .ZN(n7316) );
  NAND2_X1 U8267 ( .A1(n7326), .A2(n7318), .ZN(n7317) );
  AND2_X1 U8268 ( .A1(n7618), .A2(n7019), .ZN(n7018) );
  INV_X1 U8269 ( .A(n8049), .ZN(n7019) );
  AND2_X1 U8270 ( .A1(n7307), .A2(n7308), .ZN(n7306) );
  INV_X1 U8271 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7308) );
  AND2_X1 U8272 ( .A1(n7593), .A2(n7592), .ZN(n7893) );
  AOI21_X1 U8273 ( .B1(n7331), .B2(n7333), .A(n6664), .ZN(n7329) );
  NOR2_X1 U8274 ( .A1(n7580), .A2(n7335), .ZN(n7334) );
  NAND2_X1 U8275 ( .A1(n7552), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U8276 ( .A1(n7021), .A2(n7312), .ZN(n7311) );
  NAND2_X1 U8277 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7052), .ZN(n7051) );
  INV_X1 U8278 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7052) );
  INV_X1 U8279 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U8280 ( .A1(n6818), .A2(n6726), .ZN(n6817) );
  INV_X1 U8281 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U8282 ( .A1(n6589), .A2(n7422), .ZN(n6819) );
  NAND2_X1 U8283 ( .A1(n6828), .A2(n7408), .ZN(n12480) );
  NAND2_X1 U8284 ( .A1(n7404), .A2(n11497), .ZN(n11509) );
  INV_X1 U8285 ( .A(n11511), .ZN(n7404) );
  AND2_X1 U8286 ( .A1(n12270), .A2(n10795), .ZN(n15038) );
  INV_X1 U8287 ( .A(n6856), .ZN(n6855) );
  OAI22_X1 U8288 ( .A1(n12061), .A2(n9162), .B1(n12062), .B2(n11146), .ZN(
        n6856) );
  NAND2_X1 U8289 ( .A1(n10965), .A2(n10670), .ZN(n10671) );
  NAND2_X1 U8290 ( .A1(n7255), .A2(n7256), .ZN(n10754) );
  NAND2_X1 U8291 ( .A1(n10753), .A2(n10752), .ZN(n7251) );
  XNOR2_X1 U8292 ( .A(n11214), .B(n11198), .ZN(n11166) );
  XNOR2_X1 U8293 ( .A(n11197), .B(n11198), .ZN(n11160) );
  NOR2_X1 U8294 ( .A1(n6903), .A2(n11203), .ZN(n6900) );
  XNOR2_X1 U8295 ( .A(n11472), .B(n11464), .ZN(n11218) );
  NAND2_X1 U8296 ( .A1(n11218), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11474) );
  NOR2_X1 U8297 ( .A1(n15073), .A2(n7258), .ZN(n11463) );
  NOR2_X1 U8298 ( .A1(n15081), .A2(n9196), .ZN(n7258) );
  NAND2_X1 U8299 ( .A1(n6871), .A2(n6626), .ZN(n6870) );
  NAND2_X1 U8300 ( .A1(n11546), .A2(n11547), .ZN(n11549) );
  OR2_X1 U8301 ( .A1(n12639), .A2(n12640), .ZN(n6882) );
  NAND2_X1 U8302 ( .A1(n12678), .A2(n12677), .ZN(n12701) );
  XNOR2_X1 U8303 ( .A(n12738), .B(n12730), .ZN(n12740) );
  NOR2_X1 U8304 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7407) );
  INV_X1 U8305 ( .A(n12747), .ZN(n6878) );
  NOR2_X1 U8306 ( .A1(n12734), .A2(n6909), .ZN(n6908) );
  NOR2_X1 U8307 ( .A1(n6910), .A2(n12730), .ZN(n6909) );
  INV_X1 U8308 ( .A(n12735), .ZN(n6910) );
  AOI21_X1 U8309 ( .B1(n12740), .B2(P3_REG1_REG_17__SCAN_IN), .A(n6773), .ZN(
        n12760) );
  AND2_X1 U8310 ( .A1(n12738), .A2(n12739), .ZN(n6773) );
  NAND2_X1 U8311 ( .A1(n7236), .A2(n12786), .ZN(n6860) );
  AOI22_X1 U8312 ( .A1(n7241), .A2(n7237), .B1(n7239), .B2(n12801), .ZN(n7236)
         );
  AND2_X1 U8313 ( .A1(n7239), .A2(n7240), .ZN(n7237) );
  OR2_X1 U8314 ( .A1(n9486), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9502) );
  OR2_X1 U8315 ( .A1(n13119), .A2(n12847), .ZN(n7530) );
  AOI21_X1 U8316 ( .B1(n12861), .B2(n12252), .A(n6841), .ZN(n12846) );
  AND2_X1 U8317 ( .A1(n12872), .A2(n12627), .ZN(n6841) );
  XNOR2_X1 U8318 ( .A(n12872), .B(n12627), .ZN(n12860) );
  INV_X1 U8319 ( .A(n9434), .ZN(n9433) );
  NAND2_X1 U8320 ( .A1(n9407), .A2(n9406), .ZN(n9419) );
  NAND2_X1 U8321 ( .A1(n9622), .A2(n9621), .ZN(n12948) );
  AND2_X1 U8322 ( .A1(n9302), .A2(n9301), .ZN(n9322) );
  AND2_X1 U8323 ( .A1(n12141), .A2(n12142), .ZN(n12999) );
  OR2_X1 U8324 ( .A1(n9262), .A2(n9261), .ZN(n9287) );
  OR2_X1 U8325 ( .A1(n9228), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9262) );
  AND2_X1 U8326 ( .A1(n12115), .A2(n12116), .ZN(n12234) );
  AOI21_X1 U8327 ( .B1(n12233), .B2(n7169), .A(n7167), .ZN(n7166) );
  NOR2_X1 U8328 ( .A1(n9171), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9194) );
  INV_X1 U8329 ( .A(n12633), .ZN(n11502) );
  INV_X1 U8330 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U8331 ( .A1(n10810), .A2(n6565), .ZN(n13013) );
  NAND2_X1 U8332 ( .A1(n9536), .A2(n9535), .ZN(n13101) );
  INV_X1 U8333 ( .A(n12901), .ZN(n12880) );
  NAND2_X1 U8334 ( .A1(n7228), .A2(n7231), .ZN(n12788) );
  AND2_X1 U8335 ( .A1(n7238), .A2(n7232), .ZN(n7231) );
  NAND2_X1 U8336 ( .A1(n12799), .A2(n7233), .ZN(n7232) );
  NAND2_X1 U8337 ( .A1(n13101), .A2(n13148), .ZN(n7247) );
  NAND2_X1 U8338 ( .A1(n9527), .A2(n9526), .ZN(n13033) );
  NAND2_X1 U8339 ( .A1(n7172), .A2(n6663), .ZN(n7171) );
  AOI21_X1 U8340 ( .B1(n6844), .B2(n6847), .A(n6588), .ZN(n6843) );
  NAND2_X1 U8341 ( .A1(n12954), .A2(n12956), .ZN(n12955) );
  AND2_X1 U8342 ( .A1(n12146), .A2(n12153), .ZN(n12965) );
  AND2_X1 U8343 ( .A1(n10936), .A2(n10777), .ZN(n15155) );
  NOR2_X1 U8344 ( .A1(n9076), .A2(n6862), .ZN(n9060) );
  INV_X1 U8345 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6863) );
  INV_X1 U8346 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U8347 ( .A1(n9523), .A2(n9522), .ZN(n9530) );
  NAND2_X1 U8348 ( .A1(n9521), .A2(n9520), .ZN(n9523) );
  XNOR2_X1 U8349 ( .A(n9556), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U8350 ( .A1(n7075), .A2(n9482), .ZN(n9496) );
  NAND2_X1 U8351 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n6837) );
  NAND2_X1 U8352 ( .A1(n9469), .A2(n9456), .ZN(n9468) );
  XNOR2_X1 U8353 ( .A(n9577), .B(n9576), .ZN(n10781) );
  NAND2_X1 U8354 ( .A1(n9550), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7424) );
  NAND2_X1 U8355 ( .A1(n9382), .A2(n9381), .ZN(n9402) );
  NAND2_X1 U8356 ( .A1(n9380), .A2(n9379), .ZN(n9382) );
  AOI21_X1 U8357 ( .B1(n7087), .B2(n7089), .A(n6722), .ZN(n7085) );
  NAND2_X1 U8358 ( .A1(n7526), .A2(n9334), .ZN(n9349) );
  NAND2_X1 U8359 ( .A1(n9218), .A2(n7192), .ZN(n9297) );
  NOR2_X1 U8360 ( .A1(n7418), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7192) );
  XNOR2_X1 U8361 ( .A(n9294), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9293) );
  AND2_X1 U8362 ( .A1(n9250), .A2(n9240), .ZN(n9241) );
  NAND2_X1 U8363 ( .A1(n9222), .A2(n9221), .ZN(n9237) );
  INV_X1 U8364 ( .A(n7105), .ZN(n7104) );
  AOI21_X1 U8365 ( .B1(n7103), .B2(n7105), .A(n7102), .ZN(n7101) );
  INV_X1 U8366 ( .A(n9203), .ZN(n7102) );
  AND2_X1 U8367 ( .A1(n9221), .A2(n9205), .ZN(n9206) );
  NAND2_X1 U8368 ( .A1(n9207), .A2(n9206), .ZN(n9222) );
  OR2_X1 U8369 ( .A1(n9185), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n9201) );
  NOR2_X1 U8370 ( .A1(n10681), .A2(n9056), .ZN(n7264) );
  XNOR2_X1 U8371 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n7073) );
  OR2_X1 U8372 ( .A1(n11866), .A2(n7521), .ZN(n7520) );
  INV_X1 U8373 ( .A(n11447), .ZN(n7521) );
  INV_X1 U8374 ( .A(n11425), .ZN(n7522) );
  OR2_X1 U8375 ( .A1(n8482), .A2(n8481), .ZN(n8498) );
  OR2_X1 U8376 ( .A1(n11940), .A2(n11941), .ZN(n7499) );
  XNOR2_X1 U8377 ( .A(n10386), .B(n13217), .ZN(n10432) );
  XNOR2_X1 U8378 ( .A(n14598), .B(n13255), .ZN(n11868) );
  OR2_X1 U8379 ( .A1(n8556), .A2(n15325), .ZN(n8570) );
  NOR2_X1 U8380 ( .A1(n8570), .A2(n13317), .ZN(n8579) );
  NAND2_X1 U8381 ( .A1(n11184), .A2(n7505), .ZN(n11229) );
  INV_X1 U8382 ( .A(n7501), .ZN(n7505) );
  NAND2_X1 U8383 ( .A1(n10328), .A2(n9905), .ZN(n10316) );
  XNOR2_X1 U8384 ( .A(n13674), .B(n13217), .ZN(n13193) );
  INV_X1 U8385 ( .A(n10658), .ZN(n10656) );
  AND2_X1 U8386 ( .A1(n8988), .A2(n7345), .ZN(n7542) );
  AND2_X1 U8387 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  NAND2_X1 U8388 ( .A1(n8974), .A2(n7346), .ZN(n7345) );
  OR2_X1 U8389 ( .A1(n8985), .A2(n8984), .ZN(n8986) );
  NAND2_X1 U8390 ( .A1(n8974), .A2(n8973), .ZN(n8989) );
  AND4_X1 U8391 ( .A1(n8595), .A2(n8594), .A3(n8593), .A4(n8592), .ZN(n13282)
         );
  OR2_X1 U8392 ( .A1(n8291), .A2(n8287), .ZN(n8293) );
  OR2_X1 U8393 ( .A1(n14844), .A2(n14843), .ZN(n14845) );
  AND2_X1 U8394 ( .A1(n14870), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n14872) );
  NAND2_X1 U8395 ( .A1(n8703), .A2(n7466), .ZN(n7465) );
  INV_X1 U8396 ( .A(n6619), .ZN(n7466) );
  AOI21_X1 U8397 ( .B1(n13456), .B2(n13466), .A(n6753), .ZN(n13439) );
  AND2_X1 U8398 ( .A1(n13228), .A2(n13343), .ZN(n6753) );
  NOR2_X1 U8399 ( .A1(n13466), .A2(n7468), .ZN(n7467) );
  OAI21_X1 U8400 ( .B1(n13497), .B2(n13499), .A(n8699), .ZN(n13482) );
  OR2_X1 U8401 ( .A1(n13528), .A2(n6628), .ZN(n7153) );
  NAND2_X1 U8402 ( .A1(n7153), .A2(n6590), .ZN(n13498) );
  NAND2_X1 U8403 ( .A1(n13547), .A2(n13709), .ZN(n13534) );
  AOI21_X1 U8404 ( .B1(n7474), .B2(n7472), .A(n6653), .ZN(n7471) );
  INV_X1 U8405 ( .A(n7474), .ZN(n7473) );
  INV_X1 U8406 ( .A(n8697), .ZN(n7472) );
  AND2_X1 U8407 ( .A1(n8999), .A2(n8998), .ZN(n13551) );
  NOR2_X1 U8408 ( .A1(n7457), .A2(n6668), .ZN(n7454) );
  INV_X1 U8409 ( .A(n11400), .ZN(n8459) );
  NOR2_X1 U8410 ( .A1(n14938), .A2(n11431), .ZN(n6916) );
  NAND2_X1 U8411 ( .A1(n14942), .A2(n15019), .ZN(n14941) );
  NAND2_X1 U8412 ( .A1(n10845), .A2(n8401), .ZN(n11002) );
  NAND2_X1 U8413 ( .A1(n7209), .A2(n15201), .ZN(n14996) );
  NAND2_X1 U8414 ( .A1(n7453), .A2(n8673), .ZN(n10729) );
  AOI21_X1 U8415 ( .B1(n7450), .B2(n7452), .A(n6635), .ZN(n7448) );
  AOI21_X1 U8416 ( .B1(n9003), .B2(n7133), .A(n6649), .ZN(n7134) );
  NAND2_X1 U8417 ( .A1(n10599), .A2(n14978), .ZN(n10598) );
  CLKBUF_X1 U8418 ( .A(n10191), .Z(n6757) );
  OR3_X1 U8419 ( .A1(n13507), .A2(n13506), .A3(n13202), .ZN(n13639) );
  OR2_X1 U8420 ( .A1(n11616), .A2(n8274), .ZN(n8569) );
  NAND2_X1 U8421 ( .A1(n8555), .A2(n8554), .ZN(n13657) );
  OR2_X1 U8422 ( .A1(n11642), .A2(n8274), .ZN(n8555) );
  OR2_X1 U8423 ( .A1(n14968), .A2(n9933), .ZN(n15018) );
  AND2_X1 U8424 ( .A1(n8230), .A2(n7482), .ZN(n7481) );
  AND2_X1 U8425 ( .A1(n7484), .A2(n8236), .ZN(n7482) );
  OR2_X1 U8426 ( .A1(n8712), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8715) );
  OR2_X1 U8427 ( .A1(n8346), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8359) );
  OR2_X1 U8428 ( .A1(n8375), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8322) );
  INV_X1 U8429 ( .A(n8018), .ZN(n8032) );
  NOR2_X1 U8430 ( .A1(n7971), .A2(n13759), .ZN(n7986) );
  AOI21_X1 U8431 ( .B1(n6987), .B2(n6989), .A(n6652), .ZN(n6985) );
  NAND2_X1 U8432 ( .A1(n11568), .A2(n6651), .ZN(n11713) );
  AND2_X1 U8433 ( .A1(n10366), .A2(n10367), .ZN(n10368) );
  NAND2_X1 U8434 ( .A1(n10372), .A2(n10371), .ZN(n13764) );
  OR2_X1 U8435 ( .A1(n10370), .A2(n8097), .ZN(n10371) );
  AND2_X1 U8436 ( .A1(n7986), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8004) );
  AOI21_X1 U8437 ( .B1(n6993), .B2(n6995), .A(n6645), .ZN(n6991) );
  INV_X1 U8438 ( .A(n10913), .ZN(n12418) );
  AND2_X1 U8439 ( .A1(n7295), .A2(n7294), .ZN(n7293) );
  NAND2_X1 U8440 ( .A1(n12422), .A2(n6758), .ZN(n7295) );
  AOI22_X1 U8441 ( .A1(n10264), .A2(P1_IR_REG_0__SCAN_IN), .B1(n12423), .B2(
        n10263), .ZN(n7294) );
  NAND2_X1 U8442 ( .A1(n7293), .A2(n10370), .ZN(n10372) );
  NOR2_X1 U8443 ( .A1(n7852), .A2(n11996), .ZN(n7867) );
  NAND2_X1 U8444 ( .A1(n7292), .A2(n12325), .ZN(n7291) );
  NAND2_X1 U8445 ( .A1(n13847), .A2(n13848), .ZN(n13846) );
  NAND2_X1 U8446 ( .A1(n13857), .A2(n13858), .ZN(n13856) );
  AND2_X1 U8447 ( .A1(n7770), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7785) );
  NOR2_X1 U8448 ( .A1(n7905), .A2(n7904), .ZN(n7926) );
  AND4_X1 U8449 ( .A1(n7891), .A2(n7890), .A3(n7889), .A4(n7888), .ZN(n13885)
         );
  INV_X1 U8450 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U8451 ( .A1(n14113), .A2(n6591), .ZN(n8200) );
  AND2_X1 U8452 ( .A1(n6591), .A2(n7064), .ZN(n7063) );
  NAND2_X1 U8453 ( .A1(n14089), .A2(n14099), .ZN(n14090) );
  NAND2_X1 U8454 ( .A1(n6611), .A2(n6977), .ZN(n6772) );
  NAND2_X1 U8455 ( .A1(n6611), .A2(n7119), .ZN(n14139) );
  NAND2_X1 U8456 ( .A1(n8013), .A2(n6979), .ZN(n7119) );
  NAND2_X1 U8457 ( .A1(n14160), .A2(n8131), .ZN(n14146) );
  NAND2_X1 U8458 ( .A1(n14162), .A2(n14161), .ZN(n14160) );
  NAND2_X1 U8459 ( .A1(n7048), .A2(n8129), .ZN(n14177) );
  OAI211_X1 U8460 ( .C1(n8125), .C2(n7272), .A(n7049), .B(n14191), .ZN(n7048)
         );
  NAND2_X1 U8461 ( .A1(n14205), .A2(n7995), .ZN(n14192) );
  NAND2_X1 U8462 ( .A1(n7068), .A2(n7067), .ZN(n14218) );
  NAND2_X1 U8463 ( .A1(n12019), .A2(n8122), .ZN(n14233) );
  AND2_X1 U8464 ( .A1(n14344), .A2(n11971), .ZN(n12023) );
  INV_X1 U8465 ( .A(n14344), .ZN(n11975) );
  AND3_X1 U8466 ( .A1(n7942), .A2(n7941), .A3(n7940), .ZN(n13862) );
  NOR2_X1 U8467 ( .A1(n14351), .A2(n11842), .ZN(n11971) );
  NAND2_X1 U8468 ( .A1(n7072), .A2(n7071), .ZN(n11842) );
  AOI21_X1 U8469 ( .B1(n8115), .B2(n6932), .A(n6657), .ZN(n6931) );
  INV_X1 U8470 ( .A(n8113), .ZN(n6932) );
  INV_X1 U8471 ( .A(n13906), .ZN(n11998) );
  NAND2_X1 U8472 ( .A1(n7266), .A2(n7267), .ZN(n11340) );
  NOR2_X1 U8473 ( .A1(n7800), .A2(n7799), .ZN(n7815) );
  NAND2_X1 U8474 ( .A1(n8106), .A2(n8105), .ZN(n10696) );
  NAND2_X1 U8475 ( .A1(n6971), .A2(n6970), .ZN(n10691) );
  AOI21_X1 U8476 ( .B1(n7124), .B2(n6972), .A(n6634), .ZN(n6970) );
  NAND2_X1 U8477 ( .A1(n10558), .A2(n10921), .ZN(n10692) );
  AND2_X1 U8478 ( .A1(n12459), .A2(n8098), .ZN(n10513) );
  INV_X1 U8479 ( .A(n10452), .ZN(n10466) );
  NAND2_X1 U8480 ( .A1(n8099), .A2(n7716), .ZN(n10452) );
  AND2_X1 U8481 ( .A1(n9691), .A2(n9690), .ZN(n10497) );
  INV_X1 U8482 ( .A(n14140), .ZN(n14234) );
  INV_X1 U8483 ( .A(n14142), .ZN(n14236) );
  OR3_X1 U8484 ( .A1(n10456), .A2(n10455), .A3(n10454), .ZN(n14063) );
  AND4_X1 U8485 ( .A1(n7667), .A2(n7666), .A3(n7665), .A4(n7664), .ZN(n12457)
         );
  OAI211_X1 U8486 ( .C1(n8190), .C2(n8171), .A(n8170), .B(n8169), .ZN(n9987)
         );
  NAND2_X1 U8487 ( .A1(n7432), .A2(n7648), .ZN(n7431) );
  INV_X1 U8488 ( .A(n7433), .ZN(n7432) );
  NAND2_X1 U8489 ( .A1(n8957), .A2(n8956), .ZN(n13722) );
  OR3_X1 U8490 ( .A1(n8948), .A2(n8943), .A3(n8950), .ZN(n8957) );
  NAND2_X1 U8491 ( .A1(n7434), .A2(n7646), .ZN(n7433) );
  NAND2_X1 U8492 ( .A1(n7964), .A2(n7640), .ZN(n8163) );
  XNOR2_X1 U8493 ( .A(n8920), .B(n8919), .ZN(n13728) );
  NAND2_X1 U8494 ( .A1(n7324), .A2(n7630), .ZN(n8920) );
  NAND2_X1 U8495 ( .A1(n7964), .A2(n7004), .ZN(n8161) );
  NAND2_X1 U8496 ( .A1(n7608), .A2(n7607), .ZN(n8000) );
  INV_X1 U8497 ( .A(n8091), .ZN(n8156) );
  NAND2_X1 U8498 ( .A1(n7598), .A2(n7597), .ZN(n7934) );
  NAND2_X1 U8499 ( .A1(n7588), .A2(n7340), .ZN(n7877) );
  NAND2_X1 U8500 ( .A1(n7586), .A2(n7588), .ZN(n7875) );
  INV_X1 U8501 ( .A(n7964), .ZN(n7963) );
  OAI21_X1 U8502 ( .B1(n7726), .B2(n6935), .A(n6933), .ZN(n7747) );
  AOI21_X1 U8503 ( .B1(n7731), .B2(n6934), .A(n6936), .ZN(n6933) );
  INV_X1 U8504 ( .A(n7560), .ZN(n6936) );
  OR2_X1 U8505 ( .A1(n7737), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7751) );
  AND2_X1 U8506 ( .A1(n7734), .A2(n7733), .ZN(n9943) );
  NAND2_X1 U8507 ( .A1(n7732), .A2(n7731), .ZN(n7734) );
  NAND2_X1 U8508 ( .A1(n7726), .A2(n7556), .ZN(n7732) );
  INV_X1 U8509 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7631) );
  INV_X1 U8510 ( .A(n7548), .ZN(n7309) );
  NAND2_X1 U8511 ( .A1(n7311), .A2(n7548), .ZN(n7679) );
  NAND2_X1 U8512 ( .A1(n14427), .A2(n14426), .ZN(n14473) );
  NAND2_X1 U8513 ( .A1(n7058), .A2(n14477), .ZN(n14478) );
  AOI21_X1 U8514 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14436), .A(n14435), .ZN(
        n14446) );
  AOI21_X1 U8515 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14441), .A(n14440), .ZN(
        n14491) );
  NOR2_X1 U8516 ( .A1(n14487), .A2(n14486), .ZN(n14440) );
  AND2_X1 U8517 ( .A1(n6889), .A2(n7056), .ZN(n14500) );
  NAND2_X1 U8518 ( .A1(n7400), .A2(n7401), .ZN(n11597) );
  INV_X1 U8519 ( .A(n7402), .ZN(n7401) );
  OAI21_X1 U8520 ( .B1(n11497), .B2(n7403), .A(n11594), .ZN(n7402) );
  NAND2_X1 U8521 ( .A1(n11509), .A2(n11500), .ZN(n11501) );
  NAND2_X1 U8522 ( .A1(n9500), .A2(n9499), .ZN(n13037) );
  NAND2_X1 U8523 ( .A1(n6813), .A2(n6817), .ZN(n12488) );
  NAND2_X1 U8524 ( .A1(n6819), .A2(n6710), .ZN(n6813) );
  AND2_X1 U8525 ( .A1(n11819), .A2(n11817), .ZN(n7415) );
  INV_X1 U8526 ( .A(n15138), .ZN(n11302) );
  OR2_X1 U8527 ( .A1(n7395), .A2(n7396), .ZN(n11025) );
  INV_X1 U8528 ( .A(n7399), .ZN(n7395) );
  NAND2_X1 U8529 ( .A1(n12560), .A2(n12308), .ZN(n12518) );
  NAND2_X1 U8530 ( .A1(n7422), .A2(n12285), .ZN(n12528) );
  NAND2_X1 U8531 ( .A1(n6826), .A2(n6825), .ZN(n12539) );
  NAND2_X1 U8532 ( .A1(n6827), .A2(n6620), .ZN(n6826) );
  INV_X1 U8533 ( .A(n12501), .ZN(n6827) );
  AND2_X1 U8534 ( .A1(n10994), .A2(n10993), .ZN(n10995) );
  NAND2_X1 U8535 ( .A1(n11731), .A2(n11730), .ZN(n11733) );
  NAND2_X1 U8536 ( .A1(n12562), .A2(n12561), .ZN(n12560) );
  NAND2_X1 U8537 ( .A1(n12501), .A2(n12305), .ZN(n12562) );
  INV_X1 U8538 ( .A(n12628), .ZN(n13001) );
  NAND2_X1 U8539 ( .A1(n6819), .A2(n12287), .ZN(n12570) );
  INV_X1 U8540 ( .A(n12790), .ZN(n12815) );
  NAND2_X1 U8541 ( .A1(n6820), .A2(n6821), .ZN(n12604) );
  AOI21_X1 U8542 ( .B1(n6823), .B2(n6822), .A(n6665), .ZN(n6821) );
  INV_X1 U8543 ( .A(n15040), .ZN(n12623) );
  INV_X1 U8544 ( .A(n12969), .ZN(n13002) );
  NAND2_X1 U8545 ( .A1(n12270), .A2(n10798), .ZN(n12618) );
  OR2_X1 U8546 ( .A1(n6814), .A2(n6723), .ZN(n6811) );
  INV_X1 U8547 ( .A(n15043), .ZN(n12613) );
  NAND2_X1 U8548 ( .A1(n10792), .A2(n10791), .ZN(n12620) );
  NOR2_X1 U8549 ( .A1(n12256), .A2(n12070), .ZN(n7179) );
  NAND2_X1 U8550 ( .A1(n7099), .A2(n7178), .ZN(n7177) );
  AND4_X1 U8551 ( .A1(n12066), .A2(n9540), .A3(n9539), .A4(n9538), .ZN(n12792)
         );
  NAND2_X1 U8552 ( .A1(n6855), .A2(n6629), .ZN(n12633) );
  OR2_X1 U8553 ( .A1(n12062), .A2(n11093), .ZN(n9122) );
  NAND4_X2 U8554 ( .A1(n9091), .A2(n9090), .A3(n9089), .A4(n9088), .ZN(n15116)
         );
  NAND2_X1 U8555 ( .A1(n9117), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U8556 ( .A1(n9117), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9067) );
  OR2_X1 U8557 ( .A1(n10964), .A2(n10669), .ZN(n10965) );
  NAND2_X1 U8558 ( .A1(n6737), .A2(n7255), .ZN(n11091) );
  AND2_X1 U8559 ( .A1(n9130), .A2(n9129), .ZN(n11127) );
  INV_X1 U8560 ( .A(n7263), .ZN(n15051) );
  OAI21_X1 U8561 ( .B1(n15060), .B2(n15059), .A(n15058), .ZN(n15062) );
  NAND2_X1 U8562 ( .A1(n15060), .A2(n6615), .ZN(n6901) );
  XNOR2_X1 U8563 ( .A(n11463), .B(n11464), .ZN(n11201) );
  NOR2_X1 U8564 ( .A1(n11201), .A2(n11207), .ZN(n11465) );
  INV_X1 U8565 ( .A(n7249), .ZN(n11886) );
  INV_X1 U8566 ( .A(n6870), .ZN(n11536) );
  AOI21_X1 U8567 ( .B1(n11541), .B2(n11540), .A(n6896), .ZN(n11543) );
  AND2_X1 U8568 ( .A1(n11538), .A2(n11539), .ZN(n6896) );
  XNOR2_X1 U8569 ( .A(n12638), .B(n12647), .ZN(n11888) );
  NOR2_X1 U8570 ( .A1(n11888), .A2(n13007), .ZN(n12639) );
  INV_X1 U8571 ( .A(n7260), .ZN(n12668) );
  INV_X1 U8572 ( .A(n6882), .ZN(n12643) );
  NOR2_X1 U8573 ( .A1(n12645), .A2(n6911), .ZN(n12653) );
  AND2_X1 U8574 ( .A1(n12646), .A2(n12647), .ZN(n6911) );
  NAND2_X1 U8575 ( .A1(n12653), .A2(n12652), .ZN(n12678) );
  XNOR2_X1 U8576 ( .A(n12701), .B(n14528), .ZN(n12682) );
  NOR2_X1 U8577 ( .A1(n12689), .A2(n12690), .ZN(n12692) );
  INV_X1 U8578 ( .A(n7259), .ZN(n12687) );
  NOR2_X1 U8579 ( .A1(n12692), .A2(n12691), .ZN(n12711) );
  NAND2_X1 U8580 ( .A1(n6876), .A2(n6874), .ZN(n12771) );
  OR2_X1 U8581 ( .A1(n12748), .A2(n12747), .ZN(n6876) );
  NAND2_X1 U8582 ( .A1(n6877), .A2(n6875), .ZN(n6874) );
  AND2_X1 U8583 ( .A1(n6878), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8584 ( .A1(n7241), .A2(n7240), .ZN(n12802) );
  NAND2_X1 U8585 ( .A1(n12822), .A2(n12192), .ZN(n12811) );
  OR2_X1 U8586 ( .A1(n12056), .A2(n11562), .ZN(n9471) );
  NAND2_X1 U8587 ( .A1(n7227), .A2(n9624), .ZN(n12923) );
  NAND2_X1 U8588 ( .A1(n11362), .A2(n9608), .ZN(n11365) );
  OR2_X1 U8589 ( .A1(n9583), .A2(n15172), .ZN(n15123) );
  INV_X1 U8590 ( .A(n13004), .ZN(n12991) );
  AND2_X2 U8591 ( .A1(n9652), .A2(n9651), .ZN(n15192) );
  INV_X1 U8592 ( .A(n12779), .ZN(n13097) );
  NAND2_X1 U8593 ( .A1(n9431), .A2(n9430), .ZN(n13130) );
  NAND2_X1 U8594 ( .A1(n9418), .A2(n9417), .ZN(n13136) );
  NAND2_X1 U8595 ( .A1(n9405), .A2(n9404), .ZN(n13142) );
  OAI21_X1 U8596 ( .B1(n9378), .B2(n7186), .A(n7184), .ZN(n12897) );
  OAI21_X1 U8597 ( .B1(n9622), .B2(n6847), .A(n6844), .ZN(n12911) );
  NAND2_X1 U8598 ( .A1(n12927), .A2(n12166), .ZN(n12907) );
  AND2_X1 U8599 ( .A1(n15177), .A2(n15155), .ZN(n13148) );
  NAND2_X1 U8600 ( .A1(n9275), .A2(n9274), .ZN(n12531) );
  NAND2_X1 U8601 ( .A1(n7221), .A2(n7220), .ZN(n11905) );
  OAI21_X1 U8602 ( .B1(n12270), .B2(n11071), .A(n11070), .ZN(n11076) );
  AND2_X1 U8603 ( .A1(n10781), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10016) );
  INV_X1 U8604 ( .A(n9063), .ZN(n13186) );
  XNOR2_X1 U8605 ( .A(n9554), .B(n9553), .ZN(n11560) );
  OAI21_X1 U8606 ( .B1(n9552), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9554) );
  NAND4_X1 U8607 ( .A1(n6834), .A2(n6833), .A3(n6835), .A4(n6836), .ZN(n11387)
         );
  NAND2_X1 U8608 ( .A1(n9551), .A2(n9056), .ZN(n6836) );
  OR2_X1 U8609 ( .A1(n6838), .A2(n6837), .ZN(n6835) );
  OR2_X1 U8610 ( .A1(n9317), .A2(n6837), .ZN(n6834) );
  NAND2_X1 U8611 ( .A1(n9444), .A2(n9443), .ZN(n9454) );
  AND2_X1 U8612 ( .A1(n7046), .A2(P3_U3151), .ZN(n13179) );
  NAND2_X1 U8613 ( .A1(n6623), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9543) );
  INV_X1 U8614 ( .A(SI_16_), .ZN(n15328) );
  NAND2_X1 U8615 ( .A1(n7086), .A2(n9333), .ZN(n9347) );
  NAND2_X1 U8616 ( .A1(n9332), .A2(n9331), .ZN(n7086) );
  INV_X1 U8617 ( .A(SI_11_), .ZN(n15425) );
  NAND2_X1 U8618 ( .A1(n9251), .A2(n9250), .ZN(n9269) );
  INV_X1 U8619 ( .A(SI_10_), .ZN(n9982) );
  NAND2_X1 U8620 ( .A1(n7107), .A2(n7105), .ZN(n9204) );
  NAND2_X1 U8621 ( .A1(n7107), .A2(n7108), .ZN(n9183) );
  NAND2_X1 U8622 ( .A1(n9168), .A2(n9167), .ZN(n9180) );
  INV_X1 U8623 ( .A(n9156), .ZN(n9153) );
  NAND2_X1 U8624 ( .A1(n7095), .A2(n9133), .ZN(n9136) );
  NAND2_X1 U8625 ( .A1(n9099), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8626 ( .A1(n9105), .A2(n9104), .ZN(n9132) );
  AND2_X1 U8627 ( .A1(n9934), .A2(n9933), .ZN(n14576) );
  NAND2_X1 U8628 ( .A1(n8578), .A2(n8577), .ZN(n13647) );
  NAND2_X1 U8629 ( .A1(n11184), .A2(n11183), .ZN(n11231) );
  AOI21_X1 U8630 ( .B1(n7501), .B2(n11189), .A(n7500), .ZN(n7503) );
  INV_X1 U8631 ( .A(n7495), .ZN(n7490) );
  NAND2_X1 U8632 ( .A1(n7493), .A2(n7489), .ZN(n7488) );
  INV_X1 U8633 ( .A(n7498), .ZN(n7489) );
  AOI21_X1 U8634 ( .B1(n11939), .B2(n7499), .A(n7498), .ZN(n11943) );
  AND2_X1 U8635 ( .A1(n7485), .A2(n7486), .ZN(n13293) );
  INV_X1 U8636 ( .A(n9924), .ZN(n7516) );
  INV_X1 U8637 ( .A(n9925), .ZN(n7517) );
  AND2_X1 U8638 ( .A1(n7513), .A2(n7512), .ZN(n13309) );
  NAND2_X1 U8639 ( .A1(n11448), .A2(n11447), .ZN(n11867) );
  NAND2_X1 U8640 ( .A1(n11229), .A2(n11189), .ZN(n11420) );
  NOR2_X1 U8641 ( .A1(n13191), .A2(n13190), .ZN(n13327) );
  NAND2_X1 U8642 ( .A1(n10655), .A2(n10654), .ZN(n10657) );
  AND2_X1 U8643 ( .A1(n9020), .A2(n6750), .ZN(n6749) );
  INV_X1 U8644 ( .A(n13282), .ZN(n13358) );
  AND2_X1 U8645 ( .A1(n8267), .A2(n8266), .ZN(n8269) );
  NAND2_X1 U8646 ( .A1(n8928), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8270) );
  OR2_X1 U8647 ( .A1(n14835), .A2(n14834), .ZN(n14837) );
  NOR2_X1 U8648 ( .A1(n6598), .A2(n6655), .ZN(n7197) );
  OR2_X1 U8649 ( .A1(n13472), .A2(n13425), .ZN(n7196) );
  NAND2_X1 U8650 ( .A1(n7469), .A2(n8703), .ZN(n13465) );
  NAND2_X1 U8651 ( .A1(n7469), .A2(n7467), .ZN(n13625) );
  NAND2_X1 U8652 ( .A1(n13488), .A2(n8607), .ZN(n13469) );
  AND2_X1 U8653 ( .A1(n8600), .A2(n8599), .ZN(n13487) );
  NAND2_X1 U8654 ( .A1(n7158), .A2(n6613), .ZN(n13567) );
  NAND2_X1 U8655 ( .A1(n11954), .A2(n8689), .ZN(n13602) );
  NAND2_X1 U8656 ( .A1(n14588), .A2(n7478), .ZN(n11678) );
  NAND2_X1 U8657 ( .A1(n7480), .A2(n9010), .ZN(n14588) );
  INV_X1 U8658 ( .A(n11590), .ZN(n7480) );
  NAND2_X1 U8659 ( .A1(n7455), .A2(n7456), .ZN(n11396) );
  NAND2_X1 U8660 ( .A1(n7461), .A2(n8680), .ZN(n11242) );
  NAND2_X1 U8661 ( .A1(n7463), .A2(n7462), .ZN(n7461) );
  NAND2_X1 U8662 ( .A1(n10382), .A2(n8668), .ZN(n10597) );
  NAND2_X1 U8663 ( .A1(n8320), .A2(n8319), .ZN(n10387) );
  NAND2_X1 U8664 ( .A1(n7194), .A2(n10340), .ZN(n10304) );
  INV_X1 U8665 ( .A(n10230), .ZN(n7194) );
  INV_X1 U8666 ( .A(n13604), .ZN(n15196) );
  NAND2_X1 U8667 ( .A1(n14963), .A2(n9931), .ZN(n15200) );
  OAI22_X1 U8668 ( .A1(n8273), .A2(n15286), .B1(n8277), .B2(n14771), .ZN(n6748) );
  INV_X1 U8669 ( .A(n8991), .ZN(n13694) );
  AND2_X1 U8670 ( .A1(n13613), .A2(n13612), .ZN(n13695) );
  OR2_X1 U8671 ( .A1(n13620), .A2(n13682), .ZN(n6752) );
  OR2_X1 U8672 ( .A1(n11530), .A2(n8274), .ZN(n8542) );
  AND2_X1 U8673 ( .A1(n9927), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14963) );
  NAND2_X1 U8674 ( .A1(n8740), .A2(n8739), .ZN(n14962) );
  NAND2_X1 U8675 ( .A1(n8648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7487) );
  INV_X1 U8676 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11520) );
  INV_X1 U8677 ( .A(n11409), .ZN(n13581) );
  INV_X1 U8678 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11081) );
  INV_X1 U8679 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n15492) );
  INV_X1 U8680 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10842) );
  INV_X1 U8681 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10224) );
  INV_X1 U8682 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10150) );
  INV_X1 U8683 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10011) );
  INV_X1 U8684 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9992) );
  INV_X1 U8685 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9986) );
  INV_X1 U8686 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9952) );
  INV_X1 U8687 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9942) );
  INV_X1 U8688 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9940) );
  INV_X1 U8689 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U8690 ( .A1(n7047), .A2(SI_0_), .ZN(n8276) );
  NOR2_X1 U8691 ( .A1(n11932), .A2(n14414), .ZN(n8183) );
  NAND2_X1 U8692 ( .A1(n11253), .A2(n11252), .ZN(n11568) );
  NAND2_X1 U8693 ( .A1(n13846), .A2(n12387), .ZN(n13745) );
  NAND2_X1 U8694 ( .A1(n10898), .A2(n10897), .ZN(n10899) );
  INV_X1 U8695 ( .A(n12434), .ZN(n10897) );
  INV_X1 U8696 ( .A(n12435), .ZN(n10898) );
  NAND2_X1 U8697 ( .A1(n13856), .A2(n7304), .ZN(n13755) );
  NOR2_X1 U8698 ( .A1(n13753), .A2(n7305), .ZN(n7304) );
  INV_X1 U8699 ( .A(n12360), .ZN(n7305) );
  NAND2_X1 U8700 ( .A1(n11568), .A2(n11567), .ZN(n11571) );
  AND2_X1 U8701 ( .A1(n13763), .A2(n13764), .ZN(n13765) );
  NAND2_X1 U8702 ( .A1(n13825), .A2(n12375), .ZN(n13776) );
  NAND2_X1 U8703 ( .A1(n13877), .A2(n13880), .ZN(n13794) );
  OAI21_X1 U8704 ( .B1(n12338), .B2(n6995), .A(n6993), .ZN(n13792) );
  AND2_X1 U8705 ( .A1(n10926), .A2(n10927), .ZN(n6983) );
  INV_X1 U8706 ( .A(n14338), .ZN(n13815) );
  AOI21_X1 U8707 ( .B1(n6998), .B2(n7000), .A(n6672), .ZN(n6997) );
  OAI21_X1 U8708 ( .B1(n10370), .B2(n7293), .A(n10372), .ZN(n13932) );
  NAND2_X1 U8709 ( .A1(n12326), .A2(n7291), .ZN(n13837) );
  AND2_X1 U8710 ( .A1(n7300), .A2(n7297), .ZN(n12006) );
  AND2_X1 U8711 ( .A1(n7299), .A2(n6636), .ZN(n7297) );
  NOR2_X1 U8712 ( .A1(n13765), .A2(n10373), .ZN(n10377) );
  NAND2_X1 U8713 ( .A1(n10909), .A2(n6736), .ZN(n6982) );
  NAND2_X1 U8714 ( .A1(n6986), .A2(n12410), .ZN(n13869) );
  NAND2_X1 U8715 ( .A1(n13784), .A2(n13785), .ZN(n6986) );
  OR2_X1 U8716 ( .A1(n10269), .A2(n10268), .ZN(n13889) );
  AOI21_X1 U8717 ( .B1(n9887), .B2(n9886), .A(n9888), .ZN(n9889) );
  INV_X1 U8718 ( .A(n12457), .ZN(n14092) );
  CLKBUF_X1 U8719 ( .A(n13918), .Z(n6758) );
  CLKBUF_X1 U8720 ( .A(P1_ADDR_REG_19__SCAN_IN), .Z(n14554) );
  INV_X1 U8721 ( .A(n9880), .ZN(n6802) );
  AOI21_X1 U8722 ( .B1(n7127), .B2(n7130), .A(n7126), .ZN(n8090) );
  NAND2_X1 U8723 ( .A1(n6942), .A2(n6944), .ZN(n14110) );
  NAND2_X1 U8724 ( .A1(n6943), .A2(n8134), .ZN(n14111) );
  NAND2_X1 U8725 ( .A1(n14144), .A2(n8133), .ZN(n14124) );
  NAND2_X1 U8726 ( .A1(n14178), .A2(n8026), .ZN(n14174) );
  INV_X1 U8727 ( .A(n14380), .ZN(n14186) );
  NAND2_X1 U8728 ( .A1(n14204), .A2(n8127), .ZN(n14190) );
  NAND2_X1 U8729 ( .A1(n7979), .A2(n7978), .ZN(n14207) );
  NAND2_X1 U8730 ( .A1(n7113), .A2(n7957), .ZN(n14228) );
  NAND2_X1 U8731 ( .A1(n6958), .A2(n6962), .ZN(n14247) );
  OR2_X1 U8732 ( .A1(n11970), .A2(n6963), .ZN(n6958) );
  NAND2_X1 U8733 ( .A1(n8120), .A2(n8119), .ZN(n12021) );
  NAND2_X1 U8734 ( .A1(n11968), .A2(n7931), .ZN(n12018) );
  NAND2_X1 U8735 ( .A1(n11837), .A2(n7892), .ZN(n11785) );
  NAND2_X1 U8736 ( .A1(n8114), .A2(n8113), .ZN(n11628) );
  INV_X1 U8737 ( .A(n14536), .ZN(n12001) );
  NAND2_X1 U8738 ( .A1(n11278), .A2(n8112), .ZN(n11435) );
  NAND2_X1 U8739 ( .A1(n11290), .A2(n11289), .ZN(n11288) );
  NAND2_X1 U8740 ( .A1(n11336), .A2(n7821), .ZN(n11290) );
  INV_X1 U8741 ( .A(n14251), .ZN(n14706) );
  NAND2_X1 U8742 ( .A1(n7125), .A2(n9860), .ZN(n10555) );
  OR2_X1 U8743 ( .A1(n10512), .A2(n6972), .ZN(n7125) );
  INV_X1 U8744 ( .A(n14248), .ZN(n14229) );
  INV_X1 U8745 ( .A(n14047), .ZN(n14358) );
  AND2_X1 U8746 ( .A1(n9665), .A2(n9664), .ZN(n14360) );
  INV_X1 U8747 ( .A(n14101), .ZN(n14366) );
  INV_X1 U8748 ( .A(n14135), .ZN(n14371) );
  INV_X1 U8749 ( .A(n6770), .ZN(n14376) );
  NAND2_X1 U8750 ( .A1(n14415), .A2(n8016), .ZN(n14380) );
  NAND2_X1 U8751 ( .A1(n7839), .A2(n7838), .ZN(n11525) );
  NAND2_X1 U8752 ( .A1(n10149), .A2(n9675), .ZN(n7827) );
  NAND2_X1 U8753 ( .A1(n7062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7641) );
  XNOR2_X1 U8754 ( .A(n8076), .B(n8078), .ZN(n14406) );
  NAND2_X1 U8755 ( .A1(n8063), .A2(n8062), .ZN(n14412) );
  NAND2_X1 U8756 ( .A1(n7342), .A2(n7623), .ZN(n8063) );
  INV_X1 U8757 ( .A(n7343), .ZN(n7342) );
  OR2_X1 U8758 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  NAND2_X1 U8759 ( .A1(n8091), .A2(n7307), .ZN(n8152) );
  INV_X1 U8760 ( .A(n8150), .ZN(n11644) );
  INV_X1 U8761 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11531) );
  INV_X1 U8762 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10941) );
  INV_X1 U8763 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10844) );
  INV_X1 U8764 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10592) );
  NOR2_X1 U8765 ( .A1(n7046), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14395) );
  INV_X1 U8766 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10151) );
  INV_X1 U8767 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9994) );
  INV_X1 U8768 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9984) );
  INV_X1 U8769 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9954) );
  AND2_X1 U8770 ( .A1(n9945), .A2(SI_0_), .ZN(n7697) );
  INV_X1 U8771 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14455) );
  XNOR2_X1 U8772 ( .A(n14456), .B(n6789), .ZN(n15524) );
  INV_X1 U8773 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6789) );
  AOI21_X1 U8774 ( .B1(n14521), .B2(n14459), .A(n14518), .ZN(n15521) );
  XNOR2_X1 U8775 ( .A(n14450), .B(n14787), .ZN(n15514) );
  XNOR2_X1 U8776 ( .A(n14476), .B(n6892), .ZN(n15518) );
  INV_X1 U8777 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8778 ( .A1(n14484), .A2(n14485), .ZN(n14533) );
  NAND2_X1 U8779 ( .A1(n14530), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n14484) );
  OAI21_X2 U8780 ( .B1(n14489), .B2(n14488), .A(n14633), .ZN(n14638) );
  NOR2_X1 U8781 ( .A1(n14634), .A2(n14635), .ZN(n14489) );
  AND2_X1 U8782 ( .A1(n14500), .A2(n14501), .ZN(n14645) );
  XNOR2_X1 U8783 ( .A(n12314), .B(n7413), .ZN(n12500) );
  INV_X1 U8784 ( .A(n6871), .ZN(n11534) );
  NAND2_X1 U8785 ( .A1(n6877), .A2(n12748), .ZN(n12714) );
  AOI211_X1 U8786 ( .C1(n15080), .C2(n12768), .A(n12767), .B(n12766), .ZN(
        n12777) );
  INV_X1 U8787 ( .A(n9655), .ZN(n9656) );
  MUX2_X1 U8788 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n13098), .S(n15192), .Z(
        n9653) );
  MUX2_X1 U8789 ( .A(n13034), .B(n13104), .S(n15192), .Z(n13035) );
  INV_X1 U8790 ( .A(n7242), .ZN(n13102) );
  OAI21_X1 U8791 ( .B1(n9645), .B2(n7245), .A(n7243), .ZN(n7242) );
  NAND2_X1 U8792 ( .A1(n15177), .A2(n15114), .ZN(n7245) );
  MUX2_X1 U8793 ( .A(n13105), .B(n13104), .S(n15177), .Z(n13106) );
  OAI222_X1 U8794 ( .A1(n14525), .A2(n10216), .B1(n12642), .B2(P3_U3151), .C1(
        n11389), .C2(n10215), .ZN(P3_U3281) );
  INV_X1 U8795 ( .A(n13233), .ZN(n6761) );
  INV_X1 U8796 ( .A(n6797), .ZN(n6796) );
  OAI211_X1 U8797 ( .C1(n8663), .C2(n7143), .A(n6924), .B(n8744), .ZN(n6786)
         );
  NOR2_X1 U8798 ( .A1(n7537), .A2(n9640), .ZN(n9641) );
  NAND2_X1 U8799 ( .A1(n7283), .A2(n7287), .ZN(n14612) );
  NAND2_X1 U8800 ( .A1(n6975), .A2(n6974), .ZN(n14087) );
  AOI21_X1 U8801 ( .B1(n6953), .B2(n14752), .A(n6603), .ZN(n6951) );
  NOR2_X1 U8802 ( .A1(n14751), .A2(n14329), .ZN(n6952) );
  INV_X1 U8803 ( .A(n6885), .ZN(n14629) );
  INV_X1 U8804 ( .A(n6889), .ZN(n14641) );
  INV_X1 U8805 ( .A(n6746), .ZN(n14648) );
  NOR2_X1 U8806 ( .A1(n14550), .A2(n14549), .ZN(n14559) );
  INV_X1 U8807 ( .A(n7507), .ZN(n13300) );
  NOR2_X1 U8808 ( .A1(n12478), .A2(n12477), .ZN(n6587) );
  INV_X2 U8809 ( .A(n8747), .ZN(n8968) );
  INV_X1 U8810 ( .A(n8968), .ZN(n8992) );
  INV_X2 U8811 ( .A(n8968), .ZN(n8993) );
  INV_X1 U8812 ( .A(n12898), .ZN(n12896) );
  AND2_X1 U8813 ( .A1(n6854), .A2(n12900), .ZN(n6588) );
  INV_X1 U8814 ( .A(n11341), .ZN(n7265) );
  NAND2_X1 U8815 ( .A1(n6872), .A2(n12730), .ZN(n6877) );
  AND2_X1 U8816 ( .A1(n12285), .A2(n6717), .ZN(n6589) );
  AND2_X1 U8817 ( .A1(n13516), .A2(n6616), .ZN(n6590) );
  INV_X1 U8818 ( .A(n12110), .ZN(n7167) );
  AND2_X1 U8819 ( .A1(n7065), .A2(n14081), .ZN(n6591) );
  AND2_X1 U8820 ( .A1(n7337), .A2(n6715), .ZN(n6592) );
  AND2_X1 U8821 ( .A1(n10921), .A2(n7070), .ZN(n6593) );
  INV_X1 U8822 ( .A(n9873), .ZN(n11969) );
  XOR2_X1 U8823 ( .A(n8937), .B(n8639), .Z(n6594) );
  AND2_X1 U8824 ( .A1(n8842), .A2(n8841), .ZN(n6595) );
  AND2_X1 U8825 ( .A1(n7584), .A2(n7848), .ZN(n6596) );
  INV_X1 U8826 ( .A(n8875), .ZN(n7381) );
  AND2_X1 U8827 ( .A1(n7184), .A2(n7186), .ZN(n6597) );
  AND2_X1 U8828 ( .A1(n7201), .A2(n7203), .ZN(n6598) );
  OR2_X1 U8829 ( .A1(n8016), .A2(n6954), .ZN(n6599) );
  NAND2_X1 U8830 ( .A1(n11158), .A2(n11159), .ZN(n6600) );
  NAND2_X1 U8831 ( .A1(n12479), .A2(n6829), .ZN(n6601) );
  INV_X1 U8832 ( .A(n7457), .ZN(n7456) );
  NAND2_X1 U8833 ( .A1(n6673), .A2(n7458), .ZN(n7457) );
  INV_X1 U8834 ( .A(n8903), .ZN(n7357) );
  INV_X1 U8835 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8095) );
  INV_X1 U8836 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9334) );
  AND4_X1 U8837 ( .A1(n9334), .A2(n7406), .A3(n9051), .A4(n9054), .ZN(n6602)
         );
  NAND2_X1 U8838 ( .A1(n7535), .A2(n7532), .ZN(n6603) );
  AND2_X1 U8839 ( .A1(n14978), .A2(n7208), .ZN(n6604) );
  AND2_X1 U8840 ( .A1(n6736), .A2(n10927), .ZN(n6605) );
  AND2_X1 U8841 ( .A1(n12225), .A2(n12224), .ZN(n6606) );
  AOI21_X1 U8842 ( .B1(n7410), .B2(n7409), .A(n6667), .ZN(n7408) );
  NOR2_X1 U8843 ( .A1(n14376), .A2(n14141), .ZN(n6607) );
  OR2_X1 U8844 ( .A1(n12313), .A2(n12627), .ZN(n6608) );
  NAND2_X1 U8845 ( .A1(n7205), .A2(n7206), .ZN(n13573) );
  INV_X1 U8846 ( .A(n13573), .ZN(n6914) );
  NAND2_X1 U8847 ( .A1(n8480), .A2(n8479), .ZN(n11878) );
  INV_X1 U8848 ( .A(n11878), .ZN(n7210) );
  INV_X1 U8849 ( .A(n14617), .ZN(n7071) );
  AND2_X1 U8850 ( .A1(n7621), .A2(SI_26_), .ZN(n6609) );
  AND2_X1 U8851 ( .A1(n8037), .A2(n7621), .ZN(n6610) );
  NAND2_X1 U8852 ( .A1(n7251), .A2(n11099), .ZN(n7255) );
  INV_X1 U8853 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7918) );
  INV_X1 U8854 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13724) );
  AND2_X1 U8855 ( .A1(n7120), .A2(n14147), .ZN(n6611) );
  OR2_X1 U8856 ( .A1(n14218), .A2(n14315), .ZN(n6612) );
  INV_X1 U8857 ( .A(n13950), .ZN(n6954) );
  XNOR2_X1 U8858 ( .A(n6883), .B(n9046), .ZN(n11099) );
  AND2_X1 U8859 ( .A1(n7157), .A2(n8540), .ZN(n6613) );
  AND4_X1 U8860 ( .A1(n9048), .A2(n9165), .A3(n9186), .A4(n9047), .ZN(n6614)
         );
  AND2_X1 U8861 ( .A1(n6907), .A2(n15058), .ZN(n6615) );
  OR2_X1 U8862 ( .A1(n13537), .A2(n13274), .ZN(n6616) );
  AND2_X1 U8863 ( .A1(n14113), .A2(n7065), .ZN(n6617) );
  NOR2_X1 U8864 ( .A1(n8893), .A2(n8892), .ZN(n6618) );
  NAND2_X1 U8865 ( .A1(n13630), .A2(n13356), .ZN(n6619) );
  AND2_X1 U8866 ( .A1(n6587), .A2(n7408), .ZN(n6620) );
  AND2_X1 U8867 ( .A1(n8690), .A2(n8689), .ZN(n6621) );
  INV_X1 U8868 ( .A(n7186), .ZN(n7185) );
  OR2_X1 U8869 ( .A1(n12162), .A2(n7187), .ZN(n7186) );
  OR2_X1 U8870 ( .A1(n12332), .A2(n12331), .ZN(n6622) );
  NAND2_X1 U8871 ( .A1(n9542), .A2(n9541), .ZN(n6623) );
  OR2_X1 U8872 ( .A1(n9076), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n6624) );
  AND2_X1 U8873 ( .A1(n7417), .A2(n9283), .ZN(n6625) );
  INV_X1 U8874 ( .A(n15065), .ZN(n11161) );
  OR2_X1 U8875 ( .A1(n11539), .A2(n11533), .ZN(n6626) );
  AND2_X1 U8876 ( .A1(n6908), .A2(n12758), .ZN(n6627) );
  AND2_X1 U8877 ( .A1(n13537), .A2(n13274), .ZN(n6628) );
  XNOR2_X1 U8878 ( .A(n7424), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10803) );
  AND2_X1 U8879 ( .A1(n9164), .A2(n9163), .ZN(n6629) );
  AND2_X1 U8880 ( .A1(n7686), .A2(n7631), .ZN(n7706) );
  INV_X1 U8881 ( .A(n13617), .ZN(n7202) );
  INV_X1 U8882 ( .A(n13705), .ZN(n8905) );
  NAND2_X1 U8883 ( .A1(n11871), .A2(n11870), .ZN(n6630) );
  AND2_X1 U8884 ( .A1(n13227), .A2(n13223), .ZN(n6631) );
  INV_X1 U8885 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9046) );
  INV_X1 U8886 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9045) );
  INV_X1 U8887 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n6864) );
  AND4_X1 U8888 ( .A1(n9551), .A2(n9576), .A3(n9283), .A4(n9553), .ZN(n6632)
         );
  INV_X1 U8889 ( .A(n13228), .ZN(n13623) );
  NAND2_X1 U8890 ( .A1(n7025), .A2(n8235), .ZN(n13228) );
  NAND2_X1 U8891 ( .A1(n12214), .A2(n12215), .ZN(n12799) );
  OR2_X1 U8892 ( .A1(n7183), .A2(n12896), .ZN(n6633) );
  AND2_X1 U8893 ( .A1(n10921), .A2(n8104), .ZN(n6634) );
  AND2_X1 U8894 ( .A1(n14978), .A2(n8670), .ZN(n6635) );
  NAND2_X1 U8895 ( .A1(n12218), .A2(n12221), .ZN(n12789) );
  INV_X1 U8896 ( .A(n12789), .ZN(n12786) );
  NAND2_X1 U8897 ( .A1(n11983), .A2(n11982), .ZN(n6636) );
  AND2_X1 U8898 ( .A1(n13630), .A2(n8997), .ZN(n6637) );
  AND2_X1 U8899 ( .A1(n7267), .A2(n7265), .ZN(n6638) );
  AND2_X1 U8900 ( .A1(n12335), .A2(n12334), .ZN(n6639) );
  AND2_X1 U8901 ( .A1(n7119), .A2(n7120), .ZN(n6640) );
  AND2_X1 U8902 ( .A1(n13446), .A2(n7467), .ZN(n6641) );
  AND3_X1 U8903 ( .A1(n7691), .A2(n7690), .A3(n7689), .ZN(n10631) );
  AND2_X1 U8904 ( .A1(n8800), .A2(n8795), .ZN(n6642) );
  AND2_X1 U8905 ( .A1(n8800), .A2(n8791), .ZN(n6643) );
  NAND2_X1 U8906 ( .A1(n7414), .A2(n9046), .ZN(n9126) );
  AND2_X1 U8907 ( .A1(n12017), .A2(n8119), .ZN(n6644) );
  NOR2_X1 U8908 ( .A1(n8203), .A2(n7131), .ZN(n7130) );
  AND2_X1 U8909 ( .A1(n12346), .A2(n12345), .ZN(n6645) );
  AND2_X1 U8910 ( .A1(n10996), .A2(n10993), .ZN(n6646) );
  INV_X1 U8911 ( .A(n10340), .ZN(n7193) );
  INV_X1 U8912 ( .A(n11189), .ZN(n7504) );
  INV_X1 U8913 ( .A(n15070), .ZN(n6906) );
  INV_X1 U8914 ( .A(n8937), .ZN(n6921) );
  INV_X1 U8915 ( .A(n13537), .ZN(n13709) );
  NAND2_X1 U8916 ( .A1(n9317), .A2(n9547), .ZN(n6647) );
  AND2_X1 U8917 ( .A1(n10386), .A2(n10429), .ZN(n6649) );
  AND2_X1 U8918 ( .A1(n7416), .A2(n11730), .ZN(n6650) );
  INV_X1 U8919 ( .A(n9804), .ZN(n7447) );
  INV_X1 U8920 ( .A(n12160), .ZN(n12937) );
  AND2_X1 U8921 ( .A1(n12163), .A2(n12169), .ZN(n12160) );
  AND2_X1 U8922 ( .A1(n11569), .A2(n11567), .ZN(n6651) );
  NAND2_X1 U8923 ( .A1(n8135), .A2(n8075), .ZN(n14108) );
  INV_X1 U8924 ( .A(n6903), .ZN(n6902) );
  NOR2_X1 U8925 ( .A1(n6904), .A2(n11155), .ZN(n6903) );
  AND2_X1 U8926 ( .A1(n12416), .A2(n12415), .ZN(n6652) );
  AND2_X1 U8927 ( .A1(n13537), .A2(n13360), .ZN(n6653) );
  AND2_X1 U8928 ( .A1(n12560), .A2(n7410), .ZN(n6654) );
  AND2_X1 U8929 ( .A1(n7203), .A2(n13228), .ZN(n6655) );
  MUX2_X1 U8930 ( .A(n13935), .B(n14416), .S(n8016), .Z(n10771) );
  INV_X1 U8931 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7648) );
  OR2_X1 U8932 ( .A1(n13066), .A2(n12900), .ZN(n12172) );
  INV_X1 U8933 ( .A(n8679), .ZN(n7462) );
  NOR2_X1 U8934 ( .A1(n11863), .A2(n13907), .ZN(n6656) );
  NOR2_X1 U8935 ( .A1(n13843), .A2(n12328), .ZN(n6657) );
  NOR2_X1 U8936 ( .A1(n11525), .A2(n11998), .ZN(n6658) );
  NOR2_X1 U8937 ( .A1(n14351), .A2(n13902), .ZN(n6659) );
  NOR2_X1 U8938 ( .A1(n14745), .A2(n11721), .ZN(n6660) );
  NOR2_X1 U8939 ( .A1(n9768), .A2(n6578), .ZN(n6661) );
  NOR2_X1 U8940 ( .A1(n13142), .A2(n12522), .ZN(n6662) );
  INV_X1 U8941 ( .A(n7290), .ZN(n7289) );
  NAND2_X1 U8942 ( .A1(n6622), .A2(n7291), .ZN(n7290) );
  INV_X1 U8943 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9944) );
  INV_X1 U8944 ( .A(n7411), .ZN(n7410) );
  OR2_X1 U8945 ( .A1(n12519), .A2(n7412), .ZN(n7411) );
  INV_X1 U8946 ( .A(n11155), .ZN(n6907) );
  INV_X1 U8947 ( .A(n6851), .ZN(n6850) );
  NOR2_X1 U8948 ( .A1(n12959), .A2(n12940), .ZN(n6851) );
  NAND2_X1 U8949 ( .A1(n12823), .A2(n12205), .ZN(n6663) );
  AND2_X1 U8950 ( .A1(n7581), .A2(n15425), .ZN(n6664) );
  NOR2_X1 U8951 ( .A1(n12481), .A2(n12626), .ZN(n6665) );
  OR2_X1 U8952 ( .A1(n9297), .A2(n7528), .ZN(n6666) );
  AND2_X1 U8953 ( .A1(n12310), .A2(n12880), .ZN(n6667) );
  AND2_X1 U8954 ( .A1(n14598), .A2(n13369), .ZN(n6668) );
  INV_X1 U8955 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9350) );
  NAND2_X1 U8956 ( .A1(n8687), .A2(n9010), .ZN(n6669) );
  INV_X1 U8957 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U8958 ( .A1(n9239), .A2(n9238), .ZN(n6670) );
  OR2_X1 U8959 ( .A1(n14286), .A2(n13895), .ZN(n6671) );
  AND2_X1 U8960 ( .A1(n12394), .A2(n12393), .ZN(n6672) );
  OR2_X1 U8961 ( .A1(n11356), .A2(n11191), .ZN(n6673) );
  INV_X1 U8962 ( .A(n8703), .ZN(n7468) );
  AND2_X1 U8963 ( .A1(n13815), .A2(n14235), .ZN(n9772) );
  AND2_X1 U8964 ( .A1(n12633), .A2(n11496), .ZN(n6674) );
  INV_X1 U8965 ( .A(n7584), .ZN(n7031) );
  NOR2_X1 U8966 ( .A1(n14161), .A2(n7123), .ZN(n7122) );
  AND2_X1 U8967 ( .A1(n8874), .A2(n8873), .ZN(n6675) );
  INV_X1 U8968 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U8969 ( .A1(n7597), .A2(SI_17_), .ZN(n6676) );
  INV_X1 U8970 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9551) );
  INV_X1 U8971 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9980) );
  AND2_X1 U8972 ( .A1(n6696), .A2(n8907), .ZN(n6677) );
  NAND2_X1 U8973 ( .A1(n7645), .A2(n7644), .ZN(n14067) );
  INV_X1 U8974 ( .A(n14067), .ZN(n7064) );
  OR2_X1 U8975 ( .A1(n14479), .A2(n14478), .ZN(n6678) );
  OR2_X1 U8976 ( .A1(n7509), .A2(n13195), .ZN(n6679) );
  OR2_X1 U8977 ( .A1(n14969), .A2(n8968), .ZN(n6680) );
  AND3_X1 U8978 ( .A1(n9053), .A2(n9350), .A3(n9544), .ZN(n6681) );
  AND2_X1 U8979 ( .A1(n9601), .A2(n10807), .ZN(n6682) );
  AND2_X1 U8980 ( .A1(n13618), .A2(n6752), .ZN(n6683) );
  AND2_X1 U8981 ( .A1(n7486), .A2(n13292), .ZN(n6684) );
  INV_X1 U8982 ( .A(n13425), .ZN(n7203) );
  NAND2_X1 U8983 ( .A1(n8926), .A2(n8925), .ZN(n13425) );
  AND2_X1 U8984 ( .A1(n10732), .A2(n8673), .ZN(n6685) );
  AND2_X1 U8985 ( .A1(n8587), .A2(n8586), .ZN(n13705) );
  AND2_X1 U8986 ( .A1(n12205), .A2(n7176), .ZN(n6686) );
  OR2_X1 U8987 ( .A1(n6900), .A2(n15070), .ZN(n6687) );
  INV_X1 U8988 ( .A(n11500), .ZN(n7403) );
  NOR2_X1 U8989 ( .A1(n8118), .A2(n7117), .ZN(n7116) );
  NOR2_X1 U8990 ( .A1(n8681), .A2(n7460), .ZN(n7459) );
  AND2_X1 U8991 ( .A1(n7977), .A2(n7957), .ZN(n6688) );
  AND2_X1 U8992 ( .A1(n12779), .A2(n12780), .ZN(n12257) );
  INV_X1 U8993 ( .A(n12257), .ZN(n7099) );
  AND2_X1 U8994 ( .A1(n8784), .A2(n8783), .ZN(n6689) );
  AND2_X1 U8995 ( .A1(n10656), .A2(n10654), .ZN(n6690) );
  AND2_X1 U8996 ( .A1(n12377), .A2(n12375), .ZN(n6691) );
  OR2_X1 U8997 ( .A1(n9733), .A2(n9731), .ZN(n6692) );
  OR2_X1 U8998 ( .A1(n9724), .A2(n9722), .ZN(n6693) );
  OR2_X1 U8999 ( .A1(n9715), .A2(n9713), .ZN(n6694) );
  AND2_X1 U9000 ( .A1(n7066), .A2(n14092), .ZN(n6695) );
  NAND2_X1 U9001 ( .A1(n8904), .A2(n7357), .ZN(n6696) );
  OR2_X1 U9002 ( .A1(n9805), .A2(n7447), .ZN(n6697) );
  OR2_X1 U9003 ( .A1(n9815), .A2(n7429), .ZN(n6698) );
  AND2_X1 U9004 ( .A1(n6838), .A2(n9551), .ZN(n6699) );
  AND2_X1 U9005 ( .A1(n9626), .A2(n7224), .ZN(n6700) );
  AND2_X1 U9006 ( .A1(n13425), .A2(n7202), .ZN(n6701) );
  AND2_X1 U9007 ( .A1(n8908), .A2(n7355), .ZN(n6702) );
  AND2_X1 U9008 ( .A1(n6906), .A2(n6615), .ZN(n6703) );
  INV_X1 U9009 ( .A(n7270), .ZN(n7269) );
  AND2_X1 U9010 ( .A1(n6631), .A2(n14574), .ZN(n6704) );
  NAND2_X1 U9011 ( .A1(n7375), .A2(n7376), .ZN(n6705) );
  AND2_X1 U9012 ( .A1(n7153), .A2(n6616), .ZN(n6706) );
  OR2_X1 U9013 ( .A1(n13623), .A2(n13343), .ZN(n6707) );
  AND2_X1 U9014 ( .A1(n6825), .A2(n6824), .ZN(n6823) );
  AND2_X1 U9015 ( .A1(n8166), .A2(n7642), .ZN(n7434) );
  INV_X1 U9016 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8166) );
  INV_X1 U9017 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6928) );
  INV_X1 U9018 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7406) );
  NAND2_X1 U9019 ( .A1(n6625), .A2(n6839), .ZN(n9546) );
  INV_X1 U9020 ( .A(n9546), .ZN(n9317) );
  OR2_X1 U9021 ( .A1(n14362), .A2(n14361), .ZN(P1_U3526) );
  OR2_X1 U9022 ( .A1(n14262), .A2(n14261), .ZN(P1_U3558) );
  NAND2_X1 U9024 ( .A1(n9378), .A2(n9377), .ZN(n12927) );
  INV_X1 U9025 ( .A(SI_1_), .ZN(n7312) );
  AND2_X1 U9026 ( .A1(n6818), .A2(n12287), .ZN(n6710) );
  INV_X1 U9027 ( .A(n12625), .ZN(n12804) );
  NAND2_X1 U9028 ( .A1(n12955), .A2(n12152), .ZN(n12936) );
  INV_X1 U9029 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7421) );
  XNOR2_X1 U9030 ( .A(n11939), .B(n11940), .ZN(n11942) );
  OR2_X1 U9031 ( .A1(n9245), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U9032 ( .A1(n9218), .A2(n9219), .ZN(n9245) );
  AND2_X1 U9033 ( .A1(n8834), .A2(n8833), .ZN(n6712) );
  INV_X1 U9034 ( .A(n7206), .ZN(n13594) );
  INV_X1 U9035 ( .A(n7068), .ZN(n14239) );
  AND2_X1 U9036 ( .A1(n14588), .A2(n8685), .ZN(n6713) );
  OR2_X1 U9037 ( .A1(n12792), .A2(n13016), .ZN(n6714) );
  OR2_X1 U9038 ( .A1(n7946), .A2(SI_18_), .ZN(n6715) );
  AOI21_X1 U9039 ( .B1(n13354), .B2(n13316), .A(n8661), .ZN(n8662) );
  AND2_X1 U9040 ( .A1(n12791), .A2(n6714), .ZN(n6716) );
  NAND2_X1 U9041 ( .A1(n12526), .A2(n13001), .ZN(n6717) );
  AND2_X1 U9042 ( .A1(n12313), .A2(n12627), .ZN(n6718) );
  NAND2_X1 U9043 ( .A1(n12290), .A2(n13002), .ZN(n6719) );
  OR2_X1 U9044 ( .A1(n7961), .A2(n7599), .ZN(n6720) );
  AND2_X1 U9045 ( .A1(n7490), .A2(n7488), .ZN(n6721) );
  AND2_X1 U9046 ( .A1(n10941), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6722) );
  AND2_X1 U9047 ( .A1(n6710), .A2(n12489), .ZN(n6723) );
  AND2_X1 U9048 ( .A1(n8125), .A2(n8124), .ZN(n6724) );
  INV_X1 U9049 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9949) );
  INV_X1 U9050 ( .A(n13583), .ZN(n7205) );
  NAND2_X1 U9051 ( .A1(n9389), .A2(n9388), .ZN(n13066) );
  NAND2_X2 U9052 ( .A1(n11076), .A2(n11075), .ZN(n15177) );
  NOR2_X1 U9053 ( .A1(n11607), .A2(n12234), .ZN(n6725) );
  NAND2_X1 U9054 ( .A1(n7327), .A2(n8919), .ZN(n7326) );
  INV_X1 U9055 ( .A(n14325), .ZN(n7067) );
  AND2_X1 U9056 ( .A1(n12288), .A2(n12491), .ZN(n6726) );
  NOR2_X1 U9057 ( .A1(n11465), .A2(n11466), .ZN(n6727) );
  INV_X1 U9058 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7148) );
  AND2_X1 U9059 ( .A1(n6901), .A2(n6900), .ZN(n6728) );
  INV_X1 U9060 ( .A(n7621), .ZN(n7017) );
  AND2_X1 U9061 ( .A1(n6901), .A2(n6902), .ZN(n6729) );
  INV_X1 U9062 ( .A(n7213), .ZN(n11407) );
  AND2_X1 U9063 ( .A1(n6916), .A2(n14942), .ZN(n7213) );
  OR2_X1 U9064 ( .A1(n11209), .A2(n11210), .ZN(n6898) );
  AND2_X1 U9065 ( .A1(n7125), .A2(n7124), .ZN(n6730) );
  AND2_X1 U9066 ( .A1(n11697), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6731) );
  INV_X1 U9067 ( .A(n7072), .ZN(n11841) );
  NOR2_X1 U9068 ( .A1(n11654), .A2(n13843), .ZN(n7072) );
  INV_X1 U9069 ( .A(n7211), .ZN(n11680) );
  AND3_X1 U9070 ( .A1(n7212), .A2(n7213), .A3(n6915), .ZN(n7211) );
  INV_X1 U9071 ( .A(n7326), .ZN(n7325) );
  AND2_X1 U9072 ( .A1(n11818), .A2(n11817), .ZN(n6732) );
  INV_X1 U9073 ( .A(n14741), .ZN(n14329) );
  INV_X1 U9074 ( .A(n11036), .ZN(n7070) );
  NAND2_X1 U9075 ( .A1(n9934), .A2(n9922), .ZN(n13350) );
  INV_X1 U9076 ( .A(n15003), .ZN(n7207) );
  INV_X1 U9077 ( .A(n14983), .ZN(n7208) );
  INV_X1 U9078 ( .A(n14745), .ZN(n7069) );
  AND2_X1 U9079 ( .A1(n6593), .A2(n10558), .ZN(n6733) );
  NAND2_X1 U9080 ( .A1(n11096), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6734) );
  AND2_X1 U9081 ( .A1(n7399), .A2(n7397), .ZN(n6735) );
  NAND2_X1 U9082 ( .A1(n10916), .A2(n10915), .ZN(n6736) );
  INV_X1 U9083 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7112) );
  INV_X1 U9084 ( .A(n9941), .ZN(n6956) );
  INV_X1 U9085 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7050) );
  AND2_X1 U9086 ( .A1(n7256), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6737) );
  INV_X1 U9087 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7023) );
  INV_X1 U9088 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6745) );
  INV_X1 U9089 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7057) );
  XNOR2_X1 U9090 ( .A(n6908), .B(n12758), .ZN(n12736) );
  XNOR2_X2 U9091 ( .A(n14548), .B(n14547), .ZN(n14546) );
  NAND2_X1 U9092 ( .A1(n15514), .A2(n15513), .ZN(n6788) );
  AOI21_X1 U9093 ( .B1(n14638), .B2(n14639), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n6890) );
  INV_X1 U9094 ( .A(n14630), .ZN(n6755) );
  OAI21_X1 U9095 ( .B1(n14543), .B2(n14544), .A(P2_ADDR_REG_17__SCAN_IN), .ZN(
        n6740) );
  INV_X1 U9096 ( .A(n14642), .ZN(n6739) );
  NAND2_X2 U9097 ( .A1(n14542), .A2(n6740), .ZN(n14548) );
  OAI21_X1 U9098 ( .B1(n13200), .B2(n13199), .A(n13270), .ZN(n13204) );
  NOR2_X1 U9099 ( .A1(n13309), .A2(n6769), .ZN(n13272) );
  NAND2_X1 U9100 ( .A1(n13225), .A2(n13226), .ZN(n6744) );
  NAND3_X1 U9101 ( .A1(n6744), .A2(n13267), .A3(n14574), .ZN(n6762) );
  NAND2_X1 U9102 ( .A1(n7485), .A2(n6684), .ZN(n13279) );
  NAND2_X1 U9103 ( .A1(n10655), .A2(n6690), .ZN(n10708) );
  OAI21_X1 U9104 ( .B1(n11184), .B2(n7504), .A(n7503), .ZN(n11422) );
  NAND2_X1 U9105 ( .A1(n6887), .A2(n14842), .ZN(n6886) );
  NAND2_X1 U9106 ( .A1(n14507), .A2(n14506), .ZN(n6746) );
  NAND2_X1 U9107 ( .A1(n9666), .A2(n11644), .ZN(n9670) );
  AND2_X4 U9108 ( .A1(n7795), .A2(n7632), .ZN(n7964) );
  OAI22_X1 U9109 ( .A1(n9825), .A2(n7425), .B1(n9826), .B2(n7426), .ZN(n9832)
         );
  INV_X1 U9110 ( .A(n7332), .ZN(n7331) );
  NAND2_X1 U9111 ( .A1(n8014), .A2(n8565), .ZN(n8567) );
  OR2_X1 U9112 ( .A1(n9903), .A2(n10584), .ZN(n8298) );
  INV_X2 U9113 ( .A(n10463), .ZN(n14716) );
  NAND2_X1 U9114 ( .A1(n14071), .A2(n7045), .ZN(n7044) );
  NAND2_X4 U9115 ( .A1(n8016), .A2(n9945), .ZN(n8064) );
  NOR2_X4 U9116 ( .A1(n10613), .A2(n10929), .ZN(n10558) );
  INV_X1 U9117 ( .A(n7043), .ZN(n6953) );
  NAND2_X1 U9118 ( .A1(n7615), .A2(n7614), .ZN(n8038) );
  NAND4_X1 U9119 ( .A1(n6594), .A2(n8977), .A3(n6749), .A4(n9019), .ZN(n9030)
         );
  OR2_X1 U9120 ( .A1(n9032), .A2(n9031), .ZN(n9033) );
  NAND2_X1 U9121 ( .A1(n13619), .A2(n6683), .ZN(n13698) );
  NAND2_X1 U9122 ( .A1(n8040), .A2(n7618), .ZN(n8050) );
  NAND2_X1 U9123 ( .A1(n13445), .A2(n13446), .ZN(n13444) );
  NAND2_X1 U9124 ( .A1(n7467), .A2(n13478), .ZN(n7011) );
  NAND2_X1 U9125 ( .A1(n10233), .A2(n10232), .ZN(n6795) );
  XNOR2_X2 U9126 ( .A(n10343), .B(n13381), .ZN(n10232) );
  BUF_X4 U9127 ( .A(n8273), .Z(n8960) );
  NAND2_X1 U9128 ( .A1(n7328), .A2(n7329), .ZN(n7849) );
  NAND2_X1 U9129 ( .A1(n7896), .A2(n7593), .ZN(n7914) );
  NAND2_X1 U9130 ( .A1(n7026), .A2(SI_20_), .ZN(n7997) );
  NAND2_X1 U9131 ( .A1(n7311), .A2(n7677), .ZN(n7310) );
  AND2_X1 U9132 ( .A1(n9783), .A2(n6801), .ZN(n6800) );
  NAND2_X1 U9133 ( .A1(n10875), .A2(n10881), .ZN(n11184) );
  NAND2_X1 U9134 ( .A1(n14452), .A2(n14451), .ZN(n7053) );
  NAND2_X1 U9135 ( .A1(n10708), .A2(n10707), .ZN(n10713) );
  XNOR2_X1 U9136 ( .A(n14471), .B(n7057), .ZN(n14524) );
  OAI21_X1 U9137 ( .B1(n7510), .B2(n13191), .A(n7506), .ZN(n13302) );
  NAND2_X1 U9138 ( .A1(n9741), .A2(n9740), .ZN(n9748) );
  NAND2_X1 U9139 ( .A1(n7494), .A2(n7491), .ZN(n12036) );
  INV_X1 U9140 ( .A(n13195), .ZN(n7511) );
  NAND2_X1 U9141 ( .A1(n8234), .A2(n8233), .ZN(n8659) );
  NAND2_X1 U9142 ( .A1(n13591), .A2(n13603), .ZN(n6756) );
  OAI21_X2 U9143 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9698) );
  NAND2_X1 U9144 ( .A1(n8707), .A2(n8230), .ZN(n8717) );
  AOI22_X1 U9145 ( .A1(n9841), .A2(n9840), .B1(n9839), .B2(n9838), .ZN(n9846)
         );
  NAND2_X1 U9146 ( .A1(n9846), .A2(n6763), .ZN(n9890) );
  NOR2_X1 U9147 ( .A1(n9846), .A2(n6804), .ZN(n6803) );
  NAND2_X1 U9148 ( .A1(n7427), .A2(n7428), .ZN(n9818) );
  NAND2_X1 U9149 ( .A1(n9795), .A2(n9794), .ZN(n9798) );
  INV_X1 U9150 ( .A(n14179), .ZN(n7121) );
  INV_X1 U9151 ( .A(n7980), .ZN(n7026) );
  NAND2_X1 U9152 ( .A1(n7794), .A2(n7574), .ZN(n7808) );
  NAND2_X1 U9153 ( .A1(n7981), .A2(n7997), .ZN(n7983) );
  NAND2_X1 U9154 ( .A1(n7712), .A2(n7551), .ZN(n7724) );
  NAND2_X1 U9155 ( .A1(n7766), .A2(n7567), .ZN(n7778) );
  OAI21_X1 U9156 ( .B1(n8761), .B2(n8760), .A(n8759), .ZN(n8763) );
  AOI21_X1 U9157 ( .B1(n8768), .B2(n8767), .A(n8766), .ZN(n8770) );
  NAND2_X1 U9158 ( .A1(n7354), .A2(n7350), .ZN(n8911) );
  NAND2_X1 U9159 ( .A1(n6782), .A2(n6781), .ZN(n8782) );
  OAI21_X1 U9160 ( .B1(n8837), .B2(n7383), .A(n7382), .ZN(n8842) );
  NAND2_X1 U9161 ( .A1(n8812), .A2(n8811), .ZN(n8818) );
  OAI22_X1 U9162 ( .A1(n8825), .A2(n7385), .B1(n8826), .B2(n7384), .ZN(n8832)
         );
  OAI22_X1 U9163 ( .A1(n8847), .A2(n7393), .B1(n8846), .B2(n8845), .ZN(n8855)
         );
  OAI21_X1 U9164 ( .B1(n8990), .B2(n8989), .A(n7542), .ZN(n8995) );
  OAI211_X1 U9165 ( .C1(n7366), .C2(n8870), .A(n8872), .B(n7378), .ZN(n7377)
         );
  NAND2_X1 U9166 ( .A1(n9818), .A2(n9819), .ZN(n9817) );
  NAND2_X1 U9167 ( .A1(n6762), .A2(n6761), .ZN(P2_U3186) );
  NAND3_X1 U9168 ( .A1(n9712), .A2(n9711), .A3(n6694), .ZN(n7437) );
  NAND2_X1 U9169 ( .A1(n6764), .A2(n9779), .ZN(n9780) );
  OAI21_X1 U9170 ( .B1(n9776), .B2(n9775), .A(n6765), .ZN(n6764) );
  OR2_X1 U9171 ( .A1(n9778), .A2(n9777), .ZN(n6765) );
  NAND2_X1 U9172 ( .A1(n6768), .A2(n6767), .ZN(n6766) );
  NAND2_X1 U9173 ( .A1(n9767), .A2(n9766), .ZN(n6768) );
  NAND2_X1 U9174 ( .A1(n7349), .A2(n6702), .ZN(n8910) );
  NOR2_X1 U9175 ( .A1(n8918), .A2(n8917), .ZN(n8990) );
  NAND3_X1 U9176 ( .A1(n6982), .A2(n6981), .A3(n11032), .ZN(n11039) );
  INV_X4 U9177 ( .A(n10375), .ZN(n12422) );
  INV_X1 U9178 ( .A(n11848), .ZN(n11850) );
  NOR2_X1 U9179 ( .A1(n10401), .A2(n9685), .ZN(n10260) );
  INV_X1 U9180 ( .A(n11851), .ZN(n7296) );
  NAND2_X1 U9181 ( .A1(n7168), .A2(n7166), .ZN(n11374) );
  AOI21_X2 U9182 ( .B1(n12859), .B2(n12860), .A(n12196), .ZN(n12843) );
  OAI21_X2 U9183 ( .B1(n12876), .B2(n9440), .A(n12187), .ZN(n12859) );
  INV_X1 U9184 ( .A(n7420), .ZN(n7419) );
  NAND2_X1 U9185 ( .A1(n12071), .A2(n12224), .ZN(n7180) );
  NOR2_X1 U9186 ( .A1(n7418), .A2(n7190), .ZN(n7191) );
  AND3_X2 U9187 ( .A1(n8229), .A2(n8252), .A3(n8228), .ZN(n8707) );
  NAND2_X1 U9188 ( .A1(n11811), .A2(n11810), .ZN(n13684) );
  NAND2_X1 U9189 ( .A1(n6926), .A2(n15037), .ZN(n6924) );
  INV_X1 U9190 ( .A(n6786), .ZN(n6923) );
  INV_X1 U9191 ( .A(n7451), .ZN(n7450) );
  NAND2_X1 U9192 ( .A1(n7449), .A2(n7448), .ZN(n10539) );
  NAND2_X1 U9193 ( .A1(n14267), .A2(n7531), .ZN(n14268) );
  OAI21_X1 U9194 ( .B1(n7334), .B2(n7333), .A(n7835), .ZN(n7332) );
  INV_X1 U9195 ( .A(n7577), .ZN(n7335) );
  NAND2_X1 U9196 ( .A1(n7027), .A2(n7029), .ZN(n7586) );
  XNOR2_X1 U9197 ( .A(n8090), .B(n6802), .ZN(n14060) );
  INV_X1 U9198 ( .A(n7128), .ZN(n7126) );
  INV_X1 U9199 ( .A(n6611), .ZN(n6978) );
  NAND2_X1 U9200 ( .A1(n7310), .A2(n7548), .ZN(n7709) );
  NAND2_X1 U9201 ( .A1(n9429), .A2(n9428), .ZN(n9442) );
  NAND2_X1 U9202 ( .A1(n9314), .A2(n9313), .ZN(n9316) );
  NAND2_X1 U9203 ( .A1(n9271), .A2(n9270), .ZN(n9279) );
  NAND2_X1 U9204 ( .A1(n7077), .A2(n9403), .ZN(n9415) );
  NAND2_X1 U9205 ( .A1(n7076), .A2(n9416), .ZN(n9427) );
  NAND2_X1 U9206 ( .A1(n9293), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9296) );
  OAI21_X1 U9207 ( .B1(n9468), .B2(n11795), .A(n9469), .ZN(n9481) );
  INV_X1 U9208 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9069) );
  NAND4_X1 U9209 ( .A1(n7040), .A2(n7041), .A3(n7042), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7039) );
  NAND3_X1 U9210 ( .A1(n6771), .A2(n6973), .A3(n8205), .ZN(n8210) );
  NAND2_X1 U9211 ( .A1(n14084), .A2(n14741), .ZN(n6771) );
  NAND2_X1 U9212 ( .A1(n7724), .A2(n7723), .ZN(n7726) );
  AOI21_X1 U9213 ( .B1(n7122), .B2(n7121), .A(n6607), .ZN(n7120) );
  NAND2_X1 U9214 ( .A1(n7034), .A2(n7032), .ZN(n7028) );
  NAND2_X1 U9215 ( .A1(n14363), .A2(n14759), .ZN(n14267) );
  NAND2_X1 U9216 ( .A1(n6941), .A2(n6939), .ZN(n14088) );
  NAND2_X1 U9217 ( .A1(n11477), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11546) );
  NAND4_X1 U9218 ( .A1(n9882), .A2(n9881), .A3(n9880), .A4(n9883), .ZN(n9884)
         );
  NAND2_X1 U9219 ( .A1(n7623), .A2(n7622), .ZN(n8060) );
  NAND2_X1 U9220 ( .A1(n8040), .A2(n7018), .ZN(n7014) );
  NAND2_X1 U9221 ( .A1(n9784), .A2(n6800), .ZN(n6799) );
  NAND2_X1 U9222 ( .A1(n6808), .A2(n7446), .ZN(n9808) );
  OAI21_X1 U9223 ( .B1(n9893), .B2(n6803), .A(n9892), .ZN(n6807) );
  NAND2_X1 U9224 ( .A1(n9808), .A2(n9809), .ZN(n9807) );
  NAND3_X1 U9225 ( .A1(n6776), .A2(n6775), .A3(n6692), .ZN(n7440) );
  NAND2_X1 U9226 ( .A1(n9730), .A2(n9729), .ZN(n6775) );
  NAND2_X1 U9227 ( .A1(n9726), .A2(n9725), .ZN(n6776) );
  NAND3_X1 U9228 ( .A1(n6778), .A2(n6777), .A3(n6693), .ZN(n7443) );
  NAND2_X1 U9229 ( .A1(n9721), .A2(n9720), .ZN(n6777) );
  NAND2_X1 U9230 ( .A1(n9717), .A2(n9716), .ZN(n6778) );
  NAND2_X1 U9231 ( .A1(n9682), .A2(n10460), .ZN(n9661) );
  OR2_X1 U9232 ( .A1(n8842), .A2(n8841), .ZN(n6783) );
  OR2_X1 U9233 ( .A1(n8770), .A2(n8769), .ZN(n8775) );
  INV_X1 U9234 ( .A(n8781), .ZN(n6782) );
  AOI21_X1 U9235 ( .B1(n8865), .B2(n7369), .A(n7367), .ZN(n7366) );
  NAND3_X1 U9236 ( .A1(n9044), .A2(n9043), .A3(n6779), .ZN(P2_U3328) );
  OAI21_X2 U9237 ( .B1(n8320), .B2(n7135), .A(n7134), .ZN(n10593) );
  NAND2_X1 U9238 ( .A1(n10847), .A2(n10846), .ZN(n10845) );
  OAI21_X1 U9239 ( .B1(n11676), .B2(n8488), .A(n8489), .ZN(n11797) );
  NAND2_X1 U9240 ( .A1(n13544), .A2(n8999), .ZN(n8564) );
  NAND3_X1 U9242 ( .A1(n8756), .A2(n6780), .A3(n6680), .ZN(n8761) );
  OAI21_X1 U9243 ( .B1(n6595), .B2(n8840), .A(n6783), .ZN(n8847) );
  NAND2_X1 U9244 ( .A1(n6648), .A2(n6784), .ZN(n8837) );
  INV_X1 U9245 ( .A(n6785), .ZN(n6784) );
  AOI21_X1 U9246 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n6785) );
  NAND2_X1 U9247 ( .A1(n11402), .A2(n8460), .ZN(n11580) );
  NAND2_X1 U9248 ( .A1(n8416), .A2(n8415), .ZN(n14932) );
  NAND2_X1 U9249 ( .A1(n6795), .A2(n8310), .ZN(n10307) );
  INV_X1 U9250 ( .A(n10733), .ZN(n7136) );
  OAI21_X1 U9251 ( .B1(n8865), .B2(n7372), .A(n6790), .ZN(n8872) );
  NAND2_X1 U9252 ( .A1(n7493), .A2(n7492), .ZN(n7491) );
  NAND2_X1 U9253 ( .A1(n7034), .A2(n7583), .ZN(n7861) );
  NAND2_X1 U9254 ( .A1(n7709), .A2(n7550), .ZN(n7712) );
  NAND2_X1 U9255 ( .A1(n7746), .A2(n7747), .ZN(n7749) );
  NAND2_X1 U9256 ( .A1(n14449), .A2(n14423), .ZN(n7060) );
  NAND2_X1 U9257 ( .A1(n14524), .A2(n14523), .ZN(n6893) );
  NAND2_X1 U9258 ( .A1(n14460), .A2(n14461), .ZN(n6891) );
  NAND2_X1 U9259 ( .A1(n14630), .A2(n14631), .ZN(n6887) );
  NAND2_X1 U9260 ( .A1(n14453), .A2(n14454), .ZN(n14419) );
  AOI21_X1 U9261 ( .B1(n8911), .B2(n8910), .A(n8909), .ZN(n8918) );
  OAI21_X1 U9262 ( .B1(n8775), .B2(n8774), .A(n6792), .ZN(n8781) );
  NAND2_X1 U9263 ( .A1(n6794), .A2(n6793), .ZN(n6792) );
  NAND2_X1 U9264 ( .A1(n8775), .A2(n8774), .ZN(n6794) );
  NAND2_X1 U9265 ( .A1(n6798), .A2(n6796), .ZN(P2_U3236) );
  NAND2_X1 U9266 ( .A1(n13431), .A2(n13512), .ZN(n6798) );
  NAND2_X1 U9267 ( .A1(n7136), .A2(n10728), .ZN(n10735) );
  NAND2_X1 U9268 ( .A1(n7152), .A2(n7150), .ZN(n8597) );
  NAND2_X1 U9269 ( .A1(n7749), .A2(n7564), .ZN(n7764) );
  NAND2_X1 U9270 ( .A1(n7894), .A2(n7893), .ZN(n7896) );
  NAND2_X1 U9271 ( .A1(n7598), .A2(n6592), .ZN(n7008) );
  NAND2_X1 U9272 ( .A1(n7588), .A2(n7341), .ZN(n7894) );
  INV_X1 U9273 ( .A(n7546), .ZN(n7021) );
  NAND2_X1 U9274 ( .A1(n6807), .A2(n9896), .ZN(P1_U3242) );
  NAND3_X1 U9275 ( .A1(n9803), .A2(n9802), .A3(n6697), .ZN(n6808) );
  NAND2_X1 U9276 ( .A1(n6810), .A2(n6811), .ZN(n12616) );
  NAND3_X1 U9277 ( .A1(n6589), .A2(n7422), .A3(n6812), .ZN(n6810) );
  NAND2_X1 U9278 ( .A1(n12501), .A2(n6823), .ZN(n6820) );
  NAND2_X1 U9279 ( .A1(n12501), .A2(n6831), .ZN(n6828) );
  NAND2_X1 U9280 ( .A1(n9317), .A2(n6699), .ZN(n6833) );
  NAND2_X1 U9281 ( .A1(n9317), .A2(n6838), .ZN(n9552) );
  AND2_X2 U9282 ( .A1(n9128), .A2(n6614), .ZN(n9218) );
  NAND2_X1 U9283 ( .A1(n9622), .A2(n6844), .ZN(n6842) );
  NAND2_X1 U9284 ( .A1(n6842), .A2(n6843), .ZN(n12899) );
  INV_X1 U9285 ( .A(n13066), .ZN(n6854) );
  NAND3_X1 U9286 ( .A1(n6855), .A2(n11496), .A3(n6629), .ZN(n12110) );
  NAND3_X1 U9287 ( .A1(n9074), .A2(n6864), .A3(n6863), .ZN(n6862) );
  NAND2_X1 U9288 ( .A1(n6867), .A2(n6865), .ZN(n6868) );
  NAND2_X1 U9289 ( .A1(n6873), .A2(n6877), .ZN(n12749) );
  OAI21_X1 U9290 ( .B1(n11201), .B2(n6880), .A(n6879), .ZN(n15101) );
  INV_X1 U9291 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U9292 ( .A1(n14642), .A2(n14643), .ZN(n14494) );
  NAND2_X2 U9293 ( .A1(n6891), .A2(n14421), .ZN(n14422) );
  XNOR2_X2 U9294 ( .A(n14482), .B(n6894), .ZN(n14530) );
  AND2_X2 U9295 ( .A1(n6895), .A2(n6678), .ZN(n14482) );
  NAND2_X1 U9296 ( .A1(n15060), .A2(n6703), .ZN(n6899) );
  NAND2_X1 U9297 ( .A1(n6899), .A2(n6687), .ZN(n15069) );
  AND3_X2 U9298 ( .A1(n10681), .A2(n6912), .A3(n9045), .ZN(n9128) );
  NOR2_X2 U9299 ( .A1(n13595), .A2(n13674), .ZN(n7206) );
  NAND2_X1 U9300 ( .A1(n13472), .A2(n6922), .ZN(n13447) );
  OR2_X1 U9301 ( .A1(n13472), .A2(n6921), .ZN(n6920) );
  INV_X1 U9302 ( .A(n7146), .ZN(n13436) );
  NAND2_X1 U9303 ( .A1(n7020), .A2(n15037), .ZN(n6925) );
  NOR2_X1 U9304 ( .A1(n7020), .A2(n6926), .ZN(n7144) );
  NAND2_X1 U9305 ( .A1(n6925), .A2(n6923), .ZN(P2_U3528) );
  INV_X2 U9306 ( .A(n7552), .ZN(n9945) );
  NAND4_X1 U9307 ( .A1(n13705), .A2(n13547), .A3(n6929), .A4(n13487), .ZN(
        n13484) );
  INV_X1 U9308 ( .A(n6930), .ZN(n13521) );
  OAI21_X1 U9309 ( .B1(n8114), .B2(n11630), .A(n6931), .ZN(n11831) );
  NAND2_X1 U9310 ( .A1(n11831), .A2(n11840), .ZN(n8116) );
  INV_X1 U9311 ( .A(n7731), .ZN(n6935) );
  INV_X1 U9312 ( .A(n6937), .ZN(n7276) );
  NAND2_X1 U9313 ( .A1(n6938), .A2(n11434), .ZN(n6937) );
  NAND2_X1 U9314 ( .A1(n11289), .A2(n8112), .ZN(n6938) );
  NAND2_X1 U9315 ( .A1(n14144), .A2(n6944), .ZN(n6941) );
  NAND2_X1 U9316 ( .A1(n14073), .A2(n6952), .ZN(n6950) );
  NAND2_X1 U9317 ( .A1(n6950), .A2(n6951), .ZN(P1_U3525) );
  AOI21_X1 U9318 ( .B1(n14073), .B2(n14741), .A(n6953), .ZN(n8199) );
  MUX2_X1 U9319 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7552), .Z(n7553) );
  INV_X1 U9320 ( .A(n8064), .ZN(n9675) );
  XNOR2_X2 U9321 ( .A(n13914), .B(n10892), .ZN(n10608) );
  NAND3_X1 U9322 ( .A1(n7964), .A2(n7640), .A3(n8166), .ZN(n7280) );
  AND3_X2 U9323 ( .A1(n7540), .A2(n7639), .A3(n8154), .ZN(n7640) );
  AND4_X2 U9324 ( .A1(n7634), .A2(n7633), .A3(n7635), .A4(n7898), .ZN(n7540)
         );
  NAND2_X1 U9325 ( .A1(n7979), .A2(n6957), .ZN(n14205) );
  NAND2_X1 U9326 ( .A1(n11970), .A2(n6962), .ZN(n6961) );
  NAND2_X1 U9327 ( .A1(n6966), .A2(n6968), .ZN(n11439) );
  NAND2_X1 U9328 ( .A1(n11337), .A2(n6967), .ZN(n6966) );
  NAND2_X1 U9329 ( .A1(n10512), .A2(n7124), .ZN(n6971) );
  INV_X1 U9330 ( .A(n9861), .ZN(n6972) );
  NAND3_X1 U9331 ( .A1(n6975), .A2(n6974), .A3(n14626), .ZN(n6973) );
  NAND2_X1 U9332 ( .A1(n14098), .A2(n7130), .ZN(n6974) );
  NAND2_X1 U9333 ( .A1(n6976), .A2(n8203), .ZN(n6975) );
  XNOR2_X2 U9334 ( .A(n7647), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9335 ( .A1(n7296), .A2(n11984), .ZN(n7299) );
  NAND2_X1 U9336 ( .A1(n10926), .A2(n6605), .ZN(n6981) );
  XNOR2_X2 U9337 ( .A(n10908), .B(n10904), .ZN(n10926) );
  NOR2_X1 U9338 ( .A1(n6983), .A2(n10909), .ZN(n11033) );
  NOR2_X2 U9339 ( .A1(n12443), .A2(n10903), .ZN(n10908) );
  NAND2_X1 U9340 ( .A1(n13784), .A2(n6987), .ZN(n6984) );
  NAND2_X1 U9341 ( .A1(n6984), .A2(n6985), .ZN(n12454) );
  NAND2_X1 U9342 ( .A1(n12338), .A2(n6993), .ZN(n6990) );
  NAND2_X1 U9343 ( .A1(n6990), .A2(n6991), .ZN(n13806) );
  NAND2_X1 U9344 ( .A1(n13847), .A2(n6998), .ZN(n6996) );
  NAND2_X1 U9345 ( .A1(n6996), .A2(n6997), .ZN(n13818) );
  INV_X1 U9346 ( .A(n7005), .ZN(n7003) );
  NOR2_X1 U9347 ( .A1(n7005), .A2(n8155), .ZN(n7004) );
  NAND2_X1 U9348 ( .A1(n7964), .A2(n7540), .ZN(n7966) );
  NAND2_X1 U9349 ( .A1(n7980), .A2(n7603), .ZN(n7608) );
  NAND2_X1 U9350 ( .A1(n7008), .A2(n7336), .ZN(n7007) );
  NAND2_X1 U9351 ( .A1(n7464), .A2(n13446), .ZN(n7010) );
  NAND3_X1 U9352 ( .A1(n7010), .A2(n7009), .A3(n8704), .ZN(n8705) );
  NAND2_X1 U9353 ( .A1(n7012), .A2(n7011), .ZN(n13445) );
  INV_X1 U9354 ( .A(n7464), .ZN(n7012) );
  NAND2_X1 U9355 ( .A1(n8038), .A2(n8037), .ZN(n8040) );
  OAI21_X1 U9356 ( .B1(n7552), .B2(n7023), .A(n7022), .ZN(n7546) );
  NAND2_X1 U9357 ( .A1(n7552), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U9358 ( .A1(n7849), .A2(n6596), .ZN(n7027) );
  NAND2_X2 U9359 ( .A1(n7036), .A2(n7035), .ZN(n14144) );
  NAND4_X1 U9360 ( .A1(n7545), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n7038), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7037) );
  INV_X2 U9361 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7545) );
  NAND2_X4 U9362 ( .A1(n8016), .A2(n7047), .ZN(n9677) );
  MUX2_X1 U9363 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n9945), .Z(n7565) );
  MUX2_X1 U9364 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7046), .Z(n7575) );
  MUX2_X1 U9365 ( .A(n15492), .B(n10941), .S(n7046), .Z(n7594) );
  MUX2_X1 U9366 ( .A(n10842), .B(n10844), .S(n7046), .Z(n7590) );
  MUX2_X1 U9367 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7046), .Z(n7600) );
  MUX2_X1 U9368 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7046), .Z(n7946) );
  MUX2_X1 U9369 ( .A(n11081), .B(n15367), .S(n7046), .Z(n7932) );
  MUX2_X1 U9370 ( .A(n11529), .B(n11531), .S(n7046), .Z(n7982) );
  MUX2_X1 U9371 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7046), .Z(n7616) );
  MUX2_X1 U9372 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7046), .Z(n7628) );
  MUX2_X1 U9373 ( .A(n13740), .B(n14411), .S(n7046), .Z(n8061) );
  MUX2_X1 U9374 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7046), .Z(n8942) );
  INV_X2 U9375 ( .A(n9945), .ZN(n7047) );
  OAI21_X4 U9376 ( .B1(n11530), .B2(n8064), .A(n7985), .ZN(n14315) );
  NAND2_X1 U9377 ( .A1(n14494), .A2(n14869), .ZN(n7056) );
  XNOR2_X1 U9378 ( .A(n14478), .B(n14479), .ZN(n14529) );
  NAND2_X1 U9379 ( .A1(n15518), .A2(n15519), .ZN(n7058) );
  NAND3_X1 U9380 ( .A1(n7964), .A2(n7640), .A3(n7434), .ZN(n7062) );
  AND2_X2 U9381 ( .A1(n14113), .A2(n7063), .ZN(n14054) );
  NOR2_X2 U9382 ( .A1(n6612), .A2(n14384), .ZN(n14195) );
  NAND3_X1 U9383 ( .A1(n6593), .A2(n10558), .A3(n11249), .ZN(n11055) );
  NAND4_X1 U9384 ( .A1(n6593), .A2(n10558), .A3(n11249), .A4(n7069), .ZN(
        n11346) );
  NOR2_X2 U9385 ( .A1(n11440), .A2(n11525), .ZN(n11655) );
  NAND2_X1 U9386 ( .A1(n9093), .A2(n7073), .ZN(n9095) );
  XNOR2_X1 U9387 ( .A(n9092), .B(n7073), .ZN(n9962) );
  NAND2_X1 U9388 ( .A1(n9496), .A2(n9495), .ZN(n7074) );
  NAND2_X1 U9389 ( .A1(n9481), .A2(n9480), .ZN(n7075) );
  NAND2_X1 U9390 ( .A1(n9415), .A2(n9414), .ZN(n7076) );
  NAND2_X1 U9391 ( .A1(n9402), .A2(n9401), .ZN(n7077) );
  INV_X1 U9392 ( .A(n9444), .ZN(n7078) );
  NAND2_X1 U9393 ( .A1(n7078), .A2(n9453), .ZN(n7081) );
  NAND2_X1 U9394 ( .A1(n7081), .A2(n7082), .ZN(n9455) );
  NAND2_X1 U9395 ( .A1(n9332), .A2(n7087), .ZN(n7084) );
  NAND2_X1 U9396 ( .A1(n7084), .A2(n7085), .ZN(n9363) );
  NAND2_X1 U9397 ( .A1(n9105), .A2(n7096), .ZN(n7095) );
  OAI21_X1 U9398 ( .B1(n9168), .B2(n7104), .A(n7101), .ZN(n9207) );
  NAND2_X1 U9399 ( .A1(n7113), .A2(n6688), .ZN(n7979) );
  NAND2_X1 U9400 ( .A1(n11839), .A2(n7116), .ZN(n7114) );
  INV_X1 U9401 ( .A(n14100), .ZN(n7127) );
  AOI21_X1 U9402 ( .B1(n7130), .B2(n7129), .A(n6695), .ZN(n7128) );
  INV_X1 U9403 ( .A(n14099), .ZN(n7129) );
  INV_X1 U9404 ( .A(n8319), .ZN(n7133) );
  NAND2_X1 U9405 ( .A1(n10593), .A2(n10596), .ZN(n8345) );
  NAND2_X1 U9406 ( .A1(n13490), .A2(n7139), .ZN(n7137) );
  OR2_X2 U9407 ( .A1(n8663), .A2(n13530), .ZN(n7145) );
  NAND2_X1 U9408 ( .A1(n7145), .A2(n8662), .ZN(n13431) );
  NAND2_X1 U9409 ( .A1(n13528), .A2(n6590), .ZN(n7152) );
  OR2_X2 U9410 ( .A1(n11797), .A2(n11810), .ZN(n11798) );
  NAND2_X1 U9411 ( .A1(n13577), .A2(n6613), .ZN(n7154) );
  NAND2_X1 U9412 ( .A1(n7154), .A2(n7155), .ZN(n13544) );
  NAND2_X1 U9413 ( .A1(n8520), .A2(n8519), .ZN(n13591) );
  NAND2_X1 U9414 ( .A1(n8459), .A2(n8458), .ZN(n11402) );
  XNOR2_X1 U9415 ( .A(n8640), .B(n6594), .ZN(n8663) );
  NAND2_X2 U9416 ( .A1(n11798), .A2(n8504), .ZN(n11951) );
  NAND2_X1 U9417 ( .A1(n13442), .A2(n8631), .ZN(n8640) );
  AOI22_X1 U9418 ( .A1(n8530), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8529), .B2(
        n10106), .ZN(n8317) );
  NAND2_X1 U9419 ( .A1(n7730), .A2(n7729), .ZN(n10512) );
  NAND2_X1 U9420 ( .A1(n11437), .A2(n7847), .ZN(n11647) );
  NAND2_X1 U9421 ( .A1(n11047), .A2(n7790), .ZN(n10981) );
  OR2_X2 U9422 ( .A1(n9946), .A2(n8064), .ZN(n7715) );
  OR2_X2 U9423 ( .A1(n14181), .A2(n6770), .ZN(n14168) );
  NAND2_X1 U9424 ( .A1(n13025), .A2(n7159), .ZN(n12081) );
  NAND2_X1 U9425 ( .A1(n10814), .A2(n7159), .ZN(n10815) );
  XNOR2_X1 U9426 ( .A(n10813), .B(n7159), .ZN(n11019) );
  OAI22_X1 U9427 ( .A1(n12609), .A2(n11266), .B1(n12618), .B2(n7159), .ZN(
        n10799) );
  OAI22_X1 U9428 ( .A1(n12623), .A2(n15122), .B1(n12609), .B2(n7159), .ZN(
        n11023) );
  NAND2_X1 U9429 ( .A1(n12954), .A2(n7163), .ZN(n7162) );
  NAND3_X1 U9430 ( .A1(n11259), .A2(n12233), .A3(n12237), .ZN(n7168) );
  INV_X1 U9431 ( .A(n12100), .ZN(n7169) );
  NAND2_X1 U9432 ( .A1(n11261), .A2(n12100), .ZN(n11361) );
  NAND2_X1 U9433 ( .A1(n11259), .A2(n12237), .ZN(n11261) );
  NAND2_X1 U9434 ( .A1(n12841), .A2(n7173), .ZN(n7170) );
  NAND2_X1 U9435 ( .A1(n7170), .A2(n7171), .ZN(n12800) );
  AOI21_X2 U9436 ( .B1(n7180), .B2(n7179), .A(n7177), .ZN(n12072) );
  OAI21_X2 U9437 ( .B1(n12787), .B2(n12789), .A(n12221), .ZN(n12071) );
  NOR2_X2 U9438 ( .A1(n12798), .A2(n9509), .ZN(n12787) );
  INV_X1 U9439 ( .A(n7528), .ZN(n7189) );
  AND2_X1 U9440 ( .A1(n10230), .A2(n7193), .ZN(n10384) );
  AND2_X1 U9441 ( .A1(n7195), .A2(n14952), .ZN(n10230) );
  NAND3_X1 U9442 ( .A1(n7198), .A2(n7197), .A3(n7196), .ZN(n13426) );
  OAI21_X1 U9443 ( .B1(n7552), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7204), .ZN(
        n7547) );
  NAND2_X1 U9444 ( .A1(n7552), .A2(n9069), .ZN(n7204) );
  NAND3_X1 U9445 ( .A1(n7209), .A2(n15201), .A3(n7207), .ZN(n10852) );
  INV_X1 U9446 ( .A(n10807), .ZN(n15122) );
  OAI211_X2 U9447 ( .C1(n10662), .C2(n10979), .A(n7215), .B(n7214), .ZN(n10807) );
  OR2_X1 U9448 ( .A1(n9100), .A2(n9962), .ZN(n7214) );
  OR2_X1 U9449 ( .A1(n9138), .A2(n7312), .ZN(n7215) );
  NAND2_X1 U9450 ( .A1(n7223), .A2(n7222), .ZN(n11375) );
  AOI21_X1 U9451 ( .B1(n9608), .B2(n12237), .A(n6674), .ZN(n7222) );
  NAND2_X1 U9452 ( .A1(n11263), .A2(n9608), .ZN(n7223) );
  NAND2_X1 U9453 ( .A1(n12828), .A2(n7229), .ZN(n7228) );
  NAND2_X1 U9454 ( .A1(n12828), .A2(n7530), .ZN(n12812) );
  OAI21_X1 U9455 ( .B1(n9645), .B2(n13019), .A(n9644), .ZN(n13098) );
  OAI211_X1 U9456 ( .C1(n10753), .C2(n7253), .A(n7252), .B(n7250), .ZN(n11115)
         );
  INV_X1 U9457 ( .A(n11099), .ZN(n7257) );
  XNOR2_X2 U9458 ( .A(n7264), .B(n9045), .ZN(n10749) );
  OAI21_X1 U9459 ( .B1(n11052), .B2(n8110), .A(n8109), .ZN(n10984) );
  NAND2_X1 U9460 ( .A1(n9868), .A2(n7271), .ZN(n7270) );
  OAI21_X1 U9461 ( .B1(n11277), .B2(n6937), .A(n7274), .ZN(n11649) );
  NOR2_X4 U9462 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7686) );
  NAND3_X1 U9463 ( .A1(n8099), .A2(n7716), .A3(n10465), .ZN(n10464) );
  NAND2_X2 U9464 ( .A1(n7282), .A2(n7281), .ZN(n12338) );
  INV_X1 U9465 ( .A(n12327), .ZN(n7292) );
  INV_X1 U9466 ( .A(n11984), .ZN(n7302) );
  NAND2_X1 U9467 ( .A1(n11852), .A2(n11851), .ZN(n11985) );
  NAND2_X1 U9468 ( .A1(n11719), .A2(n11718), .ZN(n11852) );
  NAND2_X1 U9469 ( .A1(n13825), .A2(n6691), .ZN(n13774) );
  NAND2_X1 U9470 ( .A1(n8091), .A2(n7306), .ZN(n7538) );
  NAND2_X1 U9471 ( .A1(n8091), .A2(n8095), .ZN(n8093) );
  OR2_X1 U9472 ( .A1(n7310), .A2(n7309), .ZN(n7681) );
  NAND2_X1 U9473 ( .A1(n7668), .A2(n7314), .ZN(n7313) );
  NAND2_X1 U9474 ( .A1(n7668), .A2(n7630), .ZN(n7320) );
  OR2_X1 U9475 ( .A1(n7668), .A2(n7669), .ZN(n7324) );
  NAND2_X1 U9476 ( .A1(n7810), .A2(n7331), .ZN(n7328) );
  NAND2_X1 U9477 ( .A1(n7586), .A2(n7587), .ZN(n7341) );
  INV_X1 U9478 ( .A(n8061), .ZN(n7344) );
  NAND2_X1 U9479 ( .A1(n8900), .A2(n8899), .ZN(n7347) );
  NAND2_X1 U9480 ( .A1(n8902), .A2(n8901), .ZN(n7348) );
  NAND3_X1 U9481 ( .A1(n7348), .A2(n7347), .A3(n6696), .ZN(n7349) );
  NAND3_X1 U9482 ( .A1(n7348), .A2(n7347), .A3(n6677), .ZN(n7354) );
  INV_X1 U9483 ( .A(n8904), .ZN(n7356) );
  NAND2_X1 U9484 ( .A1(n8796), .A2(n8795), .ZN(n7359) );
  NAND2_X1 U9485 ( .A1(n8792), .A2(n8791), .ZN(n7360) );
  NAND2_X1 U9486 ( .A1(n7361), .A2(n7358), .ZN(n8807) );
  NAND3_X1 U9487 ( .A1(n7360), .A2(n7359), .A3(n7364), .ZN(n7358) );
  NAND3_X1 U9488 ( .A1(n7363), .A2(n7362), .A3(n7365), .ZN(n7361) );
  NAND2_X1 U9489 ( .A1(n8782), .A2(n6705), .ZN(n7373) );
  INV_X1 U9490 ( .A(n8787), .ZN(n7376) );
  NAND2_X1 U9491 ( .A1(n7377), .A2(n7380), .ZN(n8880) );
  NOR2_X1 U9492 ( .A1(n8880), .A2(n8879), .ZN(n8881) );
  NAND2_X1 U9493 ( .A1(n6675), .A2(n7381), .ZN(n7380) );
  NAND2_X1 U9494 ( .A1(n8855), .A2(n8856), .ZN(n8854) );
  NOR2_X2 U9495 ( .A1(n8722), .A2(n8217), .ZN(n8229) );
  NAND2_X1 U9496 ( .A1(n7396), .A2(n7399), .ZN(n11018) );
  INV_X1 U9497 ( .A(n10812), .ZN(n7394) );
  NAND2_X1 U9498 ( .A1(n10808), .A2(n13014), .ZN(n7399) );
  NAND2_X1 U9499 ( .A1(n11511), .A2(n11500), .ZN(n7400) );
  NAND2_X2 U9500 ( .A1(n12584), .A2(n12583), .ZN(n7422) );
  NAND2_X1 U9501 ( .A1(n9542), .A2(n7423), .ZN(n9550) );
  NAND2_X2 U9502 ( .A1(n7649), .A2(n7650), .ZN(n8149) );
  NAND3_X1 U9503 ( .A1(n7649), .A2(n7650), .A3(P1_REG1_REG_1__SCAN_IN), .ZN(
        n7673) );
  INV_X1 U9504 ( .A(n9832), .ZN(n9829) );
  NAND3_X1 U9505 ( .A1(n9813), .A2(n9812), .A3(n6698), .ZN(n7427) );
  INV_X1 U9506 ( .A(n9814), .ZN(n7429) );
  NAND2_X1 U9507 ( .A1(n9787), .A2(n9785), .ZN(n7430) );
  NAND2_X1 U9508 ( .A1(n7437), .A2(n7438), .ZN(n9718) );
  NAND2_X1 U9509 ( .A1(n7440), .A2(n7441), .ZN(n9736) );
  NAND2_X1 U9510 ( .A1(n7443), .A2(n7444), .ZN(n9727) );
  NAND2_X1 U9511 ( .A1(n10383), .A2(n7450), .ZN(n7449) );
  NAND2_X1 U9512 ( .A1(n7453), .A2(n6685), .ZN(n10731) );
  NAND2_X1 U9513 ( .A1(n14940), .A2(n7459), .ZN(n7455) );
  NAND2_X1 U9514 ( .A1(n7455), .A2(n7454), .ZN(n8683) );
  INV_X1 U9515 ( .A(n13478), .ZN(n7470) );
  OAI21_X1 U9516 ( .B1(n13466), .B2(n7465), .A(n6707), .ZN(n7464) );
  OAI21_X1 U9517 ( .B1(n13552), .B2(n7473), .A(n7471), .ZN(n13515) );
  OAI21_X1 U9518 ( .B1(n13552), .B2(n8696), .A(n8697), .ZN(n13533) );
  NAND4_X1 U9519 ( .A1(n8229), .A2(n8252), .A3(n8228), .A4(n7481), .ZN(n8238)
         );
  NAND2_X1 U9520 ( .A1(n13279), .A2(n13211), .ZN(n13216) );
  NAND2_X1 U9521 ( .A1(n13235), .A2(n13234), .ZN(n7485) );
  NAND2_X1 U9522 ( .A1(n13208), .A2(n13207), .ZN(n7486) );
  XNOR2_X2 U9523 ( .A(n13208), .B(n13206), .ZN(n13235) );
  XNOR2_X2 U9524 ( .A(n8650), .B(P2_IR_REG_20__SCAN_IN), .ZN(n9024) );
  XNOR2_X1 U9525 ( .A(n9035), .B(n6577), .ZN(n8706) );
  NAND2_X1 U9526 ( .A1(n13326), .A2(n13189), .ZN(n7508) );
  NAND3_X1 U9527 ( .A1(n7511), .A2(n13326), .A3(n13189), .ZN(n7510) );
  NAND2_X1 U9528 ( .A1(n7507), .A2(n13245), .ZN(n7512) );
  NOR2_X1 U9529 ( .A1(n13302), .A2(n13303), .ZN(n7513) );
  NAND2_X1 U9530 ( .A1(n13193), .A2(n13194), .ZN(n7509) );
  NAND2_X1 U9531 ( .A1(n13351), .A2(n6704), .ZN(n7514) );
  NAND2_X1 U9532 ( .A1(n13351), .A2(n6631), .ZN(n13267) );
  NAND2_X1 U9533 ( .A1(n13351), .A2(n13223), .ZN(n13225) );
  NAND2_X1 U9534 ( .A1(n7514), .A2(n13254), .ZN(n13258) );
  OAI21_X1 U9535 ( .B1(n9925), .B2(n9924), .A(n10349), .ZN(n7515) );
  NAND2_X1 U9536 ( .A1(n7515), .A2(n10424), .ZN(n10426) );
  NAND2_X1 U9537 ( .A1(n10350), .A2(n10349), .ZN(n10431) );
  NAND2_X1 U9538 ( .A1(n7517), .A2(n7516), .ZN(n10350) );
  NAND2_X1 U9539 ( .A1(n7520), .A2(n6630), .ZN(n7518) );
  NAND2_X1 U9540 ( .A1(n8527), .A2(n8252), .ZN(n8641) );
  OR2_X1 U9541 ( .A1(n9661), .A2(n9685), .ZN(n14723) );
  NAND2_X1 U9542 ( .A1(n9634), .A2(n6576), .ZN(n9636) );
  INV_X1 U9543 ( .A(n9653), .ZN(n9657) );
  NAND2_X1 U9544 ( .A1(n10607), .A2(n8100), .ZN(n10522) );
  OAI211_X2 U9545 ( .C1(n8016), .C2(n13944), .A(n7715), .B(n7714), .ZN(n10463)
         );
  NAND2_X1 U9546 ( .A1(n14091), .A2(n8137), .ZN(n8204) );
  CLKBUF_X1 U9547 ( .A(n10900), .Z(n12436) );
  INV_X1 U9548 ( .A(n8807), .ZN(n8810) );
  NAND2_X1 U9549 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  NAND4_X2 U9550 ( .A1(n7703), .A2(n7702), .A3(n7701), .A4(n7700), .ZN(n13915)
         );
  OAI22_X1 U9551 ( .A1(n10610), .A2(n10913), .B1(n14716), .B2(n12458), .ZN(
        n10374) );
  NAND4_X2 U9552 ( .A1(n9068), .A2(n9067), .A3(n9066), .A4(n9065), .ZN(n15110)
         );
  NAND2_X1 U9553 ( .A1(n8664), .A2(n10329), .ZN(n10188) );
  INV_X1 U9554 ( .A(n6757), .ZN(n8664) );
  NAND4_X2 U9555 ( .A1(n9085), .A2(n9084), .A3(n9083), .A4(n9082), .ZN(n9601)
         );
  NAND2_X1 U9556 ( .A1(n13600), .A2(n8691), .ZN(n13575) );
  XNOR2_X2 U9557 ( .A(n9079), .B(n9078), .ZN(n10979) );
  INV_X1 U9558 ( .A(n8246), .ZN(n12277) );
  AND2_X1 U9559 ( .A1(n9035), .A2(n11409), .ZN(n10409) );
  INV_X1 U9560 ( .A(n9064), .ZN(n12447) );
  CLKBUF_X1 U9561 ( .A(n9902), .Z(n14974) );
  NAND2_X1 U9562 ( .A1(n8299), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8268) );
  INV_X1 U9563 ( .A(n6579), .ZN(n8931) );
  NAND4_X4 U9564 ( .A1(n7676), .A2(n7675), .A3(n7674), .A4(n7673), .ZN(n13917)
         );
  NAND2_X1 U9565 ( .A1(n13204), .A2(n13203), .ZN(n13205) );
  INV_X1 U9566 ( .A(n11399), .ZN(n8458) );
  OR2_X1 U9567 ( .A1(n8818), .A2(n8817), .ZN(n7524) );
  OR2_X1 U9568 ( .A1(n6576), .A2(n9635), .ZN(n7525) );
  AND2_X1 U9569 ( .A1(n9317), .A2(n9051), .ZN(n7526) );
  CLKBUF_X3 U9570 ( .A(n9121), .Z(n12062) );
  OR3_X1 U9571 ( .A1(n10272), .A2(n14140), .A3(n14407), .ZN(n7527) );
  INV_X2 U9572 ( .A(n14757), .ZN(n14759) );
  AND2_X1 U9573 ( .A1(n13360), .A2(n13202), .ZN(n7529) );
  OR2_X1 U9574 ( .A1(n14759), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7531) );
  OR2_X1 U9575 ( .A1(n14752), .A2(n8198), .ZN(n7532) );
  NOR3_X1 U9576 ( .A1(n13694), .A2(n8969), .A3(n13421), .ZN(n7533) );
  AND3_X1 U9577 ( .A1(n13694), .A2(n8993), .A3(n13421), .ZN(n7534) );
  OR2_X1 U9578 ( .A1(n11712), .A2(n11711), .ZN(n7536) );
  AND2_X1 U9579 ( .A1(n8937), .A2(n9638), .ZN(n7537) );
  OR2_X1 U9580 ( .A1(n10019), .A2(n10026), .ZN(n13340) );
  NAND2_X1 U9581 ( .A1(n13512), .A2(n10414), .ZN(n14951) );
  INV_X1 U9582 ( .A(n14304), .ZN(n8207) );
  AND2_X2 U9583 ( .A1(n9590), .A2(n15123), .ZN(n15129) );
  AND2_X1 U9584 ( .A1(n14270), .A2(n14093), .ZN(n7539) );
  NAND2_X1 U9585 ( .A1(n14752), .A2(n14744), .ZN(n14381) );
  NOR2_X1 U9586 ( .A1(n7064), .A2(n14304), .ZN(n8193) );
  NAND2_X1 U9587 ( .A1(n9852), .A2(n9853), .ZN(n7541) );
  INV_X1 U9588 ( .A(n13360), .ZN(n13274) );
  AND2_X1 U9589 ( .A1(n9594), .A2(n9593), .ZN(n7543) );
  AND2_X1 U9590 ( .A1(n10413), .A2(n15200), .ZN(n10410) );
  INV_X1 U9591 ( .A(n13718), .ZN(n9638) );
  AND2_X2 U9592 ( .A1(n9637), .A2(n14962), .ZN(n15027) );
  INV_X1 U9593 ( .A(n13672), .ZN(n8743) );
  AND2_X2 U9594 ( .A1(n9637), .A2(n9920), .ZN(n15037) );
  OAI21_X1 U9595 ( .B1(n9835), .B2(n14716), .A(n10610), .ZN(n9697) );
  NAND2_X1 U9596 ( .A1(n10337), .A2(n8992), .ZN(n8757) );
  INV_X1 U9597 ( .A(n8808), .ZN(n8809) );
  AOI21_X1 U9598 ( .B1(n8818), .B2(n8817), .A(n8815), .ZN(n8816) );
  AND2_X1 U9599 ( .A1(n9760), .A2(n9759), .ZN(n9761) );
  NAND2_X1 U9600 ( .A1(n8819), .A2(n7524), .ZN(n8825) );
  INV_X1 U9601 ( .A(n8826), .ZN(n8827) );
  INV_X1 U9602 ( .A(n8856), .ZN(n8857) );
  NAND2_X1 U9603 ( .A1(n8860), .A2(n8859), .ZN(n8865) );
  INV_X1 U9604 ( .A(n8869), .ZN(n8870) );
  AND2_X1 U9605 ( .A1(n10804), .A2(n12229), .ZN(n10805) );
  INV_X1 U9606 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9053) );
  INV_X1 U9607 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7636) );
  AND2_X1 U9608 ( .A1(n14900), .A2(n11755), .ZN(n11757) );
  INV_X1 U9609 ( .A(n10810), .ZN(n10811) );
  INV_X1 U9610 ( .A(n9462), .ZN(n9461) );
  NOR2_X1 U9611 ( .A1(n12067), .A2(n12781), .ZN(n9643) );
  OR2_X1 U9612 ( .A1(n10010), .A2(n9572), .ZN(n10783) );
  AND2_X1 U9613 ( .A1(n8258), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8257) );
  AND3_X1 U9614 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(n8610), .ZN(n8243) );
  INV_X1 U9615 ( .A(n13603), .ZN(n8690) );
  AND2_X1 U9616 ( .A1(n10902), .A2(n10901), .ZN(n10903) );
  INV_X1 U9617 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7840) );
  INV_X1 U9618 ( .A(n14208), .ZN(n7994) );
  INV_X1 U9619 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7799) );
  INV_X1 U9620 ( .A(n14270), .ZN(n8142) );
  NAND2_X1 U9621 ( .A1(n11338), .A2(n8111), .ZN(n11277) );
  INV_X1 U9622 ( .A(n11512), .ZN(n11497) );
  INV_X1 U9623 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15488) );
  NOR2_X1 U9624 ( .A1(n9356), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U9625 ( .A1(n9461), .A2(n9460), .ZN(n9473) );
  NOR2_X1 U9626 ( .A1(n9287), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9302) );
  INV_X1 U9627 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n13099) );
  INV_X1 U9628 ( .A(n12928), .ZN(n9377) );
  OR2_X1 U9629 ( .A1(n10936), .A2(n12764), .ZN(n10779) );
  INV_X1 U9630 ( .A(n11015), .ZN(n13025) );
  OR2_X1 U9631 ( .A1(n10010), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U9632 ( .A1(n9427), .A2(n9426), .ZN(n9429) );
  NOR2_X1 U9633 ( .A1(n8588), .A2(n13295), .ZN(n8610) );
  INV_X1 U9634 ( .A(n13217), .ZN(n13255) );
  INV_X1 U9635 ( .A(n6585), .ZN(n9036) );
  AND2_X1 U9636 ( .A1(n8257), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8533) );
  OR2_X1 U9637 ( .A1(n8498), .A2(n8497), .ZN(n8510) );
  OR2_X1 U9638 ( .A1(n14819), .A2(n14818), .ZN(n14821) );
  OR2_X1 U9639 ( .A1(n14848), .A2(n14847), .ZN(n14849) );
  AND2_X1 U9640 ( .A1(n14873), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n14875) );
  AND2_X1 U9641 ( .A1(n8243), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8622) );
  OR2_X1 U9642 ( .A1(n8423), .A2(n15402), .ZN(n8449) );
  INV_X1 U9643 ( .A(n10907), .ZN(n10904) );
  INV_X1 U9644 ( .A(n8031), .ZN(n8043) );
  NAND2_X1 U9645 ( .A1(n7938), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7952) );
  OR2_X1 U9646 ( .A1(n7841), .A2(n7840), .ZN(n7852) );
  INV_X1 U9647 ( .A(n14113), .ZN(n14127) );
  OR2_X1 U9648 ( .A1(n7829), .A2(n7828), .ZN(n7841) );
  INV_X1 U9649 ( .A(n14054), .ZN(n8144) );
  NAND2_X1 U9650 ( .A1(n8567), .A2(n7611), .ZN(n8027) );
  NOR2_X1 U9651 ( .A1(n14481), .A2(n14480), .ZN(n14435) );
  INV_X1 U9652 ( .A(n12473), .ZN(n12313) );
  AND2_X1 U9653 ( .A1(n9194), .A2(n9193), .ZN(n9211) );
  INV_X1 U9654 ( .A(n12826), .ZN(n12863) );
  NAND2_X1 U9655 ( .A1(n9338), .A2(n15488), .ZN(n9356) );
  NAND2_X1 U9656 ( .A1(n9211), .A2(n11219), .ZN(n9228) );
  OR2_X1 U9657 ( .A1(n9160), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9171) );
  INV_X1 U9658 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9635) );
  INV_X1 U9659 ( .A(n12626), .ZN(n12847) );
  NAND2_X1 U9660 ( .A1(n9433), .A2(n9432), .ZN(n9447) );
  INV_X1 U9661 ( .A(n12949), .ZN(n12925) );
  AND2_X1 U9662 ( .A1(n9322), .A2(n9321), .ZN(n9338) );
  INV_X1 U9663 ( .A(n12261), .ZN(n15124) );
  NAND2_X1 U9664 ( .A1(n13101), .A2(n13068), .ZN(n9654) );
  OR2_X1 U9665 ( .A1(n9579), .A2(n9578), .ZN(n9649) );
  OR2_X1 U9666 ( .A1(n15177), .A2(n13099), .ZN(n13100) );
  INV_X1 U9667 ( .A(n15120), .ZN(n12985) );
  AND2_X1 U9668 ( .A1(n9633), .A2(n10779), .ZN(n13019) );
  AND2_X1 U9669 ( .A1(n9588), .A2(n9587), .ZN(n12867) );
  NAND2_X1 U9670 ( .A1(n9548), .A2(n6647), .ZN(n10936) );
  INV_X1 U9671 ( .A(n13340), .ZN(n13316) );
  INV_X1 U9672 ( .A(n9037), .ZN(n9933) );
  INV_X1 U9673 ( .A(n11557), .ZN(n9029) );
  OR2_X1 U9674 ( .A1(n10143), .A2(n10142), .ZN(n10279) );
  OR2_X1 U9675 ( .A1(n10136), .A2(n10137), .ZN(n10288) );
  OR2_X1 U9676 ( .A1(n10284), .A2(n10285), .ZN(n11763) );
  INV_X1 U9677 ( .A(n9010), .ZN(n11589) );
  OR2_X1 U9678 ( .A1(n10019), .A2(n8658), .ZN(n13342) );
  NAND2_X1 U9679 ( .A1(n13684), .A2(n8688), .ZN(n11956) );
  INV_X1 U9680 ( .A(n9008), .ZN(n14939) );
  NAND2_X1 U9681 ( .A1(n10857), .A2(n8675), .ZN(n11007) );
  AND2_X1 U9682 ( .A1(n8932), .A2(n8651), .ZN(n13530) );
  OR2_X1 U9683 ( .A1(n8419), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8433) );
  INV_X1 U9684 ( .A(n8252), .ZN(n8402) );
  NAND2_X1 U9685 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NOR2_X1 U9686 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  OR2_X1 U9687 ( .A1(n10269), .A2(n10255), .ZN(n13831) );
  OR2_X1 U9688 ( .A1(n8070), .A2(n14077), .ZN(n7665) );
  AND2_X1 U9689 ( .A1(n8004), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8017) );
  OR2_X1 U9690 ( .A1(n7952), .A2(n7951), .ZN(n7971) );
  NAND2_X1 U9691 ( .A1(n14093), .A2(n14234), .ZN(n14094) );
  INV_X1 U9692 ( .A(n9772), .ZN(n8121) );
  INV_X1 U9693 ( .A(n11532), .ZN(n9685) );
  INV_X1 U9694 ( .A(n13908), .ZN(n11860) );
  AND2_X1 U9695 ( .A1(n8955), .A2(n8954), .ZN(n8956) );
  AND2_X1 U9696 ( .A1(n7597), .A2(n7596), .ZN(n7913) );
  XNOR2_X1 U9697 ( .A(n7582), .B(SI_12_), .ZN(n7848) );
  AND2_X1 U9698 ( .A1(n7571), .A2(n7570), .ZN(n7777) );
  INV_X1 U9699 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U9700 ( .A1(n12599), .A2(n12598), .ZN(n12597) );
  NAND2_X1 U9701 ( .A1(n10794), .A2(n15123), .ZN(n15040) );
  OR2_X1 U9702 ( .A1(n11560), .A2(n9575), .ZN(n10782) );
  OR2_X1 U9703 ( .A1(n10674), .A2(n10665), .ZN(n10680) );
  INV_X1 U9704 ( .A(n15071), .ZN(n15099) );
  INV_X1 U9705 ( .A(n12765), .ZN(n15097) );
  NOR2_X1 U9706 ( .A1(n10680), .A2(n10679), .ZN(n12774) );
  INV_X1 U9707 ( .A(n13019), .ZN(n15114) );
  INV_X1 U9708 ( .A(n15123), .ZN(n12990) );
  AND2_X1 U9709 ( .A1(n15192), .A2(n15155), .ZN(n13068) );
  INV_X1 U9710 ( .A(n12999), .ZN(n12994) );
  NAND2_X1 U9711 ( .A1(n12867), .A2(n15166), .ZN(n15174) );
  INV_X1 U9712 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9283) );
  AND2_X1 U9713 ( .A1(n10021), .A2(n10020), .ZN(n10032) );
  INV_X1 U9714 ( .A(n13342), .ZN(n13315) );
  INV_X1 U9715 ( .A(n13350), .ZN(n14574) );
  INV_X1 U9716 ( .A(n14581), .ZN(n13322) );
  INV_X1 U9717 ( .A(n6583), .ZN(n8657) );
  AND4_X1 U9718 ( .A1(n8606), .A2(n8605), .A3(n8604), .A4(n8603), .ZN(n13341)
         );
  INV_X1 U9719 ( .A(n14883), .ZN(n14922) );
  AND2_X1 U9720 ( .A1(n10024), .A2(n10023), .ZN(n14915) );
  INV_X1 U9721 ( .A(n14951), .ZN(n14937) );
  INV_X1 U9722 ( .A(n10410), .ZN(n13512) );
  INV_X1 U9723 ( .A(n15024), .ZN(n13682) );
  NAND2_X1 U9724 ( .A1(n14974), .A2(n14970), .ZN(n15024) );
  NOR2_X1 U9725 ( .A1(n14964), .A2(n8738), .ZN(n9637) );
  INV_X1 U9726 ( .A(n13831), .ZN(n14615) );
  NAND2_X1 U9727 ( .A1(n10258), .A2(n14698), .ZN(n14618) );
  INV_X1 U9728 ( .A(n7988), .ZN(n9660) );
  INV_X1 U9729 ( .A(n14691), .ZN(n14002) );
  INV_X1 U9730 ( .A(n14687), .ZN(n14038) );
  NAND2_X1 U9731 ( .A1(n14095), .A2(n14094), .ZN(n14096) );
  NAND2_X1 U9732 ( .A1(n10257), .A2(n10256), .ZN(n14698) );
  INV_X1 U9733 ( .A(n14381), .ZN(n8212) );
  INV_X1 U9734 ( .A(n14626), .ZN(n14749) );
  NAND2_X1 U9735 ( .A1(n10501), .A2(n14723), .ZN(n14626) );
  NAND2_X1 U9736 ( .A1(n8141), .A2(n8140), .ZN(n14741) );
  XNOR2_X1 U9737 ( .A(n8186), .B(n8185), .ZN(n10000) );
  AND2_X1 U9738 ( .A1(n10674), .A2(n10673), .ZN(n15093) );
  INV_X1 U9739 ( .A(n12620), .ZN(n11826) );
  NAND2_X1 U9740 ( .A1(n10819), .A2(n11073), .ZN(n15043) );
  AND4_X1 U9741 ( .A1(n12066), .A2(n9600), .A3(n9599), .A4(n9598), .ZN(n12067)
         );
  OR2_X2 U9742 ( .A1(n10782), .A2(n9900), .ZN(n12637) );
  INV_X1 U9743 ( .A(n15093), .ZN(n15088) );
  INV_X1 U9744 ( .A(n12774), .ZN(n15103) );
  OR2_X1 U9745 ( .A1(n9590), .A2(n9589), .ZN(n13004) );
  NAND2_X1 U9746 ( .A1(n6576), .A2(n15127), .ZN(n13011) );
  AND2_X1 U9747 ( .A1(n11380), .A2(n11379), .ZN(n15159) );
  NAND2_X1 U9748 ( .A1(n15192), .A2(n15174), .ZN(n13095) );
  INV_X1 U9749 ( .A(n15192), .ZN(n15189) );
  NAND2_X1 U9750 ( .A1(n15177), .A2(n15174), .ZN(n13177) );
  INV_X1 U9751 ( .A(n15177), .ZN(n15176) );
  INV_X1 U9752 ( .A(n13148), .ZN(n13169) );
  NAND2_X1 U9753 ( .A1(n10010), .A2(n10016), .ZN(n10080) );
  INV_X1 U9754 ( .A(SI_17_), .ZN(n10451) );
  INV_X1 U9755 ( .A(SI_12_), .ZN(n10008) );
  INV_X1 U9756 ( .A(n15081), .ZN(n11213) );
  AND2_X1 U9757 ( .A1(n10032), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14760) );
  INV_X1 U9758 ( .A(n14576), .ZN(n13318) );
  INV_X1 U9759 ( .A(n13313), .ZN(n13325) );
  INV_X1 U9760 ( .A(n13343), .ZN(n13355) );
  OR2_X1 U9761 ( .A1(n10022), .A2(n10023), .ZN(n14883) );
  INV_X1 U9762 ( .A(n14760), .ZN(n14930) );
  NAND2_X1 U9763 ( .A1(n13512), .A2(n10441), .ZN(n13604) );
  AOI21_X1 U9764 ( .B1(n8937), .B2(n8743), .A(n8742), .ZN(n8744) );
  INV_X1 U9765 ( .A(n15037), .ZN(n15035) );
  AND2_X1 U9766 ( .A1(n14595), .A2(n14594), .ZN(n14608) );
  INV_X1 U9767 ( .A(n15027), .ZN(n15025) );
  INV_X1 U9768 ( .A(n14959), .ZN(n14960) );
  INV_X1 U9769 ( .A(n14963), .ZN(n14966) );
  INV_X1 U9770 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11529) );
  INV_X1 U9771 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10336) );
  INV_X1 U9772 ( .A(n11525), .ZN(n12016) );
  NAND2_X1 U9773 ( .A1(n7527), .A2(n9895), .ZN(n9896) );
  INV_X1 U9774 ( .A(n13862), .ZN(n14235) );
  OR2_X1 U9775 ( .A1(n14657), .A2(n10044), .ZN(n14687) );
  OR2_X1 U9776 ( .A1(n14657), .A2(n13934), .ZN(n14691) );
  INV_X1 U9777 ( .A(n14121), .ZN(n14232) );
  AND2_X2 U9778 ( .A1(n14063), .A2(n14698), .ZN(n14712) );
  NAND2_X1 U9779 ( .A1(n14225), .A2(n10513), .ZN(n14248) );
  NOR2_X1 U9780 ( .A1(n8193), .A2(n8194), .ZN(n8195) );
  NAND2_X1 U9781 ( .A1(n14759), .A2(n14744), .ZN(n14304) );
  OR2_X1 U9782 ( .A1(n8197), .A2(n8196), .ZN(n14757) );
  OR2_X1 U9783 ( .A1(n8197), .A2(n10455), .ZN(n14751) );
  INV_X2 U9784 ( .A(n14751), .ZN(n14752) );
  AND2_X1 U9785 ( .A1(n10000), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9989) );
  INV_X1 U9786 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n15367) );
  INV_X1 U9787 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10221) );
  INV_X1 U9788 ( .A(n12637), .ZN(P3_U3897) );
  NAND2_X1 U9789 ( .A1(n9657), .A2(n9656), .ZN(P3_U3488) );
  OAI21_X1 U9790 ( .B1(n9642), .B2(n15025), .A(n9641), .ZN(P2_U3496) );
  NOR2_X1 U9791 ( .A1(n10262), .A2(n10002), .ZN(P1_U4016) );
  NAND2_X1 U9792 ( .A1(n7546), .A2(SI_1_), .ZN(n7548) );
  INV_X1 U9793 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9070) );
  INV_X1 U9794 ( .A(SI_0_), .ZN(n9072) );
  NOR2_X1 U9795 ( .A1(n7547), .A2(n9072), .ZN(n7677) );
  NAND2_X1 U9796 ( .A1(n7549), .A2(SI_2_), .ZN(n7551) );
  OAI21_X1 U9797 ( .B1(SI_2_), .B2(n7549), .A(n7551), .ZN(n7710) );
  INV_X1 U9798 ( .A(n7710), .ZN(n7550) );
  NAND2_X1 U9799 ( .A1(n7553), .A2(SI_3_), .ZN(n7556) );
  INV_X1 U9800 ( .A(n7553), .ZN(n7554) );
  INV_X1 U9801 ( .A(SI_3_), .ZN(n15372) );
  NAND2_X1 U9802 ( .A1(n7554), .A2(n15372), .ZN(n7555) );
  AND2_X1 U9803 ( .A1(n7556), .A2(n7555), .ZN(n7723) );
  NAND2_X1 U9804 ( .A1(n7557), .A2(SI_4_), .ZN(n7560) );
  INV_X1 U9805 ( .A(n7557), .ZN(n7558) );
  INV_X1 U9806 ( .A(SI_4_), .ZN(n9971) );
  NAND2_X1 U9807 ( .A1(n7558), .A2(n9971), .ZN(n7559) );
  AND2_X1 U9808 ( .A1(n7560), .A2(n7559), .ZN(n7731) );
  MUX2_X1 U9809 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7047), .Z(n7561) );
  NAND2_X1 U9810 ( .A1(n7561), .A2(SI_5_), .ZN(n7564) );
  INV_X1 U9811 ( .A(n7561), .ZN(n7562) );
  INV_X1 U9812 ( .A(SI_5_), .ZN(n9974) );
  NAND2_X1 U9813 ( .A1(n7562), .A2(n9974), .ZN(n7563) );
  NAND2_X1 U9814 ( .A1(n7565), .A2(SI_6_), .ZN(n7567) );
  OAI21_X1 U9815 ( .B1(SI_6_), .B2(n7565), .A(n7567), .ZN(n7566) );
  INV_X1 U9816 ( .A(n7566), .ZN(n7763) );
  NAND2_X1 U9817 ( .A1(n7764), .A2(n7763), .ZN(n7766) );
  MUX2_X1 U9818 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9957), .Z(n7568) );
  NAND2_X1 U9819 ( .A1(n7568), .A2(SI_7_), .ZN(n7571) );
  INV_X1 U9820 ( .A(n7568), .ZN(n7569) );
  INV_X1 U9821 ( .A(SI_7_), .ZN(n9977) );
  NAND2_X1 U9822 ( .A1(n7569), .A2(n9977), .ZN(n7570) );
  NAND2_X1 U9823 ( .A1(n7778), .A2(n7777), .ZN(n7780) );
  NAND2_X1 U9824 ( .A1(n7780), .A2(n7571), .ZN(n7792) );
  MUX2_X1 U9825 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9957), .Z(n7572) );
  NAND2_X1 U9826 ( .A1(n7572), .A2(SI_8_), .ZN(n7574) );
  OAI21_X1 U9827 ( .B1(SI_8_), .B2(n7572), .A(n7574), .ZN(n7573) );
  INV_X1 U9828 ( .A(n7573), .ZN(n7791) );
  NAND2_X1 U9829 ( .A1(n7792), .A2(n7791), .ZN(n7794) );
  NAND2_X1 U9830 ( .A1(n7575), .A2(SI_9_), .ZN(n7577) );
  OAI21_X1 U9831 ( .B1(SI_9_), .B2(n7575), .A(n7577), .ZN(n7576) );
  INV_X1 U9832 ( .A(n7576), .ZN(n7807) );
  MUX2_X1 U9833 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9957), .Z(n7822) );
  NOR2_X1 U9834 ( .A1(n7578), .A2(n9982), .ZN(n7580) );
  NAND2_X1 U9835 ( .A1(n7578), .A2(n9982), .ZN(n7579) );
  MUX2_X1 U9836 ( .A(n10221), .B(n10224), .S(n9957), .Z(n7581) );
  MUX2_X1 U9837 ( .A(n9280), .B(n10336), .S(n9957), .Z(n7582) );
  NAND2_X1 U9838 ( .A1(n7582), .A2(n10008), .ZN(n7583) );
  MUX2_X1 U9839 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9957), .Z(n7859) );
  NOR2_X1 U9840 ( .A1(n7859), .A2(SI_13_), .ZN(n7585) );
  NAND2_X1 U9841 ( .A1(n7859), .A2(SI_13_), .ZN(n7584) );
  MUX2_X1 U9842 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9957), .Z(n7874) );
  INV_X1 U9843 ( .A(n7874), .ZN(n7587) );
  INV_X1 U9844 ( .A(SI_15_), .ZN(n7589) );
  NAND2_X1 U9845 ( .A1(n7590), .A2(n7589), .ZN(n7593) );
  INV_X1 U9846 ( .A(n7590), .ZN(n7591) );
  NAND2_X1 U9847 ( .A1(n7591), .A2(SI_15_), .ZN(n7592) );
  INV_X1 U9848 ( .A(n7594), .ZN(n7595) );
  NAND2_X1 U9849 ( .A1(n7595), .A2(SI_16_), .ZN(n7596) );
  XNOR2_X1 U9850 ( .A(n7600), .B(SI_19_), .ZN(n7961) );
  INV_X1 U9851 ( .A(n7946), .ZN(n7959) );
  INV_X1 U9852 ( .A(SI_18_), .ZN(n10511) );
  NOR2_X1 U9853 ( .A1(n7959), .A2(n10511), .ZN(n7599) );
  INV_X1 U9854 ( .A(n7600), .ZN(n7601) );
  INV_X1 U9855 ( .A(SI_19_), .ZN(n10537) );
  NAND2_X1 U9856 ( .A1(n7601), .A2(n10537), .ZN(n7602) );
  NAND2_X1 U9857 ( .A1(n7605), .A2(SI_20_), .ZN(n7603) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9957), .Z(n7604) );
  NAND2_X1 U9859 ( .A1(n7604), .A2(SI_21_), .ZN(n7609) );
  OAI21_X1 U9860 ( .B1(SI_21_), .B2(n7604), .A(n7609), .ZN(n7996) );
  NOR2_X1 U9861 ( .A1(n7605), .A2(SI_20_), .ZN(n7606) );
  NOR2_X1 U9862 ( .A1(n7996), .A2(n7606), .ZN(n7607) );
  INV_X1 U9863 ( .A(SI_22_), .ZN(n15431) );
  MUX2_X1 U9864 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9957), .Z(n8565) );
  NAND2_X1 U9865 ( .A1(n7610), .A2(SI_22_), .ZN(n7611) );
  MUX2_X1 U9866 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9957), .Z(n7612) );
  NAND2_X1 U9867 ( .A1(n7612), .A2(SI_23_), .ZN(n7614) );
  OAI21_X1 U9868 ( .B1(SI_23_), .B2(n7612), .A(n7614), .ZN(n8028) );
  INV_X1 U9869 ( .A(n8028), .ZN(n7613) );
  NAND2_X1 U9870 ( .A1(n8027), .A2(n7613), .ZN(n7615) );
  NAND2_X1 U9871 ( .A1(n7616), .A2(SI_24_), .ZN(n7618) );
  OAI21_X1 U9872 ( .B1(SI_24_), .B2(n7616), .A(n7618), .ZN(n7617) );
  INV_X1 U9873 ( .A(n7617), .ZN(n8037) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9957), .Z(n7619) );
  XNOR2_X1 U9875 ( .A(n7619), .B(SI_25_), .ZN(n8049) );
  INV_X1 U9876 ( .A(n7619), .ZN(n7620) );
  INV_X1 U9877 ( .A(SI_25_), .ZN(n11562) );
  NAND2_X1 U9878 ( .A1(n7620), .A2(n11562), .ZN(n7621) );
  INV_X1 U9879 ( .A(SI_26_), .ZN(n15326) );
  INV_X1 U9880 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14411) );
  INV_X1 U9881 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13740) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9957), .Z(n8077) );
  INV_X1 U9883 ( .A(n8077), .ZN(n7624) );
  NAND2_X1 U9884 ( .A1(n7624), .A2(n15275), .ZN(n7625) );
  NAND2_X1 U9885 ( .A1(n8077), .A2(SI_27_), .ZN(n7626) );
  XNOR2_X1 U9886 ( .A(n7628), .B(SI_28_), .ZN(n7669) );
  INV_X1 U9887 ( .A(n7628), .ZN(n7629) );
  INV_X1 U9888 ( .A(SI_28_), .ZN(n12433) );
  NAND2_X1 U9889 ( .A1(n7629), .A2(n12433), .ZN(n7630) );
  INV_X1 U9890 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14398) );
  INV_X1 U9891 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13732) );
  MUX2_X1 U9892 ( .A(n14398), .B(n13732), .S(n9957), .Z(n8921) );
  XNOR2_X1 U9893 ( .A(n8921), .B(SI_29_), .ZN(n8919) );
  NOR2_X2 U9894 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n7898) );
  NOR2_X1 U9895 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7635) );
  NOR2_X1 U9896 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7634) );
  NOR2_X1 U9897 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7633) );
  NOR2_X1 U9898 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7638) );
  NOR2_X1 U9899 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7637) );
  NOR2_X1 U9900 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n7639) );
  NAND2_X2 U9901 ( .A1(n14401), .A2(n14653), .ZN(n8016) );
  NAND2_X1 U9902 ( .A1(n13728), .A2(n9675), .ZN(n7645) );
  OR2_X1 U9903 ( .A1(n9677), .A2(n14398), .ZN(n7644) );
  INV_X1 U9904 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n15369) );
  OR2_X1 U9905 ( .A1(n8149), .A2(n15369), .ZN(n7659) );
  NAND2_X1 U9906 ( .A1(n7699), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U9907 ( .A1(n7988), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7657) );
  AND3_X1 U9908 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U9909 ( .A1(n7785), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U9910 ( .A1(n7815), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7829) );
  INV_X1 U9911 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U9912 ( .A1(n7867), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7885) );
  INV_X1 U9913 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7884) );
  INV_X1 U9914 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7904) );
  INV_X1 U9915 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7951) );
  INV_X1 U9916 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13759) );
  NAND2_X1 U9917 ( .A1(n8017), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U9918 ( .A1(n8032), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U9919 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n8043), .ZN(n8054) );
  INV_X1 U9920 ( .A(n8054), .ZN(n7652) );
  NAND2_X1 U9921 ( .A1(n7652), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8068) );
  INV_X1 U9922 ( .A(n8068), .ZN(n7653) );
  NAND2_X1 U9923 ( .A1(n7653), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8082) );
  INV_X1 U9924 ( .A(n8082), .ZN(n7654) );
  NAND2_X1 U9925 ( .A1(n7654), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8084) );
  INV_X1 U9926 ( .A(n8084), .ZN(n7655) );
  NAND2_X1 U9927 ( .A1(n7655), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14061) );
  OR2_X1 U9928 ( .A1(n8070), .A2(n14061), .ZN(n7656) );
  NAND4_X1 U9929 ( .A1(n7659), .A2(n7658), .A3(n7657), .A4(n7656), .ZN(n13892)
         );
  XNOR2_X1 U9930 ( .A(n14067), .B(n13892), .ZN(n9880) );
  NAND2_X1 U9931 ( .A1(n6584), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7667) );
  INV_X1 U9932 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7660) );
  OR2_X1 U9933 ( .A1(n8009), .A2(n7660), .ZN(n7666) );
  INV_X1 U9934 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9935 ( .A1(n8084), .A2(n7661), .ZN(n7662) );
  NAND2_X1 U9936 ( .A1(n14061), .A2(n7662), .ZN(n14077) );
  INV_X1 U9937 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7663) );
  OR2_X1 U9938 ( .A1(n9660), .A2(n7663), .ZN(n7664) );
  NAND2_X1 U9939 ( .A1(n13733), .A2(n9675), .ZN(n7671) );
  INV_X1 U9940 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14404) );
  OR2_X1 U9941 ( .A1(n9677), .A2(n14404), .ZN(n7670) );
  NAND2_X1 U9942 ( .A1(n7699), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7676) );
  INV_X1 U9943 ( .A(n7677), .ZN(n7678) );
  NAND2_X1 U9944 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  NAND2_X1 U9945 ( .A1(n7681), .A2(n7680), .ZN(n9948) );
  NAND2_X1 U9946 ( .A1(n9957), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7682) );
  OAI21_X1 U9947 ( .B1(n9948), .B2(n9957), .A(n7682), .ZN(n7683) );
  INV_X1 U9948 ( .A(n14401), .ZN(n13934) );
  NAND2_X1 U9949 ( .A1(n7683), .A2(n13934), .ZN(n7691) );
  NAND2_X1 U9950 ( .A1(n9948), .A2(n9945), .ZN(n7684) );
  INV_X1 U9951 ( .A(n6586), .ZN(n10059) );
  OAI211_X1 U9952 ( .C1(n9945), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n7684), .B(
        n10059), .ZN(n7690) );
  NAND2_X1 U9953 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7685) );
  MUX2_X1 U9954 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7685), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7688) );
  INV_X1 U9955 ( .A(n7686), .ZN(n7687) );
  NAND2_X1 U9956 ( .A1(n7688), .A2(n7687), .ZN(n13921) );
  INV_X1 U9957 ( .A(n13921), .ZN(n13926) );
  NAND3_X1 U9958 ( .A1(n14401), .A2(n13926), .A3(n6586), .ZN(n7689) );
  OR2_X2 U9959 ( .A1(n13917), .A2(n10631), .ZN(n9691) );
  NAND2_X1 U9960 ( .A1(n13917), .A2(n10631), .ZN(n9690) );
  NAND2_X1 U9961 ( .A1(n7928), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7696) );
  INV_X1 U9962 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7692) );
  OR2_X1 U9963 ( .A1(n8009), .A2(n7692), .ZN(n7695) );
  INV_X1 U9964 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10769) );
  OR2_X1 U9965 ( .A1(n8044), .A2(n10769), .ZN(n7694) );
  INV_X1 U9966 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14652) );
  INV_X1 U9967 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13935) );
  XNOR2_X1 U9968 ( .A(n7697), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14416) );
  INV_X1 U9969 ( .A(n10771), .ZN(n10263) );
  NAND2_X1 U9970 ( .A1(n13918), .A2(n10263), .ZN(n10493) );
  INV_X1 U9971 ( .A(n10493), .ZN(n7698) );
  INV_X1 U9972 ( .A(n10631), .ZN(n13770) );
  NAND2_X1 U9973 ( .A1(n7672), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U9974 ( .A1(n8020), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U9975 ( .A1(n7741), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7701) );
  NOR2_X1 U9976 ( .A1(n7686), .A2(n7918), .ZN(n7704) );
  MUX2_X1 U9977 ( .A(n7918), .B(n7704), .S(P1_IR_REG_2__SCAN_IN), .Z(n7705) );
  INV_X1 U9978 ( .A(n7705), .ZN(n7708) );
  INV_X1 U9979 ( .A(n7706), .ZN(n7707) );
  NAND2_X1 U9980 ( .A1(n7708), .A2(n7707), .ZN(n13944) );
  INV_X1 U9981 ( .A(n7709), .ZN(n7711) );
  NAND2_X1 U9982 ( .A1(n7711), .A2(n7710), .ZN(n7713) );
  NAND2_X1 U9983 ( .A1(n7713), .A2(n7712), .ZN(n9946) );
  OR2_X2 U9984 ( .A1(n9677), .A2(n9947), .ZN(n7714) );
  NAND2_X1 U9985 ( .A1(n13915), .A2(n14716), .ZN(n7716) );
  NAND2_X1 U9986 ( .A1(n10453), .A2(n10452), .ZN(n7718) );
  OR2_X1 U9987 ( .A1(n13915), .A2(n10463), .ZN(n7717) );
  NAND2_X1 U9988 ( .A1(n7718), .A2(n7717), .ZN(n10606) );
  NAND2_X1 U9989 ( .A1(n7741), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U9990 ( .A1(n7672), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7721) );
  NAND2_X1 U9991 ( .A1(n7757), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7720) );
  OR2_X1 U9992 ( .A1(n8044), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7719) );
  OR2_X1 U9993 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  AND2_X1 U9994 ( .A1(n7726), .A2(n7725), .ZN(n9941) );
  OR2_X1 U9995 ( .A1(n7706), .A2(n7918), .ZN(n7727) );
  XNOR2_X1 U9996 ( .A(n7727), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13950) );
  INV_X1 U9997 ( .A(n10608), .ZN(n7728) );
  NAND2_X1 U9998 ( .A1(n10606), .A2(n7728), .ZN(n7730) );
  INV_X1 U9999 ( .A(n10892), .ZN(n14727) );
  NAND2_X1 U10000 ( .A1(n10896), .A2(n14727), .ZN(n7729) );
  OR2_X1 U10001 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  NAND2_X1 U10002 ( .A1(n9943), .A2(n9675), .ZN(n7740) );
  NAND2_X1 U10003 ( .A1(n7706), .A2(n7735), .ZN(n7737) );
  NAND2_X1 U10004 ( .A1(n7737), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7736) );
  MUX2_X1 U10005 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7736), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7738) );
  AND2_X1 U10006 ( .A1(n7738), .A2(n7751), .ZN(n13972) );
  AOI22_X1 U10007 ( .A1(n7968), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9999), .B2(
        n13972), .ZN(n7739) );
  NAND2_X1 U10008 ( .A1(n7740), .A2(n7739), .ZN(n10929) );
  INV_X1 U10009 ( .A(n10929), .ZN(n14736) );
  NAND2_X1 U10010 ( .A1(n6584), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U10011 ( .A1(n7757), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10012 ( .A1(n7741), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7743) );
  XNOR2_X1 U10014 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10928) );
  OR2_X1 U10015 ( .A1(n8070), .A2(n10928), .ZN(n7742) );
  NAND4_X1 U10016 ( .A1(n7745), .A2(n7744), .A3(n7743), .A4(n7742), .ZN(n13913) );
  INV_X1 U10017 ( .A(n13913), .ZN(n10905) );
  NAND2_X1 U10018 ( .A1(n14736), .A2(n10905), .ZN(n9861) );
  NAND2_X1 U10019 ( .A1(n10929), .A2(n13913), .ZN(n9860) );
  OR2_X1 U10020 ( .A1(n7747), .A2(n7746), .ZN(n7748) );
  NAND2_X1 U10021 ( .A1(n7749), .A2(n7748), .ZN(n9953) );
  OR2_X1 U10022 ( .A1(n9953), .A2(n8064), .ZN(n7756) );
  NAND2_X1 U10023 ( .A1(n7751), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7750) );
  MUX2_X1 U10024 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7750), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7754) );
  INV_X1 U10025 ( .A(n7751), .ZN(n7753) );
  INV_X1 U10026 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7752) );
  NAND2_X1 U10027 ( .A1(n7753), .A2(n7752), .ZN(n7781) );
  NAND2_X1 U10028 ( .A1(n7754), .A2(n7781), .ZN(n10052) );
  INV_X1 U10029 ( .A(n10052), .ZN(n13985) );
  AOI22_X1 U10030 ( .A1(n7968), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9999), .B2(
        n13985), .ZN(n7755) );
  NAND2_X1 U10031 ( .A1(n7756), .A2(n7755), .ZN(n10914) );
  NAND2_X1 U10032 ( .A1(n6584), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U10033 ( .A1(n7757), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7761) );
  AOI21_X1 U10034 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7758) );
  NOR2_X1 U10035 ( .A1(n7758), .A2(n7770), .ZN(n10923) );
  NAND2_X1 U10036 ( .A1(n8020), .A2(n10923), .ZN(n7760) );
  NAND2_X1 U10037 ( .A1(n7741), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7759) );
  NAND4_X1 U10038 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n13912) );
  INV_X1 U10039 ( .A(n13912), .ZN(n8104) );
  XNOR2_X1 U10040 ( .A(n10914), .B(n8104), .ZN(n9864) );
  INV_X1 U10041 ( .A(n9864), .ZN(n10561) );
  INV_X1 U10042 ( .A(n10914), .ZN(n10921) );
  OR2_X1 U10043 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  NAND2_X1 U10044 ( .A1(n7766), .A2(n7765), .ZN(n9979) );
  OR2_X1 U10045 ( .A1(n9979), .A2(n8064), .ZN(n7769) );
  NAND2_X1 U10046 ( .A1(n7781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7767) );
  XNOR2_X1 U10047 ( .A(n7767), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U10048 ( .A1(n7968), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9999), .B2(
        n10122), .ZN(n7768) );
  NAND2_X1 U10049 ( .A1(n7769), .A2(n7768), .ZN(n11036) );
  NAND2_X1 U10050 ( .A1(n7757), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U10051 ( .A1(n6584), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7774) );
  NOR2_X1 U10052 ( .A1(n7770), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7771) );
  NOR2_X1 U10053 ( .A1(n7785), .A2(n7771), .ZN(n11044) );
  NAND2_X1 U10054 ( .A1(n8020), .A2(n11044), .ZN(n7773) );
  NAND2_X1 U10055 ( .A1(n7741), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7772) );
  NAND4_X1 U10056 ( .A1(n7775), .A2(n7774), .A3(n7773), .A4(n7772), .ZN(n13911) );
  XNOR2_X1 U10057 ( .A(n11036), .B(n13911), .ZN(n9865) );
  INV_X1 U10058 ( .A(n9865), .ZN(n10695) );
  NAND2_X1 U10059 ( .A1(n10691), .A2(n10695), .ZN(n10690) );
  OR2_X1 U10060 ( .A1(n11036), .A2(n13911), .ZN(n7776) );
  NAND2_X1 U10061 ( .A1(n10690), .A2(n7776), .ZN(n11048) );
  OR2_X1 U10062 ( .A1(n7778), .A2(n7777), .ZN(n7779) );
  NAND2_X1 U10063 ( .A1(n7780), .A2(n7779), .ZN(n9985) );
  OR2_X1 U10064 ( .A1(n9985), .A2(n8064), .ZN(n7784) );
  OAI21_X1 U10065 ( .B1(n7781), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7782) );
  XNOR2_X1 U10066 ( .A(n7782), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14004) );
  AOI22_X1 U10067 ( .A1(n7968), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9999), .B2(
        n14004), .ZN(n7783) );
  NAND2_X1 U10068 ( .A1(n7784), .A2(n7783), .ZN(n14702) );
  NAND2_X1 U10069 ( .A1(n6584), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10070 ( .A1(n7757), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U10071 ( .A1(n7741), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7787) );
  OAI21_X1 U10072 ( .B1(n7785), .B2(P1_REG3_REG_7__SCAN_IN), .A(n7800), .ZN(
        n14699) );
  OR2_X1 U10073 ( .A1(n8044), .A2(n14699), .ZN(n7786) );
  NAND4_X1 U10074 ( .A1(n7789), .A2(n7788), .A3(n7787), .A4(n7786), .ZN(n13910) );
  XNOR2_X1 U10075 ( .A(n14702), .B(n13910), .ZN(n9866) );
  INV_X1 U10076 ( .A(n9866), .ZN(n11051) );
  NAND2_X1 U10077 ( .A1(n11048), .A2(n11051), .ZN(n11047) );
  OR2_X1 U10078 ( .A1(n14702), .A2(n13910), .ZN(n7790) );
  OR2_X1 U10079 ( .A1(n7792), .A2(n7791), .ZN(n7793) );
  NAND2_X1 U10080 ( .A1(n7794), .A2(n7793), .ZN(n9993) );
  OR2_X1 U10081 ( .A1(n9993), .A2(n8064), .ZN(n7798) );
  OR2_X1 U10082 ( .A1(n7795), .A2(n7918), .ZN(n7796) );
  XNOR2_X1 U10083 ( .A(n7796), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U10084 ( .A1(n7968), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9999), .B2(
        n10072), .ZN(n7797) );
  NAND2_X2 U10085 ( .A1(n7798), .A2(n7797), .ZN(n14745) );
  NAND2_X1 U10086 ( .A1(n7757), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U10087 ( .A1(n6584), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U10088 ( .A1(n7741), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7803) );
  AND2_X1 U10089 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  OR2_X1 U10090 ( .A1(n7801), .A2(n7815), .ZN(n11574) );
  OR2_X1 U10091 ( .A1(n8070), .A2(n11574), .ZN(n7802) );
  NAND4_X1 U10092 ( .A1(n7805), .A2(n7804), .A3(n7803), .A4(n7802), .ZN(n13909) );
  XNOR2_X1 U10093 ( .A(n14745), .B(n13909), .ZN(n9868) );
  INV_X1 U10094 ( .A(n9868), .ZN(n10983) );
  NAND2_X1 U10095 ( .A1(n10981), .A2(n10983), .ZN(n10980) );
  OR2_X1 U10096 ( .A1(n14745), .A2(n13909), .ZN(n7806) );
  NAND2_X1 U10097 ( .A1(n10980), .A2(n7806), .ZN(n11337) );
  OR2_X1 U10098 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  NAND2_X1 U10099 ( .A1(n7810), .A2(n7809), .ZN(n10012) );
  OR2_X1 U10100 ( .A1(n10012), .A2(n8064), .ZN(n7814) );
  INV_X1 U10101 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U10102 ( .A1(n7795), .A2(n7811), .ZN(n7824) );
  NAND2_X1 U10103 ( .A1(n7824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7812) );
  XNOR2_X1 U10104 ( .A(n7812), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U10105 ( .A1(n7968), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9999), .B2(
        n10156), .ZN(n7813) );
  NAND2_X1 U10106 ( .A1(n7672), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U10107 ( .A1(n7757), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U10108 ( .A1(n7741), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7818) );
  OR2_X1 U10109 ( .A1(n7815), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U10110 ( .A1(n7829), .A2(n7816), .ZN(n11720) );
  OR2_X1 U10111 ( .A1(n8070), .A2(n11720), .ZN(n7817) );
  NAND4_X1 U10112 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n13908) );
  XNOR2_X1 U10113 ( .A(n11716), .B(n11860), .ZN(n11341) );
  OR2_X1 U10114 ( .A1(n11716), .A2(n13908), .ZN(n7821) );
  XNOR2_X1 U10115 ( .A(n7822), .B(SI_10_), .ZN(n7823) );
  OAI21_X1 U10116 ( .B1(n7824), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7825) );
  XNOR2_X1 U10117 ( .A(n7825), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U10118 ( .A1(n7968), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9999), 
        .B2(n10178), .ZN(n7826) );
  NAND2_X2 U10119 ( .A1(n7827), .A2(n7826), .ZN(n11863) );
  NAND2_X1 U10120 ( .A1(n7757), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U10121 ( .A1(n7741), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U10122 ( .A1(n6584), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7832) );
  NAND2_X1 U10123 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U10124 ( .A1(n7841), .A2(n7830), .ZN(n11859) );
  OR2_X1 U10125 ( .A1(n8044), .A2(n11859), .ZN(n7831) );
  NAND4_X1 U10126 ( .A1(n7834), .A2(n7833), .A3(n7832), .A4(n7831), .ZN(n13907) );
  XNOR2_X1 U10127 ( .A(n11863), .B(n13907), .ZN(n11279) );
  INV_X1 U10128 ( .A(n11279), .ZN(n11289) );
  XNOR2_X1 U10129 ( .A(n7836), .B(n7835), .ZN(n10220) );
  NAND2_X1 U10130 ( .A1(n10220), .A2(n9675), .ZN(n7839) );
  NAND2_X1 U10131 ( .A1(n7963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7837) );
  XNOR2_X1 U10132 ( .A(n7837), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U10133 ( .A1(n7968), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9999), 
        .B2(n10219), .ZN(n7838) );
  NAND2_X1 U10134 ( .A1(n7757), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U10135 ( .A1(n7988), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10136 ( .A1(n6584), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10137 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  NAND2_X1 U10138 ( .A1(n7852), .A2(n7842), .ZN(n11441) );
  OR2_X1 U10139 ( .A1(n8070), .A2(n11441), .ZN(n7843) );
  NAND4_X1 U10140 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n13906) );
  XNOR2_X1 U10141 ( .A(n11525), .B(n13906), .ZN(n11434) );
  INV_X1 U10142 ( .A(n11434), .ZN(n11438) );
  NAND2_X1 U10143 ( .A1(n11439), .A2(n11438), .ZN(n11437) );
  OR2_X1 U10144 ( .A1(n11525), .A2(n13906), .ZN(n7847) );
  XNOR2_X1 U10145 ( .A(n7849), .B(n7848), .ZN(n10247) );
  NAND2_X1 U10146 ( .A1(n10247), .A2(n9675), .ZN(n7851) );
  OR2_X1 U10147 ( .A1(n7963), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10148 ( .A1(n7900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7863) );
  XNOR2_X1 U10149 ( .A(n7863), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U10150 ( .A1(n7968), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9999), 
        .B2(n10482), .ZN(n7850) );
  NAND2_X1 U10151 ( .A1(n7988), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7857) );
  INV_X1 U10152 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10200) );
  OR2_X1 U10153 ( .A1(n8149), .A2(n10200), .ZN(n7856) );
  INV_X1 U10154 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11653) );
  OR2_X1 U10155 ( .A1(n8009), .A2(n11653), .ZN(n7855) );
  AND2_X1 U10156 ( .A1(n7852), .A2(n11996), .ZN(n7853) );
  OR2_X1 U10157 ( .A1(n7853), .A2(n7867), .ZN(n11997) );
  OR2_X1 U10158 ( .A1(n8070), .A2(n11997), .ZN(n7854) );
  XNOR2_X1 U10159 ( .A(n12001), .B(n13905), .ZN(n11648) );
  INV_X1 U10160 ( .A(n11648), .ZN(n11646) );
  NAND2_X1 U10161 ( .A1(n11647), .A2(n11646), .ZN(n11645) );
  NAND2_X1 U10162 ( .A1(n14536), .A2(n13840), .ZN(n7858) );
  NAND2_X1 U10163 ( .A1(n11645), .A2(n7858), .ZN(n11631) );
  INV_X1 U10164 ( .A(SI_13_), .ZN(n15411) );
  XNOR2_X1 U10165 ( .A(n7859), .B(n15411), .ZN(n7860) );
  XNOR2_X1 U10166 ( .A(n7861), .B(n7860), .ZN(n10397) );
  NAND2_X1 U10167 ( .A1(n10397), .A2(n9675), .ZN(n7866) );
  INV_X1 U10168 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10169 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  NAND2_X1 U10170 ( .A1(n7864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7879) );
  XNOR2_X1 U10171 ( .A(n7879), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U10172 ( .A1(n7968), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9999), 
        .B2(n10483), .ZN(n7865) );
  NAND2_X2 U10173 ( .A1(n7866), .A2(n7865), .ZN(n13843) );
  INV_X1 U10174 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11633) );
  OR2_X1 U10175 ( .A1(n8009), .A2(n11633), .ZN(n7872) );
  NAND2_X1 U10176 ( .A1(n6584), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10177 ( .A1(n7988), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7870) );
  OR2_X1 U10178 ( .A1(n7867), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U10179 ( .A1(n7885), .A2(n7868), .ZN(n13839) );
  OR2_X1 U10180 ( .A1(n8044), .A2(n13839), .ZN(n7869) );
  NAND4_X1 U10181 ( .A1(n7872), .A2(n7871), .A3(n7870), .A4(n7869), .ZN(n13904) );
  XNOR2_X1 U10182 ( .A(n13843), .B(n12328), .ZN(n11630) );
  NAND2_X1 U10183 ( .A1(n11631), .A2(n11630), .ZN(n11629) );
  OR2_X1 U10184 ( .A1(n13843), .A2(n13904), .ZN(n7873) );
  NAND2_X1 U10185 ( .A1(n11629), .A2(n7873), .ZN(n11839) );
  NAND2_X1 U10186 ( .A1(n7875), .A2(n7874), .ZN(n7876) );
  NAND2_X1 U10187 ( .A1(n7877), .A2(n7876), .ZN(n10589) );
  NAND2_X1 U10188 ( .A1(n10589), .A2(n9675), .ZN(n7883) );
  INV_X1 U10189 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U10190 ( .A1(n7879), .A2(n7878), .ZN(n7880) );
  NAND2_X1 U10191 ( .A1(n7880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7881) );
  XNOR2_X1 U10192 ( .A(n7881), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U10193 ( .A1(n7968), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9999), 
        .B2(n10486), .ZN(n7882) );
  NAND2_X1 U10194 ( .A1(n7988), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7891) );
  INV_X1 U10195 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10487) );
  OR2_X1 U10196 ( .A1(n8009), .A2(n10487), .ZN(n7890) );
  NAND2_X1 U10197 ( .A1(n7885), .A2(n7884), .ZN(n7886) );
  NAND2_X1 U10198 ( .A1(n7905), .A2(n7886), .ZN(n14621) );
  OR2_X1 U10199 ( .A1(n8070), .A2(n14621), .ZN(n7889) );
  INV_X1 U10200 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7887) );
  OR2_X1 U10201 ( .A1(n8149), .A2(n7887), .ZN(n7888) );
  NAND2_X1 U10202 ( .A1(n14617), .A2(n13885), .ZN(n9749) );
  INV_X1 U10203 ( .A(n11830), .ZN(n11840) );
  INV_X1 U10204 ( .A(n13885), .ZN(n13903) );
  NAND2_X1 U10205 ( .A1(n14617), .A2(n13903), .ZN(n7892) );
  OR2_X1 U10206 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  NAND2_X1 U10207 ( .A1(n7896), .A2(n7895), .ZN(n10841) );
  NAND2_X1 U10208 ( .A1(n10841), .A2(n9675), .ZN(n7903) );
  INV_X1 U10209 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10210 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  NOR2_X1 U10211 ( .A1(n7900), .A2(n7899), .ZN(n7916) );
  OR2_X1 U10212 ( .A1(n7916), .A2(n7918), .ZN(n7901) );
  XNOR2_X1 U10213 ( .A(n7901), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U10214 ( .A1(n7968), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9999), 
        .B2(n11316), .ZN(n7902) );
  AND2_X1 U10215 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  OR2_X1 U10216 ( .A1(n7906), .A2(n7926), .ZN(n13881) );
  NAND2_X1 U10217 ( .A1(n7988), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7907) );
  OAI21_X1 U10218 ( .B1(n13881), .B2(n8070), .A(n7907), .ZN(n7912) );
  INV_X1 U10219 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7910) );
  INV_X1 U10220 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7908) );
  OR2_X1 U10221 ( .A1(n8009), .A2(n7908), .ZN(n7909) );
  OAI21_X1 U10222 ( .B1(n8149), .B2(n7910), .A(n7909), .ZN(n7911) );
  NOR2_X1 U10223 ( .A1(n7912), .A2(n7911), .ZN(n13799) );
  NAND2_X1 U10224 ( .A1(n14351), .A2(n13799), .ZN(n9768) );
  NAND2_X1 U10225 ( .A1(n9766), .A2(n9768), .ZN(n11791) );
  INV_X1 U10226 ( .A(n11791), .ZN(n8118) );
  INV_X1 U10227 ( .A(n13799), .ZN(n13902) );
  XNOR2_X1 U10228 ( .A(n7914), .B(n7913), .ZN(n10940) );
  NAND2_X1 U10229 ( .A1(n10940), .A2(n9675), .ZN(n7925) );
  INV_X1 U10230 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7915) );
  AND2_X1 U10231 ( .A1(n7916), .A2(n7915), .ZN(n7921) );
  NOR2_X1 U10232 ( .A1(n7921), .A2(n7918), .ZN(n7917) );
  MUX2_X1 U10233 ( .A(n7918), .B(n7917), .S(P1_IR_REG_16__SCAN_IN), .Z(n7919)
         );
  INV_X1 U10234 ( .A(n7919), .ZN(n7922) );
  INV_X1 U10235 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10236 ( .A1(n7921), .A2(n7920), .ZN(n7947) );
  NAND2_X1 U10237 ( .A1(n7922), .A2(n7947), .ZN(n14027) );
  INV_X1 U10238 ( .A(n14027), .ZN(n7923) );
  AOI22_X1 U10239 ( .A1(n7923), .A2(n9999), .B1(n7968), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n7924) );
  NOR2_X1 U10240 ( .A1(n7926), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7927) );
  OR2_X1 U10241 ( .A1(n7938), .A2(n7927), .ZN(n13797) );
  AOI22_X1 U10242 ( .A1(n7672), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n7757), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10243 ( .A1(n7988), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7929) );
  OAI211_X1 U10244 ( .C1(n13797), .C2(n8044), .A(n7930), .B(n7929), .ZN(n13901) );
  XNOR2_X1 U10245 ( .A(n11975), .B(n13901), .ZN(n9873) );
  INV_X1 U10246 ( .A(n13901), .ZN(n13882) );
  NAND2_X1 U10247 ( .A1(n14344), .A2(n13882), .ZN(n7931) );
  XNOR2_X1 U10248 ( .A(n7932), .B(SI_17_), .ZN(n7933) );
  XNOR2_X1 U10249 ( .A(n7934), .B(n7933), .ZN(n11079) );
  NAND2_X1 U10250 ( .A1(n11079), .A2(n9675), .ZN(n7937) );
  NAND2_X1 U10251 ( .A1(n7947), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7935) );
  XNOR2_X1 U10252 ( .A(n7935), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14025) );
  AOI22_X1 U10253 ( .A1(n7968), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n14025), 
        .B2(n9999), .ZN(n7936) );
  OR2_X1 U10254 ( .A1(n7938), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7939) );
  AND2_X1 U10255 ( .A1(n7952), .A2(n7939), .ZN(n12025) );
  NAND2_X1 U10256 ( .A1(n12025), .A2(n8020), .ZN(n7942) );
  AOI22_X1 U10257 ( .A1(n6584), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n7757), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n7941) );
  NAND2_X1 U10258 ( .A1(n7988), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7940) );
  INV_X1 U10259 ( .A(n9773), .ZN(n7943) );
  NAND2_X1 U10260 ( .A1(n7944), .A2(n10511), .ZN(n7945) );
  NAND2_X1 U10261 ( .A1(n11461), .A2(n9675), .ZN(n7950) );
  OAI21_X1 U10262 ( .B1(n7947), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7948) );
  XNOR2_X1 U10263 ( .A(n7948), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U10264 ( .A1(n9999), .A2(n14030), .B1(n7968), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7949) );
  NAND2_X2 U10265 ( .A1(n7950), .A2(n7949), .ZN(n14332) );
  NAND2_X1 U10266 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  NAND2_X1 U10267 ( .A1(n7971), .A2(n7953), .ZN(n13860) );
  AOI22_X1 U10268 ( .A1(n7672), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n7757), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n7955) );
  INV_X1 U10269 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15427) );
  OR2_X1 U10270 ( .A1(n9660), .A2(n15427), .ZN(n7954) );
  OAI211_X1 U10271 ( .C1(n13860), .C2(n8070), .A(n7955), .B(n7954), .ZN(n13900) );
  OR2_X1 U10272 ( .A1(n14332), .A2(n13900), .ZN(n7956) );
  NAND2_X1 U10273 ( .A1(n14332), .A2(n13900), .ZN(n7957) );
  XNOR2_X1 U10274 ( .A(n7962), .B(n7961), .ZN(n11517) );
  NAND2_X1 U10275 ( .A1(n11517), .A2(n9675), .ZN(n7970) );
  NAND2_X1 U10276 ( .A1(n7966), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7965) );
  MUX2_X1 U10277 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7965), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n7967) );
  AOI22_X1 U10278 ( .A1(n7968), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10460), 
        .B2(n9999), .ZN(n7969) );
  AND2_X1 U10279 ( .A1(n7971), .A2(n13759), .ZN(n7972) );
  OR2_X1 U10280 ( .A1(n7972), .A2(n7986), .ZN(n14220) );
  INV_X1 U10281 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14032) );
  NAND2_X1 U10282 ( .A1(n7988), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10283 ( .A1(n7757), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7973) );
  OAI211_X1 U10284 ( .C1(n8149), .C2(n14032), .A(n7974), .B(n7973), .ZN(n7975)
         );
  INV_X1 U10285 ( .A(n7975), .ZN(n7976) );
  OAI21_X1 U10286 ( .B1(n14220), .B2(n8070), .A(n7976), .ZN(n14237) );
  INV_X1 U10287 ( .A(n14227), .ZN(n7977) );
  OR2_X1 U10288 ( .A1(n14325), .A2(n14237), .ZN(n7978) );
  INV_X1 U10289 ( .A(SI_20_), .ZN(n12324) );
  NAND2_X1 U10290 ( .A1(n7980), .A2(n12324), .ZN(n7981) );
  NAND2_X1 U10291 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  OR2_X1 U10292 ( .A1(n9677), .A2(n11531), .ZN(n7985) );
  NOR2_X1 U10293 ( .A1(n7986), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7987) );
  OR2_X1 U10294 ( .A1(n8004), .A2(n7987), .ZN(n13828) );
  INV_X1 U10295 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U10296 ( .A1(n7988), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10297 ( .A1(n7757), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7989) );
  OAI211_X1 U10298 ( .C1(n8149), .C2(n7991), .A(n7990), .B(n7989), .ZN(n7992)
         );
  INV_X1 U10299 ( .A(n7992), .ZN(n7993) );
  OAI21_X1 U10300 ( .B1(n13828), .B2(n8070), .A(n7993), .ZN(n13899) );
  NAND2_X1 U10301 ( .A1(n14315), .A2(n13899), .ZN(n7995) );
  AND2_X1 U10302 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  NAND2_X1 U10303 ( .A1(n7999), .A2(n7998), .ZN(n8001) );
  NAND2_X1 U10304 ( .A1(n8001), .A2(n8000), .ZN(n11642) );
  OR2_X1 U10305 ( .A1(n11642), .A2(n8064), .ZN(n8003) );
  INV_X1 U10306 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11643) );
  OR2_X1 U10307 ( .A1(n9677), .A2(n11643), .ZN(n8002) );
  NOR2_X1 U10308 ( .A1(n8004), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8005) );
  OR2_X1 U10309 ( .A1(n8017), .A2(n8005), .ZN(n14197) );
  INV_X1 U10310 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U10311 ( .A1(n6584), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U10312 ( .A1(n7988), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8006) );
  OAI211_X1 U10313 ( .C1(n8009), .C2(n8008), .A(n8007), .B(n8006), .ZN(n8010)
         );
  INV_X1 U10314 ( .A(n8010), .ZN(n8011) );
  OAI21_X1 U10315 ( .B1(n14197), .B2(n8070), .A(n8011), .ZN(n13898) );
  XNOR2_X1 U10316 ( .A(n14384), .B(n13898), .ZN(n14191) );
  OR2_X1 U10317 ( .A1(n14384), .A2(n13898), .ZN(n8012) );
  NAND2_X1 U10318 ( .A1(n8014), .A2(n9945), .ZN(n8015) );
  XNOR2_X1 U10319 ( .A(n8015), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14415) );
  OR2_X1 U10320 ( .A1(n8017), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8019) );
  AND2_X1 U10321 ( .A1(n8019), .A2(n8018), .ZN(n14183) );
  NAND2_X1 U10322 ( .A1(n14183), .A2(n8020), .ZN(n8025) );
  INV_X1 U10323 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n15359) );
  NAND2_X1 U10324 ( .A1(n7757), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10325 ( .A1(n7672), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8021) );
  OAI211_X1 U10326 ( .C1(n9660), .C2(n15359), .A(n8022), .B(n8021), .ZN(n8023)
         );
  INV_X1 U10327 ( .A(n8023), .ZN(n8024) );
  NAND2_X1 U10328 ( .A1(n8025), .A2(n8024), .ZN(n13897) );
  XNOR2_X1 U10329 ( .A(n14380), .B(n13897), .ZN(n14179) );
  OR2_X1 U10330 ( .A1(n14186), .A2(n13897), .ZN(n8026) );
  XNOR2_X1 U10331 ( .A(n8027), .B(n8028), .ZN(n11693) );
  NAND2_X1 U10332 ( .A1(n11693), .A2(n9675), .ZN(n8030) );
  INV_X1 U10333 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11691) );
  OR2_X1 U10334 ( .A1(n9677), .A2(n11691), .ZN(n8029) );
  NAND2_X1 U10335 ( .A1(n7757), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10336 ( .A1(n7988), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8035) );
  OAI21_X1 U10337 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8032), .A(n8031), .ZN(
        n14165) );
  OR2_X1 U10338 ( .A1(n8070), .A2(n14165), .ZN(n8034) );
  INV_X1 U10339 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15397) );
  OR2_X1 U10340 ( .A1(n8149), .A2(n15397), .ZN(n8033) );
  NAND4_X1 U10341 ( .A1(n8036), .A2(n8035), .A3(n8034), .A4(n8033), .ZN(n13896) );
  XNOR2_X1 U10342 ( .A(n14172), .B(n14141), .ZN(n14173) );
  INV_X1 U10343 ( .A(n14173), .ZN(n14161) );
  NAND2_X1 U10344 ( .A1(n8040), .A2(n8039), .ZN(n11827) );
  OR2_X1 U10345 ( .A1(n11827), .A2(n8064), .ZN(n8042) );
  INV_X1 U10346 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11828) );
  OR2_X1 U10347 ( .A1(n9677), .A2(n11828), .ZN(n8041) );
  NAND2_X2 U10348 ( .A1(n8042), .A2(n8041), .ZN(n14286) );
  NAND2_X1 U10349 ( .A1(n7757), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8048) );
  INV_X1 U10350 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15351) );
  OR2_X1 U10351 ( .A1(n9660), .A2(n15351), .ZN(n8047) );
  NAND2_X1 U10352 ( .A1(n6584), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8046) );
  OAI21_X1 U10353 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8043), .A(n8054), .ZN(
        n14152) );
  OR2_X1 U10354 ( .A1(n8044), .A2(n14152), .ZN(n8045) );
  NAND4_X1 U10355 ( .A1(n8048), .A2(n8047), .A3(n8046), .A4(n8045), .ZN(n13895) );
  INV_X1 U10356 ( .A(n13895), .ZN(n8132) );
  XNOR2_X1 U10357 ( .A(n14286), .B(n8132), .ZN(n14147) );
  XNOR2_X1 U10358 ( .A(n8050), .B(n8049), .ZN(n11931) );
  NAND2_X1 U10359 ( .A1(n11931), .A2(n9675), .ZN(n8052) );
  INV_X1 U10360 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11933) );
  OR2_X1 U10361 ( .A1(n9677), .A2(n11933), .ZN(n8051) );
  NAND2_X1 U10362 ( .A1(n7757), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10363 ( .A1(n7672), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10364 ( .A1(n7988), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8057) );
  INV_X1 U10365 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8053) );
  NAND2_X1 U10366 ( .A1(n8054), .A2(n8053), .ZN(n8055) );
  NAND2_X1 U10367 ( .A1(n8068), .A2(n8055), .ZN(n14130) );
  OR2_X1 U10368 ( .A1(n8070), .A2(n14130), .ZN(n8056) );
  NAND4_X1 U10369 ( .A1(n8059), .A2(n8058), .A3(n8057), .A4(n8056), .ZN(n13894) );
  XNOR2_X1 U10370 ( .A(n14135), .B(n14143), .ZN(n14125) );
  INV_X1 U10371 ( .A(n14125), .ZN(n14123) );
  NAND2_X1 U10372 ( .A1(n8060), .A2(n8061), .ZN(n8062) );
  OR2_X1 U10373 ( .A1(n9677), .A2(n14411), .ZN(n8065) );
  NAND2_X1 U10374 ( .A1(n7757), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10375 ( .A1(n6584), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10376 ( .A1(n7988), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8072) );
  INV_X1 U10377 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10378 ( .A1(n8068), .A2(n8067), .ZN(n8069) );
  NAND2_X1 U10379 ( .A1(n8082), .A2(n8069), .ZN(n14115) );
  OR2_X1 U10380 ( .A1(n8070), .A2(n14115), .ZN(n8071) );
  NAND4_X1 U10381 ( .A1(n8074), .A2(n8073), .A3(n8072), .A4(n8071), .ZN(n14093) );
  INV_X1 U10382 ( .A(n14093), .ZN(n12425) );
  NAND2_X1 U10383 ( .A1(n14270), .A2(n12425), .ZN(n8135) );
  OR2_X1 U10384 ( .A1(n14270), .A2(n12425), .ZN(n8075) );
  XNOR2_X1 U10385 ( .A(n8077), .B(SI_27_), .ZN(n8078) );
  NAND2_X1 U10386 ( .A1(n14406), .A2(n9675), .ZN(n8080) );
  INV_X1 U10387 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14409) );
  OR2_X1 U10388 ( .A1(n9677), .A2(n14409), .ZN(n8079) );
  NAND2_X1 U10389 ( .A1(n7757), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10390 ( .A1(n7988), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10391 ( .A1(n7672), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8086) );
  INV_X1 U10392 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10393 ( .A1(n8082), .A2(n8081), .ZN(n8083) );
  NAND2_X1 U10394 ( .A1(n8084), .A2(n8083), .ZN(n14102) );
  OR2_X1 U10395 ( .A1(n8070), .A2(n14102), .ZN(n8085) );
  NAND4_X1 U10396 ( .A1(n8088), .A2(n8087), .A3(n8086), .A4(n8085), .ZN(n13893) );
  INV_X1 U10397 ( .A(n13893), .ZN(n8136) );
  XNOR2_X1 U10398 ( .A(n14101), .B(n8136), .ZN(n14099) );
  OR2_X1 U10399 ( .A1(n14101), .A2(n13893), .ZN(n8089) );
  XNOR2_X1 U10400 ( .A(n7066), .B(n12457), .ZN(n9879) );
  NAND2_X1 U10401 ( .A1(n8143), .A2(n14040), .ZN(n9662) );
  NAND2_X1 U10402 ( .A1(n8093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10403 ( .A1(n8156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10404 ( .A1(n9662), .A2(n10259), .ZN(n10369) );
  INV_X4 U10405 ( .A(n8097), .ZN(n12459) );
  OR2_X1 U10406 ( .A1(n9662), .A2(n10259), .ZN(n8098) );
  NAND2_X1 U10407 ( .A1(n10513), .A2(n14040), .ZN(n10501) );
  INV_X1 U10408 ( .A(n8143), .ZN(n9682) );
  XNOR2_X1 U10409 ( .A(n14332), .B(n13900), .ZN(n14246) );
  NAND2_X1 U10410 ( .A1(n9686), .A2(n9690), .ZN(n9688) );
  NAND2_X1 U10411 ( .A1(n9688), .A2(n9691), .ZN(n10465) );
  NAND2_X1 U10412 ( .A1(n10464), .A2(n8099), .ZN(n10609) );
  NAND2_X1 U10413 ( .A1(n10609), .A2(n10608), .ZN(n10607) );
  NAND2_X1 U10414 ( .A1(n10896), .A2(n10892), .ZN(n8100) );
  NAND2_X1 U10415 ( .A1(n14736), .A2(n13913), .ZN(n8101) );
  NAND2_X1 U10416 ( .A1(n10522), .A2(n8101), .ZN(n8103) );
  NAND2_X1 U10417 ( .A1(n10905), .A2(n10929), .ZN(n8102) );
  NAND2_X1 U10418 ( .A1(n8103), .A2(n8102), .ZN(n10562) );
  NAND2_X1 U10419 ( .A1(n10562), .A2(n10561), .ZN(n8106) );
  NAND2_X1 U10420 ( .A1(n10914), .A2(n8104), .ZN(n8105) );
  NAND2_X1 U10421 ( .A1(n10696), .A2(n9865), .ZN(n8108) );
  INV_X1 U10422 ( .A(n13911), .ZN(n11034) );
  NAND2_X1 U10423 ( .A1(n11036), .A2(n11034), .ZN(n8107) );
  NAND2_X1 U10424 ( .A1(n8108), .A2(n8107), .ZN(n11052) );
  INV_X1 U10425 ( .A(n13910), .ZN(n11575) );
  AND2_X1 U10426 ( .A1(n14702), .A2(n11575), .ZN(n8110) );
  OR2_X1 U10427 ( .A1(n14702), .A2(n11575), .ZN(n8109) );
  INV_X1 U10428 ( .A(n13909), .ZN(n11721) );
  NAND2_X1 U10429 ( .A1(n11716), .A2(n11860), .ZN(n8111) );
  INV_X1 U10430 ( .A(n13907), .ZN(n12010) );
  OR2_X1 U10431 ( .A1(n11863), .A2(n12010), .ZN(n8112) );
  NAND2_X1 U10432 ( .A1(n11649), .A2(n11648), .ZN(n8114) );
  NAND2_X1 U10433 ( .A1(n14536), .A2(n13905), .ZN(n8113) );
  INV_X1 U10434 ( .A(n11630), .ZN(n8115) );
  NAND2_X1 U10435 ( .A1(n8116), .A2(n9764), .ZN(n11792) );
  INV_X1 U10436 ( .A(n9766), .ZN(n8117) );
  AOI21_X1 U10437 ( .B1(n11792), .B2(n8118), .A(n8117), .ZN(n11966) );
  OR2_X1 U10438 ( .A1(n14344), .A2(n13901), .ZN(n8119) );
  NAND2_X1 U10439 ( .A1(n9773), .A2(n8121), .ZN(n12017) );
  INV_X1 U10440 ( .A(n12017), .ZN(n12022) );
  NAND2_X1 U10441 ( .A1(n14338), .A2(n14235), .ZN(n8122) );
  INV_X1 U10442 ( .A(n13900), .ZN(n13812) );
  NOR2_X1 U10443 ( .A1(n14332), .A2(n13812), .ZN(n8123) );
  NAND2_X1 U10444 ( .A1(n14217), .A2(n14227), .ZN(n8125) );
  INV_X1 U10445 ( .A(n14237), .ZN(n13861) );
  NAND2_X1 U10446 ( .A1(n14325), .A2(n13861), .ZN(n8124) );
  INV_X1 U10447 ( .A(n13899), .ZN(n8126) );
  OR2_X1 U10448 ( .A1(n14315), .A2(n8126), .ZN(n8127) );
  INV_X1 U10449 ( .A(n13898), .ZN(n8128) );
  OR2_X1 U10450 ( .A1(n14384), .A2(n8128), .ZN(n8129) );
  INV_X1 U10451 ( .A(n13897), .ZN(n12381) );
  NAND2_X1 U10452 ( .A1(n14186), .A2(n12381), .ZN(n8130) );
  NAND2_X1 U10453 ( .A1(n6770), .A2(n14141), .ZN(n8131) );
  OR2_X1 U10454 ( .A1(n14286), .A2(n8132), .ZN(n8133) );
  NAND2_X1 U10455 ( .A1(n14135), .A2(n14143), .ZN(n8134) );
  INV_X1 U10456 ( .A(n14108), .ZN(n14112) );
  NAND2_X1 U10457 ( .A1(n7129), .A2(n14088), .ZN(n14091) );
  NAND2_X1 U10458 ( .A1(n14101), .A2(n8136), .ZN(n8137) );
  OAI21_X1 U10459 ( .B1(n12457), .B2(n7066), .A(n8204), .ZN(n8138) );
  OAI21_X1 U10460 ( .B1(n14081), .B2(n14092), .A(n8138), .ZN(n8139) );
  NAND2_X1 U10461 ( .A1(n8143), .A2(n10460), .ZN(n8141) );
  OR2_X1 U10462 ( .A1(n11644), .A2(n11532), .ZN(n8140) );
  INV_X1 U10463 ( .A(n14702), .ZN(n11249) );
  AND2_X1 U10464 ( .A1(n10771), .A2(n10631), .ZN(n10495) );
  NAND2_X1 U10465 ( .A1(n10495), .A2(n14716), .ZN(n10612) );
  OR2_X1 U10466 ( .A1(n10612), .A2(n10892), .ZN(n10613) );
  OR2_X2 U10467 ( .A1(n11346), .A2(n11716), .ZN(n11282) );
  OR2_X2 U10468 ( .A1(n11282), .A2(n11863), .ZN(n11440) );
  NAND2_X1 U10469 ( .A1(n14338), .A2(n12023), .ZN(n14240) );
  NAND2_X1 U10470 ( .A1(n14380), .A2(n14195), .ZN(n14181) );
  OR2_X2 U10471 ( .A1(n14168), .A2(n14286), .ZN(n14150) );
  NOR2_X2 U10472 ( .A1(n14150), .A2(n14135), .ZN(n14113) );
  INV_X1 U10473 ( .A(n8200), .ZN(n8145) );
  OAI211_X1 U10474 ( .C1(n7064), .C2(n8145), .A(n14254), .B(n8144), .ZN(n14071) );
  INV_X1 U10475 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10476 ( .A1(n7757), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10477 ( .A1(n7988), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8146) );
  OAI211_X1 U10478 ( .C1(n8149), .C2(n8148), .A(n8147), .B(n8146), .ZN(n13891)
         );
  NAND2_X1 U10479 ( .A1(n8143), .A2(n8150), .ZN(n9998) );
  INV_X1 U10480 ( .A(P1_B_REG_SCAN_IN), .ZN(n8168) );
  NOR2_X1 U10481 ( .A1(n6586), .A2(n8168), .ZN(n8151) );
  NOR2_X1 U10482 ( .A1(n14142), .A2(n8151), .ZN(n14049) );
  NAND2_X1 U10483 ( .A1(n13891), .A2(n14049), .ZN(n14062) );
  OR2_X1 U10484 ( .A1(n9998), .A2(n14401), .ZN(n14140) );
  NAND2_X1 U10485 ( .A1(n14092), .A2(n14234), .ZN(n14064) );
  INV_X1 U10486 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U10487 ( .A1(n8161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8162) );
  MUX2_X1 U10488 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8162), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8165) );
  NAND2_X1 U10489 ( .A1(n8165), .A2(n8164), .ZN(n11932) );
  NAND2_X1 U10490 ( .A1(n11932), .A2(P1_B_REG_SCAN_IN), .ZN(n8171) );
  NAND2_X1 U10491 ( .A1(n8164), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8167) );
  INV_X1 U10492 ( .A(n14414), .ZN(n8170) );
  NAND2_X1 U10493 ( .A1(n8190), .A2(n8168), .ZN(n8169) );
  NAND2_X1 U10494 ( .A1(n11932), .A2(n14414), .ZN(n9988) );
  OAI21_X1 U10495 ( .B1(n9987), .B2(P1_D_REG_1__SCAN_IN), .A(n9988), .ZN(
        n10454) );
  NAND2_X1 U10496 ( .A1(n14254), .A2(n10460), .ZN(n10270) );
  NAND2_X1 U10497 ( .A1(n10454), .A2(n10270), .ZN(n8189) );
  INV_X1 U10498 ( .A(n9987), .ZN(n8182) );
  NOR4_X1 U10499 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n8180) );
  NOR4_X1 U10500 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8179) );
  INV_X1 U10501 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15459) );
  INV_X1 U10502 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15450) );
  INV_X1 U10503 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15270) );
  INV_X1 U10504 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15311) );
  NAND4_X1 U10505 ( .A1(n15459), .A2(n15450), .A3(n15270), .A4(n15311), .ZN(
        n8177) );
  NOR4_X1 U10506 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n8175) );
  NOR4_X1 U10507 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n8174) );
  NOR4_X1 U10508 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8173) );
  NOR4_X1 U10509 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n8172) );
  NAND4_X1 U10510 ( .A1(n8175), .A2(n8174), .A3(n8173), .A4(n8172), .ZN(n8176)
         );
  NOR4_X1 U10511 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8177), .A4(n8176), .ZN(n8178) );
  NAND3_X1 U10512 ( .A1(n8180), .A2(n8179), .A3(n8178), .ZN(n8181) );
  NAND2_X1 U10513 ( .A1(n8182), .A2(n8181), .ZN(n10251) );
  AND2_X1 U10514 ( .A1(n11532), .A2(n14040), .ZN(n8184) );
  OR2_X1 U10515 ( .A1(n9998), .A2(n8184), .ZN(n10254) );
  NAND2_X1 U10516 ( .A1(n7538), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8186) );
  INV_X1 U10517 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8185) );
  AND2_X1 U10518 ( .A1(n10254), .A2(n10000), .ZN(n8187) );
  NAND2_X1 U10519 ( .A1(n10262), .A2(n8187), .ZN(n10272) );
  NOR2_X1 U10520 ( .A1(n10272), .A2(P1_U3086), .ZN(n8188) );
  NAND2_X1 U10521 ( .A1(n10251), .A2(n8188), .ZN(n10456) );
  OR2_X1 U10522 ( .A1(n8189), .A2(n10456), .ZN(n8197) );
  INV_X1 U10523 ( .A(n8190), .ZN(n11829) );
  NAND2_X1 U10524 ( .A1(n11829), .A2(n14414), .ZN(n10003) );
  OAI21_X1 U10525 ( .B1(n9987), .B2(P1_D_REG_0__SCAN_IN), .A(n10003), .ZN(
        n8196) );
  INV_X1 U10526 ( .A(n10401), .ZN(n8191) );
  NAND2_X1 U10527 ( .A1(n8191), .A2(n9685), .ZN(n10459) );
  NAND2_X1 U10528 ( .A1(n8191), .A2(n10460), .ZN(n8192) );
  NOR2_X1 U10529 ( .A1(n14759), .A2(n15369), .ZN(n8194) );
  OAI21_X1 U10530 ( .B1(n8199), .B2(n14757), .A(n8195), .ZN(P1_U3557) );
  INV_X1 U10531 ( .A(n8196), .ZN(n10455) );
  INV_X1 U10532 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8198) );
  OAI211_X1 U10533 ( .C1(n14081), .C2(n6617), .A(n14254), .B(n8200), .ZN(
        n14076) );
  NAND2_X1 U10534 ( .A1(n13892), .A2(n14236), .ZN(n8202) );
  NAND2_X1 U10535 ( .A1(n13893), .A2(n14234), .ZN(n8201) );
  AND2_X1 U10536 ( .A1(n8202), .A2(n8201), .ZN(n14078) );
  AND2_X1 U10537 ( .A1(n14076), .A2(n14078), .ZN(n8205) );
  XNOR2_X1 U10538 ( .A(n8204), .B(n8203), .ZN(n14084) );
  MUX2_X1 U10539 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n8210), .S(n14759), .Z(
        n8206) );
  INV_X1 U10540 ( .A(n8206), .ZN(n8209) );
  NAND2_X1 U10541 ( .A1(n7066), .A2(n8207), .ZN(n8208) );
  NAND2_X1 U10542 ( .A1(n8209), .A2(n8208), .ZN(P1_U3556) );
  MUX2_X1 U10543 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n8210), .S(n14752), .Z(
        n8211) );
  INV_X1 U10544 ( .A(n8211), .ZN(n8214) );
  NAND2_X1 U10545 ( .A1(n7066), .A2(n8212), .ZN(n8213) );
  NAND2_X1 U10546 ( .A1(n8214), .A2(n8213), .ZN(P1_U3524) );
  NAND4_X1 U10547 ( .A1(n8524), .A2(n8216), .A3(n8215), .A4(n8644), .ZN(n8722)
         );
  NAND2_X1 U10548 ( .A1(n8523), .A2(n8726), .ZN(n8217) );
  NOR2_X2 U10549 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8306) );
  INV_X1 U10550 ( .A(n8526), .ZN(n8228) );
  NAND2_X1 U10551 ( .A1(n8717), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8232) );
  INV_X1 U10552 ( .A(n8237), .ZN(n8233) );
  NAND2_X2 U10553 ( .A1(n6568), .A2(n9957), .ZN(n8274) );
  INV_X1 U10554 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13738) );
  OR2_X1 U10555 ( .A1(n8960), .A2(n13738), .ZN(n8235) );
  NOR2_X2 U10556 ( .A1(n8238), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n13723) );
  OR2_X2 U10557 ( .A1(n13723), .A2(n13724), .ZN(n8279) );
  AND2_X2 U10558 ( .A1(n12277), .A2(n8294), .ZN(n8339) );
  NAND2_X1 U10559 ( .A1(n8654), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8251) );
  INV_X1 U10560 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8240) );
  OR2_X1 U10561 ( .A1(n8657), .A2(n8240), .ZN(n8250) );
  AND2_X2 U10562 ( .A1(n8246), .A2(n8294), .ZN(n8571) );
  INV_X2 U10563 ( .A(n8571), .ZN(n8634) );
  NAND2_X1 U10564 ( .A1(n8335), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8365) );
  INV_X1 U10565 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8364) );
  NOR2_X1 U10566 ( .A1(n8365), .A2(n8364), .ZN(n8363) );
  AND2_X1 U10567 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n8241) );
  NAND2_X1 U10568 ( .A1(n8381), .A2(n8241), .ZN(n8423) );
  INV_X1 U10569 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n15402) );
  NAND2_X1 U10570 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n8242) );
  NAND2_X1 U10571 ( .A1(n8450), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8482) );
  INV_X1 U10572 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8481) );
  INV_X1 U10573 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8497) );
  INV_X1 U10574 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U10575 ( .A1(n8533), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8556) );
  INV_X1 U10576 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n15325) );
  INV_X1 U10577 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U10578 ( .A1(n8579), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8588) );
  INV_X1 U10579 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13295) );
  INV_X1 U10580 ( .A(n8622), .ZN(n8624) );
  INV_X1 U10581 ( .A(n8243), .ZN(n8614) );
  INV_X1 U10582 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10583 ( .A1(n8614), .A2(n8244), .ZN(n8245) );
  NAND2_X1 U10584 ( .A1(n8624), .A2(n8245), .ZN(n13460) );
  OR2_X1 U10585 ( .A1(n8634), .A2(n13460), .ZN(n8249) );
  INV_X1 U10586 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8247) );
  OR2_X1 U10587 ( .A1(n8931), .A2(n8247), .ZN(n8248) );
  XNOR2_X1 U10588 ( .A(n13228), .B(n13355), .ZN(n13466) );
  NAND2_X1 U10589 ( .A1(n11461), .A2(n8958), .ZN(n8256) );
  NOR2_X1 U10590 ( .A1(n8402), .A2(n8526), .ZN(n8475) );
  NAND2_X1 U10591 ( .A1(n8724), .A2(n8522), .ZN(n8505) );
  OAI21_X1 U10592 ( .B1(n8505), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8254) );
  INV_X1 U10593 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8253) );
  XNOR2_X1 U10594 ( .A(n8254), .B(n8253), .ZN(n14925) );
  INV_X1 U10595 ( .A(n14925), .ZN(n11756) );
  AOI22_X1 U10596 ( .A1(n8530), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n11756), 
        .B2(n8529), .ZN(n8255) );
  INV_X1 U10597 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8265) );
  INV_X1 U10598 ( .A(n8257), .ZN(n8535) );
  INV_X1 U10599 ( .A(n8258), .ZN(n8512) );
  INV_X1 U10600 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10601 ( .A1(n8512), .A2(n8259), .ZN(n8260) );
  NAND2_X1 U10602 ( .A1(n8535), .A2(n8260), .ZN(n13596) );
  OR2_X1 U10603 ( .A1(n13596), .A2(n8634), .ZN(n8264) );
  NAND2_X1 U10604 ( .A1(n6582), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8262) );
  INV_X1 U10605 ( .A(n8654), .ZN(n8513) );
  INV_X1 U10606 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14917) );
  OR2_X1 U10607 ( .A1(n8513), .A2(n14917), .ZN(n8261) );
  AND2_X1 U10608 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  OAI211_X1 U10609 ( .C1(n8931), .C2(n8265), .A(n8264), .B(n8263), .ZN(n13364)
         );
  NAND2_X1 U10610 ( .A1(n8339), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8267) );
  NAND2_X1 U10611 ( .A1(n8571), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8266) );
  NAND3_X2 U10612 ( .A1(n8269), .A2(n8270), .A3(n8268), .ZN(n9903) );
  NAND2_X1 U10613 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8271) );
  MUX2_X1 U10614 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8271), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8272) );
  INV_X1 U10615 ( .A(n8306), .ZN(n8304) );
  NAND2_X1 U10616 ( .A1(n8272), .A2(n8304), .ZN(n14771) );
  INV_X1 U10617 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8278) );
  XNOR2_X1 U10618 ( .A(n9069), .B(n8276), .ZN(n13743) );
  INV_X1 U10619 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8286) );
  AOI22_X1 U10620 ( .A1(n8286), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n8284) );
  INV_X1 U10621 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10622 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n8280) );
  OAI21_X1 U10623 ( .B1(n8281), .B2(P2_IR_REG_30__SCAN_IN), .A(n8280), .ZN(
        n8282) );
  NAND2_X1 U10624 ( .A1(n8291), .A2(n8282), .ZN(n8283) );
  OAI21_X1 U10625 ( .B1(n8291), .B2(n8284), .A(n8283), .ZN(n8285) );
  NAND2_X1 U10626 ( .A1(n8285), .A2(n13730), .ZN(n8297) );
  AOI22_X1 U10627 ( .A1(n8286), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n8287) );
  INV_X1 U10628 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10629 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .ZN(n8288) );
  OAI21_X1 U10630 ( .B1(n8289), .B2(P2_IR_REG_30__SCAN_IN), .A(n8288), .ZN(
        n8290) );
  NAND2_X1 U10631 ( .A1(n8293), .A2(n8292), .ZN(n8295) );
  NAND2_X1 U10632 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  NOR2_X1 U10633 ( .A1(n14969), .A2(n8750), .ZN(n10192) );
  NAND2_X1 U10634 ( .A1(n10191), .A2(n10192), .ZN(n10190) );
  INV_X1 U10635 ( .A(n10337), .ZN(n10584) );
  NAND2_X1 U10636 ( .A1(n10190), .A2(n8298), .ZN(n10233) );
  NAND2_X1 U10637 ( .A1(n8571), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U10638 ( .A1(n6583), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10639 ( .A1(n6580), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10640 ( .A1(n8339), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8300) );
  NAND4_X2 U10641 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n13381) );
  NOR2_X1 U10642 ( .A1(n9946), .A2(n8274), .ZN(n8309) );
  NAND2_X1 U10643 ( .A1(n8304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8305) );
  MUX2_X1 U10644 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8305), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8307) );
  NAND2_X1 U10645 ( .A1(n8306), .A2(n8223), .ZN(n8375) );
  NAND2_X1 U10646 ( .A1(n8307), .A2(n8375), .ZN(n13382) );
  OAI22_X1 U10647 ( .A1(n8960), .A2(n9940), .B1(n10017), .B2(n13382), .ZN(
        n8308) );
  INV_X1 U10648 ( .A(n10343), .ZN(n14952) );
  OR2_X1 U10649 ( .A1(n13381), .A2(n14952), .ZN(n8310) );
  NAND2_X1 U10650 ( .A1(n6583), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U10651 ( .A1(n6580), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U10652 ( .A1(n8339), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8311) );
  NAND4_X1 U10653 ( .A1(n8314), .A2(n8313), .A3(n8312), .A4(n8311), .ZN(n13380) );
  NAND2_X1 U10654 ( .A1(n9941), .A2(n8958), .ZN(n8318) );
  NAND2_X1 U10655 ( .A1(n8375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8315) );
  MUX2_X1 U10656 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8315), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8316) );
  AND2_X1 U10657 ( .A1(n8316), .A2(n8322), .ZN(n10106) );
  NAND2_X2 U10658 ( .A1(n8318), .A2(n8317), .ZN(n10340) );
  XNOR2_X1 U10659 ( .A(n13380), .B(n10340), .ZN(n9002) );
  NAND2_X1 U10660 ( .A1(n10307), .A2(n9002), .ZN(n8320) );
  INV_X1 U10661 ( .A(n13380), .ZN(n10357) );
  NAND2_X1 U10662 ( .A1(n10357), .A2(n10340), .ZN(n8319) );
  NAND2_X1 U10663 ( .A1(n9943), .A2(n8958), .ZN(n8327) );
  NAND2_X1 U10664 ( .A1(n8322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8321) );
  MUX2_X1 U10665 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8321), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8325) );
  INV_X1 U10666 ( .A(n8322), .ZN(n8324) );
  INV_X1 U10667 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10668 ( .A1(n8324), .A2(n8323), .ZN(n8346) );
  NAND2_X1 U10669 ( .A1(n8325), .A2(n8346), .ZN(n14783) );
  INV_X1 U10670 ( .A(n14783), .ZN(n10108) );
  AOI22_X1 U10671 ( .A1(n8530), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8529), .B2(
        n10108), .ZN(n8326) );
  NAND2_X2 U10672 ( .A1(n8327), .A2(n8326), .ZN(n10386) );
  NAND2_X1 U10673 ( .A1(n6582), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8331) );
  XNOR2_X1 U10674 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10570) );
  OR2_X1 U10675 ( .A1(n8634), .A2(n10570), .ZN(n8330) );
  NAND2_X1 U10676 ( .A1(n6579), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8329) );
  NAND2_X1 U10677 ( .A1(n8339), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8328) );
  INV_X1 U10678 ( .A(n13378), .ZN(n10429) );
  OR2_X1 U10679 ( .A1(n9953), .A2(n8274), .ZN(n8334) );
  NAND2_X1 U10680 ( .A1(n8346), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8332) );
  XNOR2_X1 U10681 ( .A(n8332), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U10682 ( .A1(n8530), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8529), .B2(
        n10111), .ZN(n8333) );
  NAND2_X1 U10683 ( .A1(n8334), .A2(n8333), .ZN(n10425) );
  NAND2_X1 U10684 ( .A1(n6583), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8343) );
  INV_X1 U10685 ( .A(n8335), .ZN(n8351) );
  INV_X1 U10686 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10687 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8336) );
  NAND2_X1 U10688 ( .A1(n8337), .A2(n8336), .ZN(n8338) );
  NAND2_X1 U10689 ( .A1(n8351), .A2(n8338), .ZN(n10427) );
  OR2_X1 U10690 ( .A1(n8634), .A2(n10427), .ZN(n8342) );
  NAND2_X1 U10691 ( .A1(n8654), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10692 ( .A1(n6580), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8340) );
  NAND4_X1 U10693 ( .A1(n8343), .A2(n8342), .A3(n8341), .A4(n8340), .ZN(n13377) );
  XNOR2_X1 U10694 ( .A(n10425), .B(n13377), .ZN(n10596) );
  INV_X1 U10695 ( .A(n13377), .ZN(n8670) );
  NAND2_X1 U10696 ( .A1(n10425), .A2(n8670), .ZN(n8344) );
  NAND2_X1 U10697 ( .A1(n8345), .A2(n8344), .ZN(n10542) );
  OR2_X1 U10698 ( .A1(n9979), .A2(n8274), .ZN(n8349) );
  NAND2_X1 U10699 ( .A1(n8359), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8347) );
  XNOR2_X1 U10700 ( .A(n8347), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U10701 ( .A1(n8530), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8529), .B2(
        n14801), .ZN(n8348) );
  NAND2_X1 U10702 ( .A1(n6583), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8356) );
  INV_X1 U10703 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10704 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U10705 ( .A1(n8365), .A2(n8352), .ZN(n10646) );
  OR2_X1 U10706 ( .A1(n8634), .A2(n10646), .ZN(n8355) );
  NAND2_X1 U10707 ( .A1(n8339), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10708 ( .A1(n6580), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8353) );
  NAND4_X1 U10709 ( .A1(n8356), .A2(n8355), .A3(n8354), .A4(n8353), .ZN(n13376) );
  INV_X1 U10710 ( .A(n13376), .ZN(n10428) );
  XNOR2_X1 U10711 ( .A(n14983), .B(n10428), .ZN(n10538) );
  INV_X1 U10712 ( .A(n10538), .ZN(n10541) );
  NAND2_X1 U10713 ( .A1(n10542), .A2(n10541), .ZN(n8358) );
  NAND2_X1 U10714 ( .A1(n14983), .A2(n10428), .ZN(n8357) );
  OR2_X1 U10715 ( .A1(n9985), .A2(n8274), .ZN(n8362) );
  OAI21_X1 U10716 ( .B1(n8359), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8360) );
  XNOR2_X1 U10717 ( .A(n8360), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U10718 ( .A1(n8530), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8529), .B2(
        n10115), .ZN(n8361) );
  NAND2_X1 U10719 ( .A1(n8362), .A2(n8361), .ZN(n10839) );
  NAND2_X1 U10720 ( .A1(n8654), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8370) );
  INV_X1 U10721 ( .A(n8363), .ZN(n8383) );
  NAND2_X1 U10722 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  NAND2_X1 U10723 ( .A1(n8383), .A2(n8366), .ZN(n15199) );
  OR2_X1 U10724 ( .A1(n8634), .A2(n15199), .ZN(n8369) );
  NAND2_X1 U10725 ( .A1(n6582), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10726 ( .A1(n6579), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8367) );
  NAND4_X1 U10727 ( .A1(n8370), .A2(n8369), .A3(n8368), .A4(n8367), .ZN(n13375) );
  INV_X1 U10728 ( .A(n13375), .ZN(n10722) );
  AND2_X1 U10729 ( .A1(n10839), .A2(n10722), .ZN(n8371) );
  OR2_X1 U10730 ( .A1(n10839), .A2(n10722), .ZN(n8372) );
  OR2_X1 U10731 ( .A1(n9993), .A2(n8274), .ZN(n8380) );
  INV_X1 U10732 ( .A(n8373), .ZN(n8374) );
  NOR2_X1 U10733 ( .A1(n8374), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8377) );
  INV_X1 U10734 ( .A(n8375), .ZN(n8376) );
  NAND2_X1 U10735 ( .A1(n8377), .A2(n8376), .ZN(n8391) );
  NAND2_X1 U10736 ( .A1(n8391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8378) );
  XNOR2_X1 U10737 ( .A(n8378), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U10738 ( .A1(n8530), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8529), .B2(
        n10138), .ZN(n8379) );
  NAND2_X1 U10739 ( .A1(n8654), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8388) );
  INV_X1 U10740 ( .A(n8381), .ZN(n8408) );
  INV_X1 U10741 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10742 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  NAND2_X1 U10743 ( .A1(n8408), .A2(n8384), .ZN(n10742) );
  OR2_X1 U10744 ( .A1(n8634), .A2(n10742), .ZN(n8387) );
  NAND2_X1 U10745 ( .A1(n6582), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10746 ( .A1(n6579), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8385) );
  NAND4_X1 U10747 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(n13374) );
  XNOR2_X1 U10748 ( .A(n15003), .B(n13374), .ZN(n10728) );
  INV_X1 U10749 ( .A(n10728), .ZN(n10732) );
  INV_X1 U10750 ( .A(n13374), .ZN(n8389) );
  NAND2_X1 U10751 ( .A1(n15003), .A2(n8389), .ZN(n8390) );
  NAND2_X1 U10752 ( .A1(n10735), .A2(n8390), .ZN(n10847) );
  OR2_X1 U10753 ( .A1(n10012), .A2(n8274), .ZN(n8395) );
  OAI21_X1 U10754 ( .B1(n8391), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8392) );
  MUX2_X1 U10755 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8392), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8393) );
  AND2_X1 U10756 ( .A1(n8393), .A2(n8402), .ZN(n10141) );
  AOI22_X1 U10757 ( .A1(n8530), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8529), .B2(
        n10141), .ZN(n8394) );
  INV_X1 U10758 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10277) );
  OR2_X1 U10759 ( .A1(n8513), .A2(n10277), .ZN(n8399) );
  INV_X1 U10760 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8407) );
  XNOR2_X1 U10761 ( .A(n8408), .B(n8407), .ZN(n10879) );
  OR2_X1 U10762 ( .A1(n8634), .A2(n10879), .ZN(n8398) );
  INV_X1 U10763 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10854) );
  OR2_X1 U10764 ( .A1(n8931), .A2(n10854), .ZN(n8397) );
  NAND2_X1 U10765 ( .A1(n6582), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8396) );
  NAND4_X1 U10766 ( .A1(n8399), .A2(n8398), .A3(n8397), .A4(n8396), .ZN(n13373) );
  NAND2_X1 U10767 ( .A1(n10951), .A2(n13373), .ZN(n8675) );
  OR2_X1 U10768 ( .A1(n10951), .A2(n13373), .ZN(n8400) );
  NAND2_X1 U10769 ( .A1(n8675), .A2(n8400), .ZN(n10846) );
  INV_X1 U10770 ( .A(n13373), .ZN(n11004) );
  NAND2_X1 U10771 ( .A1(n10951), .A2(n11004), .ZN(n8401) );
  NAND2_X1 U10772 ( .A1(n10149), .A2(n8958), .ZN(n8405) );
  NAND2_X1 U10773 ( .A1(n8402), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8403) );
  XNOR2_X1 U10774 ( .A(n8403), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U10775 ( .A1(n8530), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8529), 
        .B2(n10289), .ZN(n8404) );
  NAND2_X2 U10776 ( .A1(n8405), .A2(n8404), .ZN(n11235) );
  NAND2_X1 U10777 ( .A1(n8654), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8413) );
  INV_X1 U10778 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8406) );
  OAI21_X1 U10779 ( .B1(n8408), .B2(n8407), .A(n8406), .ZN(n8409) );
  NAND2_X1 U10780 ( .A1(n8409), .A2(n8423), .ZN(n11228) );
  OR2_X1 U10781 ( .A1(n8634), .A2(n11228), .ZN(n8412) );
  NAND2_X1 U10782 ( .A1(n6583), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U10783 ( .A1(n6580), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8410) );
  NAND4_X1 U10784 ( .A1(n8413), .A2(n8412), .A3(n8411), .A4(n8410), .ZN(n13372) );
  INV_X1 U10785 ( .A(n13372), .ZN(n11192) );
  OR2_X1 U10786 ( .A1(n11235), .A2(n11192), .ZN(n8414) );
  NAND2_X1 U10787 ( .A1(n11002), .A2(n8414), .ZN(n8416) );
  NAND2_X1 U10788 ( .A1(n11235), .A2(n11192), .ZN(n8415) );
  NAND2_X1 U10789 ( .A1(n10220), .A2(n8958), .ZN(n8422) );
  NAND2_X1 U10790 ( .A1(n8252), .A2(n8417), .ZN(n8419) );
  NAND2_X1 U10791 ( .A1(n8419), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8418) );
  MUX2_X1 U10792 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8418), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n8420) );
  AND2_X1 U10793 ( .A1(n8420), .A2(n8433), .ZN(n10291) );
  AOI22_X1 U10794 ( .A1(n8530), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8529), 
        .B2(n10291), .ZN(n8421) );
  NAND2_X1 U10795 ( .A1(n8654), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10796 ( .A1(n8423), .A2(n15402), .ZN(n8424) );
  NAND2_X1 U10797 ( .A1(n8449), .A2(n8424), .ZN(n14935) );
  OR2_X1 U10798 ( .A1(n8634), .A2(n14935), .ZN(n8427) );
  NAND2_X1 U10799 ( .A1(n6582), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U10800 ( .A1(n6579), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8425) );
  NAND4_X1 U10801 ( .A1(n8428), .A2(n8427), .A3(n8426), .A4(n8425), .ZN(n13371) );
  INV_X1 U10802 ( .A(n13371), .ZN(n11003) );
  XNOR2_X1 U10803 ( .A(n14938), .B(n11003), .ZN(n9008) );
  NAND2_X1 U10804 ( .A1(n14932), .A2(n14939), .ZN(n8430) );
  NAND2_X1 U10805 ( .A1(n14938), .A2(n11003), .ZN(n8429) );
  NAND2_X1 U10806 ( .A1(n10247), .A2(n8958), .ZN(n8436) );
  NAND2_X1 U10807 ( .A1(n8433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8431) );
  MUX2_X1 U10808 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8431), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8432) );
  INV_X1 U10809 ( .A(n8432), .ZN(n8434) );
  NOR2_X1 U10810 ( .A1(n8433), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8443) );
  NOR2_X1 U10811 ( .A1(n8434), .A2(n8443), .ZN(n10296) );
  AOI22_X1 U10812 ( .A1(n8530), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8529), 
        .B2(n10296), .ZN(n8435) );
  INV_X1 U10813 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11760) );
  OR2_X1 U10814 ( .A1(n8513), .A2(n11760), .ZN(n8440) );
  INV_X1 U10815 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8448) );
  XNOR2_X1 U10816 ( .A(n8449), .B(n8448), .ZN(n11426) );
  OR2_X1 U10817 ( .A1(n8634), .A2(n11426), .ZN(n8439) );
  INV_X1 U10818 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11742) );
  OR2_X1 U10819 ( .A1(n8931), .A2(n11742), .ZN(n8438) );
  NAND2_X1 U10820 ( .A1(n6582), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8437) );
  NAND4_X1 U10821 ( .A1(n8440), .A2(n8439), .A3(n8438), .A4(n8437), .ZN(n13370) );
  AND2_X1 U10822 ( .A1(n11431), .A2(n11191), .ZN(n8441) );
  OR2_X1 U10823 ( .A1(n11431), .A2(n11191), .ZN(n8442) );
  NAND2_X1 U10824 ( .A1(n10397), .A2(n8958), .ZN(n8446) );
  INV_X1 U10825 ( .A(n8443), .ZN(n8461) );
  NAND2_X1 U10826 ( .A1(n8461), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8444) );
  XNOR2_X1 U10827 ( .A(n8444), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U10828 ( .A1(n8530), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8529), 
        .B2(n11765), .ZN(n8445) );
  INV_X1 U10829 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8447) );
  OAI21_X1 U10830 ( .B1(n8449), .B2(n8448), .A(n8447), .ZN(n8451) );
  INV_X1 U10831 ( .A(n8450), .ZN(n8466) );
  NAND2_X1 U10832 ( .A1(n8451), .A2(n8466), .ZN(n11449) );
  OR2_X1 U10833 ( .A1(n8634), .A2(n11449), .ZN(n8455) );
  NAND2_X1 U10834 ( .A1(n6583), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10835 ( .A1(n6580), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10836 ( .A1(n8654), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8452) );
  NAND4_X1 U10837 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n13369) );
  INV_X1 U10838 ( .A(n13369), .ZN(n8456) );
  NAND2_X1 U10839 ( .A1(n14598), .A2(n8456), .ZN(n8460) );
  OR2_X1 U10840 ( .A1(n14598), .A2(n8456), .ZN(n8457) );
  NAND2_X1 U10841 ( .A1(n8460), .A2(n8457), .ZN(n11399) );
  NAND2_X1 U10842 ( .A1(n10589), .A2(n8958), .ZN(n8464) );
  OAI21_X1 U10843 ( .B1(n8461), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10844 ( .A(n8462), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U10845 ( .A1(n8530), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8529), 
        .B2(n11767), .ZN(n8463) );
  NAND2_X1 U10846 ( .A1(n6582), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8471) );
  INV_X1 U10847 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8465) );
  NAND2_X1 U10848 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  NAND2_X1 U10849 ( .A1(n8482), .A2(n8467), .ZN(n14580) );
  OR2_X1 U10850 ( .A1(n8634), .A2(n14580), .ZN(n8470) );
  NAND2_X1 U10851 ( .A1(n6580), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10852 ( .A1(n8654), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8468) );
  NAND4_X1 U10853 ( .A1(n8471), .A2(n8470), .A3(n8469), .A4(n8468), .ZN(n13368) );
  INV_X1 U10854 ( .A(n13368), .ZN(n8684) );
  OR2_X1 U10855 ( .A1(n14589), .A2(n8684), .ZN(n8472) );
  NAND2_X1 U10856 ( .A1(n11580), .A2(n8472), .ZN(n8474) );
  NAND2_X1 U10857 ( .A1(n14589), .A2(n8684), .ZN(n8473) );
  NAND2_X1 U10858 ( .A1(n10841), .A2(n8958), .ZN(n8480) );
  INV_X1 U10859 ( .A(n8475), .ZN(n8476) );
  NAND2_X1 U10860 ( .A1(n8476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8477) );
  MUX2_X1 U10861 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8477), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n8478) );
  INV_X1 U10862 ( .A(n8724), .ZN(n8490) );
  AND2_X1 U10863 ( .A1(n8478), .A2(n8490), .ZN(n11770) );
  AOI22_X1 U10864 ( .A1(n8530), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8529), 
        .B2(n11770), .ZN(n8479) );
  NAND2_X1 U10865 ( .A1(n6583), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U10866 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NAND2_X1 U10867 ( .A1(n8498), .A2(n8483), .ZN(n11681) );
  OR2_X1 U10868 ( .A1(n8634), .A2(n11681), .ZN(n8486) );
  NAND2_X1 U10869 ( .A1(n8654), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10870 ( .A1(n6579), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8484) );
  NAND4_X1 U10871 ( .A1(n8487), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(n13367) );
  INV_X1 U10872 ( .A(n13367), .ZN(n11801) );
  AND2_X1 U10873 ( .A1(n11878), .A2(n11801), .ZN(n8488) );
  OR2_X1 U10874 ( .A1(n11878), .A2(n11801), .ZN(n8489) );
  NAND2_X1 U10875 ( .A1(n10940), .A2(n8958), .ZN(n8496) );
  NAND2_X1 U10876 ( .A1(n8490), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8491) );
  MUX2_X1 U10877 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8491), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8492) );
  INV_X1 U10878 ( .A(n8492), .ZN(n8494) );
  INV_X1 U10879 ( .A(n8505), .ZN(n8493) );
  NOR2_X1 U10880 ( .A1(n8494), .A2(n8493), .ZN(n14893) );
  AOI22_X1 U10881 ( .A1(n8530), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8529), 
        .B2(n14893), .ZN(n8495) );
  NAND2_X1 U10882 ( .A1(n8498), .A2(n8497), .ZN(n8499) );
  NAND2_X1 U10883 ( .A1(n8510), .A2(n8499), .ZN(n11947) );
  OR2_X1 U10884 ( .A1(n8634), .A2(n11947), .ZN(n8503) );
  NAND2_X1 U10885 ( .A1(n8654), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U10886 ( .A1(n6583), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10887 ( .A1(n6579), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8500) );
  NAND4_X1 U10888 ( .A1(n8503), .A2(n8502), .A3(n8501), .A4(n8500), .ZN(n13366) );
  INV_X1 U10889 ( .A(n13366), .ZN(n11952) );
  XNOR2_X1 U10890 ( .A(n13687), .B(n11952), .ZN(n11810) );
  NAND2_X1 U10891 ( .A1(n13687), .A2(n11952), .ZN(n8504) );
  NAND2_X1 U10892 ( .A1(n11079), .A2(n8958), .ZN(n8508) );
  NAND2_X1 U10893 ( .A1(n8505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8506) );
  XNOR2_X1 U10894 ( .A(n8506), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U10895 ( .A1(n8530), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8529), 
        .B2(n11773), .ZN(n8507) );
  NAND2_X1 U10896 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U10897 ( .A1(n8512), .A2(n8511), .ZN(n12039) );
  OR2_X1 U10898 ( .A1(n12039), .A2(n8634), .ZN(n8517) );
  INV_X1 U10899 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n15357) );
  OR2_X1 U10900 ( .A1(n8513), .A2(n15357), .ZN(n8516) );
  NAND2_X1 U10901 ( .A1(n6583), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10902 ( .A1(n6580), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8514) );
  NAND4_X1 U10903 ( .A1(n8517), .A2(n8516), .A3(n8515), .A4(n8514), .ZN(n13365) );
  INV_X1 U10904 ( .A(n13365), .ZN(n13328) );
  OR2_X1 U10905 ( .A1(n13679), .A2(n13328), .ZN(n8518) );
  NAND2_X1 U10906 ( .A1(n11951), .A2(n8518), .ZN(n8520) );
  NAND2_X1 U10907 ( .A1(n13679), .A2(n13328), .ZN(n8519) );
  INV_X1 U10908 ( .A(n13364), .ZN(n13247) );
  NAND2_X1 U10909 ( .A1(n13674), .A2(n13247), .ZN(n8521) );
  NAND2_X1 U10910 ( .A1(n11517), .A2(n8958), .ZN(n8532) );
  NAND3_X1 U10911 ( .A1(n8524), .A2(n8523), .A3(n8522), .ZN(n8525) );
  NOR2_X1 U10912 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  NAND2_X1 U10913 ( .A1(n8641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8528) );
  AOI22_X1 U10914 ( .A1(n8530), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11409), 
        .B2(n8529), .ZN(n8531) );
  INV_X1 U10915 ( .A(n8533), .ZN(n8544) );
  INV_X1 U10916 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U10917 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  NAND2_X1 U10918 ( .A1(n8544), .A2(n8536), .ZN(n13584) );
  AOI22_X1 U10919 ( .A1(n6582), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n8654), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10920 ( .A1(n6579), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8537) );
  OAI211_X1 U10921 ( .C1(n13584), .C2(n8634), .A(n8538), .B(n8537), .ZN(n13363) );
  INV_X1 U10922 ( .A(n13363), .ZN(n13329) );
  AND2_X1 U10923 ( .A1(n13583), .A2(n13329), .ZN(n8539) );
  OR2_X1 U10924 ( .A1(n13583), .A2(n13329), .ZN(n8540) );
  OR2_X1 U10925 ( .A1(n8960), .A2(n11529), .ZN(n8541) );
  NAND2_X2 U10926 ( .A1(n8542), .A2(n8541), .ZN(n13713) );
  INV_X1 U10927 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U10928 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  NAND2_X1 U10929 ( .A1(n8556), .A2(n8545), .ZN(n13560) );
  OR2_X1 U10930 ( .A1(n13560), .A2(n8634), .ZN(n8551) );
  INV_X1 U10931 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10932 ( .A1(n8654), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10933 ( .A1(n6579), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8546) );
  OAI211_X1 U10934 ( .C1(n8657), .C2(n8548), .A(n8547), .B(n8546), .ZN(n8549)
         );
  INV_X1 U10935 ( .A(n8549), .ZN(n8550) );
  NAND2_X1 U10936 ( .A1(n8551), .A2(n8550), .ZN(n13362) );
  INV_X1 U10937 ( .A(n13362), .ZN(n13273) );
  NAND2_X1 U10938 ( .A1(n13713), .A2(n13273), .ZN(n8553) );
  OR2_X1 U10939 ( .A1(n13713), .A2(n13273), .ZN(n8552) );
  NAND2_X1 U10940 ( .A1(n8553), .A2(n8552), .ZN(n13564) );
  INV_X1 U10941 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11558) );
  OR2_X1 U10942 ( .A1(n8960), .A2(n11558), .ZN(n8554) );
  NAND2_X1 U10943 ( .A1(n8556), .A2(n15325), .ZN(n8557) );
  AND2_X1 U10944 ( .A1(n8570), .A2(n8557), .ZN(n13548) );
  NAND2_X1 U10945 ( .A1(n13548), .A2(n8571), .ZN(n8563) );
  INV_X1 U10946 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10947 ( .A1(n8654), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10948 ( .A1(n6580), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8558) );
  OAI211_X1 U10949 ( .C1(n8657), .C2(n8560), .A(n8559), .B(n8558), .ZN(n8561)
         );
  INV_X1 U10950 ( .A(n8561), .ZN(n8562) );
  NAND2_X1 U10951 ( .A1(n8563), .A2(n8562), .ZN(n13361) );
  INV_X1 U10952 ( .A(n13361), .ZN(n8885) );
  OR2_X1 U10953 ( .A1(n13657), .A2(n8885), .ZN(n8999) );
  NAND2_X1 U10954 ( .A1(n13657), .A2(n8885), .ZN(n8998) );
  OR2_X1 U10955 ( .A1(n8014), .A2(n8565), .ZN(n8566) );
  NAND2_X1 U10956 ( .A1(n8567), .A2(n8566), .ZN(n11616) );
  INV_X1 U10957 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11617) );
  OR2_X1 U10958 ( .A1(n8960), .A2(n11617), .ZN(n8568) );
  AOI21_X1 U10959 ( .B1(n8570), .B2(n13317), .A(n8579), .ZN(n13538) );
  NAND2_X1 U10960 ( .A1(n13538), .A2(n8571), .ZN(n8576) );
  INV_X1 U10961 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n15354) );
  NAND2_X1 U10962 ( .A1(n8654), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U10963 ( .A1(n6580), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8572) );
  OAI211_X1 U10964 ( .C1(n8657), .C2(n15354), .A(n8573), .B(n8572), .ZN(n8574)
         );
  INV_X1 U10965 ( .A(n8574), .ZN(n8575) );
  NAND2_X1 U10966 ( .A1(n8576), .A2(n8575), .ZN(n13360) );
  NAND2_X1 U10967 ( .A1(n11693), .A2(n8958), .ZN(n8578) );
  INV_X1 U10968 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11697) );
  OR2_X1 U10969 ( .A1(n8960), .A2(n11697), .ZN(n8577) );
  NAND2_X1 U10970 ( .A1(n8654), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8583) );
  OAI21_X1 U10971 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8579), .A(n8588), .ZN(
        n13238) );
  OR2_X1 U10972 ( .A1(n8634), .A2(n13238), .ZN(n8582) );
  NAND2_X1 U10973 ( .A1(n6582), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10974 ( .A1(n6579), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8580) );
  NAND4_X1 U10975 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n13359) );
  INV_X1 U10976 ( .A(n13359), .ZN(n8584) );
  NAND2_X1 U10977 ( .A1(n13647), .A2(n8584), .ZN(n13500) );
  OR2_X1 U10978 ( .A1(n13647), .A2(n8584), .ZN(n8585) );
  OR2_X1 U10979 ( .A1(n11827), .A2(n8274), .ZN(n8587) );
  INV_X1 U10980 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11795) );
  OR2_X1 U10981 ( .A1(n8960), .A2(n11795), .ZN(n8586) );
  NAND2_X1 U10982 ( .A1(n8654), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8595) );
  INV_X1 U10983 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13703) );
  OR2_X1 U10984 ( .A1(n8657), .A2(n13703), .ZN(n8594) );
  INV_X1 U10985 ( .A(n8588), .ZN(n8590) );
  INV_X1 U10986 ( .A(n8610), .ZN(n8589) );
  OAI21_X1 U10987 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8590), .A(n8589), .ZN(
        n13294) );
  OR2_X1 U10988 ( .A1(n8634), .A2(n13294), .ZN(n8593) );
  INV_X1 U10989 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8591) );
  OR2_X1 U10990 ( .A1(n8931), .A2(n8591), .ZN(n8592) );
  NAND2_X1 U10991 ( .A1(n8905), .A2(n13358), .ZN(n8699) );
  OR2_X1 U10992 ( .A1(n8905), .A2(n13358), .ZN(n8596) );
  NAND2_X1 U10993 ( .A1(n8699), .A2(n8596), .ZN(n13499) );
  NAND2_X1 U10994 ( .A1(n8597), .A2(n13499), .ZN(n13503) );
  OR2_X1 U10995 ( .A1(n13705), .A2(n13358), .ZN(n8598) );
  NAND2_X1 U10996 ( .A1(n11931), .A2(n8958), .ZN(n8600) );
  INV_X1 U10997 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11936) );
  OR2_X1 U10998 ( .A1(n8960), .A2(n11936), .ZN(n8599) );
  NAND2_X1 U10999 ( .A1(n8654), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8606) );
  INV_X1 U11000 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8601) );
  OR2_X1 U11001 ( .A1(n8657), .A2(n8601), .ZN(n8605) );
  XNOR2_X1 U11002 ( .A(P2_REG3_REG_25__SCAN_IN), .B(n8610), .ZN(n13287) );
  OR2_X1 U11003 ( .A1(n8634), .A2(n13287), .ZN(n8604) );
  INV_X1 U11004 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8602) );
  OR2_X1 U11005 ( .A1(n8931), .A2(n8602), .ZN(n8603) );
  OR2_X1 U11006 ( .A1(n13487), .A2(n13357), .ZN(n8607) );
  OR2_X1 U11007 ( .A1(n8960), .A2(n13740), .ZN(n8608) );
  NAND2_X1 U11008 ( .A1(n8654), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8618) );
  INV_X1 U11009 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U11010 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(n8610), .ZN(n8611) );
  NAND2_X1 U11011 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  NAND2_X1 U11012 ( .A1(n8614), .A2(n8613), .ZN(n13473) );
  OR2_X1 U11013 ( .A1(n8634), .A2(n13473), .ZN(n8617) );
  NAND2_X1 U11014 ( .A1(n6583), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U11015 ( .A1(n6580), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8615) );
  NAND4_X1 U11016 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), .ZN(n13356) );
  INV_X1 U11017 ( .A(n13356), .ZN(n8997) );
  OR2_X1 U11018 ( .A1(n13630), .A2(n8997), .ZN(n8619) );
  NAND2_X1 U11019 ( .A1(n13733), .A2(n8958), .ZN(n8621) );
  INV_X1 U11020 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9524) );
  OR2_X1 U11021 ( .A1(n8960), .A2(n9524), .ZN(n8620) );
  NAND2_X1 U11022 ( .A1(n6582), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11023 ( .A1(n8622), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13432) );
  INV_X1 U11024 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U11025 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  NAND2_X1 U11026 ( .A1(n13432), .A2(n8625), .ZN(n13449) );
  OR2_X1 U11027 ( .A1(n8634), .A2(n13449), .ZN(n8628) );
  NAND2_X1 U11028 ( .A1(n8654), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11029 ( .A1(n6579), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8626) );
  NAND4_X1 U11030 ( .A1(n8629), .A2(n8628), .A3(n8627), .A4(n8626), .ZN(n13354) );
  NAND2_X1 U11031 ( .A1(n13617), .A2(n13354), .ZN(n8704) );
  OR2_X1 U11032 ( .A1(n13617), .A2(n13354), .ZN(n8630) );
  NAND2_X1 U11033 ( .A1(n8704), .A2(n8630), .ZN(n9020) );
  NAND2_X1 U11034 ( .A1(n13439), .A2(n9020), .ZN(n13442) );
  INV_X1 U11035 ( .A(n13354), .ZN(n8652) );
  NAND2_X1 U11036 ( .A1(n13728), .A2(n8958), .ZN(n8633) );
  OR2_X1 U11037 ( .A1(n8960), .A2(n13732), .ZN(n8632) );
  NAND2_X1 U11038 ( .A1(n6583), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8638) );
  OR2_X1 U11039 ( .A1(n8634), .A2(n13432), .ZN(n8637) );
  NAND2_X1 U11040 ( .A1(n8654), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U11041 ( .A1(n6580), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8635) );
  NAND4_X1 U11042 ( .A1(n8638), .A2(n8637), .A3(n8636), .A4(n8635), .ZN(n13353) );
  INV_X1 U11043 ( .A(n13353), .ZN(n8639) );
  INV_X1 U11044 ( .A(n8641), .ZN(n8643) );
  INV_X1 U11045 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11046 ( .A1(n8643), .A2(n8642), .ZN(n8649) );
  OAI21_X2 U11047 ( .B1(n8649), .B2(P2_IR_REG_20__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U11048 ( .A1(n8646), .A2(n8645), .ZN(n8648) );
  NAND2_X1 U11049 ( .A1(n9036), .A2(n11409), .ZN(n8932) );
  NAND2_X1 U11050 ( .A1(n8649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11051 ( .A1(n9029), .A2(n9024), .ZN(n8651) );
  NAND2_X1 U11052 ( .A1(n9036), .A2(n9029), .ZN(n10019) );
  CLKBUF_X1 U11053 ( .A(n8653), .Z(n10026) );
  INV_X1 U11054 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13696) );
  NAND2_X1 U11055 ( .A1(n6579), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11056 ( .A1(n8654), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8655) );
  OAI211_X1 U11057 ( .C1(n8657), .C2(n13696), .A(n8656), .B(n8655), .ZN(n13352) );
  INV_X1 U11058 ( .A(n13352), .ZN(n8996) );
  INV_X1 U11059 ( .A(n10026), .ZN(n8658) );
  INV_X1 U11060 ( .A(n8659), .ZN(n10023) );
  NAND2_X1 U11061 ( .A1(n10023), .A2(P2_B_REG_SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11062 ( .A1(n13315), .A2(n8660), .ZN(n13419) );
  NOR2_X1 U11063 ( .A1(n8996), .A2(n13419), .ZN(n8661) );
  INV_X1 U11064 ( .A(n13679), .ZN(n11962) );
  INV_X1 U11065 ( .A(n14938), .ZN(n15019) );
  INV_X1 U11066 ( .A(n10839), .ZN(n15201) );
  NAND2_X1 U11067 ( .A1(n10584), .A2(n14969), .ZN(n10231) );
  INV_X1 U11068 ( .A(n10386), .ZN(n10574) );
  AND2_X1 U11069 ( .A1(n10384), .A2(n10574), .ZN(n10599) );
  INV_X1 U11070 ( .A(n10425), .ZN(n14978) );
  OR2_X1 U11071 ( .A1(n10852), .A2(n10951), .ZN(n10851) );
  NOR2_X1 U11072 ( .A1(n11235), .A2(n10851), .ZN(n14942) );
  NOR2_X1 U11073 ( .A1(n13687), .A2(n11803), .ZN(n11957) );
  NAND2_X1 U11074 ( .A1(n11962), .A2(n11957), .ZN(n13595) );
  NAND2_X1 U11075 ( .A1(n6585), .A2(n11557), .ZN(n14968) );
  OR2_X2 U11076 ( .A1(n14968), .A2(n9024), .ZN(n13574) );
  INV_X1 U11077 ( .A(n14969), .ZN(n10241) );
  NAND2_X1 U11078 ( .A1(n10241), .A2(n8750), .ZN(n10329) );
  INV_X1 U11079 ( .A(n10329), .ZN(n10186) );
  OR2_X1 U11080 ( .A1(n9903), .A2(n10337), .ZN(n8665) );
  INV_X1 U11081 ( .A(n10232), .ZN(n10228) );
  NAND2_X1 U11082 ( .A1(n10229), .A2(n10228), .ZN(n10227) );
  OR2_X1 U11083 ( .A1(n13381), .A2(n10343), .ZN(n8666) );
  NAND2_X1 U11084 ( .A1(n10227), .A2(n8666), .ZN(n10303) );
  INV_X1 U11085 ( .A(n9002), .ZN(n10306) );
  NAND2_X1 U11086 ( .A1(n10303), .A2(n10306), .ZN(n10302) );
  NAND2_X1 U11087 ( .A1(n10357), .A2(n7193), .ZN(n8667) );
  NAND2_X1 U11088 ( .A1(n10302), .A2(n8667), .ZN(n10383) );
  OR2_X1 U11089 ( .A1(n10386), .A2(n13378), .ZN(n8668) );
  NAND2_X1 U11090 ( .A1(n10425), .A2(n13377), .ZN(n8669) );
  NAND2_X1 U11091 ( .A1(n10539), .A2(n10538), .ZN(n8672) );
  OR2_X1 U11092 ( .A1(n14983), .A2(n13376), .ZN(n8671) );
  NAND2_X1 U11093 ( .A1(n8672), .A2(n8671), .ZN(n15000) );
  XNOR2_X1 U11094 ( .A(n10839), .B(n13375), .ZN(n14990) );
  INV_X1 U11095 ( .A(n14990), .ZN(n14999) );
  OR2_X1 U11096 ( .A1(n10839), .A2(n13375), .ZN(n8673) );
  NAND2_X1 U11097 ( .A1(n15003), .A2(n13374), .ZN(n8674) );
  NAND2_X1 U11098 ( .A1(n10731), .A2(n8674), .ZN(n10859) );
  INV_X1 U11099 ( .A(n10846), .ZN(n10858) );
  NAND2_X1 U11100 ( .A1(n10859), .A2(n10858), .ZN(n10857) );
  OR2_X1 U11101 ( .A1(n11235), .A2(n13372), .ZN(n8676) );
  NAND2_X1 U11102 ( .A1(n11007), .A2(n8676), .ZN(n8678) );
  NAND2_X1 U11103 ( .A1(n11235), .A2(n13372), .ZN(n8677) );
  NAND2_X1 U11104 ( .A1(n8678), .A2(n8677), .ZN(n14940) );
  AND2_X1 U11105 ( .A1(n14938), .A2(n13371), .ZN(n8679) );
  OR2_X1 U11106 ( .A1(n14938), .A2(n13371), .ZN(n8680) );
  NOR2_X1 U11107 ( .A1(n11431), .A2(n13370), .ZN(n8681) );
  INV_X1 U11108 ( .A(n11431), .ZN(n11356) );
  OR2_X1 U11109 ( .A1(n14598), .A2(n13369), .ZN(n8682) );
  NAND2_X1 U11110 ( .A1(n8683), .A2(n8682), .ZN(n11590) );
  XNOR2_X1 U11111 ( .A(n14589), .B(n8684), .ZN(n9010) );
  NAND2_X1 U11112 ( .A1(n14589), .A2(n13368), .ZN(n8685) );
  XNOR2_X1 U11113 ( .A(n11878), .B(n11801), .ZN(n11679) );
  INV_X1 U11114 ( .A(n11679), .ZN(n8686) );
  OR2_X1 U11115 ( .A1(n11878), .A2(n13367), .ZN(n8687) );
  NAND2_X1 U11116 ( .A1(n13687), .A2(n13366), .ZN(n8688) );
  XNOR2_X1 U11117 ( .A(n13679), .B(n13328), .ZN(n11955) );
  NAND2_X1 U11118 ( .A1(n13679), .A2(n13365), .ZN(n8689) );
  OR2_X1 U11119 ( .A1(n13674), .A2(n13364), .ZN(n8691) );
  NAND2_X1 U11120 ( .A1(n13583), .A2(n13363), .ZN(n9013) );
  NAND2_X1 U11121 ( .A1(n13575), .A2(n9013), .ZN(n8692) );
  OR2_X1 U11122 ( .A1(n13583), .A2(n13363), .ZN(n9014) );
  NAND2_X1 U11123 ( .A1(n8692), .A2(n9014), .ZN(n13556) );
  NAND2_X1 U11124 ( .A1(n13713), .A2(n13362), .ZN(n8693) );
  NAND2_X1 U11125 ( .A1(n13556), .A2(n8693), .ZN(n8695) );
  OR2_X1 U11126 ( .A1(n13713), .A2(n13362), .ZN(n8694) );
  NAND2_X1 U11127 ( .A1(n8695), .A2(n8694), .ZN(n13552) );
  NOR2_X1 U11128 ( .A1(n13657), .A2(n13361), .ZN(n8696) );
  NAND2_X1 U11129 ( .A1(n13657), .A2(n13361), .ZN(n8697) );
  XNOR2_X1 U11130 ( .A(n13537), .B(n13274), .ZN(n13532) );
  AND2_X1 U11131 ( .A1(n13647), .A2(n13359), .ZN(n8698) );
  OAI22_X1 U11132 ( .A1(n13515), .A2(n8698), .B1(n13359), .B2(n13647), .ZN(
        n13497) );
  NAND2_X1 U11133 ( .A1(n13487), .A2(n13341), .ZN(n8700) );
  NAND2_X1 U11134 ( .A1(n13482), .A2(n8700), .ZN(n8702) );
  OR2_X1 U11135 ( .A1(n13487), .A2(n13341), .ZN(n8701) );
  NAND2_X1 U11136 ( .A1(n8702), .A2(n8701), .ZN(n13478) );
  OR2_X1 U11137 ( .A1(n13630), .A2(n13356), .ZN(n8703) );
  INV_X1 U11138 ( .A(n9020), .ZN(n13446) );
  XNOR2_X1 U11139 ( .A(n8705), .B(n6594), .ZN(n13430) );
  NAND2_X1 U11140 ( .A1(n8706), .A2(n13581), .ZN(n9902) );
  NAND2_X1 U11141 ( .A1(n6577), .A2(n11409), .ZN(n8753) );
  OR2_X1 U11142 ( .A1(n8753), .A2(n9024), .ZN(n14970) );
  NAND2_X1 U11143 ( .A1(n8707), .A2(n7148), .ZN(n8712) );
  NAND2_X1 U11144 ( .A1(n8712), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8708) );
  MUX2_X1 U11145 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8708), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8709) );
  NAND2_X1 U11146 ( .A1(n8709), .A2(n8715), .ZN(n11934) );
  INV_X1 U11147 ( .A(P2_B_REG_SCAN_IN), .ZN(n9028) );
  NOR2_X1 U11148 ( .A1(n8707), .A2(n13724), .ZN(n8710) );
  MUX2_X1 U11149 ( .A(n13724), .B(n8710), .S(P2_IR_REG_24__SCAN_IN), .Z(n8711)
         );
  INV_X1 U11150 ( .A(n8711), .ZN(n8713) );
  NAND2_X1 U11151 ( .A1(n8713), .A2(n8712), .ZN(n11796) );
  XOR2_X1 U11152 ( .A(n9028), .B(n11796), .Z(n8714) );
  AND2_X1 U11153 ( .A1(n11934), .A2(n8714), .ZN(n8719) );
  NAND2_X1 U11154 ( .A1(n8715), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8716) );
  MUX2_X1 U11155 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8716), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8718) );
  NAND2_X1 U11156 ( .A1(n8718), .A2(n8717), .ZN(n13742) );
  INV_X1 U11157 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15487) );
  AOI22_X1 U11158 ( .A1(n14958), .A2(n15487), .B1(n13742), .B2(n11934), .ZN(
        n9919) );
  INV_X1 U11159 ( .A(n13742), .ZN(n8721) );
  NOR2_X1 U11160 ( .A1(n11796), .A2(n11934), .ZN(n8720) );
  NAND2_X1 U11161 ( .A1(n8721), .A2(n8720), .ZN(n9897) );
  INV_X1 U11162 ( .A(n8722), .ZN(n8723) );
  NAND2_X1 U11163 ( .A1(n8724), .A2(n8723), .ZN(n8725) );
  NAND2_X1 U11164 ( .A1(n8725), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8727) );
  XNOR2_X1 U11165 ( .A(n8727), .B(n8726), .ZN(n9898) );
  AND2_X1 U11166 ( .A1(n9897), .A2(n9898), .ZN(n9927) );
  OR2_X1 U11167 ( .A1(n9919), .A2(n14966), .ZN(n14964) );
  NOR4_X1 U11168 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8731) );
  NOR4_X1 U11169 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8730) );
  NOR4_X1 U11170 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8729) );
  NOR4_X1 U11171 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n8728) );
  NAND4_X1 U11172 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n8737)
         );
  NOR2_X1 U11173 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n8735) );
  NOR4_X1 U11174 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8734) );
  NOR4_X1 U11175 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n8733) );
  NOR4_X1 U11176 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8732) );
  NAND4_X1 U11177 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n8736)
         );
  OAI21_X1 U11178 ( .B1(n8737), .B2(n8736), .A(n14958), .ZN(n9918) );
  INV_X1 U11179 ( .A(n9024), .ZN(n11528) );
  NAND2_X1 U11180 ( .A1(n11528), .A2(n13581), .ZN(n9037) );
  OR2_X1 U11181 ( .A1(n10019), .A2(n9933), .ZN(n10404) );
  NAND3_X1 U11182 ( .A1(n9918), .A2(n9930), .A3(n10404), .ZN(n8738) );
  INV_X1 U11183 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U11184 ( .A1(n14958), .A2(n14961), .ZN(n8740) );
  NAND2_X1 U11185 ( .A1(n13742), .A2(n11796), .ZN(n8739) );
  INV_X1 U11186 ( .A(n14962), .ZN(n9920) );
  NAND2_X1 U11187 ( .A1(n15037), .A2(n14597), .ZN(n13672) );
  INV_X1 U11188 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8741) );
  NOR2_X1 U11189 ( .A1(n15037), .A2(n8741), .ZN(n8742) );
  AND2_X2 U11190 ( .A1(n10409), .A2(n6577), .ZN(n8747) );
  NAND2_X1 U11191 ( .A1(n8750), .A2(n8747), .ZN(n8748) );
  INV_X1 U11192 ( .A(n8751), .ZN(n8749) );
  INV_X1 U11193 ( .A(n8750), .ZN(n9000) );
  NAND2_X1 U11194 ( .A1(n8968), .A2(n8750), .ZN(n8752) );
  NAND2_X1 U11195 ( .A1(n8752), .A2(n8751), .ZN(n8755) );
  NAND2_X1 U11196 ( .A1(n8753), .A2(n9035), .ZN(n8754) );
  NAND2_X1 U11197 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  NAND2_X1 U11198 ( .A1(n9903), .A2(n8968), .ZN(n8758) );
  NAND2_X1 U11199 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  NAND2_X1 U11200 ( .A1(n8761), .A2(n8760), .ZN(n8762) );
  NAND2_X1 U11201 ( .A1(n8763), .A2(n8762), .ZN(n8768) );
  NAND2_X1 U11202 ( .A1(n13381), .A2(n8848), .ZN(n8765) );
  NAND2_X1 U11203 ( .A1(n10343), .A2(n8993), .ZN(n8764) );
  NAND2_X1 U11204 ( .A1(n8765), .A2(n8764), .ZN(n8767) );
  AOI22_X1 U11205 ( .A1(n13381), .A2(n8992), .B1(n10343), .B2(n8848), .ZN(
        n8766) );
  NOR2_X1 U11206 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  INV_X2 U11207 ( .A(n8968), .ZN(n8969) );
  NAND2_X1 U11208 ( .A1(n13380), .A2(n8969), .ZN(n8772) );
  NAND2_X1 U11209 ( .A1(n10340), .A2(n8848), .ZN(n8771) );
  NAND2_X1 U11210 ( .A1(n8772), .A2(n8771), .ZN(n8774) );
  AOI22_X1 U11211 ( .A1(n13380), .A2(n8848), .B1(n10340), .B2(n8969), .ZN(
        n8773) );
  NAND2_X1 U11212 ( .A1(n10386), .A2(n8969), .ZN(n8777) );
  NAND2_X1 U11213 ( .A1(n13378), .A2(n8848), .ZN(n8776) );
  NAND2_X1 U11214 ( .A1(n8777), .A2(n8776), .ZN(n8780) );
  INV_X2 U11215 ( .A(n8993), .ZN(n8970) );
  AOI22_X1 U11216 ( .A1(n10386), .A2(n8970), .B1(n8969), .B2(n13378), .ZN(
        n8778) );
  AOI21_X1 U11217 ( .B1(n8781), .B2(n8780), .A(n8778), .ZN(n8779) );
  NAND2_X1 U11218 ( .A1(n10425), .A2(n8848), .ZN(n8784) );
  NAND2_X1 U11219 ( .A1(n13377), .A2(n8969), .ZN(n8783) );
  NAND2_X1 U11220 ( .A1(n10425), .A2(n8969), .ZN(n8786) );
  NAND2_X1 U11221 ( .A1(n13377), .A2(n8970), .ZN(n8785) );
  NAND2_X1 U11222 ( .A1(n8786), .A2(n8785), .ZN(n8787) );
  NAND2_X1 U11223 ( .A1(n14983), .A2(n8969), .ZN(n8789) );
  NAND2_X1 U11224 ( .A1(n13376), .A2(n8970), .ZN(n8788) );
  NAND2_X1 U11225 ( .A1(n8789), .A2(n8788), .ZN(n8794) );
  NAND2_X1 U11226 ( .A1(n8793), .A2(n8794), .ZN(n8792) );
  AOI22_X1 U11227 ( .A1(n14983), .A2(n8970), .B1(n8969), .B2(n13376), .ZN(
        n8790) );
  INV_X1 U11228 ( .A(n8790), .ZN(n8791) );
  INV_X1 U11229 ( .A(n8793), .ZN(n8796) );
  INV_X1 U11230 ( .A(n8794), .ZN(n8795) );
  NAND2_X1 U11231 ( .A1(n10839), .A2(n8970), .ZN(n8798) );
  NAND2_X1 U11232 ( .A1(n13375), .A2(n8969), .ZN(n8797) );
  NAND2_X1 U11233 ( .A1(n8798), .A2(n8797), .ZN(n8800) );
  AOI22_X1 U11234 ( .A1(n10839), .A2(n8969), .B1(n13375), .B2(n8970), .ZN(
        n8799) );
  NAND2_X1 U11235 ( .A1(n15003), .A2(n8969), .ZN(n8802) );
  NAND2_X1 U11236 ( .A1(n13374), .A2(n8848), .ZN(n8801) );
  NAND2_X1 U11237 ( .A1(n8802), .A2(n8801), .ZN(n8808) );
  NAND2_X1 U11238 ( .A1(n8807), .A2(n8808), .ZN(n8806) );
  NAND2_X1 U11239 ( .A1(n15003), .A2(n8970), .ZN(n8804) );
  NAND2_X1 U11240 ( .A1(n13374), .A2(n8969), .ZN(n8803) );
  NAND2_X1 U11241 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  NAND2_X1 U11242 ( .A1(n8806), .A2(n8805), .ZN(n8812) );
  NAND2_X1 U11243 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  NAND2_X1 U11244 ( .A1(n10951), .A2(n8970), .ZN(n8814) );
  NAND2_X1 U11245 ( .A1(n13373), .A2(n8969), .ZN(n8813) );
  NAND2_X1 U11246 ( .A1(n8814), .A2(n8813), .ZN(n8817) );
  AOI22_X1 U11247 ( .A1(n10951), .A2(n8969), .B1(n13373), .B2(n8970), .ZN(
        n8815) );
  INV_X1 U11248 ( .A(n8816), .ZN(n8819) );
  NAND2_X1 U11249 ( .A1(n11235), .A2(n8969), .ZN(n8821) );
  NAND2_X1 U11250 ( .A1(n13372), .A2(n8848), .ZN(n8820) );
  NAND2_X1 U11251 ( .A1(n8821), .A2(n8820), .ZN(n8826) );
  NAND2_X1 U11252 ( .A1(n11235), .A2(n8970), .ZN(n8823) );
  NAND2_X1 U11253 ( .A1(n13372), .A2(n8969), .ZN(n8822) );
  NAND2_X1 U11254 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  NAND2_X1 U11255 ( .A1(n14938), .A2(n8970), .ZN(n8829) );
  NAND2_X1 U11256 ( .A1(n13371), .A2(n8969), .ZN(n8828) );
  NAND2_X1 U11257 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  AOI22_X1 U11258 ( .A1(n14938), .A2(n8969), .B1(n13371), .B2(n8970), .ZN(
        n8830) );
  NAND2_X1 U11259 ( .A1(n11431), .A2(n8969), .ZN(n8834) );
  NAND2_X1 U11260 ( .A1(n13370), .A2(n8848), .ZN(n8833) );
  NAND2_X1 U11261 ( .A1(n11431), .A2(n8970), .ZN(n8835) );
  OAI21_X1 U11262 ( .B1(n11191), .B2(n8970), .A(n8835), .ZN(n8836) );
  NAND2_X1 U11263 ( .A1(n14598), .A2(n8970), .ZN(n8839) );
  NAND2_X1 U11264 ( .A1(n13369), .A2(n8969), .ZN(n8838) );
  NAND2_X1 U11265 ( .A1(n8839), .A2(n8838), .ZN(n8841) );
  AOI22_X1 U11266 ( .A1(n14598), .A2(n8969), .B1(n13369), .B2(n8848), .ZN(
        n8840) );
  NAND2_X1 U11267 ( .A1(n14589), .A2(n8969), .ZN(n8844) );
  NAND2_X1 U11268 ( .A1(n13368), .A2(n8970), .ZN(n8843) );
  NAND2_X1 U11269 ( .A1(n8844), .A2(n8843), .ZN(n8846) );
  AOI22_X1 U11270 ( .A1(n14589), .A2(n8970), .B1(n8969), .B2(n13368), .ZN(
        n8845) );
  NAND2_X1 U11271 ( .A1(n11878), .A2(n8848), .ZN(n8850) );
  NAND2_X1 U11272 ( .A1(n13367), .A2(n8993), .ZN(n8849) );
  NAND2_X1 U11273 ( .A1(n8850), .A2(n8849), .ZN(n8856) );
  NAND2_X1 U11274 ( .A1(n11878), .A2(n8969), .ZN(n8852) );
  NAND2_X1 U11275 ( .A1(n13367), .A2(n8970), .ZN(n8851) );
  NAND2_X1 U11276 ( .A1(n8852), .A2(n8851), .ZN(n8853) );
  NAND2_X1 U11277 ( .A1(n8854), .A2(n8853), .ZN(n8860) );
  INV_X1 U11278 ( .A(n8855), .ZN(n8858) );
  NAND2_X1 U11279 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  NAND2_X1 U11280 ( .A1(n13687), .A2(n8969), .ZN(n8862) );
  NAND2_X1 U11281 ( .A1(n13366), .A2(n8970), .ZN(n8861) );
  NAND2_X1 U11282 ( .A1(n8862), .A2(n8861), .ZN(n8864) );
  AOI22_X1 U11283 ( .A1(n13687), .A2(n8970), .B1(n8969), .B2(n13366), .ZN(
        n8863) );
  NAND2_X1 U11284 ( .A1(n13679), .A2(n8970), .ZN(n8867) );
  NAND2_X1 U11285 ( .A1(n13365), .A2(n8992), .ZN(n8866) );
  NAND2_X1 U11286 ( .A1(n8867), .A2(n8866), .ZN(n8871) );
  NAND2_X1 U11287 ( .A1(n13679), .A2(n8969), .ZN(n8868) );
  OAI21_X1 U11288 ( .B1(n13328), .B2(n8993), .A(n8868), .ZN(n8869) );
  NAND2_X1 U11289 ( .A1(n13674), .A2(n8969), .ZN(n8874) );
  NAND2_X1 U11290 ( .A1(n13364), .A2(n8970), .ZN(n8873) );
  AOI22_X1 U11291 ( .A1(n13674), .A2(n8970), .B1(n8969), .B2(n13364), .ZN(
        n8875) );
  NAND2_X1 U11292 ( .A1(n13583), .A2(n8970), .ZN(n8877) );
  NAND2_X1 U11293 ( .A1(n13363), .A2(n8969), .ZN(n8876) );
  NAND2_X1 U11294 ( .A1(n8877), .A2(n8876), .ZN(n8879) );
  AOI22_X1 U11295 ( .A1(n13583), .A2(n8992), .B1(n13363), .B2(n8970), .ZN(
        n8878) );
  AOI21_X1 U11296 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8882) );
  AND2_X1 U11297 ( .A1(n13362), .A2(n8970), .ZN(n8883) );
  AOI21_X1 U11298 ( .B1(n13713), .B2(n8969), .A(n8883), .ZN(n8888) );
  NAND2_X1 U11299 ( .A1(n13657), .A2(n8993), .ZN(n8884) );
  OAI21_X1 U11300 ( .B1(n8885), .B2(n8993), .A(n8884), .ZN(n8890) );
  NAND2_X1 U11301 ( .A1(n13713), .A2(n8970), .ZN(n8886) );
  OAI21_X1 U11302 ( .B1(n13273), .B2(n8970), .A(n8886), .ZN(n8887) );
  INV_X1 U11303 ( .A(n8890), .ZN(n8893) );
  AND2_X1 U11304 ( .A1(n13361), .A2(n8969), .ZN(n8891) );
  AOI21_X1 U11305 ( .B1(n13657), .B2(n8970), .A(n8891), .ZN(n8894) );
  INV_X1 U11306 ( .A(n8894), .ZN(n8892) );
  NAND2_X1 U11307 ( .A1(n13537), .A2(n8969), .ZN(n8896) );
  NAND2_X1 U11308 ( .A1(n13360), .A2(n8970), .ZN(n8895) );
  NAND2_X1 U11309 ( .A1(n8896), .A2(n8895), .ZN(n8898) );
  NAND2_X1 U11310 ( .A1(n8897), .A2(n8898), .ZN(n8902) );
  OAI22_X1 U11311 ( .A1(n13709), .A2(n8993), .B1(n13274), .B2(n8970), .ZN(
        n8901) );
  INV_X1 U11312 ( .A(n8897), .ZN(n8900) );
  INV_X1 U11313 ( .A(n8898), .ZN(n8899) );
  AOI22_X1 U11314 ( .A1(n13647), .A2(n8970), .B1(n8969), .B2(n13359), .ZN(
        n8903) );
  AOI22_X1 U11315 ( .A1(n13647), .A2(n8969), .B1(n13359), .B2(n8970), .ZN(
        n8904) );
  OAI22_X1 U11316 ( .A1(n13705), .A2(n8970), .B1(n13282), .B2(n8993), .ZN(
        n8907) );
  AOI22_X1 U11317 ( .A1(n8905), .A2(n8970), .B1(n8969), .B2(n13358), .ZN(n8906) );
  INV_X1 U11318 ( .A(n8907), .ZN(n8908) );
  AOI22_X1 U11319 ( .A1(n13635), .A2(n8970), .B1(n8969), .B2(n13357), .ZN(
        n8916) );
  OAI22_X1 U11320 ( .A1(n13487), .A2(n8970), .B1(n13341), .B2(n8993), .ZN(
        n8915) );
  AND2_X1 U11321 ( .A1(n8916), .A2(n8915), .ZN(n8909) );
  AND2_X1 U11322 ( .A1(n13356), .A2(n8969), .ZN(n8912) );
  AOI21_X1 U11323 ( .B1(n13630), .B2(n8970), .A(n8912), .ZN(n8972) );
  NAND2_X1 U11324 ( .A1(n13630), .A2(n8992), .ZN(n8914) );
  NAND2_X1 U11325 ( .A1(n13356), .A2(n8970), .ZN(n8913) );
  NAND2_X1 U11326 ( .A1(n8914), .A2(n8913), .ZN(n8971) );
  OAI22_X1 U11327 ( .A1(n8972), .A2(n8971), .B1(n8916), .B2(n8915), .ZN(n8917)
         );
  INV_X1 U11328 ( .A(SI_29_), .ZN(n13188) );
  NAND2_X1 U11329 ( .A1(n8921), .A2(n13188), .ZN(n8944) );
  MUX2_X1 U11330 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9957), .Z(n8922) );
  NAND2_X1 U11331 ( .A1(n8922), .A2(SI_30_), .ZN(n8949) );
  INV_X1 U11332 ( .A(n8922), .ZN(n8923) );
  INV_X1 U11333 ( .A(SI_30_), .ZN(n12449) );
  NAND2_X1 U11334 ( .A1(n8923), .A2(n12449), .ZN(n8945) );
  AND2_X1 U11335 ( .A1(n8949), .A2(n8945), .ZN(n8924) );
  NAND2_X1 U11336 ( .A1(n12276), .A2(n8958), .ZN(n8926) );
  INV_X1 U11337 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12278) );
  OR2_X1 U11338 ( .A1(n8960), .A2(n12278), .ZN(n8925) );
  AND2_X1 U11339 ( .A1(n13352), .A2(n8969), .ZN(n8927) );
  AOI21_X1 U11340 ( .B1(n13425), .B2(n8970), .A(n8927), .ZN(n8985) );
  INV_X1 U11341 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U11342 ( .A1(n6582), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U11343 ( .A1(n8654), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8929) );
  OAI211_X1 U11344 ( .C1(n8931), .C2(n15449), .A(n8930), .B(n8929), .ZN(n13421) );
  OAI211_X1 U11345 ( .C1(n8932), .C2(n9024), .A(n9029), .B(n9037), .ZN(n8933)
         );
  AOI21_X1 U11346 ( .B1(n13421), .B2(n8970), .A(n8933), .ZN(n8935) );
  NAND2_X1 U11347 ( .A1(n13425), .A2(n8969), .ZN(n8934) );
  OAI21_X1 U11348 ( .B1(n8996), .B2(n8935), .A(n8934), .ZN(n8984) );
  NAND2_X1 U11349 ( .A1(n8985), .A2(n8984), .ZN(n8941) );
  AND2_X1 U11350 ( .A1(n13353), .A2(n8969), .ZN(n8936) );
  AOI21_X1 U11351 ( .B1(n8937), .B2(n8970), .A(n8936), .ZN(n8981) );
  NAND2_X1 U11352 ( .A1(n8937), .A2(n8969), .ZN(n8939) );
  NAND2_X1 U11353 ( .A1(n13353), .A2(n8848), .ZN(n8938) );
  NAND2_X1 U11354 ( .A1(n8939), .A2(n8938), .ZN(n8980) );
  NAND2_X1 U11355 ( .A1(n8981), .A2(n8980), .ZN(n8940) );
  NAND2_X1 U11356 ( .A1(n8941), .A2(n8940), .ZN(n8963) );
  INV_X1 U11357 ( .A(n8949), .ZN(n8943) );
  XNOR2_X1 U11358 ( .A(n8942), .B(SI_31_), .ZN(n8950) );
  NAND2_X1 U11359 ( .A1(n8945), .A2(n8944), .ZN(n8951) );
  INV_X1 U11360 ( .A(n8950), .ZN(n8946) );
  NOR2_X1 U11361 ( .A1(n8951), .A2(n8946), .ZN(n8947) );
  NAND2_X1 U11362 ( .A1(n8948), .A2(n8947), .ZN(n8955) );
  XNOR2_X1 U11363 ( .A(n8950), .B(n8949), .ZN(n8953) );
  NOR2_X1 U11364 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  OR2_X1 U11365 ( .A1(n8953), .A2(n8952), .ZN(n8954) );
  NAND2_X1 U11366 ( .A1(n13722), .A2(n8958), .ZN(n8962) );
  INV_X1 U11367 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8959) );
  OR2_X1 U11368 ( .A1(n8960), .A2(n8959), .ZN(n8961) );
  NAND2_X1 U11369 ( .A1(n8962), .A2(n8961), .ZN(n8991) );
  XNOR2_X1 U11370 ( .A(n8991), .B(n13421), .ZN(n8977) );
  NAND2_X1 U11371 ( .A1(n8963), .A2(n8977), .ZN(n8982) );
  AND2_X1 U11372 ( .A1(n13354), .A2(n8969), .ZN(n8964) );
  AOI21_X1 U11373 ( .B1(n13617), .B2(n8970), .A(n8964), .ZN(n8979) );
  NAND2_X1 U11374 ( .A1(n13617), .A2(n8969), .ZN(n8966) );
  NAND2_X1 U11375 ( .A1(n13354), .A2(n8970), .ZN(n8965) );
  NAND2_X1 U11376 ( .A1(n8966), .A2(n8965), .ZN(n8978) );
  NAND2_X1 U11377 ( .A1(n8979), .A2(n8978), .ZN(n8967) );
  OAI22_X1 U11378 ( .A1(n13623), .A2(n8970), .B1(n13343), .B2(n8993), .ZN(
        n8975) );
  AOI22_X1 U11379 ( .A1(n13228), .A2(n8970), .B1(n8969), .B2(n13355), .ZN(
        n8976) );
  AOI22_X1 U11380 ( .A1(n8975), .A2(n8976), .B1(n8972), .B2(n8971), .ZN(n8973)
         );
  INV_X1 U11381 ( .A(n8977), .ZN(n9021) );
  OAI22_X1 U11382 ( .A1(n8981), .A2(n8980), .B1(n8979), .B2(n8978), .ZN(n8983)
         );
  OAI21_X1 U11383 ( .B1(n9021), .B2(n8983), .A(n8982), .ZN(n8987) );
  NOR2_X1 U11384 ( .A1(n7533), .A2(n7534), .ZN(n8994) );
  NAND2_X1 U11385 ( .A1(n8995), .A2(n8994), .ZN(n9042) );
  INV_X1 U11386 ( .A(n9898), .ZN(n10018) );
  NAND2_X1 U11387 ( .A1(n10018), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11694) );
  OR2_X1 U11388 ( .A1(n11694), .A2(n13581), .ZN(n9025) );
  NOR2_X1 U11389 ( .A1(n9025), .A2(n9029), .ZN(n9023) );
  XNOR2_X1 U11390 ( .A(n13425), .B(n8996), .ZN(n9022) );
  XNOR2_X1 U11391 ( .A(n13630), .B(n8997), .ZN(n13477) );
  XNOR2_X1 U11392 ( .A(n11431), .B(n11191), .ZN(n11241) );
  XNOR2_X1 U11393 ( .A(n11235), .B(n11192), .ZN(n11006) );
  NAND2_X1 U11394 ( .A1(n9000), .A2(n14969), .ZN(n9001) );
  NAND2_X1 U11395 ( .A1(n10329), .A2(n9001), .ZN(n14971) );
  AND4_X1 U11396 ( .A1(n6757), .A2(n10232), .A3(n9024), .A4(n14971), .ZN(n9004) );
  NAND4_X1 U11397 ( .A1(n10596), .A2(n9004), .A3(n9003), .A4(n9002), .ZN(n9005) );
  NOR2_X1 U11398 ( .A1(n10538), .A2(n9005), .ZN(n9006) );
  NAND4_X1 U11399 ( .A1(n10846), .A2(n9006), .A3(n10728), .A4(n14990), .ZN(
        n9007) );
  OR4_X1 U11400 ( .A1(n11399), .A2(n11006), .A3(n9008), .A4(n9007), .ZN(n9009)
         );
  OR3_X1 U11401 ( .A1(n9010), .A2(n11241), .A3(n9009), .ZN(n9011) );
  OR4_X1 U11402 ( .A1(n11955), .A2(n11810), .A3(n11679), .A4(n9011), .ZN(n9012) );
  NOR2_X1 U11403 ( .A1(n13564), .A2(n9012), .ZN(n9015) );
  NAND2_X1 U11404 ( .A1(n9014), .A2(n9013), .ZN(n13576) );
  NAND4_X1 U11405 ( .A1(n13551), .A2(n9015), .A3(n13603), .A4(n13576), .ZN(
        n9016) );
  NOR2_X1 U11406 ( .A1(n13532), .A2(n9016), .ZN(n9017) );
  NAND4_X1 U11407 ( .A1(n13489), .A2(n13516), .A3(n9017), .A4(n13499), .ZN(
        n9018) );
  NOR2_X1 U11408 ( .A1(n13477), .A2(n9018), .ZN(n9019) );
  OAI211_X1 U11409 ( .C1(n9042), .C2(n9024), .A(n9023), .B(n9030), .ZN(n9044)
         );
  MUX2_X1 U11410 ( .A(n6577), .B(n11557), .S(n9024), .Z(n9026) );
  NOR2_X1 U11411 ( .A1(n9026), .A2(n9025), .ZN(n9034) );
  INV_X1 U11412 ( .A(n11694), .ZN(n9038) );
  NOR4_X1 U11413 ( .A1(n14966), .A2(n8659), .A3(n13340), .A4(n9037), .ZN(n9027) );
  AOI211_X1 U11414 ( .C1(n9038), .C2(n6577), .A(n9028), .B(n9027), .ZN(n9032)
         );
  AOI21_X1 U11415 ( .B1(n9042), .B2(n9034), .A(n9033), .ZN(n9043) );
  INV_X1 U11416 ( .A(n9035), .ZN(n9901) );
  NOR2_X1 U11417 ( .A1(n9036), .A2(n9901), .ZN(n9040) );
  OAI21_X1 U11418 ( .B1(n11557), .B2(n11409), .A(n9037), .ZN(n9039) );
  OAI21_X1 U11419 ( .B1(n9040), .B2(n9039), .A(n9038), .ZN(n9041) );
  NOR2_X1 U11420 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n9052) );
  NAND2_X1 U11421 ( .A1(n9058), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9059) );
  INV_X1 U11422 ( .A(n9060), .ZN(n13181) );
  INV_X1 U11423 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9062) );
  OR2_X1 U11424 ( .A1(n9119), .A2(n9062), .ZN(n9068) );
  AND2_X2 U11425 ( .A1(n12447), .A2(n9063), .ZN(n9117) );
  AND2_X2 U11426 ( .A1(n9064), .A2(n9063), .ZN(n9141) );
  NAND2_X1 U11427 ( .A1(n9141), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9066) );
  INV_X1 U11428 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11131) );
  OR2_X1 U11429 ( .A1(n9121), .A2(n11131), .ZN(n9065) );
  INV_X1 U11430 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U11431 ( .A1(n9069), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U11432 ( .A1(n9070), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9071) );
  AND2_X1 U11433 ( .A1(n9092), .A2(n9071), .ZN(n9073) );
  MUX2_X1 U11434 ( .A(n9073), .B(n9072), .S(n9957), .Z(n9939) );
  XNOR2_X2 U11435 ( .A(n9075), .B(n9074), .ZN(n12431) );
  NAND2_X1 U11436 ( .A1(n9076), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9077) );
  XNOR2_X2 U11437 ( .A(n9077), .B(n6864), .ZN(n12733) );
  MUX2_X1 U11438 ( .A(n10667), .B(n9939), .S(n6567), .Z(n11078) );
  NOR2_X2 U11439 ( .A1(n15110), .A2(n11078), .ZN(n12075) );
  INV_X1 U11440 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U11441 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9078) );
  NAND2_X1 U11442 ( .A1(n9141), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9085) );
  INV_X1 U11443 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9080) );
  OR2_X1 U11444 ( .A1(n9119), .A2(n9080), .ZN(n9083) );
  INV_X1 U11445 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9081) );
  OR2_X1 U11446 ( .A1(n9121), .A2(n9081), .ZN(n9082) );
  NAND2_X1 U11447 ( .A1(n15122), .A2(n9601), .ZN(n12077) );
  NAND2_X1 U11448 ( .A1(n9141), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U11449 ( .A1(n9117), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9090) );
  INV_X1 U11450 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9086) );
  OR2_X1 U11451 ( .A1(n9119), .A2(n9086), .ZN(n9089) );
  INV_X1 U11452 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9087) );
  OR2_X1 U11453 ( .A1(n9121), .A2(n9087), .ZN(n9088) );
  INV_X1 U11454 ( .A(n9092), .ZN(n9093) );
  NAND2_X1 U11455 ( .A1(n15286), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11456 ( .A1(n9095), .A2(n9094), .ZN(n9101) );
  XNOR2_X1 U11457 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9096) );
  XNOR2_X1 U11458 ( .A(n9101), .B(n9096), .ZN(n9963) );
  OR2_X1 U11459 ( .A1(n9100), .A2(n9963), .ZN(n9098) );
  OR2_X1 U11460 ( .A1(n9138), .A2(SI_2_), .ZN(n9097) );
  NAND2_X1 U11461 ( .A1(n15116), .A2(n11015), .ZN(n12086) );
  NAND2_X1 U11462 ( .A1(n13013), .A2(n13018), .ZN(n13012) );
  NAND2_X1 U11463 ( .A1(n13012), .A2(n12081), .ZN(n11294) );
  INV_X1 U11464 ( .A(n9101), .ZN(n9103) );
  NAND2_X1 U11465 ( .A1(n9940), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U11466 ( .A1(n9947), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9104) );
  XNOR2_X1 U11467 ( .A(n9942), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n9106) );
  XNOR2_X1 U11468 ( .A(n9132), .B(n9106), .ZN(n9968) );
  OR2_X1 U11469 ( .A1(n9100), .A2(n9968), .ZN(n9108) );
  OR2_X1 U11470 ( .A1(n9138), .A2(SI_3_), .ZN(n9107) );
  OAI211_X1 U11471 ( .C1(n7257), .C2(n10662), .A(n9108), .B(n9107), .ZN(n15138) );
  INV_X1 U11472 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11473 ( .A1(n9141), .A2(n9109), .ZN(n9115) );
  NAND2_X1 U11474 ( .A1(n9117), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9114) );
  INV_X1 U11475 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9110) );
  OR2_X1 U11476 ( .A1(n9119), .A2(n9110), .ZN(n9113) );
  INV_X1 U11477 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9111) );
  OR2_X1 U11478 ( .A1(n9121), .A2(n9111), .ZN(n9112) );
  NAND4_X1 U11479 ( .A1(n9115), .A2(n9114), .A3(n9113), .A4(n9112), .ZN(n12636) );
  NAND2_X1 U11480 ( .A1(n12636), .A2(n15138), .ZN(n12087) );
  AND2_X1 U11481 ( .A1(n12094), .A2(n12087), .ZN(n11295) );
  NAND2_X1 U11482 ( .A1(n11294), .A2(n11295), .ZN(n9116) );
  NAND2_X1 U11483 ( .A1(n9116), .A2(n12094), .ZN(n11325) );
  NAND2_X1 U11484 ( .A1(n6573), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9125) );
  AND2_X1 U11485 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9118) );
  OR2_X1 U11486 ( .A1(n9118), .A2(n9142), .ZN(n10991) );
  NAND2_X1 U11487 ( .A1(n9141), .A2(n10991), .ZN(n9124) );
  INV_X1 U11488 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9120) );
  OR2_X1 U11489 ( .A1(n12061), .A2(n9120), .ZN(n9123) );
  INV_X1 U11490 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U11491 ( .A1(n9126), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9127) );
  MUX2_X1 U11492 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9127), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9130) );
  INV_X1 U11493 ( .A(n9128), .ZN(n9129) );
  NAND2_X1 U11494 ( .A1(n9942), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11495 ( .A1(n6928), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11496 ( .A1(n9944), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U11497 ( .A1(n9150), .A2(n9134), .ZN(n9135) );
  NAND2_X1 U11498 ( .A1(n9136), .A2(n9135), .ZN(n9137) );
  AND2_X1 U11499 ( .A1(n9151), .A2(n9137), .ZN(n9970) );
  OR2_X1 U11500 ( .A1(n9244), .A2(n9970), .ZN(n9140) );
  OR2_X1 U11501 ( .A1(n12056), .A2(SI_4_), .ZN(n9139) );
  OAI211_X1 U11502 ( .C1(n11127), .C2(n10662), .A(n9140), .B(n9139), .ZN(
        n15142) );
  NAND2_X1 U11503 ( .A1(n11266), .A2(n10999), .ZN(n12091) );
  NAND2_X1 U11504 ( .A1(n12635), .A2(n15142), .ZN(n12092) );
  NAND2_X1 U11505 ( .A1(n11325), .A2(n9605), .ZN(n11326) );
  NAND2_X1 U11506 ( .A1(n11326), .A2(n12091), .ZN(n11259) );
  NAND2_X1 U11507 ( .A1(n6575), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U11508 ( .A1(n9142), .A2(n11105), .ZN(n9160) );
  OR2_X1 U11509 ( .A1(n9142), .A2(n11105), .ZN(n9143) );
  NAND2_X1 U11510 ( .A1(n9160), .A2(n9143), .ZN(n11273) );
  NAND2_X1 U11511 ( .A1(n6571), .A2(n11273), .ZN(n9147) );
  INV_X1 U11512 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n9144) );
  OR2_X1 U11513 ( .A1(n12061), .A2(n9144), .ZN(n9146) );
  INV_X1 U11514 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11087) );
  OR2_X1 U11515 ( .A1(n12062), .A2(n11087), .ZN(n9145) );
  OR2_X1 U11516 ( .A1(n9128), .A2(n9056), .ZN(n9149) );
  XNOR2_X1 U11517 ( .A(n9149), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U11518 ( .A1(n9954), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11519 ( .A1(n9952), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U11520 ( .A1(n9167), .A2(n9152), .ZN(n9154) );
  NAND2_X1 U11521 ( .A1(n9153), .A2(n9154), .ZN(n9157) );
  INV_X1 U11522 ( .A(n9154), .ZN(n9155) );
  AND2_X1 U11523 ( .A1(n9157), .A2(n9168), .ZN(n9973) );
  OR2_X1 U11524 ( .A1(n9244), .A2(n9973), .ZN(n9159) );
  OR2_X1 U11525 ( .A1(n12056), .A2(SI_5_), .ZN(n9158) );
  OAI211_X1 U11526 ( .C1(n11164), .C2(n10662), .A(n9159), .B(n9158), .ZN(
        n15146) );
  INV_X1 U11527 ( .A(n15146), .ZN(n11274) );
  NAND2_X1 U11528 ( .A1(n11492), .A2(n11274), .ZN(n12100) );
  NAND2_X1 U11529 ( .A1(n12634), .A2(n15146), .ZN(n12104) );
  NAND2_X1 U11530 ( .A1(n6575), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U11531 ( .A1(n9160), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11532 ( .A1(n9171), .A2(n9161), .ZN(n11515) );
  NAND2_X1 U11533 ( .A1(n6571), .A2(n11515), .ZN(n9163) );
  INV_X1 U11534 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9162) );
  INV_X1 U11535 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U11536 ( .A1(n9128), .A2(n9165), .ZN(n9185) );
  NAND2_X1 U11537 ( .A1(n9185), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U11538 ( .A(n9166), .B(P3_IR_REG_6__SCAN_IN), .ZN(n15065) );
  INV_X1 U11539 ( .A(SI_6_), .ZN(n9961) );
  OR2_X1 U11540 ( .A1(n12056), .A2(n9961), .ZN(n9170) );
  XNOR2_X1 U11541 ( .A(n9180), .B(n9178), .ZN(n9960) );
  OR2_X1 U11542 ( .A1(n9244), .A2(n9960), .ZN(n9169) );
  OAI211_X1 U11543 ( .C1(n10662), .C2(n11161), .A(n9170), .B(n9169), .ZN(
        n11496) );
  INV_X1 U11544 ( .A(n11496), .ZN(n15150) );
  NAND2_X1 U11545 ( .A1(n12633), .A2(n15150), .ZN(n12105) );
  AND2_X1 U11546 ( .A1(n9171), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9172) );
  OR2_X1 U11547 ( .A1(n9172), .A2(n9194), .ZN(n11488) );
  NAND2_X1 U11548 ( .A1(n6571), .A2(n11488), .ZN(n9177) );
  NAND2_X1 U11549 ( .A1(n6575), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9176) );
  INV_X1 U11550 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n9173) );
  OR2_X1 U11551 ( .A1(n12061), .A2(n9173), .ZN(n9175) );
  INV_X1 U11552 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11151) );
  OR2_X1 U11553 ( .A1(n12062), .A2(n11151), .ZN(n9174) );
  NAND4_X1 U11554 ( .A1(n9177), .A2(n9176), .A3(n9175), .A4(n9174), .ZN(n12632) );
  INV_X1 U11555 ( .A(n12632), .ZN(n11600) );
  OR2_X1 U11556 ( .A1(n12056), .A2(SI_7_), .ZN(n9190) );
  INV_X1 U11557 ( .A(n9178), .ZN(n9179) );
  NAND2_X1 U11558 ( .A1(n9984), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11559 ( .A1(n9986), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11560 ( .A1(n9203), .A2(n9181), .ZN(n9182) );
  NAND2_X1 U11561 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  AND2_X1 U11562 ( .A1(n9204), .A2(n9184), .ZN(n9976) );
  OR2_X1 U11563 ( .A1(n9244), .A2(n9976), .ZN(n9189) );
  NAND2_X1 U11564 ( .A1(n9201), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9187) );
  XNOR2_X1 U11565 ( .A(n9187), .B(n9186), .ZN(n11215) );
  NAND2_X1 U11566 ( .A1(n9387), .A2(n11215), .ZN(n9188) );
  NAND2_X1 U11567 ( .A1(n11600), .A2(n15154), .ZN(n12112) );
  INV_X1 U11568 ( .A(n15154), .ZN(n9191) );
  NAND2_X1 U11569 ( .A1(n12632), .A2(n9191), .ZN(n12111) );
  NAND2_X1 U11570 ( .A1(n11374), .A2(n12235), .ZN(n9192) );
  NAND2_X1 U11571 ( .A1(n9192), .A2(n12112), .ZN(n11606) );
  NAND2_X1 U11572 ( .A1(n6574), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9200) );
  NOR2_X1 U11573 ( .A1(n9194), .A2(n9193), .ZN(n9195) );
  OR2_X1 U11574 ( .A1(n9211), .A2(n9195), .ZN(n11593) );
  NAND2_X1 U11575 ( .A1(n6571), .A2(n11593), .ZN(n9199) );
  OR2_X1 U11576 ( .A1(n12061), .A2(n15164), .ZN(n9198) );
  INV_X1 U11577 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n9196) );
  OR2_X1 U11578 ( .A1(n12062), .A2(n9196), .ZN(n9197) );
  NAND4_X1 U11579 ( .A1(n9200), .A2(n9199), .A3(n9198), .A4(n9197), .ZN(n11728) );
  INV_X1 U11580 ( .A(n11728), .ZN(n11735) );
  OAI21_X1 U11581 ( .B1(n9201), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9202) );
  XNOR2_X1 U11582 ( .A(n9202), .B(P3_IR_REG_8__SCAN_IN), .ZN(n15081) );
  INV_X1 U11583 ( .A(SI_8_), .ZN(n15360) );
  OR2_X1 U11584 ( .A1(n12056), .A2(n15360), .ZN(n9209) );
  NAND2_X1 U11585 ( .A1(n9994), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11586 ( .A1(n9992), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9205) );
  OAI21_X1 U11587 ( .B1(n9207), .B2(n9206), .A(n9222), .ZN(n9966) );
  OR2_X1 U11588 ( .A1(n9244), .A2(n9966), .ZN(n9208) );
  OAI211_X1 U11589 ( .C1(n10662), .C2(n11213), .A(n9209), .B(n9208), .ZN(
        n11603) );
  NAND2_X1 U11590 ( .A1(n11735), .A2(n11603), .ZN(n12115) );
  INV_X1 U11591 ( .A(n11603), .ZN(n15160) );
  NAND2_X1 U11592 ( .A1(n11728), .A2(n15160), .ZN(n12116) );
  NAND2_X1 U11593 ( .A1(n11606), .A2(n12234), .ZN(n9210) );
  NAND2_X1 U11594 ( .A1(n9210), .A2(n12115), .ZN(n11618) );
  OR2_X1 U11595 ( .A1(n9211), .A2(n11219), .ZN(n9212) );
  NAND2_X1 U11596 ( .A1(n9228), .A2(n9212), .ZN(n11738) );
  NAND2_X1 U11597 ( .A1(n6571), .A2(n11738), .ZN(n9217) );
  NAND2_X1 U11598 ( .A1(n6574), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9216) );
  INV_X1 U11599 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n9213) );
  OR2_X1 U11600 ( .A1(n12061), .A2(n9213), .ZN(n9215) );
  INV_X1 U11601 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11207) );
  OR2_X1 U11602 ( .A1(n12062), .A2(n11207), .ZN(n9214) );
  NAND4_X1 U11603 ( .A1(n9217), .A2(n9216), .A3(n9215), .A4(n9214), .ZN(n12631) );
  OR2_X1 U11604 ( .A1(n9218), .A2(n9056), .ZN(n9220) );
  XNOR2_X1 U11605 ( .A(n9220), .B(n9219), .ZN(n11473) );
  INV_X1 U11606 ( .A(n11473), .ZN(n11464) );
  OR2_X1 U11607 ( .A1(n12056), .A2(SI_9_), .ZN(n9224) );
  XNOR2_X1 U11608 ( .A(n10011), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n9236) );
  XNOR2_X1 U11609 ( .A(n9237), .B(n9236), .ZN(n9955) );
  OR2_X1 U11610 ( .A1(n9244), .A2(n9955), .ZN(n9223) );
  OAI211_X1 U11611 ( .C1(n11464), .C2(n10662), .A(n9224), .B(n9223), .ZN(
        n15165) );
  NAND2_X1 U11612 ( .A1(n12631), .A2(n15165), .ZN(n9225) );
  NAND2_X1 U11613 ( .A1(n11618), .A2(n9225), .ZN(n9227) );
  INV_X1 U11614 ( .A(n12631), .ZN(n11820) );
  INV_X1 U11615 ( .A(n15165), .ZN(n12119) );
  NAND2_X1 U11616 ( .A1(n11820), .A2(n12119), .ZN(n9226) );
  NAND2_X1 U11617 ( .A1(n9227), .A2(n9226), .ZN(n11917) );
  NAND2_X1 U11618 ( .A1(n6574), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U11619 ( .A1(n9228), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11620 ( .A1(n9262), .A2(n9229), .ZN(n11814) );
  NAND2_X1 U11621 ( .A1(n6571), .A2(n11814), .ZN(n9234) );
  INV_X1 U11622 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9230) );
  OR2_X1 U11623 ( .A1(n12061), .A2(n9230), .ZN(n9233) );
  INV_X1 U11624 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9231) );
  OR2_X1 U11625 ( .A1(n12062), .A2(n9231), .ZN(n9232) );
  NAND4_X1 U11626 ( .A1(n9235), .A2(n9234), .A3(n9233), .A4(n9232), .ZN(n12630) );
  NAND2_X1 U11627 ( .A1(n10011), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11628 ( .A1(n10151), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U11629 ( .A1(n10150), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9240) );
  INV_X1 U11630 ( .A(n9241), .ZN(n9242) );
  NAND2_X1 U11631 ( .A1(n6670), .A2(n9242), .ZN(n9243) );
  NAND2_X1 U11632 ( .A1(n9251), .A2(n9243), .ZN(n9983) );
  NAND2_X1 U11633 ( .A1(n9983), .A2(n12055), .ZN(n9248) );
  NAND2_X1 U11634 ( .A1(n9245), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9246) );
  XNOR2_X1 U11635 ( .A(n9246), .B(n7421), .ZN(n11471) );
  NAND2_X1 U11636 ( .A1(n9387), .A2(n11471), .ZN(n9247) );
  OAI211_X1 U11637 ( .C1(SI_10_), .C2(n12056), .A(n9248), .B(n9247), .ZN(
        n15171) );
  NAND2_X1 U11638 ( .A1(n12630), .A2(n15171), .ZN(n12125) );
  NAND2_X1 U11639 ( .A1(n11917), .A2(n12125), .ZN(n9249) );
  INV_X1 U11640 ( .A(n12630), .ZN(n12588) );
  INV_X1 U11641 ( .A(n15171), .ZN(n11823) );
  NAND2_X1 U11642 ( .A1(n12588), .A2(n11823), .ZN(n12126) );
  NAND2_X1 U11643 ( .A1(n9249), .A2(n12126), .ZN(n11668) );
  XNOR2_X1 U11644 ( .A(n10224), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n9252) );
  XNOR2_X1 U11645 ( .A(n9269), .B(n9252), .ZN(n9996) );
  NAND2_X1 U11646 ( .A1(n9996), .A2(n12055), .ZN(n9255) );
  NAND2_X1 U11647 ( .A1(n6711), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9253) );
  XNOR2_X1 U11648 ( .A(n9253), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U11649 ( .A1(n9457), .A2(SI_11_), .B1(n9387), .B2(n11539), .ZN(
        n9254) );
  NAND2_X1 U11650 ( .A1(n9255), .A2(n9254), .ZN(n12587) );
  NAND2_X1 U11651 ( .A1(n6575), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9260) );
  XNOR2_X1 U11652 ( .A(n9262), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U11653 ( .A1(n6571), .A2(n12586), .ZN(n9259) );
  INV_X1 U11654 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9256) );
  OR2_X1 U11655 ( .A1(n12061), .A2(n9256), .ZN(n9258) );
  INV_X1 U11656 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11670) );
  OR2_X1 U11657 ( .A1(n12062), .A2(n11670), .ZN(n9257) );
  NAND4_X1 U11658 ( .A1(n9260), .A2(n9259), .A3(n9258), .A4(n9257), .ZN(n12629) );
  XNOR2_X1 U11659 ( .A(n12587), .B(n12629), .ZN(n12243) );
  NAND2_X1 U11660 ( .A1(n11668), .A2(n12243), .ZN(n11669) );
  NAND2_X1 U11661 ( .A1(n12583), .A2(n12587), .ZN(n12128) );
  NAND2_X1 U11662 ( .A1(n11669), .A2(n12128), .ZN(n11911) );
  NAND2_X1 U11663 ( .A1(n6574), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9267) );
  OAI21_X1 U11664 ( .B1(n9262), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n9263) );
  INV_X1 U11665 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11479) );
  INV_X1 U11666 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U11667 ( .A1(n11479), .A2(n11550), .ZN(n9261) );
  NAND2_X1 U11668 ( .A1(n9263), .A2(n9287), .ZN(n12530) );
  NAND2_X1 U11669 ( .A1(n6571), .A2(n12530), .ZN(n9266) );
  INV_X1 U11670 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n11910) );
  OR2_X1 U11671 ( .A1(n12061), .A2(n11910), .ZN(n9265) );
  INV_X1 U11672 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11926) );
  OR2_X1 U11673 ( .A1(n12062), .A2(n11926), .ZN(n9264) );
  NAND4_X1 U11674 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n12628) );
  NAND2_X1 U11675 ( .A1(n10224), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11676 ( .A1(n10221), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9270) );
  XNOR2_X1 U11677 ( .A(n9280), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n9277) );
  XNOR2_X1 U11678 ( .A(n9279), .B(n9277), .ZN(n10007) );
  NAND2_X1 U11679 ( .A1(n10007), .A2(n12055), .ZN(n9275) );
  OR2_X1 U11680 ( .A1(n9272), .A2(n9056), .ZN(n9273) );
  XNOR2_X1 U11681 ( .A(n9273), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U11682 ( .A1(n9457), .A2(SI_12_), .B1(n9387), .B2(n11897), .ZN(
        n9274) );
  OR2_X1 U11683 ( .A1(n13001), .A2(n12531), .ZN(n12132) );
  NAND2_X1 U11684 ( .A1(n12531), .A2(n13001), .ZN(n12137) );
  NAND2_X1 U11685 ( .A1(n11911), .A2(n12244), .ZN(n9276) );
  INV_X1 U11686 ( .A(n9277), .ZN(n9278) );
  NAND2_X1 U11687 ( .A1(n9280), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9281) );
  XNOR2_X1 U11688 ( .A(n9293), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10154) );
  NAND2_X1 U11689 ( .A1(n10154), .A2(n12055), .ZN(n9286) );
  NAND2_X1 U11690 ( .A1(n9297), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9284) );
  XNOR2_X1 U11691 ( .A(n9284), .B(n9283), .ZN(n12655) );
  AOI22_X1 U11692 ( .A1(n9457), .A2(n15411), .B1(n9387), .B2(n12655), .ZN(
        n9285) );
  NAND2_X1 U11693 ( .A1(n9286), .A2(n9285), .ZN(n13003) );
  NAND2_X1 U11694 ( .A1(n6574), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9292) );
  AND2_X1 U11695 ( .A1(n9287), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9288) );
  OR2_X1 U11696 ( .A1(n9288), .A2(n9302), .ZN(n13005) );
  NAND2_X1 U11697 ( .A1(n6571), .A2(n13005), .ZN(n9291) );
  INV_X1 U11698 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13175) );
  OR2_X1 U11699 ( .A1(n12061), .A2(n13175), .ZN(n9290) );
  INV_X1 U11700 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13007) );
  OR2_X1 U11701 ( .A1(n12062), .A2(n13007), .ZN(n9289) );
  NAND4_X1 U11702 ( .A1(n9292), .A2(n9291), .A3(n9290), .A4(n9289), .ZN(n12984) );
  NOR2_X1 U11703 ( .A1(n13003), .A2(n12984), .ZN(n9617) );
  NAND2_X1 U11704 ( .A1(n13003), .A2(n12984), .ZN(n12142) );
  INV_X1 U11705 ( .A(n12977), .ZN(n9310) );
  INV_X1 U11706 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U11707 ( .A1(n9294), .A2(n10398), .ZN(n9295) );
  XNOR2_X1 U11708 ( .A(n10592), .B(P1_DATAO_REG_14__SCAN_IN), .ZN(n9312) );
  XNOR2_X1 U11709 ( .A(n9314), .B(n9312), .ZN(n10214) );
  NAND2_X1 U11710 ( .A1(n10214), .A2(n12055), .ZN(n9300) );
  NAND2_X1 U11711 ( .A1(n9546), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9298) );
  XNOR2_X1 U11712 ( .A(n9298), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U11713 ( .A1(n9457), .A2(SI_14_), .B1(n9387), .B2(n12660), .ZN(
        n9299) );
  NAND2_X1 U11714 ( .A1(n9300), .A2(n9299), .ZN(n13087) );
  NAND2_X1 U11715 ( .A1(n6574), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9308) );
  INV_X1 U11716 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n9301) );
  NOR2_X1 U11717 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  OR2_X1 U11718 ( .A1(n9322), .A2(n9303), .ZN(n12989) );
  NAND2_X1 U11719 ( .A1(n9141), .A2(n12989), .ZN(n9307) );
  INV_X1 U11720 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n9304) );
  OR2_X1 U11721 ( .A1(n12061), .A2(n9304), .ZN(n9306) );
  INV_X1 U11722 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12641) );
  OR2_X1 U11723 ( .A1(n12062), .A2(n12641), .ZN(n9305) );
  NAND4_X1 U11724 ( .A1(n9308), .A2(n9307), .A3(n9306), .A4(n9305), .ZN(n12969) );
  OR2_X1 U11725 ( .A1(n13087), .A2(n13002), .ZN(n12147) );
  NAND2_X1 U11726 ( .A1(n13087), .A2(n13002), .ZN(n12154) );
  NAND2_X1 U11727 ( .A1(n12147), .A2(n12154), .ZN(n12247) );
  INV_X1 U11728 ( .A(n12247), .ZN(n9309) );
  NAND2_X1 U11729 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  NAND2_X1 U11730 ( .A1(n9311), .A2(n12154), .ZN(n12964) );
  INV_X1 U11731 ( .A(n9312), .ZN(n9313) );
  NAND2_X1 U11732 ( .A1(n10592), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9315) );
  XNOR2_X1 U11733 ( .A(n10844), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n9330) );
  XNOR2_X1 U11734 ( .A(n9332), .B(n9330), .ZN(n14526) );
  NAND2_X1 U11735 ( .A1(n14526), .A2(n12055), .ZN(n9320) );
  OR2_X1 U11736 ( .A1(n7526), .A2(n9056), .ZN(n9318) );
  XNOR2_X1 U11737 ( .A(n9318), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U11738 ( .A1(n9457), .A2(SI_15_), .B1(n9387), .B2(n12688), .ZN(
        n9319) );
  NAND2_X1 U11739 ( .A1(n9320), .A2(n9319), .ZN(n12974) );
  NAND2_X1 U11740 ( .A1(n6575), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9328) );
  INV_X1 U11741 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n9321) );
  NOR2_X1 U11742 ( .A1(n9322), .A2(n9321), .ZN(n9323) );
  OR2_X1 U11743 ( .A1(n9338), .A2(n9323), .ZN(n12973) );
  NAND2_X1 U11744 ( .A1(n6571), .A2(n12973), .ZN(n9327) );
  INV_X1 U11745 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n9324) );
  OR2_X1 U11746 ( .A1(n12061), .A2(n9324), .ZN(n9326) );
  INV_X1 U11747 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12680) );
  OR2_X1 U11748 ( .A1(n12062), .A2(n12680), .ZN(n9325) );
  NAND4_X1 U11749 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(n12983) );
  INV_X1 U11750 ( .A(n12983), .ZN(n12951) );
  OR2_X1 U11751 ( .A1(n12974), .A2(n12951), .ZN(n12146) );
  NAND2_X1 U11752 ( .A1(n12974), .A2(n12951), .ZN(n12153) );
  NAND2_X1 U11753 ( .A1(n12964), .A2(n12965), .ZN(n9329) );
  NAND2_X1 U11754 ( .A1(n9329), .A2(n12153), .ZN(n12954) );
  INV_X1 U11755 ( .A(n9330), .ZN(n9331) );
  NAND2_X1 U11756 ( .A1(n10844), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9333) );
  XNOR2_X1 U11757 ( .A(n10941), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n9345) );
  XNOR2_X1 U11758 ( .A(n9347), .B(n9345), .ZN(n10346) );
  NAND2_X1 U11759 ( .A1(n10346), .A2(n12055), .ZN(n9337) );
  NAND2_X1 U11760 ( .A1(n9349), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9335) );
  XNOR2_X1 U11761 ( .A(n9335), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U11762 ( .A1(n9457), .A2(SI_16_), .B1(n9387), .B2(n12718), .ZN(
        n9336) );
  NAND2_X1 U11763 ( .A1(n6575), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9344) );
  OR2_X1 U11764 ( .A1(n9338), .A2(n15488), .ZN(n9339) );
  NAND2_X1 U11765 ( .A1(n9356), .A2(n9339), .ZN(n12957) );
  NAND2_X1 U11766 ( .A1(n6571), .A2(n12957), .ZN(n9343) );
  INV_X1 U11767 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n9340) );
  OR2_X1 U11768 ( .A1(n12061), .A2(n9340), .ZN(n9342) );
  INV_X1 U11769 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12709) );
  OR2_X1 U11770 ( .A1(n12062), .A2(n12709), .ZN(n9341) );
  NAND4_X1 U11771 ( .A1(n9344), .A2(n9343), .A3(n9342), .A4(n9341), .ZN(n12968) );
  XNOR2_X1 U11772 ( .A(n13079), .B(n12968), .ZN(n12956) );
  INV_X1 U11773 ( .A(n12968), .ZN(n12940) );
  NAND2_X1 U11774 ( .A1(n13079), .A2(n12940), .ZN(n12152) );
  INV_X1 U11775 ( .A(n9345), .ZN(n9346) );
  XNOR2_X1 U11776 ( .A(n15367), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n9348) );
  XNOR2_X1 U11777 ( .A(n9363), .B(n9348), .ZN(n10449) );
  NAND2_X1 U11778 ( .A1(n10449), .A2(n12055), .ZN(n9355) );
  INV_X1 U11779 ( .A(n9383), .ZN(n9365) );
  NAND2_X1 U11780 ( .A1(n9351), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9352) );
  MUX2_X1 U11781 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9352), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9353) );
  AND2_X1 U11782 ( .A1(n9365), .A2(n9353), .ZN(n12730) );
  AOI22_X1 U11783 ( .A1(n9457), .A2(SI_17_), .B1(n12730), .B2(n9387), .ZN(
        n9354) );
  NAND2_X1 U11784 ( .A1(n6574), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11785 ( .A1(n9356), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9357) );
  INV_X1 U11786 ( .A(n9370), .ZN(n9369) );
  NAND2_X1 U11787 ( .A1(n9357), .A2(n9369), .ZN(n12942) );
  NAND2_X1 U11788 ( .A1(n6571), .A2(n12942), .ZN(n9360) );
  INV_X1 U11789 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n15298) );
  OR2_X1 U11790 ( .A1(n12061), .A2(n15298), .ZN(n9359) );
  INV_X1 U11791 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12715) );
  OR2_X1 U11792 ( .A1(n12062), .A2(n12715), .ZN(n9358) );
  NAND4_X1 U11793 ( .A1(n9361), .A2(n9360), .A3(n9359), .A4(n9358), .ZN(n12949) );
  OR2_X1 U11794 ( .A1(n13076), .A2(n12925), .ZN(n12163) );
  NAND2_X1 U11795 ( .A1(n13076), .A2(n12925), .ZN(n12169) );
  INV_X1 U11796 ( .A(n12929), .ZN(n9378) );
  AND2_X1 U11797 ( .A1(n15367), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11798 ( .A1(n11081), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9364) );
  XNOR2_X1 U11799 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .ZN(n9379) );
  XNOR2_X1 U11800 ( .A(n9380), .B(n9379), .ZN(n10508) );
  NAND2_X1 U11801 ( .A1(n10508), .A2(n12055), .ZN(n9368) );
  NAND2_X1 U11802 ( .A1(n9365), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9366) );
  XNOR2_X1 U11803 ( .A(n9366), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U11804 ( .A1(n9387), .A2(n12758), .B1(n9457), .B2(SI_18_), .ZN(
        n9367) );
  NAND2_X1 U11805 ( .A1(n9368), .A2(n9367), .ZN(n12596) );
  NAND2_X1 U11806 ( .A1(n6575), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11807 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(n9369), .ZN(n9372) );
  INV_X1 U11808 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U11809 ( .A1(n9371), .A2(n9370), .ZN(n9392) );
  NAND2_X1 U11810 ( .A1(n9372), .A2(n9392), .ZN(n12931) );
  NAND2_X1 U11811 ( .A1(n6571), .A2(n12931), .ZN(n9375) );
  INV_X1 U11812 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13152) );
  OR2_X1 U11813 ( .A1(n12061), .A2(n13152), .ZN(n9374) );
  INV_X1 U11814 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n15465) );
  OR2_X1 U11815 ( .A1(n12062), .A2(n15465), .ZN(n9373) );
  NAND4_X1 U11816 ( .A1(n9376), .A2(n9375), .A3(n9374), .A4(n9373), .ZN(n12914) );
  NAND2_X1 U11817 ( .A1(n12596), .A2(n12941), .ZN(n12171) );
  NAND2_X1 U11818 ( .A1(n12166), .A2(n12171), .ZN(n12928) );
  INV_X1 U11819 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U11820 ( .A1(n11462), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9381) );
  XNOR2_X1 U11821 ( .A(n11520), .B(P2_DATAO_REG_19__SCAN_IN), .ZN(n9400) );
  XNOR2_X1 U11822 ( .A(n9402), .B(n9400), .ZN(n10536) );
  NAND2_X1 U11823 ( .A1(n10536), .A2(n12055), .ZN(n9389) );
  INV_X1 U11824 ( .A(n9542), .ZN(n9384) );
  NAND2_X1 U11825 ( .A1(n9384), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9385) );
  XNOR2_X2 U11826 ( .A(n9385), .B(n9541), .ZN(n12764) );
  NOR2_X1 U11827 ( .A1(n12056), .A2(SI_19_), .ZN(n9386) );
  AOI21_X1 U11828 ( .B1(n12764), .B2(n9387), .A(n9386), .ZN(n9388) );
  NAND2_X1 U11829 ( .A1(n6575), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9399) );
  INV_X1 U11830 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9391) );
  INV_X1 U11831 ( .A(n9392), .ZN(n9390) );
  NAND2_X1 U11832 ( .A1(n9391), .A2(n9390), .ZN(n9408) );
  NAND2_X1 U11833 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n9392), .ZN(n9393) );
  NAND2_X1 U11834 ( .A1(n9408), .A2(n9393), .ZN(n12919) );
  NAND2_X1 U11835 ( .A1(n9141), .A2(n12919), .ZN(n9398) );
  INV_X1 U11836 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n9394) );
  OR2_X1 U11837 ( .A1(n12061), .A2(n9394), .ZN(n9397) );
  INV_X1 U11838 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n9395) );
  OR2_X1 U11839 ( .A1(n12062), .A2(n9395), .ZN(n9396) );
  NAND4_X1 U11840 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n12900) );
  AND2_X1 U11841 ( .A1(n13066), .A2(n12900), .ZN(n12162) );
  INV_X1 U11842 ( .A(n9400), .ZN(n9401) );
  NAND2_X1 U11843 ( .A1(n11520), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9403) );
  XNOR2_X1 U11844 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .ZN(n9414) );
  XNOR2_X1 U11845 ( .A(n9415), .B(n9414), .ZN(n12322) );
  NAND2_X1 U11846 ( .A1(n12322), .A2(n12055), .ZN(n9405) );
  NAND2_X1 U11847 ( .A1(n9457), .A2(SI_20_), .ZN(n9404) );
  NAND2_X1 U11848 ( .A1(n6574), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9413) );
  INV_X1 U11849 ( .A(n9408), .ZN(n9407) );
  INV_X1 U11850 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U11851 ( .A1(n9408), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U11852 ( .A1(n9419), .A2(n9409), .ZN(n12904) );
  NAND2_X1 U11853 ( .A1(n6571), .A2(n12904), .ZN(n9412) );
  INV_X1 U11854 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13141) );
  OR2_X1 U11855 ( .A1(n12061), .A2(n13141), .ZN(n9411) );
  INV_X1 U11856 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12903) );
  OR2_X1 U11857 ( .A1(n12062), .A2(n12903), .ZN(n9410) );
  NAND4_X1 U11858 ( .A1(n9413), .A2(n9412), .A3(n9411), .A4(n9410), .ZN(n12913) );
  XNOR2_X1 U11859 ( .A(n13142), .B(n12913), .ZN(n12898) );
  INV_X1 U11860 ( .A(n12913), .ZN(n12522) );
  NAND2_X1 U11861 ( .A1(n11529), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9416) );
  XNOR2_X1 U11862 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .ZN(n9426) );
  XNOR2_X1 U11863 ( .A(n9427), .B(n9426), .ZN(n10887) );
  NAND2_X1 U11864 ( .A1(n10887), .A2(n12055), .ZN(n9418) );
  NAND2_X1 U11865 ( .A1(n9457), .A2(SI_21_), .ZN(n9417) );
  NAND2_X1 U11866 ( .A1(n6575), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U11867 ( .A1(n9419), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U11868 ( .A1(n9434), .A2(n9420), .ZN(n12893) );
  NAND2_X1 U11869 ( .A1(n6571), .A2(n12893), .ZN(n9423) );
  INV_X1 U11870 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13135) );
  OR2_X1 U11871 ( .A1(n12061), .A2(n13135), .ZN(n9422) );
  INV_X1 U11872 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12892) );
  OR2_X1 U11873 ( .A1(n12062), .A2(n12892), .ZN(n9421) );
  NAND4_X1 U11874 ( .A1(n9424), .A2(n9423), .A3(n9422), .A4(n9421), .ZN(n12901) );
  INV_X1 U11875 ( .A(n12182), .ZN(n9425) );
  NAND2_X1 U11876 ( .A1(n13136), .A2(n12880), .ZN(n12183) );
  OAI21_X2 U11877 ( .B1(n12887), .B2(n9425), .A(n12183), .ZN(n12876) );
  NAND2_X1 U11878 ( .A1(n11558), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9428) );
  XNOR2_X1 U11879 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .ZN(n9441) );
  XNOR2_X1 U11880 ( .A(n9442), .B(n9441), .ZN(n10938) );
  NAND2_X1 U11881 ( .A1(n10938), .A2(n12055), .ZN(n9431) );
  OR2_X1 U11882 ( .A1(n12056), .A2(n15431), .ZN(n9430) );
  NAND2_X1 U11883 ( .A1(n6574), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9439) );
  INV_X1 U11884 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11885 ( .A1(n9434), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9435) );
  NAND2_X1 U11886 ( .A1(n9447), .A2(n9435), .ZN(n12883) );
  NAND2_X1 U11887 ( .A1(n9141), .A2(n12883), .ZN(n9438) );
  INV_X1 U11888 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13129) );
  OR2_X1 U11889 ( .A1(n12061), .A2(n13129), .ZN(n9437) );
  INV_X1 U11890 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12882) );
  OR2_X1 U11891 ( .A1(n12062), .A2(n12882), .ZN(n9436) );
  NAND4_X1 U11892 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(n12890) );
  NAND2_X1 U11893 ( .A1(n13130), .A2(n12862), .ZN(n12188) );
  INV_X1 U11894 ( .A(n12188), .ZN(n9440) );
  NAND2_X1 U11895 ( .A1(n11617), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9443) );
  XNOR2_X1 U11896 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .ZN(n9453) );
  XNOR2_X1 U11897 ( .A(n9454), .B(n9453), .ZN(n11029) );
  NAND2_X1 U11898 ( .A1(n11029), .A2(n12055), .ZN(n9446) );
  NAND2_X1 U11899 ( .A1(n9457), .A2(SI_23_), .ZN(n9445) );
  NAND2_X1 U11900 ( .A1(n9117), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U11901 ( .A1(n9447), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U11902 ( .A1(n9462), .A2(n9448), .ZN(n12868) );
  NAND2_X1 U11903 ( .A1(n9141), .A2(n12868), .ZN(n9451) );
  INV_X1 U11904 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13125) );
  OR2_X1 U11905 ( .A1(n12061), .A2(n13125), .ZN(n9450) );
  INV_X1 U11906 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12870) );
  OR2_X1 U11907 ( .A1(n12062), .A2(n12870), .ZN(n9449) );
  NAND4_X1 U11908 ( .A1(n9452), .A2(n9451), .A3(n9450), .A4(n9449), .ZN(n12627) );
  NOR2_X1 U11909 ( .A1(n12872), .A2(n12881), .ZN(n12196) );
  NAND2_X1 U11910 ( .A1(n9455), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9456) );
  XNOR2_X1 U11911 ( .A(n9468), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U11912 ( .A1(n11385), .A2(n12055), .ZN(n9459) );
  NAND2_X1 U11913 ( .A1(n9457), .A2(SI_24_), .ZN(n9458) );
  NAND2_X2 U11914 ( .A1(n9459), .A2(n9458), .ZN(n12855) );
  INV_X1 U11915 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U11916 ( .A1(n9462), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11917 ( .A1(n9473), .A2(n9463), .ZN(n12851) );
  NAND2_X1 U11918 ( .A1(n6571), .A2(n12851), .ZN(n9467) );
  NAND2_X1 U11919 ( .A1(n6575), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9466) );
  INV_X1 U11920 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13121) );
  OR2_X1 U11921 ( .A1(n12061), .A2(n13121), .ZN(n9465) );
  INV_X1 U11922 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12853) );
  OR2_X1 U11923 ( .A1(n12062), .A2(n12853), .ZN(n9464) );
  NAND4_X1 U11924 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(n12826) );
  OR2_X1 U11925 ( .A1(n12855), .A2(n12863), .ZN(n12197) );
  NAND2_X1 U11926 ( .A1(n12843), .A2(n12842), .ZN(n12841) );
  NAND2_X1 U11927 ( .A1(n11933), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U11928 ( .A1(n11936), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U11929 ( .A1(n9482), .A2(n9470), .ZN(n9479) );
  XNOR2_X1 U11930 ( .A(n9481), .B(n9479), .ZN(n11559) );
  NAND2_X1 U11931 ( .A1(n11559), .A2(n12055), .ZN(n9472) );
  NAND2_X1 U11932 ( .A1(n9473), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U11933 ( .A1(n9486), .A2(n9474), .ZN(n12833) );
  NAND2_X1 U11934 ( .A1(n6571), .A2(n12833), .ZN(n9478) );
  NAND2_X1 U11935 ( .A1(n9117), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9477) );
  INV_X1 U11936 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13117) );
  OR2_X1 U11937 ( .A1(n12061), .A2(n13117), .ZN(n9476) );
  INV_X1 U11938 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12835) );
  OR2_X1 U11939 ( .A1(n12062), .A2(n12835), .ZN(n9475) );
  NAND4_X1 U11940 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), .ZN(n12626) );
  NAND2_X1 U11941 ( .A1(n12837), .A2(n12847), .ZN(n12192) );
  INV_X1 U11942 ( .A(n9479), .ZN(n9480) );
  NAND2_X1 U11943 ( .A1(n14411), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11944 ( .A1(n13740), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U11945 ( .A1(n9497), .A2(n9483), .ZN(n9494) );
  XNOR2_X1 U11946 ( .A(n9496), .B(n9494), .ZN(n11661) );
  NAND2_X1 U11947 ( .A1(n11661), .A2(n12055), .ZN(n9485) );
  NAND2_X1 U11948 ( .A1(n6574), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9492) );
  NAND2_X1 U11949 ( .A1(n9486), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U11950 ( .A1(n9502), .A2(n9487), .ZN(n12817) );
  NAND2_X1 U11951 ( .A1(n6571), .A2(n12817), .ZN(n9491) );
  INV_X1 U11952 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13113) );
  OR2_X1 U11953 ( .A1(n12061), .A2(n13113), .ZN(n9490) );
  INV_X1 U11954 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n9488) );
  OR2_X1 U11955 ( .A1(n12062), .A2(n9488), .ZN(n9489) );
  NAND2_X1 U11956 ( .A1(n12816), .A2(n12805), .ZN(n12206) );
  INV_X1 U11957 ( .A(n12206), .ZN(n9493) );
  INV_X1 U11958 ( .A(n9494), .ZN(n9495) );
  NAND2_X1 U11959 ( .A1(n14409), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U11960 ( .A1(n13738), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U11961 ( .A1(n9522), .A2(n9498), .ZN(n9519) );
  XNOR2_X1 U11962 ( .A(n9521), .B(n9519), .ZN(n11687) );
  NAND2_X1 U11963 ( .A1(n11687), .A2(n12055), .ZN(n9500) );
  OR2_X1 U11964 ( .A1(n12056), .A2(n15275), .ZN(n9499) );
  NAND2_X1 U11965 ( .A1(n9117), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9508) );
  INV_X1 U11966 ( .A(n9502), .ZN(n9501) );
  INV_X1 U11967 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U11968 ( .A1(n9501), .A2(n15285), .ZN(n9512) );
  NAND2_X1 U11969 ( .A1(n9502), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U11970 ( .A1(n9512), .A2(n9503), .ZN(n12806) );
  NAND2_X1 U11971 ( .A1(n6571), .A2(n12806), .ZN(n9507) );
  INV_X1 U11972 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13109) );
  OR2_X1 U11973 ( .A1(n12061), .A2(n13109), .ZN(n9506) );
  INV_X1 U11974 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9504) );
  OR2_X1 U11975 ( .A1(n12062), .A2(n9504), .ZN(n9505) );
  NAND4_X1 U11976 ( .A1(n9508), .A2(n9507), .A3(n9506), .A4(n9505), .ZN(n12790) );
  NAND2_X1 U11977 ( .A1(n13037), .A2(n12815), .ZN(n12215) );
  INV_X1 U11978 ( .A(n12215), .ZN(n9509) );
  NAND2_X1 U11979 ( .A1(n6575), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9518) );
  INV_X1 U11980 ( .A(n9512), .ZN(n9511) );
  INV_X1 U11981 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U11982 ( .A1(n9511), .A2(n9510), .ZN(n9537) );
  NAND2_X1 U11983 ( .A1(n9512), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9513) );
  NAND2_X1 U11984 ( .A1(n9537), .A2(n9513), .ZN(n12793) );
  NAND2_X1 U11985 ( .A1(n9141), .A2(n12793), .ZN(n9517) );
  INV_X1 U11986 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13105) );
  OR2_X1 U11987 ( .A1(n12061), .A2(n13105), .ZN(n9516) );
  INV_X1 U11988 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9514) );
  OR2_X1 U11989 ( .A1(n9121), .A2(n9514), .ZN(n9515) );
  NAND4_X1 U11990 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n12625) );
  INV_X1 U11991 ( .A(n9519), .ZN(n9520) );
  NAND2_X1 U11992 ( .A1(n14404), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9531) );
  NAND2_X1 U11993 ( .A1(n9524), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U11994 ( .A1(n9531), .A2(n9525), .ZN(n9528) );
  XNOR2_X1 U11995 ( .A(n9530), .B(n9528), .ZN(n12430) );
  NAND2_X1 U11996 ( .A1(n12430), .A2(n12055), .ZN(n9527) );
  OR2_X1 U11997 ( .A1(n12056), .A2(n12433), .ZN(n9526) );
  NAND2_X1 U11998 ( .A1(n13033), .A2(n12804), .ZN(n12221) );
  INV_X1 U11999 ( .A(n9528), .ZN(n9529) );
  NAND2_X1 U12000 ( .A1(n9530), .A2(n9529), .ZN(n9532) );
  AOI22_X1 U12001 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13732), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n14398), .ZN(n9533) );
  INV_X1 U12002 ( .A(n9533), .ZN(n9534) );
  XNOR2_X1 U12003 ( .A(n12044), .B(n9534), .ZN(n13185) );
  NAND2_X1 U12004 ( .A1(n13185), .A2(n12055), .ZN(n9536) );
  OR2_X1 U12005 ( .A1(n12056), .A2(n13188), .ZN(n9535) );
  INV_X1 U12006 ( .A(n9537), .ZN(n9591) );
  NAND2_X1 U12007 ( .A1(n6571), .A2(n9591), .ZN(n12066) );
  OR2_X1 U12008 ( .A1(n12061), .A2(n13099), .ZN(n9540) );
  NAND2_X1 U12009 ( .A1(n9117), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9539) );
  OR2_X1 U12010 ( .A1(n9121), .A2(n9635), .ZN(n9538) );
  NAND2_X1 U12011 ( .A1(n13101), .A2(n12792), .ZN(n12254) );
  NAND2_X1 U12012 ( .A1(n12224), .A2(n12254), .ZN(n9631) );
  XNOR2_X1 U12013 ( .A(n12071), .B(n9631), .ZN(n13103) );
  INV_X1 U12014 ( .A(n12764), .ZN(n12259) );
  OR2_X1 U12015 ( .A1(n10802), .A2(n12259), .ZN(n9549) );
  OAI21_X1 U12016 ( .B1(n9550), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9545) );
  MUX2_X1 U12017 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9545), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9548) );
  OR2_X1 U12018 ( .A1(n9549), .A2(n10936), .ZN(n9587) );
  NAND2_X1 U12019 ( .A1(n9587), .A2(n12213), .ZN(n9560) );
  INV_X1 U12020 ( .A(n9560), .ZN(n9582) );
  XNOR2_X1 U12021 ( .A(n11387), .B(P3_B_REG_SCAN_IN), .ZN(n9555) );
  NAND2_X1 U12022 ( .A1(n9555), .A2(n11560), .ZN(n9557) );
  NAND2_X1 U12023 ( .A1(n6666), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9556) );
  INV_X1 U12024 ( .A(n9573), .ZN(n11662) );
  NAND2_X1 U12025 ( .A1(n11560), .A2(n11662), .ZN(n9558) );
  NAND2_X1 U12026 ( .A1(n12211), .A2(n12229), .ZN(n10786) );
  NAND2_X1 U12027 ( .A1(n10786), .A2(n9560), .ZN(n9650) );
  NAND2_X1 U12028 ( .A1(n9650), .A2(n10780), .ZN(n9581) );
  NAND2_X1 U12029 ( .A1(n11387), .A2(n11662), .ZN(n9561) );
  XNOR2_X1 U12030 ( .A(n10801), .B(n10780), .ZN(n9579) );
  NOR2_X1 U12031 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .ZN(
        n9565) );
  NOR4_X1 U12032 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n9564) );
  NOR4_X1 U12033 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n9563) );
  NOR4_X1 U12034 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n9562) );
  NAND4_X1 U12035 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(n9571)
         );
  NOR4_X1 U12036 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n9569) );
  NOR4_X1 U12037 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9568) );
  NOR4_X1 U12038 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9567) );
  NOR4_X1 U12039 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9566) );
  NAND4_X1 U12040 ( .A1(n9569), .A2(n9568), .A3(n9567), .A4(n9566), .ZN(n9570)
         );
  NOR2_X1 U12041 ( .A1(n9571), .A2(n9570), .ZN(n9572) );
  INV_X1 U12042 ( .A(n11387), .ZN(n9574) );
  NAND2_X1 U12043 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  NAND2_X1 U12044 ( .A1(n6647), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U12045 ( .A1(n10783), .A2(n11073), .ZN(n9578) );
  INV_X1 U12046 ( .A(n9649), .ZN(n9580) );
  OAI211_X1 U12047 ( .C1(n9582), .C2(n10780), .A(n9581), .B(n9580), .ZN(n9590)
         );
  NAND2_X1 U12048 ( .A1(n10802), .A2(n12259), .ZN(n12261) );
  INV_X1 U12049 ( .A(n11073), .ZN(n10664) );
  OR2_X1 U12050 ( .A1(n12261), .A2(n10664), .ZN(n9583) );
  NAND2_X1 U12051 ( .A1(n10777), .A2(n10802), .ZN(n9584) );
  XNOR2_X1 U12052 ( .A(n10936), .B(n9584), .ZN(n9586) );
  AND2_X1 U12053 ( .A1(n10777), .A2(n12764), .ZN(n9585) );
  OR2_X1 U12054 ( .A1(n9586), .A2(n9585), .ZN(n11074) );
  INV_X1 U12055 ( .A(n12229), .ZN(n9646) );
  NAND3_X1 U12056 ( .A1(n11074), .A2(n9646), .A3(n15172), .ZN(n9588) );
  NAND2_X1 U12057 ( .A1(n15124), .A2(n10803), .ZN(n11262) );
  NAND2_X1 U12058 ( .A1(n12867), .A2(n11262), .ZN(n15127) );
  NAND2_X1 U12059 ( .A1(n15155), .A2(n12261), .ZN(n9589) );
  NAND2_X1 U12060 ( .A1(n12990), .A2(n9591), .ZN(n12782) );
  INV_X1 U12061 ( .A(n12782), .ZN(n9592) );
  AOI21_X1 U12062 ( .B1(n13101), .B2(n12991), .A(n9592), .ZN(n9593) );
  INV_X1 U12063 ( .A(n12431), .ZN(n12269) );
  INV_X1 U12064 ( .A(n12733), .ZN(n12754) );
  NAND2_X1 U12065 ( .A1(n12269), .A2(n12754), .ZN(n10679) );
  INV_X1 U12066 ( .A(P3_B_REG_SCAN_IN), .ZN(n9595) );
  NOR2_X2 U12067 ( .A1(n12213), .A2(n10796), .ZN(n15117) );
  OAI21_X1 U12068 ( .B1(n12431), .B2(n9595), .A(n15117), .ZN(n12781) );
  INV_X1 U12069 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n9596) );
  OR2_X1 U12070 ( .A1(n12061), .A2(n9596), .ZN(n9600) );
  NAND2_X1 U12071 ( .A1(n9117), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9599) );
  INV_X1 U12072 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9597) );
  OR2_X1 U12073 ( .A1(n12062), .A2(n9597), .ZN(n9598) );
  INV_X1 U12074 ( .A(n13033), .ZN(n12795) );
  INV_X1 U12075 ( .A(n13130), .ZN(n13057) );
  INV_X1 U12076 ( .A(n12900), .ZN(n12926) );
  NAND2_X1 U12077 ( .A1(n12077), .A2(n6565), .ZN(n15113) );
  INV_X1 U12078 ( .A(n11078), .ZN(n15039) );
  NAND2_X1 U12079 ( .A1(n15110), .A2(n15039), .ZN(n15112) );
  INV_X1 U12080 ( .A(n9601), .ZN(n13014) );
  NAND2_X1 U12081 ( .A1(n13014), .A2(n15122), .ZN(n13017) );
  NAND2_X1 U12082 ( .A1(n15111), .A2(n13017), .ZN(n9602) );
  INV_X1 U12083 ( .A(n13018), .ZN(n12083) );
  NAND2_X1 U12084 ( .A1(n9602), .A2(n12083), .ZN(n13021) );
  NOR2_X1 U12085 ( .A1(n15116), .A2(n13025), .ZN(n11296) );
  NOR2_X1 U12086 ( .A1(n11295), .A2(n11296), .ZN(n9603) );
  NAND2_X1 U12087 ( .A1(n13021), .A2(n9603), .ZN(n11298) );
  NAND2_X1 U12088 ( .A1(n12636), .A2(n11302), .ZN(n9604) );
  NAND2_X1 U12089 ( .A1(n11298), .A2(n9604), .ZN(n11329) );
  INV_X1 U12090 ( .A(n9605), .ZN(n12096) );
  NAND2_X1 U12091 ( .A1(n11329), .A2(n12096), .ZN(n9607) );
  NAND2_X1 U12092 ( .A1(n12635), .A2(n10999), .ZN(n9606) );
  NAND2_X1 U12093 ( .A1(n9607), .A2(n9606), .ZN(n11263) );
  NOR2_X1 U12094 ( .A1(n12634), .A2(n11274), .ZN(n11363) );
  NOR2_X1 U12095 ( .A1(n12233), .A2(n11363), .ZN(n9608) );
  INV_X1 U12096 ( .A(n12235), .ZN(n9609) );
  NAND2_X1 U12097 ( .A1(n11375), .A2(n9609), .ZN(n9611) );
  NAND2_X1 U12098 ( .A1(n12632), .A2(n15154), .ZN(n9610) );
  NAND2_X1 U12099 ( .A1(n9611), .A2(n9610), .ZN(n11607) );
  NAND2_X1 U12100 ( .A1(n12631), .A2(n12119), .ZN(n12120) );
  OAI21_X1 U12101 ( .B1(n12631), .B2(n12119), .A(n12120), .ZN(n12238) );
  NOR2_X1 U12102 ( .A1(n11728), .A2(n11603), .ZN(n11619) );
  NOR2_X1 U12103 ( .A1(n12238), .A2(n11619), .ZN(n9612) );
  OAI21_X1 U12104 ( .B1(n11607), .B2(n12234), .A(n9612), .ZN(n11620) );
  NAND2_X1 U12105 ( .A1(n11620), .A2(n12120), .ZN(n11919) );
  NAND2_X1 U12106 ( .A1(n12126), .A2(n12125), .ZN(n12239) );
  NAND2_X1 U12107 ( .A1(n12630), .A2(n11823), .ZN(n9613) );
  AND2_X1 U12108 ( .A1(n12587), .A2(n12629), .ZN(n9615) );
  INV_X1 U12109 ( .A(n12587), .ZN(n14563) );
  NAND2_X1 U12110 ( .A1(n14563), .A2(n12583), .ZN(n9614) );
  INV_X1 U12111 ( .A(n12244), .ZN(n11906) );
  NAND2_X1 U12112 ( .A1(n12531), .A2(n12628), .ZN(n9616) );
  INV_X1 U12113 ( .A(n9617), .ZN(n12141) );
  NAND2_X1 U12114 ( .A1(n12996), .A2(n12994), .ZN(n12978) );
  INV_X1 U12115 ( .A(n12984), .ZN(n12491) );
  NAND2_X1 U12116 ( .A1(n13003), .A2(n12491), .ZN(n12979) );
  AND2_X1 U12117 ( .A1(n12247), .A2(n12979), .ZN(n9618) );
  NAND2_X1 U12118 ( .A1(n12978), .A2(n9618), .ZN(n12981) );
  NAND2_X1 U12119 ( .A1(n13087), .A2(n12969), .ZN(n9619) );
  NAND2_X1 U12120 ( .A1(n12981), .A2(n9619), .ZN(n12966) );
  AND2_X1 U12121 ( .A1(n12974), .A2(n12983), .ZN(n9620) );
  OR2_X1 U12122 ( .A1(n12974), .A2(n12983), .ZN(n9621) );
  NOR2_X1 U12123 ( .A1(n13079), .A2(n12968), .ZN(n9623) );
  INV_X1 U12124 ( .A(n13079), .ZN(n12959) );
  NAND2_X1 U12125 ( .A1(n13076), .A2(n12949), .ZN(n9624) );
  INV_X1 U12126 ( .A(n12172), .ZN(n9625) );
  OR2_X1 U12127 ( .A1(n12596), .A2(n12914), .ZN(n12908) );
  AND2_X1 U12128 ( .A1(n12231), .A2(n12908), .ZN(n9626) );
  AOI22_X2 U12129 ( .A1(n12899), .A2(n12896), .B1(n12913), .B2(n13142), .ZN(
        n12889) );
  NAND2_X1 U12130 ( .A1(n13136), .A2(n12901), .ZN(n9628) );
  INV_X1 U12131 ( .A(n13136), .ZN(n9627) );
  OAI21_X1 U12132 ( .B1(n12890), .B2(n13130), .A(n12878), .ZN(n9629) );
  OAI21_X1 U12133 ( .B1(n12862), .B2(n13057), .A(n9629), .ZN(n12861) );
  INV_X1 U12134 ( .A(n12860), .ZN(n12252) );
  INV_X1 U12135 ( .A(n12855), .ZN(n13123) );
  NAND2_X1 U12136 ( .A1(n13123), .A2(n12863), .ZN(n12827) );
  AND2_X1 U12137 ( .A1(n12829), .A2(n12827), .ZN(n9630) );
  INV_X1 U12138 ( .A(n12837), .ZN(n13119) );
  INV_X1 U12139 ( .A(n13037), .ZN(n12808) );
  OAI21_X1 U12140 ( .B1(n12804), .B2(n12795), .A(n12788), .ZN(n9632) );
  INV_X1 U12141 ( .A(n10802), .ZN(n10778) );
  AND2_X1 U12142 ( .A1(n10803), .A2(n10778), .ZN(n12267) );
  INV_X1 U12143 ( .A(n12267), .ZN(n9633) );
  OAI222_X1 U12144 ( .A1(n15120), .A2(n12804), .B1(n12781), .B2(n12067), .C1(
        n9645), .C2(n13019), .ZN(n9634) );
  NAND3_X1 U12145 ( .A1(n7543), .A2(n9636), .A3(n7525), .ZN(P3_U3204) );
  NAND2_X1 U12146 ( .A1(n15027), .A2(n14597), .ZN(n13718) );
  INV_X1 U12147 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9639) );
  NOR2_X1 U12148 ( .A1(n15027), .A2(n9639), .ZN(n9640) );
  INV_X1 U12149 ( .A(n10936), .ZN(n12272) );
  AOI22_X1 U12150 ( .A1(n15155), .A2(n10802), .B1(n12272), .B2(n12764), .ZN(
        n9647) );
  OAI21_X1 U12151 ( .B1(n9647), .B2(n9646), .A(n12213), .ZN(n9648) );
  NAND2_X1 U12152 ( .A1(n9648), .A2(n10780), .ZN(n9652) );
  INV_X1 U12153 ( .A(n10780), .ZN(n10785) );
  AOI21_X1 U12154 ( .B1(n9650), .B2(n10785), .A(n9649), .ZN(n9651) );
  NAND2_X1 U12155 ( .A1(n10936), .A2(n15124), .ZN(n15166) );
  INV_X1 U12156 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15464) );
  NAND2_X1 U12157 ( .A1(n7757), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U12158 ( .A1(n7672), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9658) );
  OAI211_X1 U12159 ( .C1(n9660), .C2(n15464), .A(n9659), .B(n9658), .ZN(n14050) );
  NAND2_X1 U12160 ( .A1(n9662), .A2(n9661), .ZN(n9666) );
  INV_X1 U12161 ( .A(n9668), .ZN(n9663) );
  OAI21_X1 U12162 ( .B1(n14050), .B2(n9663), .A(n13891), .ZN(n9669) );
  NAND2_X1 U12163 ( .A1(n12276), .A2(n9675), .ZN(n9665) );
  INV_X1 U12164 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12444) );
  OR2_X1 U12165 ( .A1(n9677), .A2(n12444), .ZN(n9664) );
  NAND2_X1 U12166 ( .A1(n9666), .A2(n9685), .ZN(n9667) );
  MUX2_X1 U12167 ( .A(n9669), .B(n14360), .S(n6578), .Z(n9842) );
  INV_X1 U12168 ( .A(n14360), .ZN(n9858) );
  NAND2_X1 U12169 ( .A1(n9858), .A2(n9835), .ZN(n9674) );
  INV_X1 U12170 ( .A(n14050), .ZN(n9671) );
  OAI21_X1 U12171 ( .B1(n9671), .B2(n9835), .A(n9670), .ZN(n9672) );
  NAND2_X1 U12172 ( .A1(n9672), .A2(n13891), .ZN(n9673) );
  NAND2_X1 U12173 ( .A1(n9674), .A2(n9673), .ZN(n9843) );
  NAND2_X1 U12174 ( .A1(n13722), .A2(n9675), .ZN(n9679) );
  INV_X1 U12175 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9676) );
  OR2_X1 U12176 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  MUX2_X1 U12177 ( .A(n14050), .B(n14047), .S(n9835), .Z(n9681) );
  NOR2_X1 U12178 ( .A1(n14047), .A2(n14050), .ZN(n9680) );
  NAND2_X1 U12179 ( .A1(n9682), .A2(n11532), .ZN(n9683) );
  NAND2_X1 U12180 ( .A1(n9998), .A2(n9683), .ZN(n9684) );
  OR2_X1 U12181 ( .A1(n10259), .A2(n14040), .ZN(n10457) );
  NAND2_X1 U12182 ( .A1(n9684), .A2(n10457), .ZN(n9851) );
  NAND2_X1 U12183 ( .A1(n11644), .A2(n9685), .ZN(n9885) );
  AND2_X1 U12184 ( .A1(n9851), .A2(n9885), .ZN(n9847) );
  NAND2_X1 U12185 ( .A1(n9849), .A2(n9847), .ZN(n9857) );
  INV_X1 U12186 ( .A(n9686), .ZN(n9687) );
  NAND2_X1 U12187 ( .A1(n9691), .A2(n9687), .ZN(n9689) );
  AND2_X1 U12188 ( .A1(n9859), .A2(n10261), .ZN(n9693) );
  MUX2_X1 U12189 ( .A(n9691), .B(n9690), .S(n9835), .Z(n9692) );
  MUX2_X1 U12190 ( .A(n13915), .B(n10463), .S(n9835), .Z(n9695) );
  INV_X1 U12191 ( .A(n9695), .ZN(n9696) );
  NAND3_X1 U12192 ( .A1(n9698), .A2(n10463), .A3(n9697), .ZN(n9699) );
  NAND3_X1 U12193 ( .A1(n9700), .A2(n9699), .A3(n10608), .ZN(n9704) );
  NAND2_X1 U12194 ( .A1(n9827), .A2(n13914), .ZN(n9702) );
  NAND2_X1 U12195 ( .A1(n10896), .A2(n9835), .ZN(n9701) );
  MUX2_X1 U12196 ( .A(n9702), .B(n9701), .S(n10892), .Z(n9703) );
  NAND2_X1 U12197 ( .A1(n9704), .A2(n9703), .ZN(n9707) );
  MUX2_X1 U12198 ( .A(n13913), .B(n10929), .S(n6809), .Z(n9708) );
  NAND2_X1 U12199 ( .A1(n9707), .A2(n9708), .ZN(n9706) );
  MUX2_X1 U12200 ( .A(n10929), .B(n13913), .S(n9835), .Z(n9705) );
  NAND2_X1 U12201 ( .A1(n9706), .A2(n9705), .ZN(n9712) );
  INV_X1 U12202 ( .A(n9707), .ZN(n9710) );
  INV_X1 U12203 ( .A(n9708), .ZN(n9709) );
  NAND2_X1 U12204 ( .A1(n9710), .A2(n9709), .ZN(n9711) );
  MUX2_X1 U12205 ( .A(n10914), .B(n13912), .S(n9835), .Z(n9714) );
  MUX2_X1 U12206 ( .A(n10914), .B(n13912), .S(n6578), .Z(n9713) );
  INV_X1 U12207 ( .A(n9714), .ZN(n9715) );
  MUX2_X1 U12208 ( .A(n13911), .B(n11036), .S(n9835), .Z(n9719) );
  NAND2_X1 U12209 ( .A1(n9718), .A2(n9719), .ZN(n9717) );
  MUX2_X1 U12210 ( .A(n11036), .B(n13911), .S(n9835), .Z(n9716) );
  INV_X1 U12211 ( .A(n9718), .ZN(n9721) );
  INV_X1 U12212 ( .A(n9719), .ZN(n9720) );
  MUX2_X1 U12213 ( .A(n13910), .B(n14702), .S(n6578), .Z(n9723) );
  MUX2_X1 U12214 ( .A(n13910), .B(n14702), .S(n6809), .Z(n9722) );
  INV_X1 U12215 ( .A(n9723), .ZN(n9724) );
  MUX2_X1 U12216 ( .A(n13909), .B(n14745), .S(n6809), .Z(n9728) );
  NAND2_X1 U12217 ( .A1(n9727), .A2(n9728), .ZN(n9726) );
  MUX2_X1 U12218 ( .A(n13909), .B(n14745), .S(n6578), .Z(n9725) );
  INV_X1 U12219 ( .A(n9727), .ZN(n9730) );
  INV_X1 U12220 ( .A(n9728), .ZN(n9729) );
  MUX2_X1 U12221 ( .A(n13908), .B(n11716), .S(n6578), .Z(n9732) );
  MUX2_X1 U12222 ( .A(n13908), .B(n11716), .S(n6809), .Z(n9731) );
  INV_X1 U12223 ( .A(n9732), .ZN(n9733) );
  MUX2_X1 U12224 ( .A(n13907), .B(n11863), .S(n6809), .Z(n9737) );
  NAND2_X1 U12225 ( .A1(n9736), .A2(n9737), .ZN(n9735) );
  MUX2_X1 U12226 ( .A(n13907), .B(n11863), .S(n6578), .Z(n9734) );
  NAND2_X1 U12227 ( .A1(n9735), .A2(n9734), .ZN(n9741) );
  INV_X1 U12228 ( .A(n9736), .ZN(n9739) );
  INV_X1 U12229 ( .A(n9737), .ZN(n9738) );
  NAND2_X1 U12230 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  MUX2_X1 U12231 ( .A(n13906), .B(n11525), .S(n6578), .Z(n9747) );
  MUX2_X1 U12232 ( .A(n13904), .B(n13843), .S(n6578), .Z(n9751) );
  NAND2_X1 U12233 ( .A1(n12328), .A2(n6578), .ZN(n9742) );
  OAI21_X1 U12234 ( .B1(n13843), .B2(n6578), .A(n9742), .ZN(n9743) );
  NOR2_X1 U12235 ( .A1(n9751), .A2(n9743), .ZN(n9744) );
  NOR2_X1 U12236 ( .A1(n11830), .A2(n9744), .ZN(n9758) );
  MUX2_X1 U12237 ( .A(n13840), .B(n14536), .S(n6578), .Z(n9755) );
  MUX2_X1 U12238 ( .A(n13905), .B(n12001), .S(n6809), .Z(n9754) );
  NAND2_X1 U12239 ( .A1(n9755), .A2(n9754), .ZN(n9745) );
  OAI211_X1 U12240 ( .C1(n9748), .C2(n9747), .A(n9758), .B(n9745), .ZN(n9763)
         );
  MUX2_X1 U12241 ( .A(n11998), .B(n12016), .S(n6809), .Z(n9746) );
  AOI21_X1 U12242 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(n9762) );
  NAND2_X1 U12243 ( .A1(n9768), .A2(n9749), .ZN(n9753) );
  MUX2_X1 U12244 ( .A(n13904), .B(n13843), .S(n6809), .Z(n9750) );
  NOR2_X1 U12245 ( .A1(n11830), .A2(n9750), .ZN(n9752) );
  AOI22_X1 U12246 ( .A1(n6578), .A2(n9753), .B1(n9752), .B2(n9751), .ZN(n9760)
         );
  INV_X1 U12247 ( .A(n9754), .ZN(n9757) );
  INV_X1 U12248 ( .A(n9755), .ZN(n9756) );
  NAND3_X1 U12249 ( .A1(n9758), .A2(n9757), .A3(n9756), .ZN(n9759) );
  OAI21_X1 U12250 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9767) );
  AOI21_X1 U12251 ( .B1(n9766), .B2(n9764), .A(n6578), .ZN(n9765) );
  MUX2_X1 U12252 ( .A(n13882), .B(n14344), .S(n6578), .Z(n9770) );
  MUX2_X1 U12253 ( .A(n13901), .B(n11975), .S(n6809), .Z(n9769) );
  MUX2_X1 U12254 ( .A(n13862), .B(n14338), .S(n6578), .Z(n9771) );
  AOI21_X1 U12255 ( .B1(n9774), .B2(n9772), .A(n9771), .ZN(n9776) );
  NOR2_X1 U12256 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  XNOR2_X1 U12257 ( .A(n14332), .B(n6578), .ZN(n9778) );
  XNOR2_X1 U12258 ( .A(n13900), .B(n9835), .ZN(n9777) );
  NAND2_X1 U12259 ( .A1(n9778), .A2(n9777), .ZN(n9779) );
  NAND2_X1 U12260 ( .A1(n9780), .A2(n14227), .ZN(n9784) );
  NAND2_X1 U12261 ( .A1(n14325), .A2(n6578), .ZN(n9782) );
  OR2_X1 U12262 ( .A1(n14325), .A2(n6578), .ZN(n9781) );
  MUX2_X1 U12263 ( .A(n9782), .B(n9781), .S(n14237), .Z(n9783) );
  MUX2_X1 U12264 ( .A(n13899), .B(n14315), .S(n6578), .Z(n9786) );
  MUX2_X1 U12265 ( .A(n13899), .B(n14315), .S(n6809), .Z(n9785) );
  INV_X1 U12266 ( .A(n9786), .ZN(n9787) );
  MUX2_X1 U12267 ( .A(n13898), .B(n14384), .S(n6809), .Z(n9791) );
  NAND2_X1 U12268 ( .A1(n9790), .A2(n9791), .ZN(n9789) );
  MUX2_X1 U12269 ( .A(n13898), .B(n14384), .S(n6578), .Z(n9788) );
  NAND2_X1 U12270 ( .A1(n9789), .A2(n9788), .ZN(n9795) );
  INV_X1 U12271 ( .A(n9790), .ZN(n9793) );
  INV_X1 U12272 ( .A(n9791), .ZN(n9792) );
  NAND2_X1 U12273 ( .A1(n9793), .A2(n9792), .ZN(n9794) );
  MUX2_X1 U12274 ( .A(n13897), .B(n14186), .S(n6578), .Z(n9799) );
  NAND2_X1 U12275 ( .A1(n9798), .A2(n9799), .ZN(n9797) );
  MUX2_X1 U12276 ( .A(n13897), .B(n14186), .S(n6809), .Z(n9796) );
  NAND2_X1 U12277 ( .A1(n9797), .A2(n9796), .ZN(n9803) );
  INV_X1 U12278 ( .A(n9798), .ZN(n9801) );
  INV_X1 U12279 ( .A(n9799), .ZN(n9800) );
  NAND2_X1 U12280 ( .A1(n9801), .A2(n9800), .ZN(n9802) );
  MUX2_X1 U12281 ( .A(n13896), .B(n14172), .S(n6809), .Z(n9804) );
  MUX2_X1 U12282 ( .A(n13896), .B(n14172), .S(n6578), .Z(n9805) );
  MUX2_X1 U12283 ( .A(n13895), .B(n14286), .S(n6578), .Z(n9809) );
  MUX2_X1 U12284 ( .A(n13895), .B(n14286), .S(n6809), .Z(n9806) );
  NAND2_X1 U12285 ( .A1(n9807), .A2(n9806), .ZN(n9813) );
  INV_X1 U12286 ( .A(n9808), .ZN(n9811) );
  INV_X1 U12287 ( .A(n9809), .ZN(n9810) );
  NAND2_X1 U12288 ( .A1(n9811), .A2(n9810), .ZN(n9812) );
  MUX2_X1 U12289 ( .A(n13894), .B(n14135), .S(n6809), .Z(n9814) );
  MUX2_X1 U12290 ( .A(n13894), .B(n14135), .S(n6578), .Z(n9815) );
  MUX2_X1 U12291 ( .A(n14093), .B(n14270), .S(n6578), .Z(n9819) );
  MUX2_X1 U12292 ( .A(n14093), .B(n14270), .S(n6809), .Z(n9816) );
  NAND2_X1 U12293 ( .A1(n9817), .A2(n9816), .ZN(n9823) );
  INV_X1 U12294 ( .A(n9818), .ZN(n9821) );
  INV_X1 U12295 ( .A(n9819), .ZN(n9820) );
  NAND2_X1 U12296 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U12297 ( .A1(n9823), .A2(n9822), .ZN(n9825) );
  MUX2_X1 U12298 ( .A(n13893), .B(n14101), .S(n6809), .Z(n9826) );
  MUX2_X1 U12299 ( .A(n13893), .B(n14101), .S(n6578), .Z(n9824) );
  MUX2_X1 U12300 ( .A(n12457), .B(n14081), .S(n6578), .Z(n9830) );
  MUX2_X1 U12301 ( .A(n14092), .B(n7066), .S(n6809), .Z(n9828) );
  INV_X1 U12302 ( .A(n9830), .ZN(n9831) );
  OR2_X2 U12303 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  MUX2_X1 U12304 ( .A(n13892), .B(n14067), .S(n6809), .Z(n9837) );
  NAND2_X1 U12305 ( .A1(n9836), .A2(n9837), .ZN(n9841) );
  MUX2_X1 U12306 ( .A(n14067), .B(n13892), .S(n9835), .Z(n9840) );
  INV_X1 U12307 ( .A(n9836), .ZN(n9839) );
  INV_X1 U12308 ( .A(n9837), .ZN(n9838) );
  INV_X1 U12309 ( .A(n9842), .ZN(n9852) );
  INV_X1 U12310 ( .A(n9843), .ZN(n9853) );
  XNOR2_X1 U12311 ( .A(n14047), .B(n14050), .ZN(n9881) );
  INV_X1 U12312 ( .A(n9851), .ZN(n9844) );
  NAND2_X1 U12313 ( .A1(n9881), .A2(n9844), .ZN(n9854) );
  INV_X1 U12314 ( .A(n9854), .ZN(n9845) );
  INV_X1 U12315 ( .A(n9881), .ZN(n9848) );
  NAND2_X1 U12316 ( .A1(n9848), .A2(n9847), .ZN(n9850) );
  MUX2_X1 U12317 ( .A(n9851), .B(n9850), .S(n9849), .Z(n9856) );
  OR3_X1 U12318 ( .A1(n9854), .A2(n9853), .A3(n9852), .ZN(n9855) );
  OAI211_X1 U12319 ( .C1(n9857), .C2(n7541), .A(n9856), .B(n9855), .ZN(n9888)
         );
  XNOR2_X1 U12320 ( .A(n9858), .B(n13891), .ZN(n9883) );
  INV_X1 U12321 ( .A(n9859), .ZN(n10774) );
  NOR2_X1 U12322 ( .A1(n10774), .A2(n10452), .ZN(n9862) );
  NAND2_X1 U12323 ( .A1(n9861), .A2(n9860), .ZN(n10521) );
  NAND4_X1 U12324 ( .A1(n9862), .A2(n10497), .A3(n10608), .A4(n10521), .ZN(
        n9863) );
  NOR2_X1 U12325 ( .A1(n9864), .A2(n9863), .ZN(n9867) );
  NAND4_X1 U12326 ( .A1(n9868), .A2(n9867), .A3(n9866), .A4(n9865), .ZN(n9869)
         );
  NOR2_X1 U12327 ( .A1(n11341), .A2(n9869), .ZN(n9870) );
  NAND4_X1 U12328 ( .A1(n11648), .A2(n9870), .A3(n11434), .A4(n11279), .ZN(
        n9871) );
  OR3_X1 U12329 ( .A1(n11830), .A2(n11630), .A3(n9871), .ZN(n9872) );
  NOR2_X1 U12330 ( .A1(n11791), .A2(n9872), .ZN(n9874) );
  AND4_X1 U12331 ( .A1(n14246), .A2(n9874), .A3(n9873), .A4(n12017), .ZN(n9875) );
  NAND4_X1 U12332 ( .A1(n14191), .A2(n9875), .A3(n14208), .A4(n14227), .ZN(
        n9876) );
  NOR2_X1 U12333 ( .A1(n9879), .A2(n9878), .ZN(n9882) );
  XNOR2_X1 U12334 ( .A(n9884), .B(n10460), .ZN(n9887) );
  INV_X1 U12335 ( .A(n9885), .ZN(n9886) );
  NAND2_X1 U12336 ( .A1(n9890), .A2(n9889), .ZN(n9893) );
  INV_X1 U12337 ( .A(n10000), .ZN(n9891) );
  NAND2_X1 U12338 ( .A1(n9891), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11689) );
  INV_X1 U12339 ( .A(n11689), .ZN(n9892) );
  NAND2_X1 U12340 ( .A1(n10059), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14407) );
  OAI21_X1 U12341 ( .B1(n11689), .B2(n8143), .A(P1_B_REG_SCAN_IN), .ZN(n9894)
         );
  INV_X1 U12342 ( .A(n9894), .ZN(n9895) );
  INV_X1 U12343 ( .A(n9989), .ZN(n10002) );
  INV_X1 U12344 ( .A(n9897), .ZN(n9899) );
  NAND2_X1 U12345 ( .A1(n9899), .A2(n9898), .ZN(n10021) );
  INV_X1 U12346 ( .A(n13379), .ZN(P2_U3947) );
  INV_X1 U12347 ( .A(n10016), .ZN(n9900) );
  NAND2_X1 U12348 ( .A1(n9903), .A2(n13574), .ZN(n9907) );
  OR2_X1 U12349 ( .A1(n10241), .A2(n13217), .ZN(n10323) );
  OAI21_X1 U12350 ( .B1(n14997), .B2(n10329), .A(n10323), .ZN(n9904) );
  INV_X1 U12351 ( .A(n9904), .ZN(n9905) );
  INV_X1 U12352 ( .A(n10315), .ZN(n9906) );
  NAND2_X1 U12353 ( .A1(n9907), .A2(n9906), .ZN(n9908) );
  NAND2_X1 U12354 ( .A1(n10316), .A2(n9908), .ZN(n9909) );
  NAND2_X1 U12355 ( .A1(n13381), .A2(n13574), .ZN(n9911) );
  XNOR2_X1 U12356 ( .A(n13217), .B(n10343), .ZN(n9910) );
  XNOR2_X1 U12357 ( .A(n9911), .B(n9910), .ZN(n10317) );
  NAND2_X1 U12358 ( .A1(n9909), .A2(n10317), .ZN(n10322) );
  INV_X1 U12359 ( .A(n9910), .ZN(n9912) );
  NAND2_X1 U12360 ( .A1(n9912), .A2(n9911), .ZN(n9913) );
  XNOR2_X1 U12361 ( .A(n10340), .B(n13217), .ZN(n9914) );
  AND2_X1 U12362 ( .A1(n13380), .A2(n13574), .ZN(n9915) );
  NAND2_X1 U12363 ( .A1(n9914), .A2(n9915), .ZN(n10348) );
  INV_X1 U12364 ( .A(n9914), .ZN(n10356) );
  INV_X1 U12365 ( .A(n9915), .ZN(n9916) );
  NAND2_X1 U12366 ( .A1(n10356), .A2(n9916), .ZN(n9917) );
  NAND2_X1 U12367 ( .A1(n10348), .A2(n9917), .ZN(n9924) );
  NAND2_X1 U12368 ( .A1(n9919), .A2(n9918), .ZN(n9926) );
  INV_X1 U12369 ( .A(n9926), .ZN(n10403) );
  AND2_X1 U12370 ( .A1(n9920), .A2(n14963), .ZN(n9921) );
  AND2_X1 U12371 ( .A1(n10403), .A2(n9921), .ZN(n9934) );
  AND2_X1 U12372 ( .A1(n15018), .A2(n10019), .ZN(n9922) );
  INV_X1 U12373 ( .A(n10350), .ZN(n9923) );
  AOI211_X1 U12374 ( .C1(n9925), .C2(n9924), .A(n13350), .B(n9923), .ZN(n9937)
         );
  OAI21_X1 U12375 ( .B1(n9926), .B2(n14962), .A(n9930), .ZN(n9929) );
  AND2_X1 U12376 ( .A1(n9927), .A2(n10404), .ZN(n9928) );
  NAND2_X1 U12377 ( .A1(n9929), .A2(n9928), .ZN(n10244) );
  MUX2_X1 U12378 ( .A(n13322), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n9936) );
  NOR2_X1 U12379 ( .A1(n14968), .A2(n11528), .ZN(n10414) );
  NAND2_X1 U12380 ( .A1(n9934), .A2(n10414), .ZN(n9932) );
  INV_X1 U12381 ( .A(n9930), .ZN(n9931) );
  INV_X1 U12382 ( .A(n14578), .ZN(n13319) );
  AOI22_X1 U12383 ( .A1(n13316), .A2(n13381), .B1(n13378), .B2(n13315), .ZN(
        n10308) );
  OAI22_X1 U12384 ( .A1(n7193), .A2(n13319), .B1(n13318), .B2(n10308), .ZN(
        n9935) );
  OR3_X1 U12385 ( .A1(n9937), .A2(n9936), .A3(n9935), .ZN(P2_U3190) );
  NAND2_X1 U12386 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), .ZN(
        n9938) );
  OAI21_X1 U12387 ( .B1(n9939), .B2(P3_STATE_REG_SCAN_IN), .A(n9938), .ZN(
        P3_U3295) );
  NAND2_X1 U12388 ( .A1(n9945), .A2(P2_U3088), .ZN(n11696) );
  NAND2_X1 U12389 ( .A1(n9957), .A2(P2_U3088), .ZN(n13729) );
  OAI222_X1 U12390 ( .A1(P2_U3088), .A2(n13382), .B1(n11696), .B2(n9940), .C1(
        n13729), .C2(n9946), .ZN(P2_U3325) );
  OAI222_X1 U12391 ( .A1(P2_U3088), .A2(n14771), .B1(n11696), .B2(n15286), 
        .C1(n13729), .C2(n9948), .ZN(P2_U3326) );
  INV_X1 U12392 ( .A(n10106), .ZN(n13394) );
  OAI222_X1 U12393 ( .A1(P2_U3088), .A2(n13394), .B1(n11696), .B2(n9942), .C1(
        n13729), .C2(n6956), .ZN(P2_U3324) );
  INV_X1 U12394 ( .A(n9943), .ZN(n9950) );
  OAI222_X1 U12395 ( .A1(P2_U3088), .A2(n14783), .B1(n11696), .B2(n9944), .C1(
        n13729), .C2(n9950), .ZN(P2_U3323) );
  INV_X2 U12396 ( .A(n14395), .ZN(n14410) );
  NAND2_X1 U12397 ( .A1(n9945), .A2(P1_U3086), .ZN(n14403) );
  INV_X1 U12398 ( .A(n14403), .ZN(n14405) );
  INV_X1 U12399 ( .A(n14405), .ZN(n14413) );
  OAI222_X1 U12400 ( .A1(P1_U3086), .A2(n13944), .B1(n14410), .B2(n9947), .C1(
        n14413), .C2(n9946), .ZN(P1_U3353) );
  OAI222_X1 U12401 ( .A1(P1_U3086), .A2(n13921), .B1(n14410), .B2(n7023), .C1(
        n14413), .C2(n9948), .ZN(P1_U3354) );
  OAI222_X1 U12402 ( .A1(P1_U3086), .A2(n6954), .B1(n14410), .B2(n9949), .C1(
        n14413), .C2(n6956), .ZN(P1_U3352) );
  INV_X1 U12403 ( .A(n13972), .ZN(n9951) );
  OAI222_X1 U12404 ( .A1(P1_U3086), .A2(n9951), .B1(n14410), .B2(n6928), .C1(
        n14413), .C2(n9950), .ZN(P1_U3351) );
  INV_X1 U12405 ( .A(n10111), .ZN(n14796) );
  OAI222_X1 U12406 ( .A1(P2_U3088), .A2(n14796), .B1(n11696), .B2(n9952), .C1(
        n13729), .C2(n9953), .ZN(P2_U3322) );
  OAI222_X1 U12407 ( .A1(P1_U3086), .A2(n10052), .B1(n14410), .B2(n9954), .C1(
        n14403), .C2(n9953), .ZN(P1_U3350) );
  INV_X2 U12408 ( .A(n13179), .ZN(n11389) );
  INV_X1 U12409 ( .A(n9955), .ZN(n9959) );
  INV_X1 U12410 ( .A(SI_9_), .ZN(n9958) );
  OAI222_X1 U12411 ( .A1(n11389), .A2(n9959), .B1(n11473), .B2(P3_U3151), .C1(
        n9958), .C2(n14525), .ZN(P3_U3286) );
  OAI222_X1 U12412 ( .A1(n14525), .A2(n9961), .B1(n11161), .B2(P3_U3151), .C1(
        n11389), .C2(n9960), .ZN(P3_U3289) );
  OAI222_X1 U12413 ( .A1(n14525), .A2(n7312), .B1(n10979), .B2(P3_U3151), .C1(
        n11389), .C2(n9962), .ZN(P3_U3294) );
  INV_X1 U12414 ( .A(SI_2_), .ZN(n9965) );
  INV_X1 U12415 ( .A(n9963), .ZN(n9964) );
  INV_X1 U12416 ( .A(n10749), .ZN(n10757) );
  OAI222_X1 U12417 ( .A1(n14525), .A2(n9965), .B1(n11389), .B2(n9964), .C1(
        P3_U3151), .C2(n10757), .ZN(P3_U3293) );
  OAI222_X1 U12418 ( .A1(n14525), .A2(n15360), .B1(n11213), .B2(P3_U3151), 
        .C1(n11389), .C2(n9966), .ZN(P3_U3287) );
  INV_X1 U12419 ( .A(n13729), .ZN(n11692) );
  INV_X1 U12420 ( .A(n11692), .ZN(n13741) );
  INV_X1 U12421 ( .A(n11696), .ZN(n13735) );
  AOI22_X1 U12422 ( .A1(n14801), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n13735), .ZN(n9967) );
  OAI21_X1 U12423 ( .B1(n9979), .B2(n13741), .A(n9967), .ZN(P2_U3321) );
  INV_X1 U12424 ( .A(n9968), .ZN(n9969) );
  OAI222_X1 U12425 ( .A1(n11389), .A2(n9969), .B1(n11099), .B2(P3_U3151), .C1(
        n15372), .C2(n14525), .ZN(P3_U3292) );
  INV_X1 U12426 ( .A(n9970), .ZN(n9972) );
  INV_X1 U12427 ( .A(n11127), .ZN(n11092) );
  OAI222_X1 U12428 ( .A1(n11389), .A2(n9972), .B1(n11092), .B2(P3_U3151), .C1(
        n9971), .C2(n14525), .ZN(P3_U3291) );
  INV_X1 U12429 ( .A(n9973), .ZN(n9975) );
  INV_X1 U12430 ( .A(n11164), .ZN(n11159) );
  OAI222_X1 U12431 ( .A1(n11389), .A2(n9975), .B1(n11159), .B2(P3_U3151), .C1(
        n9974), .C2(n14525), .ZN(P3_U3290) );
  INV_X1 U12432 ( .A(n9976), .ZN(n9978) );
  OAI222_X1 U12433 ( .A1(n11389), .A2(n9978), .B1(n11215), .B2(P3_U3151), .C1(
        n9977), .C2(n14525), .ZN(P3_U3288) );
  INV_X1 U12434 ( .A(n10122), .ZN(n10053) );
  OAI222_X1 U12435 ( .A1(P1_U3086), .A2(n10053), .B1(n14410), .B2(n9980), .C1(
        n14403), .C2(n9979), .ZN(P1_U3349) );
  OAI222_X1 U12436 ( .A1(n11389), .A2(n9983), .B1(n11471), .B2(P3_U3151), .C1(
        n9982), .C2(n14525), .ZN(P3_U3285) );
  INV_X1 U12437 ( .A(n14004), .ZN(n10055) );
  OAI222_X1 U12438 ( .A1(P1_U3086), .A2(n10055), .B1(n14410), .B2(n9984), .C1(
        n14403), .C2(n9985), .ZN(P1_U3348) );
  INV_X1 U12439 ( .A(n10115), .ZN(n13406) );
  OAI222_X1 U12440 ( .A1(P2_U3088), .A2(n13406), .B1(n11696), .B2(n9986), .C1(
        n13729), .C2(n9985), .ZN(P2_U3320) );
  NAND2_X1 U12441 ( .A1(n10262), .A2(n9989), .ZN(n10253) );
  INV_X1 U12442 ( .A(n10253), .ZN(n10256) );
  NAND2_X1 U12443 ( .A1(n10256), .A2(n9987), .ZN(n14714) );
  INV_X1 U12444 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9991) );
  INV_X1 U12445 ( .A(n9988), .ZN(n9990) );
  AOI22_X1 U12446 ( .A1(n14714), .A2(n9991), .B1(n9990), .B2(n9989), .ZN(
        P1_U3446) );
  INV_X1 U12447 ( .A(n10138), .ZN(n10083) );
  OAI222_X1 U12448 ( .A1(P2_U3088), .A2(n10083), .B1(n11696), .B2(n9992), .C1(
        n13729), .C2(n9993), .ZN(P2_U3319) );
  INV_X1 U12449 ( .A(n10072), .ZN(n9995) );
  OAI222_X1 U12450 ( .A1(P1_U3086), .A2(n9995), .B1(n14410), .B2(n9994), .C1(
        n14403), .C2(n9993), .ZN(P1_U3347) );
  INV_X1 U12451 ( .A(n9996), .ZN(n9997) );
  INV_X1 U12452 ( .A(n11539), .ZN(n11545) );
  OAI222_X1 U12453 ( .A1(n11389), .A2(n9997), .B1(n11545), .B2(P3_U3151), .C1(
        n15425), .C2(n14525), .ZN(P3_U3284) );
  NAND2_X1 U12454 ( .A1(n10253), .A2(n11689), .ZN(n10043) );
  INV_X1 U12455 ( .A(n9998), .ZN(n10267) );
  AOI21_X1 U12456 ( .B1(n10267), .B2(n10000), .A(n9999), .ZN(n10042) );
  INV_X1 U12457 ( .A(n10042), .ZN(n10001) );
  AND2_X1 U12458 ( .A1(n10043), .A2(n10001), .ZN(n14655) );
  NOR2_X1 U12459 ( .A1(n14655), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12460 ( .A(n14714), .ZN(n14713) );
  OAI22_X1 U12461 ( .A1(n14713), .A2(P1_D_REG_0__SCAN_IN), .B1(n10003), .B2(
        n10002), .ZN(n10004) );
  INV_X1 U12462 ( .A(n10004), .ZN(P1_U3445) );
  INV_X1 U12463 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10006) );
  INV_X1 U12464 ( .A(n10801), .ZN(n10784) );
  NAND2_X1 U12465 ( .A1(n10784), .A2(n10016), .ZN(n10005) );
  OAI21_X1 U12466 ( .B1(n10016), .B2(n10006), .A(n10005), .ZN(P3_U3376) );
  INV_X1 U12467 ( .A(n10007), .ZN(n10009) );
  INV_X1 U12468 ( .A(n11897), .ZN(n11887) );
  OAI222_X1 U12469 ( .A1(n11389), .A2(n10009), .B1(n11887), .B2(P3_U3151), 
        .C1(n10008), .C2(n14525), .ZN(P3_U3283) );
  AND2_X1 U12470 ( .A1(n10080), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12471 ( .A1(n10080), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12472 ( .A1(n10080), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12473 ( .A1(n10080), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12474 ( .A1(n10080), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12475 ( .A1(n10080), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12476 ( .A1(n10080), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12477 ( .A1(n10080), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12478 ( .A1(n10080), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12479 ( .A1(n10080), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12480 ( .A1(n10080), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12481 ( .A1(n10080), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12482 ( .A1(n10080), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12483 ( .A1(n10080), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12484 ( .A1(n10080), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12485 ( .A1(n10080), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12486 ( .A1(n10080), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12487 ( .A1(n10080), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12488 ( .A1(n10080), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12489 ( .A1(n10080), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12490 ( .A1(n10080), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12491 ( .A1(n10080), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12492 ( .A1(n10080), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12493 ( .A1(n10080), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12494 ( .A1(n10080), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  INV_X1 U12495 ( .A(n13735), .ZN(n13739) );
  INV_X1 U12496 ( .A(n10141), .ZN(n10286) );
  OAI222_X1 U12497 ( .A1(n13739), .A2(n10011), .B1(n13729), .B2(n10012), .C1(
        n10286), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U12498 ( .A(n10156), .ZN(n10161) );
  INV_X1 U12499 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10013) );
  OAI222_X1 U12500 ( .A1(P1_U3086), .A2(n10161), .B1(n14410), .B2(n10013), 
        .C1(n14413), .C2(n10012), .ZN(P1_U3346) );
  INV_X1 U12501 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U12502 ( .A1(n10785), .A2(n10016), .ZN(n10014) );
  OAI21_X1 U12503 ( .B1(n10016), .B2(n10015), .A(n10014), .ZN(P3_U3377) );
  OAI21_X1 U12504 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10020) );
  INV_X1 U12505 ( .A(n10032), .ZN(n10028) );
  NOR2_X1 U12506 ( .A1(n10026), .A2(P2_U3088), .ZN(n13734) );
  NAND2_X1 U12507 ( .A1(n10028), .A2(n13734), .ZN(n10022) );
  INV_X1 U12508 ( .A(n10022), .ZN(n10024) );
  NAND2_X1 U12509 ( .A1(n14915), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10025) );
  OAI21_X1 U12510 ( .B1(n8289), .B2(n14883), .A(n10025), .ZN(n10031) );
  INV_X1 U12511 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U12512 ( .A1(n14915), .A2(n10412), .ZN(n10029) );
  AND2_X1 U12513 ( .A1(n10026), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10027) );
  NAND2_X1 U12514 ( .A1(n10028), .A2(n10027), .ZN(n14926) );
  OAI211_X1 U12515 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14883), .A(n10029), .B(
        n14926), .ZN(n10030) );
  MUX2_X1 U12516 ( .A(n10031), .B(n10030), .S(P2_IR_REG_0__SCAN_IN), .Z(n10034) );
  INV_X1 U12517 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15516) );
  INV_X1 U12518 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10411) );
  OAI22_X1 U12519 ( .A1(n14930), .A2(n15516), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10411), .ZN(n10033) );
  OR2_X1 U12520 ( .A1(n10034), .A2(n10033), .ZN(P2_U3214) );
  INV_X1 U12521 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10471) );
  MUX2_X1 U12522 ( .A(n10471), .B(P1_REG2_REG_2__SCAN_IN), .S(n13944), .Z(
        n13941) );
  INV_X1 U12523 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10035) );
  MUX2_X1 U12524 ( .A(n10035), .B(P1_REG2_REG_1__SCAN_IN), .S(n13921), .Z(
        n13920) );
  AND2_X1 U12525 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13931) );
  NAND2_X1 U12526 ( .A1(n13920), .A2(n13931), .ZN(n13919) );
  OAI21_X1 U12527 ( .B1(n10035), .B2(n13921), .A(n13919), .ZN(n13940) );
  NAND2_X1 U12528 ( .A1(n13941), .A2(n13940), .ZN(n13957) );
  INV_X1 U12529 ( .A(n13944), .ZN(n10036) );
  NAND2_X1 U12530 ( .A1(n10036), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13956) );
  INV_X1 U12531 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10618) );
  MUX2_X1 U12532 ( .A(n10618), .B(P1_REG2_REG_3__SCAN_IN), .S(n13950), .Z(
        n13955) );
  AOI21_X1 U12533 ( .B1(n13957), .B2(n13956), .A(n13955), .ZN(n13968) );
  NOR2_X1 U12534 ( .A1(n6954), .A2(n10618), .ZN(n13964) );
  INV_X1 U12535 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n13963) );
  MUX2_X1 U12536 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n13963), .S(n13972), .Z(
        n10037) );
  OAI21_X1 U12537 ( .B1(n13968), .B2(n13964), .A(n10037), .ZN(n13993) );
  NAND2_X1 U12538 ( .A1(n13972), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13992) );
  INV_X1 U12539 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10557) );
  MUX2_X1 U12540 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10557), .S(n10052), .Z(
        n13991) );
  AOI21_X1 U12541 ( .B1(n13993), .B2(n13992), .A(n13991), .ZN(n13990) );
  NOR2_X1 U12542 ( .A1(n10052), .A2(n10557), .ZN(n10127) );
  INV_X1 U12543 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10038) );
  MUX2_X1 U12544 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10038), .S(n10122), .Z(
        n10126) );
  OAI21_X1 U12545 ( .B1(n13990), .B2(n10127), .A(n10126), .ZN(n14014) );
  NAND2_X1 U12546 ( .A1(n10122), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14013) );
  MUX2_X1 U12547 ( .A(n14700), .B(P1_REG2_REG_7__SCAN_IN), .S(n14004), .Z(
        n14012) );
  AOI21_X1 U12548 ( .B1(n14014), .B2(n14013), .A(n14012), .ZN(n14011) );
  NOR2_X1 U12549 ( .A1(n10055), .A2(n14700), .ZN(n10071) );
  INV_X1 U12550 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10986) );
  MUX2_X1 U12551 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10986), .S(n10072), .Z(
        n10039) );
  OAI21_X1 U12552 ( .B1(n14011), .B2(n10071), .A(n10039), .ZN(n10075) );
  NAND2_X1 U12553 ( .A1(n10072), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10041) );
  INV_X1 U12554 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10160) );
  MUX2_X1 U12555 ( .A(n10160), .B(P1_REG2_REG_9__SCAN_IN), .S(n10156), .Z(
        n10040) );
  AOI21_X1 U12556 ( .B1(n10075), .B2(n10041), .A(n10040), .ZN(n10164) );
  NAND3_X1 U12557 ( .A1(n10075), .A2(n10041), .A3(n10040), .ZN(n10045) );
  NAND2_X1 U12558 ( .A1(n10043), .A2(n10042), .ZN(n14657) );
  OR2_X1 U12559 ( .A1(n14401), .A2(n6586), .ZN(n10044) );
  NAND2_X1 U12560 ( .A1(n10045), .A2(n14038), .ZN(n10066) );
  INV_X1 U12561 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14005) );
  INV_X1 U12562 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10046) );
  MUX2_X1 U12563 ( .A(n10046), .B(P1_REG1_REG_2__SCAN_IN), .S(n13944), .Z(
        n13939) );
  INV_X1 U12564 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n13922) );
  MUX2_X1 U12565 ( .A(n13922), .B(P1_REG1_REG_1__SCAN_IN), .S(n13921), .Z(
        n10048) );
  AND2_X1 U12566 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10047) );
  NAND2_X1 U12567 ( .A1(n10048), .A2(n10047), .ZN(n13925) );
  OAI21_X1 U12568 ( .B1(n13922), .B2(n13921), .A(n13925), .ZN(n13938) );
  NAND2_X1 U12569 ( .A1(n13939), .A2(n13938), .ZN(n13953) );
  OR2_X1 U12570 ( .A1(n13944), .A2(n10046), .ZN(n13952) );
  NAND2_X1 U12571 ( .A1(n13953), .A2(n13952), .ZN(n10051) );
  INV_X1 U12572 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10049) );
  MUX2_X1 U12573 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10049), .S(n13950), .Z(
        n10050) );
  NAND2_X1 U12574 ( .A1(n10051), .A2(n10050), .ZN(n13976) );
  NAND2_X1 U12575 ( .A1(n13950), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13975) );
  INV_X1 U12576 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14755) );
  MUX2_X1 U12577 ( .A(n14755), .B(P1_REG1_REG_4__SCAN_IN), .S(n13972), .Z(
        n13974) );
  AOI21_X1 U12578 ( .B1(n13976), .B2(n13975), .A(n13974), .ZN(n13973) );
  AOI21_X1 U12579 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n13972), .A(n13973), .ZN(
        n13987) );
  INV_X1 U12580 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15385) );
  MUX2_X1 U12581 ( .A(n15385), .B(P1_REG1_REG_5__SCAN_IN), .S(n10052), .Z(
        n13988) );
  NAND2_X1 U12582 ( .A1(n13987), .A2(n13988), .ZN(n13986) );
  OAI21_X1 U12583 ( .B1(n13985), .B2(P1_REG1_REG_5__SCAN_IN), .A(n13986), .ZN(
        n10125) );
  INV_X1 U12584 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10703) );
  MUX2_X1 U12585 ( .A(n10703), .B(P1_REG1_REG_6__SCAN_IN), .S(n10122), .Z(
        n10124) );
  NOR2_X1 U12586 ( .A1(n10125), .A2(n10124), .ZN(n14010) );
  NOR2_X1 U12587 ( .A1(n10053), .A2(n10703), .ZN(n14003) );
  MUX2_X1 U12588 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14005), .S(n14004), .Z(
        n10054) );
  OAI21_X1 U12589 ( .B1(n14010), .B2(n14003), .A(n10054), .ZN(n14008) );
  OAI21_X1 U12590 ( .B1(n14005), .B2(n10055), .A(n14008), .ZN(n10068) );
  INV_X1 U12591 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10056) );
  MUX2_X1 U12592 ( .A(n10056), .B(P1_REG1_REG_8__SCAN_IN), .S(n10072), .Z(
        n10069) );
  NOR2_X1 U12593 ( .A1(n10068), .A2(n10069), .ZN(n10067) );
  NOR2_X1 U12594 ( .A1(n10072), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10057) );
  INV_X1 U12595 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15447) );
  MUX2_X1 U12596 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15447), .S(n10156), .Z(
        n10058) );
  OAI21_X1 U12597 ( .B1(n10067), .B2(n10057), .A(n10058), .ZN(n10155) );
  INV_X1 U12598 ( .A(n10155), .ZN(n10061) );
  NOR3_X1 U12599 ( .A1(n10067), .A2(n10058), .A3(n10057), .ZN(n10060) );
  OR2_X1 U12600 ( .A1(n14657), .A2(n10059), .ZN(n14689) );
  INV_X1 U12601 ( .A(n14689), .ZN(n14037) );
  OAI21_X1 U12602 ( .B1(n10061), .B2(n10060), .A(n14037), .ZN(n10065) );
  INV_X1 U12603 ( .A(n14655), .ZN(n14695) );
  INV_X1 U12604 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14436) );
  NAND2_X1 U12605 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10062) );
  OAI21_X1 U12606 ( .B1(n14695), .B2(n14436), .A(n10062), .ZN(n10063) );
  AOI21_X1 U12607 ( .B1(n10156), .B2(n14002), .A(n10063), .ZN(n10064) );
  OAI211_X1 U12608 ( .C1(n10164), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        P1_U3252) );
  AOI21_X1 U12609 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n10079) );
  INV_X1 U12610 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15296) );
  NAND2_X1 U12611 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11573) );
  OAI21_X1 U12612 ( .B1(n14695), .B2(n15296), .A(n11573), .ZN(n10070) );
  AOI21_X1 U12613 ( .B1(n10072), .B2(n14002), .A(n10070), .ZN(n10078) );
  INV_X1 U12614 ( .A(n10071), .ZN(n10074) );
  MUX2_X1 U12615 ( .A(n10986), .B(P1_REG2_REG_8__SCAN_IN), .S(n10072), .Z(
        n10073) );
  NAND2_X1 U12616 ( .A1(n10074), .A2(n10073), .ZN(n10076) );
  OAI211_X1 U12617 ( .C1(n14011), .C2(n10076), .A(n10075), .B(n14038), .ZN(
        n10077) );
  OAI211_X1 U12618 ( .C1(n10079), .C2(n14689), .A(n10078), .B(n10077), .ZN(
        P1_U3251) );
  INV_X1 U12619 ( .A(n10080), .ZN(n10081) );
  INV_X1 U12620 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n15370) );
  NOR2_X1 U12621 ( .A1(n10081), .A2(n15370), .ZN(P3_U3244) );
  INV_X1 U12622 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U12623 ( .A1(n10081), .A2(n15341), .ZN(P3_U3242) );
  INV_X1 U12624 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15413) );
  NOR2_X1 U12625 ( .A1(n10081), .A2(n15413), .ZN(P3_U3253) );
  INV_X1 U12626 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n15366) );
  NOR2_X1 U12627 ( .A1(n10081), .A2(n15366), .ZN(P3_U3263) );
  INV_X1 U12628 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n15473) );
  NOR2_X1 U12629 ( .A1(n10081), .A2(n15473), .ZN(P3_U3252) );
  NAND2_X1 U12630 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10082) );
  OAI21_X1 U12631 ( .B1(n14926), .B2(n10083), .A(n10082), .ZN(n10099) );
  INV_X1 U12632 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U12633 ( .A(n10084), .B(P2_REG1_REG_1__SCAN_IN), .S(n14771), .Z(
        n14763) );
  AND2_X1 U12634 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14762) );
  NAND2_X1 U12635 ( .A1(n14763), .A2(n14762), .ZN(n14761) );
  INV_X1 U12636 ( .A(n14771), .ZN(n10101) );
  NAND2_X1 U12637 ( .A1(n10101), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U12638 ( .A1(n14761), .A2(n10085), .ZN(n13388) );
  INV_X1 U12639 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10086) );
  MUX2_X1 U12640 ( .A(n10086), .B(P2_REG1_REG_2__SCAN_IN), .S(n13382), .Z(
        n13389) );
  NAND2_X1 U12641 ( .A1(n13388), .A2(n13389), .ZN(n13387) );
  INV_X1 U12642 ( .A(n13382), .ZN(n10103) );
  NAND2_X1 U12643 ( .A1(n10103), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12644 ( .A1(n13387), .A2(n10087), .ZN(n13397) );
  INV_X1 U12645 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10088) );
  MUX2_X1 U12646 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10088), .S(n10106), .Z(
        n13398) );
  NAND2_X1 U12647 ( .A1(n13397), .A2(n13398), .ZN(n13396) );
  NAND2_X1 U12648 ( .A1(n10106), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U12649 ( .A1(n13396), .A2(n10089), .ZN(n14779) );
  XNOR2_X1 U12650 ( .A(n14783), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n14780) );
  NAND2_X1 U12651 ( .A1(n14779), .A2(n14780), .ZN(n14778) );
  NAND2_X1 U12652 ( .A1(n10108), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U12653 ( .A1(n14778), .A2(n10090), .ZN(n14792) );
  INV_X1 U12654 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10091) );
  XNOR2_X1 U12655 ( .A(n10111), .B(n10091), .ZN(n14793) );
  NAND2_X1 U12656 ( .A1(n14792), .A2(n14793), .ZN(n14791) );
  NAND2_X1 U12657 ( .A1(n10111), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U12658 ( .A1(n14791), .A2(n10092), .ZN(n14803) );
  INV_X1 U12659 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15443) );
  MUX2_X1 U12660 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15443), .S(n14801), .Z(
        n14804) );
  NAND2_X1 U12661 ( .A1(n14803), .A2(n14804), .ZN(n14802) );
  NAND2_X1 U12662 ( .A1(n14801), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U12663 ( .A1(n14802), .A2(n10093), .ZN(n13412) );
  INV_X1 U12664 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15444) );
  MUX2_X1 U12665 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15444), .S(n10115), .Z(
        n13413) );
  NAND2_X1 U12666 ( .A1(n13412), .A2(n13413), .ZN(n13411) );
  NAND2_X1 U12667 ( .A1(n10115), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10094) );
  NAND2_X1 U12668 ( .A1(n13411), .A2(n10094), .ZN(n10096) );
  INV_X1 U12669 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15032) );
  MUX2_X1 U12670 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15032), .S(n10138), .Z(
        n10095) );
  NAND2_X1 U12671 ( .A1(n10096), .A2(n10095), .ZN(n10140) );
  OAI211_X1 U12672 ( .C1(n10096), .C2(n10095), .A(n10140), .B(n14922), .ZN(
        n10097) );
  INV_X1 U12673 ( .A(n10097), .ZN(n10098) );
  AOI211_X1 U12674 ( .C1(n14760), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10099), .B(
        n10098), .ZN(n10121) );
  INV_X1 U12675 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10580) );
  MUX2_X1 U12676 ( .A(n10580), .B(P2_REG2_REG_1__SCAN_IN), .S(n14771), .Z(
        n14764) );
  AND2_X1 U12677 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10100) );
  NAND2_X1 U12678 ( .A1(n14764), .A2(n10100), .ZN(n14768) );
  NAND2_X1 U12679 ( .A1(n10101), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U12680 ( .A1(n14768), .A2(n10102), .ZN(n13385) );
  INV_X1 U12681 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n14947) );
  MUX2_X1 U12682 ( .A(n14947), .B(P2_REG2_REG_2__SCAN_IN), .S(n13382), .Z(
        n13386) );
  NAND2_X1 U12683 ( .A1(n13385), .A2(n13386), .ZN(n13384) );
  NAND2_X1 U12684 ( .A1(n10103), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U12685 ( .A1(n13384), .A2(n10104), .ZN(n13400) );
  INV_X1 U12686 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10105) );
  MUX2_X1 U12687 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10105), .S(n10106), .Z(
        n13401) );
  NAND2_X1 U12688 ( .A1(n13400), .A2(n13401), .ZN(n13399) );
  NAND2_X1 U12689 ( .A1(n10106), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U12690 ( .A1(n13399), .A2(n10107), .ZN(n14776) );
  XNOR2_X1 U12691 ( .A(n14783), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n14777) );
  NAND2_X1 U12692 ( .A1(n14776), .A2(n14777), .ZN(n14775) );
  NAND2_X1 U12693 ( .A1(n10108), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U12694 ( .A1(n14775), .A2(n10109), .ZN(n14789) );
  INV_X1 U12695 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10110) );
  XNOR2_X1 U12696 ( .A(n10111), .B(n10110), .ZN(n14790) );
  NAND2_X1 U12697 ( .A1(n14789), .A2(n14790), .ZN(n14788) );
  NAND2_X1 U12698 ( .A1(n10111), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10112) );
  NAND2_X1 U12699 ( .A1(n14788), .A2(n10112), .ZN(n14806) );
  INV_X1 U12700 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10549) );
  XNOR2_X1 U12701 ( .A(n14801), .B(n10549), .ZN(n14807) );
  NAND2_X1 U12702 ( .A1(n14806), .A2(n14807), .ZN(n14805) );
  NAND2_X1 U12703 ( .A1(n14801), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U12704 ( .A1(n14805), .A2(n10113), .ZN(n13409) );
  INV_X1 U12705 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10114) );
  MUX2_X1 U12706 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10114), .S(n10115), .Z(
        n13410) );
  NAND2_X1 U12707 ( .A1(n13409), .A2(n13410), .ZN(n13408) );
  NAND2_X1 U12708 ( .A1(n10115), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10116) );
  NAND2_X1 U12709 ( .A1(n13408), .A2(n10116), .ZN(n10119) );
  INV_X1 U12710 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10117) );
  MUX2_X1 U12711 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10117), .S(n10138), .Z(
        n10118) );
  NAND2_X1 U12712 ( .A1(n10119), .A2(n10118), .ZN(n10134) );
  OAI211_X1 U12713 ( .C1(n10119), .C2(n10118), .A(n10134), .B(n14915), .ZN(
        n10120) );
  NAND2_X1 U12714 ( .A1(n10121), .A2(n10120), .ZN(P2_U3222) );
  INV_X1 U12715 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14429) );
  NAND2_X1 U12716 ( .A1(n14002), .A2(n10122), .ZN(n10123) );
  NAND2_X1 U12717 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11040) );
  OAI211_X1 U12718 ( .C1(n14429), .C2(n14695), .A(n10123), .B(n11040), .ZN(
        n10132) );
  AOI211_X1 U12719 ( .C1(n10125), .C2(n10124), .A(n14010), .B(n14689), .ZN(
        n10131) );
  INV_X1 U12720 ( .A(n14014), .ZN(n10129) );
  NOR3_X1 U12721 ( .A1(n13990), .A2(n10127), .A3(n10126), .ZN(n10128) );
  NOR3_X1 U12722 ( .A1(n14687), .A2(n10129), .A3(n10128), .ZN(n10130) );
  OR3_X1 U12723 ( .A1(n10132), .A2(n10131), .A3(n10130), .ZN(P1_U3249) );
  XNOR2_X1 U12724 ( .A(n10141), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U12725 ( .A1(n10138), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U12726 ( .A1(n10134), .A2(n10133), .ZN(n10136) );
  INV_X1 U12727 ( .A(n10288), .ZN(n10135) );
  AOI21_X1 U12728 ( .B1(n10137), .B2(n10136), .A(n10135), .ZN(n10148) );
  INV_X1 U12729 ( .A(n14915), .ZN(n14887) );
  NAND2_X1 U12730 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10878) );
  OAI21_X1 U12731 ( .B1(n14926), .B2(n10286), .A(n10878), .ZN(n10146) );
  NAND2_X1 U12732 ( .A1(n10138), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U12733 ( .A1(n10140), .A2(n10139), .ZN(n10143) );
  MUX2_X1 U12734 ( .A(n10277), .B(P2_REG1_REG_9__SCAN_IN), .S(n10141), .Z(
        n10142) );
  NAND2_X1 U12735 ( .A1(n10143), .A2(n10142), .ZN(n10144) );
  AOI21_X1 U12736 ( .B1(n10279), .B2(n10144), .A(n14883), .ZN(n10145) );
  AOI211_X1 U12737 ( .C1(n14760), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10146), .B(
        n10145), .ZN(n10147) );
  OAI21_X1 U12738 ( .B1(n10148), .B2(n14887), .A(n10147), .ZN(P2_U3223) );
  INV_X1 U12739 ( .A(n10289), .ZN(n14824) );
  INV_X1 U12740 ( .A(n10149), .ZN(n10152) );
  OAI222_X1 U12741 ( .A1(n14824), .A2(P2_U3088), .B1(n13741), .B2(n10152), 
        .C1(n10150), .C2(n13739), .ZN(P2_U3317) );
  INV_X1 U12742 ( .A(n10178), .ZN(n10153) );
  OAI222_X1 U12743 ( .A1(n10153), .A2(P1_U3086), .B1(n14403), .B2(n10152), 
        .C1(n10151), .C2(n14410), .ZN(P1_U3345) );
  OAI222_X1 U12744 ( .A1(n11389), .A2(n10154), .B1(n12655), .B2(P3_U3151), 
        .C1(n15411), .C2(n14525), .ZN(P3_U3282) );
  OAI21_X1 U12745 ( .B1(n10156), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10155), .ZN(
        n10159) );
  INV_X1 U12746 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10157) );
  MUX2_X1 U12747 ( .A(n10157), .B(P1_REG1_REG_10__SCAN_IN), .S(n10178), .Z(
        n10158) );
  NOR2_X1 U12748 ( .A1(n10159), .A2(n10158), .ZN(n10177) );
  AOI211_X1 U12749 ( .C1(n10159), .C2(n10158), .A(n14689), .B(n10177), .ZN(
        n10170) );
  NOR2_X1 U12750 ( .A1(n10161), .A2(n10160), .ZN(n10163) );
  INV_X1 U12751 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11284) );
  MUX2_X1 U12752 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11284), .S(n10178), .Z(
        n10162) );
  OAI21_X1 U12753 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(n10174) );
  INV_X1 U12754 ( .A(n10174), .ZN(n10166) );
  NOR3_X1 U12755 ( .A1(n10164), .A2(n10163), .A3(n10162), .ZN(n10165) );
  NOR3_X1 U12756 ( .A1(n10166), .A2(n10165), .A3(n14687), .ZN(n10169) );
  INV_X1 U12757 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15476) );
  NAND2_X1 U12758 ( .A1(n14002), .A2(n10178), .ZN(n10167) );
  NAND2_X1 U12759 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11858)
         );
  OAI211_X1 U12760 ( .C1(n15476), .C2(n14695), .A(n10167), .B(n11858), .ZN(
        n10168) );
  OR3_X1 U12761 ( .A1(n10170), .A2(n10169), .A3(n10168), .ZN(P1_U3253) );
  NAND2_X1 U12762 ( .A1(n10178), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10173) );
  INV_X1 U12763 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10171) );
  MUX2_X1 U12764 ( .A(n10171), .B(P1_REG2_REG_11__SCAN_IN), .S(n10219), .Z(
        n10172) );
  AOI21_X1 U12765 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(n10205) );
  NAND3_X1 U12766 ( .A1(n10174), .A2(n10173), .A3(n10172), .ZN(n10175) );
  NAND2_X1 U12767 ( .A1(n10175), .A2(n14038), .ZN(n10185) );
  INV_X1 U12768 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10176) );
  MUX2_X1 U12769 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10176), .S(n10219), .Z(
        n10180) );
  AOI21_X1 U12770 ( .B1(n10178), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10177), 
        .ZN(n10179) );
  NAND2_X1 U12771 ( .A1(n10179), .A2(n10180), .ZN(n10203) );
  OAI21_X1 U12772 ( .B1(n10180), .B2(n10179), .A(n10203), .ZN(n10181) );
  NAND2_X1 U12773 ( .A1(n10181), .A2(n14037), .ZN(n10184) );
  INV_X1 U12774 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14439) );
  NAND2_X1 U12775 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12009)
         );
  OAI21_X1 U12776 ( .B1(n14695), .B2(n14439), .A(n12009), .ZN(n10182) );
  AOI21_X1 U12777 ( .B1(n10219), .B2(n14002), .A(n10182), .ZN(n10183) );
  OAI211_X1 U12778 ( .C1(n10205), .C2(n10185), .A(n10184), .B(n10183), .ZN(
        P1_U3254) );
  NAND2_X1 U12779 ( .A1(n6757), .A2(n10186), .ZN(n10187) );
  NAND2_X1 U12780 ( .A1(n10188), .A2(n10187), .ZN(n10586) );
  AOI21_X1 U12781 ( .B1(n10241), .B2(n10337), .A(n13202), .ZN(n10189) );
  AND2_X1 U12782 ( .A1(n10189), .A2(n10231), .ZN(n10581) );
  OAI21_X1 U12783 ( .B1(n10192), .B2(n6757), .A(n10190), .ZN(n10193) );
  NAND2_X1 U12784 ( .A1(n10193), .A2(n14992), .ZN(n10194) );
  AOI22_X1 U12785 ( .A1(n13381), .A2(n13315), .B1(n13316), .B2(n8750), .ZN(
        n10327) );
  NAND2_X1 U12786 ( .A1(n10194), .A2(n10327), .ZN(n10579) );
  AOI211_X1 U12787 ( .C1(n15024), .C2(n10586), .A(n10581), .B(n10579), .ZN(
        n10339) );
  INV_X1 U12788 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10195) );
  OAI22_X1 U12789 ( .A1(n13718), .A2(n10584), .B1(n15027), .B2(n10195), .ZN(
        n10196) );
  INV_X1 U12790 ( .A(n10196), .ZN(n10197) );
  OAI21_X1 U12791 ( .B1(n10339), .B2(n15025), .A(n10197), .ZN(P2_U3433) );
  INV_X1 U12792 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U12793 ( .A1(n15116), .A2(P3_U3897), .ZN(n10198) );
  OAI21_X1 U12794 ( .B1(P3_U3897), .B2(n10199), .A(n10198), .ZN(P3_U3493) );
  OR2_X1 U12795 ( .A1(n10219), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10201) );
  MUX2_X1 U12796 ( .A(n10200), .B(P1_REG1_REG_12__SCAN_IN), .S(n10482), .Z(
        n10202) );
  AOI21_X1 U12797 ( .B1(n10203), .B2(n10201), .A(n10202), .ZN(n10475) );
  AND3_X1 U12798 ( .A1(n10203), .A2(n10202), .A3(n10201), .ZN(n10204) );
  OAI21_X1 U12799 ( .B1(n10475), .B2(n10204), .A(n14037), .ZN(n10213) );
  MUX2_X1 U12800 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11653), .S(n10482), .Z(
        n10207) );
  AOI21_X1 U12801 ( .B1(n10219), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10205), 
        .ZN(n10206) );
  NAND2_X1 U12802 ( .A1(n10206), .A2(n10207), .ZN(n10481) );
  OAI21_X1 U12803 ( .B1(n10207), .B2(n10206), .A(n10481), .ZN(n10211) );
  INV_X1 U12804 ( .A(n10482), .ZN(n10476) );
  NOR2_X1 U12805 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11996), .ZN(n10208) );
  AOI21_X1 U12806 ( .B1(n14655), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10208), 
        .ZN(n10209) );
  OAI21_X1 U12807 ( .B1(n14691), .B2(n10476), .A(n10209), .ZN(n10210) );
  AOI21_X1 U12808 ( .B1(n10211), .B2(n14038), .A(n10210), .ZN(n10212) );
  NAND2_X1 U12809 ( .A1(n10213), .A2(n10212), .ZN(P1_U3255) );
  INV_X1 U12810 ( .A(SI_14_), .ZN(n10216) );
  INV_X1 U12811 ( .A(n12660), .ZN(n12642) );
  INV_X1 U12812 ( .A(n10214), .ZN(n10215) );
  INV_X1 U12813 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12814 ( .A1(n12900), .A2(P3_U3897), .ZN(n10217) );
  OAI21_X1 U12815 ( .B1(P3_U3897), .B2(n10218), .A(n10217), .ZN(P3_U3510) );
  INV_X1 U12816 ( .A(n10219), .ZN(n10222) );
  INV_X1 U12817 ( .A(n10220), .ZN(n10223) );
  OAI222_X1 U12818 ( .A1(P1_U3086), .A2(n10222), .B1(n14410), .B2(n10221), 
        .C1(n14413), .C2(n10223), .ZN(P1_U3344) );
  INV_X1 U12819 ( .A(n10291), .ZN(n14833) );
  OAI222_X1 U12820 ( .A1(P2_U3088), .A2(n14833), .B1(n11696), .B2(n10224), 
        .C1(n13729), .C2(n10223), .ZN(P2_U3316) );
  INV_X1 U12821 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U12822 ( .A1(n12890), .A2(P3_U3897), .ZN(n10225) );
  OAI21_X1 U12823 ( .B1(P3_U3897), .B2(n10226), .A(n10225), .ZN(P3_U3513) );
  OAI21_X1 U12824 ( .B1(n10229), .B2(n10228), .A(n10227), .ZN(n14954) );
  AOI211_X1 U12825 ( .C1(n10343), .C2(n10231), .A(n13574), .B(n10230), .ZN(
        n14946) );
  XNOR2_X1 U12826 ( .A(n10233), .B(n10232), .ZN(n10235) );
  INV_X1 U12827 ( .A(n9903), .ZN(n10234) );
  OAI22_X1 U12828 ( .A1(n10234), .A2(n13340), .B1(n10357), .B2(n13342), .ZN(
        n10313) );
  AOI21_X1 U12829 ( .B1(n10235), .B2(n14992), .A(n10313), .ZN(n14956) );
  INV_X1 U12830 ( .A(n14956), .ZN(n10236) );
  AOI211_X1 U12831 ( .C1(n15024), .C2(n14954), .A(n14946), .B(n10236), .ZN(
        n10345) );
  INV_X1 U12832 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10237) );
  OAI22_X1 U12833 ( .A1(n13718), .A2(n14952), .B1(n15027), .B2(n10237), .ZN(
        n10238) );
  INV_X1 U12834 ( .A(n10238), .ZN(n10239) );
  OAI21_X1 U12835 ( .B1(n10345), .B2(n15025), .A(n10239), .ZN(P2_U3436) );
  NAND2_X1 U12836 ( .A1(n9903), .A2(n13315), .ZN(n10406) );
  NOR2_X1 U12837 ( .A1(n13350), .A2(n14997), .ZN(n13334) );
  NAND2_X1 U12838 ( .A1(n13334), .A2(n8750), .ZN(n10243) );
  AOI21_X1 U12839 ( .B1(n8750), .B2(n13574), .A(n13350), .ZN(n10240) );
  NOR2_X1 U12840 ( .A1(n10240), .A2(n14578), .ZN(n10242) );
  MUX2_X1 U12841 ( .A(n10243), .B(n10242), .S(n10241), .Z(n10246) );
  OR2_X1 U12842 ( .A1(n10244), .A2(P2_U3088), .ZN(n10332) );
  NAND2_X1 U12843 ( .A1(n10332), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10245) );
  OAI211_X1 U12844 ( .C1(n13318), .C2(n10406), .A(n10246), .B(n10245), .ZN(
        P2_U3204) );
  INV_X1 U12845 ( .A(n10247), .ZN(n10335) );
  AOI22_X1 U12846 ( .A1(n10482), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14395), .ZN(n10248) );
  OAI21_X1 U12847 ( .B1(n10335), .B2(n14403), .A(n10248), .ZN(P1_U3343) );
  INV_X1 U12848 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12849 ( .A1(n11728), .A2(P3_U3897), .ZN(n10249) );
  OAI21_X1 U12850 ( .B1(P3_U3897), .B2(n10250), .A(n10249), .ZN(P3_U3499) );
  INV_X1 U12851 ( .A(n10454), .ZN(n10252) );
  NAND3_X1 U12852 ( .A1(n10455), .A2(n10252), .A3(n10251), .ZN(n10271) );
  OR2_X1 U12853 ( .A1(n10271), .A2(n10253), .ZN(n10269) );
  INV_X1 U12854 ( .A(n10254), .ZN(n10255) );
  NAND2_X1 U12855 ( .A1(n14615), .A2(n14236), .ZN(n13883) );
  INV_X1 U12856 ( .A(n13883), .ZN(n13767) );
  OR2_X1 U12857 ( .A1(n10269), .A2(n10459), .ZN(n10258) );
  INV_X1 U12858 ( .A(n10270), .ZN(n10257) );
  AOI22_X1 U12859 ( .A1(n13767), .A2(n13917), .B1(n10263), .B2(n14618), .ZN(
        n10276) );
  AND2_X4 U12860 ( .A1(n10262), .A2(n10259), .ZN(n12417) );
  INV_X2 U12861 ( .A(n10260), .ZN(n14317) );
  INV_X1 U12862 ( .A(n10262), .ZN(n10264) );
  NAND2_X1 U12863 ( .A1(n12423), .A2(n13918), .ZN(n10266) );
  NAND2_X1 U12864 ( .A1(n10264), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10265) );
  OAI211_X1 U12865 ( .C1(n12458), .C2(n10771), .A(n10266), .B(n10265), .ZN(
        n10370) );
  OR2_X1 U12866 ( .A1(n14744), .A2(n10267), .ZN(n10268) );
  NAND2_X1 U12867 ( .A1(n10271), .A2(n10270), .ZN(n10274) );
  INV_X1 U12868 ( .A(n10272), .ZN(n10273) );
  NAND2_X1 U12869 ( .A1(n10274), .A2(n10273), .ZN(n10918) );
  OR2_X1 U12870 ( .A1(n10918), .A2(P1_U3086), .ZN(n13769) );
  AOI22_X1 U12871 ( .A1(n13932), .A2(n14613), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n13769), .ZN(n10275) );
  NAND2_X1 U12872 ( .A1(n10276), .A2(n10275), .ZN(P1_U3232) );
  MUX2_X1 U12873 ( .A(n11760), .B(P2_REG1_REG_12__SCAN_IN), .S(n10296), .Z(
        n10285) );
  NAND2_X1 U12874 ( .A1(n10286), .A2(n10277), .ZN(n10278) );
  NAND2_X1 U12875 ( .A1(n10279), .A2(n10278), .ZN(n14815) );
  INV_X1 U12876 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10280) );
  MUX2_X1 U12877 ( .A(n10280), .B(P2_REG1_REG_10__SCAN_IN), .S(n10289), .Z(
        n14814) );
  OR2_X1 U12878 ( .A1(n14815), .A2(n14814), .ZN(n14817) );
  NAND2_X1 U12879 ( .A1(n10289), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10281) );
  NAND2_X1 U12880 ( .A1(n14817), .A2(n10281), .ZN(n14831) );
  INV_X1 U12881 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15387) );
  MUX2_X1 U12882 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15387), .S(n10291), .Z(
        n14830) );
  NAND2_X1 U12883 ( .A1(n14831), .A2(n14830), .ZN(n14829) );
  NAND2_X1 U12884 ( .A1(n10291), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12885 ( .A1(n14829), .A2(n10282), .ZN(n10284) );
  INV_X1 U12886 ( .A(n11763), .ZN(n10283) );
  AOI21_X1 U12887 ( .B1(n10285), .B2(n10284), .A(n10283), .ZN(n10301) );
  MUX2_X1 U12888 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11742), .S(n10296), .Z(
        n10295) );
  NAND2_X1 U12889 ( .A1(n10286), .A2(n10854), .ZN(n10287) );
  NAND2_X1 U12890 ( .A1(n10288), .A2(n10287), .ZN(n14819) );
  INV_X1 U12891 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11010) );
  MUX2_X1 U12892 ( .A(n11010), .B(P2_REG2_REG_10__SCAN_IN), .S(n10289), .Z(
        n14818) );
  NAND2_X1 U12893 ( .A1(n10289), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U12894 ( .A1(n14821), .A2(n10290), .ZN(n14835) );
  INV_X1 U12895 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10292) );
  MUX2_X1 U12896 ( .A(n10292), .B(P2_REG2_REG_11__SCAN_IN), .S(n10291), .Z(
        n14834) );
  NAND2_X1 U12897 ( .A1(n14833), .A2(n10292), .ZN(n10293) );
  NAND2_X1 U12898 ( .A1(n14837), .A2(n10293), .ZN(n10294) );
  NAND2_X1 U12899 ( .A1(n10294), .A2(n10295), .ZN(n11744) );
  OAI21_X1 U12900 ( .B1(n10295), .B2(n10294), .A(n11744), .ZN(n10299) );
  INV_X1 U12901 ( .A(n10296), .ZN(n11761) );
  NAND2_X1 U12902 ( .A1(n14760), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10297) );
  NAND2_X1 U12903 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11427)
         );
  OAI211_X1 U12904 ( .C1(n14926), .C2(n11761), .A(n10297), .B(n11427), .ZN(
        n10298) );
  AOI21_X1 U12905 ( .B1(n10299), .B2(n14915), .A(n10298), .ZN(n10300) );
  OAI21_X1 U12906 ( .B1(n10301), .B2(n14883), .A(n10300), .ZN(P2_U3226) );
  OAI21_X1 U12907 ( .B1(n10303), .B2(n10306), .A(n10302), .ZN(n10439) );
  NAND2_X1 U12908 ( .A1(n10304), .A2(n14997), .ZN(n10305) );
  NOR2_X1 U12909 ( .A1(n10384), .A2(n10305), .ZN(n10445) );
  XNOR2_X1 U12910 ( .A(n10307), .B(n10306), .ZN(n10309) );
  OAI21_X1 U12911 ( .B1(n10309), .B2(n13530), .A(n10308), .ZN(n10442) );
  AOI211_X1 U12912 ( .C1(n15024), .C2(n10439), .A(n10445), .B(n10442), .ZN(
        n10342) );
  INV_X1 U12913 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10310) );
  OAI22_X1 U12914 ( .A1(n13718), .A2(n7193), .B1(n15027), .B2(n10310), .ZN(
        n10311) );
  INV_X1 U12915 ( .A(n10311), .ZN(n10312) );
  OAI21_X1 U12916 ( .B1(n10342), .B2(n15025), .A(n10312), .ZN(P2_U3439) );
  INV_X1 U12917 ( .A(n10313), .ZN(n10314) );
  OAI22_X1 U12918 ( .A1(n14952), .A2(n13319), .B1(n13318), .B2(n10314), .ZN(
        n10320) );
  AOI22_X1 U12919 ( .A1(n13334), .A2(n9903), .B1(n14574), .B2(n10315), .ZN(
        n10318) );
  INV_X1 U12920 ( .A(n10316), .ZN(n10324) );
  NOR3_X1 U12921 ( .A1(n10318), .A2(n10324), .A3(n10317), .ZN(n10319) );
  AOI211_X1 U12922 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n10332), .A(n10320), .B(
        n10319), .ZN(n10321) );
  OAI21_X1 U12923 ( .B1(n13350), .B2(n10322), .A(n10321), .ZN(P2_U3209) );
  INV_X1 U12924 ( .A(n10323), .ZN(n10326) );
  INV_X1 U12925 ( .A(n10328), .ZN(n10325) );
  AOI21_X1 U12926 ( .B1(n10326), .B2(n10325), .A(n10324), .ZN(n10334) );
  OAI22_X1 U12927 ( .A1(n10584), .A2(n13319), .B1(n13318), .B2(n10327), .ZN(
        n10331) );
  INV_X1 U12928 ( .A(n13334), .ZN(n13299) );
  NOR3_X1 U12929 ( .A1(n13299), .A2(n10329), .A3(n10328), .ZN(n10330) );
  AOI211_X1 U12930 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n10332), .A(n10331), .B(
        n10330), .ZN(n10333) );
  OAI21_X1 U12931 ( .B1(n10334), .B2(n13350), .A(n10333), .ZN(P2_U3194) );
  OAI222_X1 U12932 ( .A1(P2_U3088), .A2(n11761), .B1(n11696), .B2(n10336), 
        .C1(n13741), .C2(n10335), .ZN(P2_U3315) );
  AOI22_X1 U12933 ( .A1(n8743), .A2(n10337), .B1(n15035), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10338) );
  OAI21_X1 U12934 ( .B1(n10339), .B2(n15035), .A(n10338), .ZN(P2_U3500) );
  AOI22_X1 U12935 ( .A1(n8743), .A2(n10340), .B1(n15035), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10341) );
  OAI21_X1 U12936 ( .B1(n10342), .B2(n15035), .A(n10341), .ZN(P2_U3502) );
  AOI22_X1 U12937 ( .A1(n8743), .A2(n10343), .B1(n15035), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10344) );
  OAI21_X1 U12938 ( .B1(n10345), .B2(n15035), .A(n10344), .ZN(P2_U3501) );
  INV_X1 U12939 ( .A(n10346), .ZN(n10347) );
  INV_X1 U12940 ( .A(n12718), .ZN(n12723) );
  OAI222_X1 U12941 ( .A1(n11389), .A2(n10347), .B1(n12723), .B2(P3_U3151), 
        .C1(n15328), .C2(n14525), .ZN(P3_U3279) );
  NAND2_X1 U12942 ( .A1(n13378), .A2(n13574), .ZN(n10422) );
  XNOR2_X1 U12943 ( .A(n10432), .B(n10422), .ZN(n10358) );
  AND2_X1 U12944 ( .A1(n10358), .A2(n10348), .ZN(n10349) );
  OAI21_X1 U12945 ( .B1(n10358), .B2(n10350), .A(n10431), .ZN(n10361) );
  NAND2_X1 U12946 ( .A1(n13380), .A2(n13316), .ZN(n10352) );
  NAND2_X1 U12947 ( .A1(n13377), .A2(n13315), .ZN(n10351) );
  AND2_X1 U12948 ( .A1(n10352), .A2(n10351), .ZN(n10388) );
  INV_X1 U12949 ( .A(n10388), .ZN(n10353) );
  AOI22_X1 U12950 ( .A1(n14576), .A2(n10353), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10355) );
  NAND2_X1 U12951 ( .A1(n14578), .A2(n10386), .ZN(n10354) );
  OAI211_X1 U12952 ( .C1(n14581), .C2(n10570), .A(n10355), .B(n10354), .ZN(
        n10360) );
  NOR4_X1 U12953 ( .A1(n13299), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10359) );
  AOI211_X1 U12954 ( .C1(n14574), .C2(n10361), .A(n10360), .B(n10359), .ZN(
        n10362) );
  INV_X1 U12955 ( .A(n10362), .ZN(P2_U3202) );
  NAND2_X1 U12956 ( .A1(n13917), .A2(n12423), .ZN(n10364) );
  NAND2_X1 U12957 ( .A1(n12417), .A2(n13770), .ZN(n10363) );
  NAND2_X1 U12958 ( .A1(n10364), .A2(n10363), .ZN(n10365) );
  XNOR2_X1 U12959 ( .A(n10365), .B(n10369), .ZN(n10366) );
  INV_X1 U12960 ( .A(n13917), .ZN(n10496) );
  NOR2_X1 U12961 ( .A1(n10366), .A2(n10367), .ZN(n10373) );
  NOR2_X1 U12962 ( .A1(n10373), .A2(n10368), .ZN(n13763) );
  XNOR2_X1 U12963 ( .A(n10374), .B(n12459), .ZN(n10891) );
  OAI22_X1 U12964 ( .A1(n12455), .A2(n10610), .B1(n14716), .B2(n12456), .ZN(
        n10890) );
  XNOR2_X1 U12965 ( .A(n10891), .B(n10890), .ZN(n10376) );
  AOI21_X1 U12966 ( .B1(n10377), .B2(n10376), .A(n12436), .ZN(n10381) );
  INV_X1 U12967 ( .A(n14618), .ZN(n13868) );
  NOR2_X1 U12968 ( .A1(n13868), .A2(n14716), .ZN(n10379) );
  NAND2_X1 U12969 ( .A1(n14615), .A2(n14234), .ZN(n13884) );
  OAI22_X1 U12970 ( .A1(n10496), .A2(n13884), .B1(n13883), .B2(n10896), .ZN(
        n10378) );
  AOI211_X1 U12971 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n13769), .A(n10379), .B(
        n10378), .ZN(n10380) );
  OAI21_X1 U12972 ( .B1(n10381), .B2(n13889), .A(n10380), .ZN(P1_U3237) );
  OAI21_X1 U12973 ( .B1(n10383), .B2(n7135), .A(n10382), .ZN(n10576) );
  INV_X1 U12974 ( .A(n10384), .ZN(n10385) );
  AOI211_X1 U12975 ( .C1(n10386), .C2(n10385), .A(n13202), .B(n10599), .ZN(
        n10569) );
  XNOR2_X1 U12976 ( .A(n10387), .B(n7135), .ZN(n10389) );
  OAI21_X1 U12977 ( .B1(n10389), .B2(n13530), .A(n10388), .ZN(n10568) );
  AOI211_X1 U12978 ( .C1(n15024), .C2(n10576), .A(n10569), .B(n10568), .ZN(
        n10396) );
  INV_X1 U12979 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10390) );
  OAI22_X1 U12980 ( .A1(n13718), .A2(n10574), .B1(n15027), .B2(n10390), .ZN(
        n10391) );
  INV_X1 U12981 ( .A(n10391), .ZN(n10392) );
  OAI21_X1 U12982 ( .B1(n10396), .B2(n15025), .A(n10392), .ZN(P2_U3442) );
  INV_X1 U12983 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10393) );
  OAI22_X1 U12984 ( .A1(n13672), .A2(n10574), .B1(n15037), .B2(n10393), .ZN(
        n10394) );
  INV_X1 U12985 ( .A(n10394), .ZN(n10395) );
  OAI21_X1 U12986 ( .B1(n10396), .B2(n15035), .A(n10395), .ZN(P2_U3503) );
  INV_X1 U12987 ( .A(n10397), .ZN(n10399) );
  INV_X1 U12988 ( .A(n10483), .ZN(n10531) );
  OAI222_X1 U12989 ( .A1(n14410), .A2(n10398), .B1(n14403), .B2(n10399), .C1(
        n10531), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12990 ( .A(n11765), .ZN(n14853) );
  INV_X1 U12991 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n15308) );
  OAI222_X1 U12992 ( .A1(P2_U3088), .A2(n14853), .B1(n11696), .B2(n15308), 
        .C1(n13741), .C2(n10399), .ZN(P2_U3314) );
  OAI21_X1 U12993 ( .B1(n14626), .B2(n14741), .A(n10774), .ZN(n10400) );
  NAND2_X1 U12994 ( .A1(n13917), .A2(n14236), .ZN(n10770) );
  OAI211_X1 U12995 ( .C1(n10401), .C2(n10771), .A(n10400), .B(n10770), .ZN(
        n10419) );
  NAND2_X1 U12996 ( .A1(n14759), .A2(n10419), .ZN(n10402) );
  OAI21_X1 U12997 ( .B1(n14759), .B2(n14652), .A(n10402), .ZN(P1_U3528) );
  AND2_X1 U12998 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  NAND3_X1 U12999 ( .A1(n14963), .A2(n10405), .A3(n14962), .ZN(n10413) );
  INV_X2 U13000 ( .A(n13512), .ZN(n14957) );
  INV_X1 U13001 ( .A(n10406), .ZN(n10408) );
  AOI21_X1 U13002 ( .B1(n13530), .B2(n14974), .A(n14971), .ZN(n10407) );
  NOR2_X1 U13003 ( .A1(n10408), .A2(n10407), .ZN(n14967) );
  INV_X1 U13004 ( .A(n10409), .ZN(n10440) );
  NOR2_X1 U13005 ( .A1(n14957), .A2(n10440), .ZN(n13588) );
  INV_X1 U13006 ( .A(n14971), .ZN(n10417) );
  OAI22_X1 U13007 ( .A1(n13512), .A2(n10412), .B1(n10411), .B2(n15200), .ZN(
        n10416) );
  NOR2_X2 U13008 ( .A1(n10413), .A2(n11409), .ZN(n15195) );
  AND2_X1 U13009 ( .A1(n15195), .A2(n14997), .ZN(n13418) );
  INV_X1 U13010 ( .A(n13418), .ZN(n10552) );
  AOI21_X1 U13011 ( .B1(n10552), .B2(n14951), .A(n14969), .ZN(n10415) );
  AOI211_X1 U13012 ( .C1(n13588), .C2(n10417), .A(n10416), .B(n10415), .ZN(
        n10418) );
  OAI21_X1 U13013 ( .B1(n14957), .B2(n14967), .A(n10418), .ZN(P2_U3265) );
  INV_X1 U13014 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U13015 ( .A1(n14752), .A2(n10419), .ZN(n10420) );
  OAI21_X1 U13016 ( .B1(n14752), .B2(n10421), .A(n10420), .ZN(P1_U3459) );
  INV_X1 U13017 ( .A(n10432), .ZN(n10423) );
  NAND2_X1 U13018 ( .A1(n10423), .A2(n10422), .ZN(n10424) );
  XNOR2_X1 U13019 ( .A(n10425), .B(n13217), .ZN(n10651) );
  NAND2_X1 U13020 ( .A1(n13377), .A2(n13574), .ZN(n10652) );
  XNOR2_X1 U13021 ( .A(n10651), .B(n10652), .ZN(n10433) );
  NAND2_X1 U13022 ( .A1(n10426), .A2(n10433), .ZN(n10655) );
  INV_X1 U13023 ( .A(n10427), .ZN(n10600) );
  OAI22_X1 U13024 ( .A1(n10429), .A2(n13340), .B1(n10428), .B2(n13342), .ZN(
        n10594) );
  AOI22_X1 U13025 ( .A1(n14576), .A2(n10594), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10430) );
  OAI21_X1 U13026 ( .B1(n13319), .B2(n14978), .A(n10430), .ZN(n10437) );
  INV_X1 U13027 ( .A(n10431), .ZN(n10435) );
  AOI22_X1 U13028 ( .A1(n13334), .A2(n13378), .B1(n14574), .B2(n10432), .ZN(
        n10434) );
  NOR3_X1 U13029 ( .A1(n10435), .A2(n10434), .A3(n10433), .ZN(n10436) );
  AOI211_X1 U13030 ( .C1(n13322), .C2(n10600), .A(n10437), .B(n10436), .ZN(
        n10438) );
  OAI21_X1 U13031 ( .B1(n13350), .B2(n10655), .A(n10438), .ZN(P2_U3199) );
  INV_X1 U13032 ( .A(n10439), .ZN(n10448) );
  NAND2_X1 U13033 ( .A1(n14974), .A2(n10440), .ZN(n10441) );
  INV_X1 U13034 ( .A(n10442), .ZN(n10443) );
  MUX2_X1 U13035 ( .A(n10105), .B(n10443), .S(n13512), .Z(n10447) );
  OAI22_X1 U13036 ( .A1(n14951), .A2(n7193), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n15200), .ZN(n10444) );
  AOI21_X1 U13037 ( .B1(n15195), .B2(n10445), .A(n10444), .ZN(n10446) );
  OAI211_X1 U13038 ( .C1(n10448), .C2(n13604), .A(n10447), .B(n10446), .ZN(
        P2_U3262) );
  INV_X1 U13039 ( .A(n12730), .ZN(n12739) );
  INV_X1 U13040 ( .A(n10449), .ZN(n10450) );
  OAI222_X1 U13041 ( .A1(n14525), .A2(n10451), .B1(n12739), .B2(P3_U3151), 
        .C1(n11389), .C2(n10450), .ZN(P3_U3278) );
  XNOR2_X1 U13042 ( .A(n10453), .B(n10452), .ZN(n14720) );
  INV_X1 U13043 ( .A(n14720), .ZN(n10474) );
  INV_X1 U13044 ( .A(n10457), .ZN(n10458) );
  NAND2_X1 U13045 ( .A1(n14225), .A2(n10458), .ZN(n14697) );
  NOR2_X2 U13046 ( .A1(n14712), .A2(n10459), .ZN(n14703) );
  NOR2_X2 U13047 ( .A1(n14063), .A2(n10460), .ZN(n14251) );
  OAI211_X1 U13048 ( .C1(n10495), .C2(n14716), .A(n14254), .B(n10612), .ZN(
        n14715) );
  INV_X1 U13049 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10461) );
  OAI22_X1 U13050 ( .A1(n14706), .A2(n14715), .B1(n10461), .B2(n14698), .ZN(
        n10462) );
  AOI21_X1 U13051 ( .B1(n14703), .B2(n10463), .A(n10462), .ZN(n10473) );
  INV_X1 U13052 ( .A(n10501), .ZN(n14730) );
  OAI21_X1 U13053 ( .B1(n10466), .B2(n10465), .A(n10464), .ZN(n10467) );
  NAND2_X1 U13054 ( .A1(n10467), .A2(n14741), .ZN(n10469) );
  AOI22_X1 U13055 ( .A1(n14234), .A2(n13917), .B1(n13914), .B2(n14236), .ZN(
        n10468) );
  NAND2_X1 U13056 ( .A1(n10469), .A2(n10468), .ZN(n10470) );
  AOI21_X1 U13057 ( .B1(n14720), .B2(n14730), .A(n10470), .ZN(n14717) );
  INV_X1 U13058 ( .A(n14712), .ZN(n14225) );
  MUX2_X1 U13059 ( .A(n10471), .B(n14717), .S(n14225), .Z(n10472) );
  OAI211_X1 U13060 ( .C1(n10474), .C2(n14697), .A(n10473), .B(n10472), .ZN(
        P1_U3291) );
  INV_X1 U13061 ( .A(n10486), .ZN(n11315) );
  AOI22_X1 U13062 ( .A1(n10486), .A2(n7887), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11315), .ZN(n10478) );
  INV_X1 U13063 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15339) );
  AOI21_X1 U13064 ( .B1(n10200), .B2(n10476), .A(n10475), .ZN(n10529) );
  MUX2_X1 U13065 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15339), .S(n10483), .Z(
        n10528) );
  NAND2_X1 U13066 ( .A1(n10529), .A2(n10528), .ZN(n10527) );
  OAI21_X1 U13067 ( .B1(n10531), .B2(n15339), .A(n10527), .ZN(n10477) );
  NOR2_X1 U13068 ( .A1(n10478), .A2(n10477), .ZN(n11314) );
  AOI21_X1 U13069 ( .B1(n10478), .B2(n10477), .A(n11314), .ZN(n10492) );
  NAND2_X1 U13070 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14619)
         );
  NAND2_X1 U13071 ( .A1(n14655), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10479) );
  OAI211_X1 U13072 ( .C1(n14691), .C2(n11315), .A(n14619), .B(n10479), .ZN(
        n10480) );
  INV_X1 U13073 ( .A(n10480), .ZN(n10491) );
  NAND2_X1 U13074 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10483), .ZN(n10485) );
  OAI21_X1 U13075 ( .B1(n10482), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10481), 
        .ZN(n10526) );
  MUX2_X1 U13076 ( .A(n11633), .B(P1_REG2_REG_13__SCAN_IN), .S(n10483), .Z(
        n10525) );
  OR2_X1 U13077 ( .A1(n10526), .A2(n10525), .ZN(n10484) );
  NAND2_X1 U13078 ( .A1(n10485), .A2(n10484), .ZN(n10489) );
  MUX2_X1 U13079 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10487), .S(n10486), .Z(
        n10488) );
  NAND2_X1 U13080 ( .A1(n10488), .A2(n10489), .ZN(n11308) );
  OAI211_X1 U13081 ( .C1(n10489), .C2(n10488), .A(n11308), .B(n14038), .ZN(
        n10490) );
  OAI211_X1 U13082 ( .C1(n10492), .C2(n14689), .A(n10491), .B(n10490), .ZN(
        P1_U3257) );
  XNOR2_X1 U13083 ( .A(n10497), .B(n10493), .ZN(n10627) );
  INV_X1 U13084 ( .A(n14698), .ZN(n14241) );
  NOR2_X1 U13085 ( .A1(n10610), .A2(n14142), .ZN(n10623) );
  NOR2_X1 U13086 ( .A1(n10771), .A2(n10631), .ZN(n10494) );
  OR2_X1 U13087 ( .A1(n10495), .A2(n10494), .ZN(n10505) );
  XNOR2_X1 U13088 ( .A(n10505), .B(n10496), .ZN(n10500) );
  INV_X1 U13089 ( .A(n10497), .ZN(n10498) );
  NOR2_X1 U13090 ( .A1(n10498), .A2(n14234), .ZN(n10499) );
  MUX2_X1 U13091 ( .A(n10500), .B(n10499), .S(n6758), .Z(n10503) );
  AOI21_X1 U13092 ( .B1(n6758), .B2(n14234), .A(n14741), .ZN(n10502) );
  OAI22_X1 U13093 ( .A1(n10503), .A2(n10502), .B1(n10627), .B2(n10501), .ZN(
        n10622) );
  AOI211_X1 U13094 ( .C1(n14241), .C2(P1_REG3_REG_1__SCAN_IN), .A(n10623), .B(
        n10622), .ZN(n10504) );
  MUX2_X1 U13095 ( .A(n10035), .B(n10504), .S(n14225), .Z(n10507) );
  AND2_X1 U13096 ( .A1(n14251), .A2(n14254), .ZN(n14048) );
  INV_X1 U13097 ( .A(n10505), .ZN(n10624) );
  AOI22_X1 U13098 ( .A1(n14703), .A2(n13770), .B1(n14048), .B2(n10624), .ZN(
        n10506) );
  OAI211_X1 U13099 ( .C1(n10627), .C2(n14697), .A(n10507), .B(n10506), .ZN(
        P1_U3292) );
  INV_X1 U13100 ( .A(n10508), .ZN(n10510) );
  INV_X1 U13101 ( .A(n12758), .ZN(n10509) );
  OAI222_X1 U13102 ( .A1(n14525), .A2(n10511), .B1(n11389), .B2(n10510), .C1(
        P3_U3151), .C2(n10509), .ZN(P3_U3277) );
  XNOR2_X1 U13103 ( .A(n10512), .B(n10521), .ZN(n14737) );
  NAND2_X1 U13104 ( .A1(n13912), .A2(n14236), .ZN(n10515) );
  NAND2_X1 U13105 ( .A1(n13914), .A2(n14234), .ZN(n10514) );
  AND2_X1 U13106 ( .A1(n10515), .A2(n10514), .ZN(n14733) );
  INV_X1 U13107 ( .A(n14733), .ZN(n10516) );
  MUX2_X1 U13108 ( .A(n10516), .B(P1_REG2_REG_4__SCAN_IN), .S(n14712), .Z(
        n10520) );
  NAND2_X1 U13109 ( .A1(n14225), .A2(n14040), .ZN(n14070) );
  NAND2_X1 U13110 ( .A1(n10613), .A2(n10929), .ZN(n10517) );
  NAND2_X1 U13111 ( .A1(n10517), .A2(n14254), .ZN(n10518) );
  OR2_X1 U13112 ( .A1(n10518), .A2(n10558), .ZN(n14734) );
  OAI22_X1 U13113 ( .A1(n14070), .A2(n14734), .B1(n10928), .B2(n14698), .ZN(
        n10519) );
  AOI211_X1 U13114 ( .C1(n14703), .C2(n10929), .A(n10520), .B(n10519), .ZN(
        n10524) );
  XNOR2_X1 U13115 ( .A(n10522), .B(n10521), .ZN(n14740) );
  NAND2_X1 U13116 ( .A1(n14740), .A2(n14121), .ZN(n10523) );
  OAI211_X1 U13117 ( .C1(n14737), .C2(n14248), .A(n10524), .B(n10523), .ZN(
        P1_U3289) );
  XNOR2_X1 U13118 ( .A(n10526), .B(n10525), .ZN(n10535) );
  NAND2_X1 U13119 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13838)
         );
  OAI211_X1 U13120 ( .C1(n10529), .C2(n10528), .A(n14037), .B(n10527), .ZN(
        n10530) );
  NAND2_X1 U13121 ( .A1(n13838), .A2(n10530), .ZN(n10533) );
  NOR2_X1 U13122 ( .A1(n14691), .A2(n10531), .ZN(n10532) );
  AOI211_X1 U13123 ( .C1(n14655), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n10533), 
        .B(n10532), .ZN(n10534) );
  OAI21_X1 U13124 ( .B1(n10535), .B2(n14687), .A(n10534), .ZN(P1_U3256) );
  OAI222_X1 U13125 ( .A1(n14525), .A2(n10537), .B1(n11389), .B2(n10536), .C1(
        P3_U3151), .C2(n12764), .ZN(P3_U3276) );
  XNOR2_X1 U13126 ( .A(n10539), .B(n10538), .ZN(n14986) );
  INV_X1 U13127 ( .A(n14974), .ZN(n10540) );
  NAND2_X1 U13128 ( .A1(n14986), .A2(n10540), .ZN(n10547) );
  XNOR2_X1 U13129 ( .A(n10542), .B(n10541), .ZN(n10545) );
  NAND2_X1 U13130 ( .A1(n13377), .A2(n13316), .ZN(n10544) );
  NAND2_X1 U13131 ( .A1(n13375), .A2(n13315), .ZN(n10543) );
  NAND2_X1 U13132 ( .A1(n10544), .A2(n10543), .ZN(n10644) );
  AOI21_X1 U13133 ( .B1(n10545), .B2(n14992), .A(n10644), .ZN(n10546) );
  AND2_X1 U13134 ( .A1(n10547), .A2(n10546), .ZN(n14988) );
  AND2_X1 U13135 ( .A1(n10598), .A2(n14983), .ZN(n10548) );
  OR2_X1 U13136 ( .A1(n7209), .A2(n10548), .ZN(n14984) );
  OAI22_X1 U13137 ( .A1(n13512), .A2(n10549), .B1(n10646), .B2(n15200), .ZN(
        n10550) );
  AOI21_X1 U13138 ( .B1(n14983), .B2(n14937), .A(n10550), .ZN(n10551) );
  OAI21_X1 U13139 ( .B1(n14984), .B2(n10552), .A(n10551), .ZN(n10553) );
  AOI21_X1 U13140 ( .B1(n14986), .B2(n13588), .A(n10553), .ZN(n10554) );
  OAI21_X1 U13141 ( .B1(n14988), .B2(n10410), .A(n10554), .ZN(P2_U3259) );
  AOI21_X1 U13142 ( .B1(n10561), .B2(n10555), .A(n6730), .ZN(n10637) );
  INV_X1 U13143 ( .A(n10923), .ZN(n10556) );
  OAI22_X1 U13144 ( .A1(n14225), .A2(n10557), .B1(n10556), .B2(n14698), .ZN(
        n10560) );
  OAI211_X1 U13145 ( .C1(n10558), .C2(n10921), .A(n14254), .B(n10692), .ZN(
        n10635) );
  NOR2_X1 U13146 ( .A1(n14706), .A2(n10635), .ZN(n10559) );
  AOI211_X1 U13147 ( .C1(n14703), .C2(n10914), .A(n10560), .B(n10559), .ZN(
        n10567) );
  XNOR2_X1 U13148 ( .A(n10562), .B(n10561), .ZN(n10565) );
  NAND2_X1 U13149 ( .A1(n13911), .A2(n14236), .ZN(n10564) );
  NAND2_X1 U13150 ( .A1(n13913), .A2(n14234), .ZN(n10563) );
  NAND2_X1 U13151 ( .A1(n10564), .A2(n10563), .ZN(n10919) );
  AOI21_X1 U13152 ( .B1(n10565), .B2(n14741), .A(n10919), .ZN(n10636) );
  OR2_X1 U13153 ( .A1(n10636), .A2(n14712), .ZN(n10566) );
  OAI211_X1 U13154 ( .C1(n10637), .C2(n14248), .A(n10567), .B(n10566), .ZN(
        P1_U3288) );
  INV_X1 U13155 ( .A(n10568), .ZN(n10578) );
  NAND2_X1 U13156 ( .A1(n10569), .A2(n15195), .ZN(n10573) );
  INV_X1 U13157 ( .A(n10570), .ZN(n10571) );
  INV_X1 U13158 ( .A(n15200), .ZN(n14948) );
  AOI22_X1 U13159 ( .A1(n14957), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n10571), 
        .B2(n14948), .ZN(n10572) );
  OAI211_X1 U13160 ( .C1(n10574), .C2(n14951), .A(n10573), .B(n10572), .ZN(
        n10575) );
  AOI21_X1 U13161 ( .B1(n15196), .B2(n10576), .A(n10575), .ZN(n10577) );
  OAI21_X1 U13162 ( .B1(n10578), .B2(n10410), .A(n10577), .ZN(P2_U3261) );
  INV_X1 U13163 ( .A(n10579), .ZN(n10588) );
  AOI22_X1 U13164 ( .A1(n14957), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n14948), .ZN(n10583) );
  NAND2_X1 U13165 ( .A1(n15195), .A2(n10581), .ZN(n10582) );
  OAI211_X1 U13166 ( .C1(n14951), .C2(n10584), .A(n10583), .B(n10582), .ZN(
        n10585) );
  AOI21_X1 U13167 ( .B1(n15196), .B2(n10586), .A(n10585), .ZN(n10587) );
  OAI21_X1 U13168 ( .B1(n10588), .B2(n10410), .A(n10587), .ZN(P2_U3264) );
  INV_X1 U13169 ( .A(n11767), .ZN(n14865) );
  INV_X1 U13170 ( .A(n10589), .ZN(n10591) );
  INV_X1 U13171 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10590) );
  OAI222_X1 U13172 ( .A1(n14865), .A2(P2_U3088), .B1(n13741), .B2(n10591), 
        .C1(n10590), .C2(n13739), .ZN(P2_U3313) );
  OAI222_X1 U13173 ( .A1(n14410), .A2(n10592), .B1(n14403), .B2(n10591), .C1(
        P1_U3086), .C2(n11315), .ZN(P1_U3341) );
  XNOR2_X1 U13174 ( .A(n10593), .B(n10596), .ZN(n10595) );
  AOI21_X1 U13175 ( .B1(n10595), .B2(n14992), .A(n10594), .ZN(n14977) );
  XOR2_X1 U13176 ( .A(n10597), .B(n10596), .Z(n14981) );
  NAND2_X1 U13177 ( .A1(n14981), .A2(n15196), .ZN(n10605) );
  OAI211_X1 U13178 ( .C1(n10599), .C2(n14978), .A(n14997), .B(n10598), .ZN(
        n14976) );
  INV_X1 U13179 ( .A(n14976), .ZN(n10603) );
  AOI22_X1 U13180 ( .A1(n14957), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n10600), 
        .B2(n14948), .ZN(n10601) );
  OAI21_X1 U13181 ( .B1(n14978), .B2(n14951), .A(n10601), .ZN(n10602) );
  AOI21_X1 U13182 ( .B1(n10603), .B2(n15195), .A(n10602), .ZN(n10604) );
  OAI211_X1 U13183 ( .C1(n14957), .C2(n14977), .A(n10605), .B(n10604), .ZN(
        P2_U3260) );
  XNOR2_X1 U13184 ( .A(n10606), .B(n10608), .ZN(n14724) );
  OAI21_X1 U13185 ( .B1(n10609), .B2(n10608), .A(n10607), .ZN(n10611) );
  OAI22_X1 U13186 ( .A1(n10610), .A2(n14140), .B1(n10905), .B2(n14142), .ZN(
        n12438) );
  AOI21_X1 U13187 ( .B1(n10611), .B2(n14741), .A(n12438), .ZN(n14726) );
  INV_X1 U13188 ( .A(n14726), .ZN(n10620) );
  NAND2_X1 U13189 ( .A1(n14703), .A2(n10892), .ZN(n10617) );
  AOI21_X1 U13190 ( .B1(n10612), .B2(n10892), .A(n14317), .ZN(n10614) );
  NAND2_X1 U13191 ( .A1(n10614), .A2(n10613), .ZN(n14725) );
  INV_X1 U13192 ( .A(n14725), .ZN(n10615) );
  INV_X1 U13193 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U13194 ( .A1(n14251), .A2(n10615), .B1(n14241), .B2(n13948), .ZN(
        n10616) );
  OAI211_X1 U13195 ( .C1(n10618), .C2(n14225), .A(n10617), .B(n10616), .ZN(
        n10619) );
  AOI21_X1 U13196 ( .B1(n10620), .B2(n14225), .A(n10619), .ZN(n10621) );
  OAI21_X1 U13197 ( .B1(n14248), .B2(n14724), .A(n10621), .ZN(P1_U3290) );
  INV_X1 U13198 ( .A(n10622), .ZN(n10626) );
  AOI21_X1 U13199 ( .B1(n10624), .B2(n14254), .A(n10623), .ZN(n10625) );
  OAI211_X1 U13200 ( .C1(n10627), .C2(n14723), .A(n10626), .B(n10625), .ZN(
        n10633) );
  INV_X1 U13201 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10628) );
  OAI22_X1 U13202 ( .A1(n14381), .A2(n10631), .B1(n14752), .B2(n10628), .ZN(
        n10629) );
  AOI21_X1 U13203 ( .B1(n10633), .B2(n14752), .A(n10629), .ZN(n10630) );
  INV_X1 U13204 ( .A(n10630), .ZN(P1_U3462) );
  OAI22_X1 U13205 ( .A1(n14304), .A2(n10631), .B1(n14759), .B2(n13922), .ZN(
        n10632) );
  AOI21_X1 U13206 ( .B1(n10633), .B2(n14759), .A(n10632), .ZN(n10634) );
  INV_X1 U13207 ( .A(n10634), .ZN(P1_U3529) );
  OAI211_X1 U13208 ( .C1(n10637), .C2(n14749), .A(n10636), .B(n10635), .ZN(
        n10642) );
  INV_X1 U13209 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10638) );
  OAI22_X1 U13210 ( .A1(n14381), .A2(n10921), .B1(n14752), .B2(n10638), .ZN(
        n10639) );
  AOI21_X1 U13211 ( .B1(n10642), .B2(n14752), .A(n10639), .ZN(n10640) );
  INV_X1 U13212 ( .A(n10640), .ZN(P1_U3474) );
  OAI22_X1 U13213 ( .A1(n14304), .A2(n10921), .B1(n14759), .B2(n15385), .ZN(
        n10641) );
  AOI21_X1 U13214 ( .B1(n10642), .B2(n14759), .A(n10641), .ZN(n10643) );
  INV_X1 U13215 ( .A(n10643), .ZN(P1_U3533) );
  NAND2_X1 U13216 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14812) );
  NAND2_X1 U13217 ( .A1(n14576), .A2(n10644), .ZN(n10645) );
  OAI211_X1 U13218 ( .C1(n14581), .C2(n10646), .A(n14812), .B(n10645), .ZN(
        n10660) );
  XNOR2_X1 U13219 ( .A(n14983), .B(n13217), .ZN(n10831) );
  AND2_X1 U13220 ( .A1(n13376), .A2(n13574), .ZN(n10647) );
  NAND2_X1 U13221 ( .A1(n10831), .A2(n10647), .ZN(n10707) );
  INV_X1 U13222 ( .A(n10831), .ZN(n10649) );
  INV_X1 U13223 ( .A(n10647), .ZN(n10648) );
  NAND2_X1 U13224 ( .A1(n10649), .A2(n10648), .ZN(n10650) );
  NAND2_X1 U13225 ( .A1(n10707), .A2(n10650), .ZN(n10658) );
  INV_X1 U13226 ( .A(n10651), .ZN(n10653) );
  NAND2_X1 U13227 ( .A1(n10653), .A2(n10652), .ZN(n10654) );
  INV_X1 U13228 ( .A(n10708), .ZN(n10833) );
  AOI211_X1 U13229 ( .C1(n10658), .C2(n10657), .A(n13350), .B(n10833), .ZN(
        n10659) );
  AOI211_X1 U13230 ( .C1(n14983), .C2(n14578), .A(n10660), .B(n10659), .ZN(
        n10661) );
  INV_X1 U13231 ( .A(n10661), .ZN(P2_U3211) );
  INV_X1 U13232 ( .A(n10781), .ZN(n10663) );
  OAI21_X1 U13233 ( .B1(n12213), .B2(n10663), .A(n10662), .ZN(n10674) );
  OR2_X1 U13234 ( .A1(n10781), .A2(P3_U3151), .ZN(n12274) );
  NAND2_X1 U13235 ( .A1(n10664), .A2(n12274), .ZN(n10673) );
  INV_X1 U13236 ( .A(n10673), .ZN(n10665) );
  MUX2_X1 U13237 ( .A(n10680), .B(n12637), .S(n12269), .Z(n12765) );
  INV_X1 U13238 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10666) );
  MUX2_X1 U13239 ( .A(n10666), .B(P3_REG1_REG_2__SCAN_IN), .S(n10749), .Z(
        n10672) );
  NAND2_X1 U13240 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10667), .ZN(n10668) );
  INV_X1 U13241 ( .A(n10668), .ZN(n10956) );
  OR2_X1 U13242 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10668), .ZN(n10670) );
  OAI21_X1 U13243 ( .B1(n10979), .B2(n10956), .A(n10670), .ZN(n10964) );
  INV_X1 U13244 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U13245 ( .A1(n10672), .A2(n10671), .ZN(n10759) );
  OAI21_X1 U13246 ( .B1(n10672), .B2(n10671), .A(n10759), .ZN(n10678) );
  INV_X1 U13247 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10676) );
  INV_X1 U13248 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10675) );
  OAI22_X1 U13249 ( .A1(n15088), .A2(n10676), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10675), .ZN(n10677) );
  AOI21_X1 U13250 ( .B1(n15080), .B2(n10678), .A(n10677), .ZN(n10689) );
  MUX2_X1 U13251 ( .A(n9087), .B(P3_REG2_REG_2__SCAN_IN), .S(n10749), .Z(
        n10684) );
  NOR2_X1 U13252 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11131), .ZN(n10960) );
  NAND2_X1 U13253 ( .A1(n10681), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10682) );
  OAI21_X1 U13254 ( .B1(n10979), .B2(n10960), .A(n10682), .ZN(n10972) );
  OR2_X1 U13255 ( .A1(n10972), .A2(n9081), .ZN(n10974) );
  NAND2_X1 U13256 ( .A1(n10974), .A2(n10682), .ZN(n10683) );
  NAND2_X1 U13257 ( .A1(n10684), .A2(n10683), .ZN(n10753) );
  OAI21_X1 U13258 ( .B1(n10684), .B2(n10683), .A(n10753), .ZN(n10687) );
  NAND2_X1 U13259 ( .A1(P3_U3897), .A2(n12431), .ZN(n15071) );
  MUX2_X1 U13260 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12725), .Z(n10685) );
  XNOR2_X1 U13261 ( .A(n10685), .B(n10979), .ZN(n10968) );
  INV_X1 U13262 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11067) );
  MUX2_X1 U13263 ( .A(n11131), .B(n11067), .S(n12733), .Z(n10954) );
  NAND2_X1 U13264 ( .A1(n10954), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10967) );
  OAI22_X1 U13265 ( .A1(n10968), .A2(n10967), .B1(n10685), .B2(n10979), .ZN(
        n10751) );
  MUX2_X1 U13266 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12725), .Z(n10747) );
  XNOR2_X1 U13267 ( .A(n10747), .B(n10749), .ZN(n10750) );
  XNOR2_X1 U13268 ( .A(n10751), .B(n10750), .ZN(n10686) );
  AOI22_X1 U13269 ( .A1(n12774), .A2(n10687), .B1(n15099), .B2(n10686), .ZN(
        n10688) );
  OAI211_X1 U13270 ( .C1(n10757), .C2(n12765), .A(n10689), .B(n10688), .ZN(
        P3_U3184) );
  OAI21_X1 U13271 ( .B1(n10691), .B2(n10695), .A(n10690), .ZN(n10869) );
  NAND2_X1 U13272 ( .A1(n10692), .A2(n11036), .ZN(n10693) );
  NAND2_X1 U13273 ( .A1(n10693), .A2(n14254), .ZN(n10694) );
  NOR2_X1 U13274 ( .A1(n6733), .A2(n10694), .ZN(n10863) );
  XNOR2_X1 U13275 ( .A(n10696), .B(n10695), .ZN(n10699) );
  NAND2_X1 U13276 ( .A1(n13912), .A2(n14234), .ZN(n10698) );
  NAND2_X1 U13277 ( .A1(n13910), .A2(n14236), .ZN(n10697) );
  AND2_X1 U13278 ( .A1(n10698), .A2(n10697), .ZN(n11041) );
  OAI21_X1 U13279 ( .B1(n10699), .B2(n14329), .A(n11041), .ZN(n10866) );
  AOI211_X1 U13280 ( .C1(n14626), .C2(n10869), .A(n10863), .B(n10866), .ZN(
        n10706) );
  INV_X1 U13281 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10700) );
  OAI22_X1 U13282 ( .A1(n14381), .A2(n7070), .B1(n14752), .B2(n10700), .ZN(
        n10701) );
  INV_X1 U13283 ( .A(n10701), .ZN(n10702) );
  OAI21_X1 U13284 ( .B1(n10706), .B2(n14751), .A(n10702), .ZN(P1_U3477) );
  OAI22_X1 U13285 ( .A1(n14304), .A2(n7070), .B1(n14759), .B2(n10703), .ZN(
        n10704) );
  INV_X1 U13286 ( .A(n10704), .ZN(n10705) );
  OAI21_X1 U13287 ( .B1(n10706), .B2(n14757), .A(n10705), .ZN(P1_U3534) );
  XNOR2_X1 U13288 ( .A(n15003), .B(n13217), .ZN(n10880) );
  NAND2_X1 U13289 ( .A1(n13374), .A2(n13574), .ZN(n10871) );
  XNOR2_X1 U13290 ( .A(n10880), .B(n10871), .ZN(n10723) );
  INV_X1 U13291 ( .A(n10723), .ZN(n10717) );
  XNOR2_X1 U13292 ( .A(n10839), .B(n13217), .ZN(n10709) );
  AND2_X1 U13293 ( .A1(n13375), .A2(n13202), .ZN(n10710) );
  NAND2_X1 U13294 ( .A1(n10709), .A2(n10710), .ZN(n10714) );
  INV_X1 U13295 ( .A(n10709), .ZN(n10721) );
  INV_X1 U13296 ( .A(n10710), .ZN(n10711) );
  NAND2_X1 U13297 ( .A1(n10721), .A2(n10711), .ZN(n10712) );
  AND2_X1 U13298 ( .A1(n10714), .A2(n10712), .ZN(n10832) );
  NAND2_X1 U13299 ( .A1(n10713), .A2(n10832), .ZN(n10716) );
  INV_X1 U13300 ( .A(n10716), .ZN(n10834) );
  AND2_X1 U13301 ( .A1(n10723), .A2(n10714), .ZN(n10715) );
  NAND2_X1 U13302 ( .A1(n10716), .A2(n10715), .ZN(n10874) );
  INV_X1 U13303 ( .A(n10874), .ZN(n10883) );
  AOI21_X1 U13304 ( .B1(n10717), .B2(n10834), .A(n10883), .ZN(n10727) );
  NAND2_X1 U13305 ( .A1(n13375), .A2(n13316), .ZN(n10719) );
  NAND2_X1 U13306 ( .A1(n13373), .A2(n13315), .ZN(n10718) );
  NAND2_X1 U13307 ( .A1(n10719), .A2(n10718), .ZN(n10736) );
  AOI22_X1 U13308 ( .A1(n14576), .A2(n10736), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10720) );
  OAI21_X1 U13309 ( .B1(n10742), .B2(n14581), .A(n10720), .ZN(n10725) );
  NOR4_X1 U13310 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n13299), .ZN(
        n10724) );
  AOI211_X1 U13311 ( .C1(n15003), .C2(n14578), .A(n10725), .B(n10724), .ZN(
        n10726) );
  OAI21_X1 U13312 ( .B1(n10727), .B2(n13350), .A(n10726), .ZN(P2_U3193) );
  NAND2_X1 U13313 ( .A1(n10729), .A2(n10728), .ZN(n10730) );
  NAND2_X1 U13314 ( .A1(n10731), .A2(n10730), .ZN(n10740) );
  OR2_X1 U13315 ( .A1(n10740), .A2(n14974), .ZN(n10739) );
  NAND2_X1 U13316 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  NAND2_X1 U13317 ( .A1(n10735), .A2(n10734), .ZN(n10737) );
  AOI21_X1 U13318 ( .B1(n10737), .B2(n14992), .A(n10736), .ZN(n10738) );
  AND2_X1 U13319 ( .A1(n10739), .A2(n10738), .ZN(n15009) );
  INV_X1 U13320 ( .A(n10740), .ZN(n15007) );
  NAND2_X1 U13321 ( .A1(n14996), .A2(n15003), .ZN(n10741) );
  NAND3_X1 U13322 ( .A1(n10852), .A2(n14997), .A3(n10741), .ZN(n15004) );
  INV_X1 U13323 ( .A(n15195), .ZN(n13563) );
  OAI22_X1 U13324 ( .A1(n13512), .A2(n10117), .B1(n10742), .B2(n15200), .ZN(
        n10743) );
  AOI21_X1 U13325 ( .B1(n15003), .B2(n14937), .A(n10743), .ZN(n10744) );
  OAI21_X1 U13326 ( .B1(n15004), .B2(n13563), .A(n10744), .ZN(n10745) );
  AOI21_X1 U13327 ( .B1(n15007), .B2(n13588), .A(n10745), .ZN(n10746) );
  OAI21_X1 U13328 ( .B1(n15009), .B2(n10410), .A(n10746), .ZN(P2_U3257) );
  INV_X1 U13329 ( .A(n10747), .ZN(n10748) );
  AOI22_X1 U13330 ( .A1(n10751), .A2(n10750), .B1(n10749), .B2(n10748), .ZN(
        n11084) );
  MUX2_X1 U13331 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12733), .Z(n11082) );
  XOR2_X1 U13332 ( .A(n7257), .B(n11082), .Z(n11083) );
  XNOR2_X1 U13333 ( .A(n11084), .B(n11083), .ZN(n10765) );
  NAND2_X1 U13334 ( .A1(n10757), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U13335 ( .A1(n10754), .A2(n9111), .ZN(n10755) );
  NAND2_X1 U13336 ( .A1(n11091), .A2(n10755), .ZN(n10756) );
  NAND2_X1 U13337 ( .A1(n12774), .A2(n10756), .ZN(n10763) );
  NAND2_X1 U13338 ( .A1(n10757), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10758) );
  XNOR2_X1 U13339 ( .A(n11100), .B(n7257), .ZN(n11098) );
  XNOR2_X1 U13340 ( .A(n11098), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n10760) );
  NAND2_X1 U13341 ( .A1(n15080), .A2(n10760), .ZN(n10762) );
  NOR2_X1 U13342 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9109), .ZN(n10800) );
  AOI21_X1 U13343 ( .B1(n15093), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10800), .ZN(
        n10761) );
  NAND3_X1 U13344 ( .A1(n10763), .A2(n10762), .A3(n10761), .ZN(n10764) );
  AOI21_X1 U13345 ( .B1(n15099), .B2(n10765), .A(n10764), .ZN(n10766) );
  OAI21_X1 U13346 ( .B1(n11099), .B2(n12765), .A(n10766), .ZN(P3_U3185) );
  NAND2_X1 U13347 ( .A1(n12637), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10767) );
  OAI21_X1 U13348 ( .B1(n12792), .B2(n12637), .A(n10767), .ZN(P3_U3520) );
  NAND2_X1 U13349 ( .A1(n12637), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10768) );
  OAI21_X1 U13350 ( .B1(n12067), .B2(n12637), .A(n10768), .ZN(P3_U3521) );
  OAI22_X1 U13351 ( .A1(n14712), .A2(n10770), .B1(n10769), .B2(n14698), .ZN(
        n10773) );
  INV_X1 U13352 ( .A(n14048), .ZN(n14214) );
  AOI21_X1 U13353 ( .B1(n14244), .B2(n14214), .A(n10771), .ZN(n10772) );
  AOI211_X1 U13354 ( .C1(n14712), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10773), .B(
        n10772), .ZN(n10776) );
  OAI21_X1 U13355 ( .B1(n14229), .B2(n14121), .A(n10774), .ZN(n10775) );
  NAND2_X1 U13356 ( .A1(n10776), .A2(n10775), .ZN(P1_U3293) );
  NOR2_X1 U13357 ( .A1(n10779), .A2(n12263), .ZN(n11069) );
  NAND3_X1 U13358 ( .A1(n10801), .A2(n10780), .A3(n10783), .ZN(n10816) );
  NAND2_X1 U13359 ( .A1(n11069), .A2(n10816), .ZN(n10789) );
  AND2_X1 U13360 ( .A1(n10782), .A2(n10781), .ZN(n10788) );
  NAND3_X1 U13361 ( .A1(n10785), .A2(n10784), .A3(n10783), .ZN(n10793) );
  NAND2_X1 U13362 ( .A1(n11074), .A2(n10793), .ZN(n10787) );
  NAND4_X1 U13363 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10790) );
  NAND2_X1 U13364 ( .A1(n10790), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10792) );
  NOR2_X1 U13365 ( .A1(n12213), .A2(n12229), .ZN(n11064) );
  NAND2_X1 U13366 ( .A1(n12270), .A2(n10816), .ZN(n10791) );
  INV_X1 U13367 ( .A(n10793), .ZN(n11070) );
  NAND3_X1 U13368 ( .A1(n15155), .A2(n11073), .A3(n11070), .ZN(n10794) );
  NOR2_X1 U13369 ( .A1(n10816), .A2(n10796), .ZN(n10795) );
  INV_X1 U13370 ( .A(n10796), .ZN(n10797) );
  NOR2_X1 U13371 ( .A1(n10816), .A2(n10797), .ZN(n10798) );
  AOI211_X1 U13372 ( .C1(n11302), .C2(n15040), .A(n10800), .B(n10799), .ZN(
        n10826) );
  NAND2_X1 U13373 ( .A1(n10803), .A2(n10802), .ZN(n10804) );
  XNOR2_X1 U13374 ( .A(n10809), .B(n10807), .ZN(n10808) );
  AOI21_X1 U13375 ( .B1(n7398), .B2(n15112), .A(n10811), .ZN(n10812) );
  XNOR2_X1 U13376 ( .A(n10809), .B(n11015), .ZN(n10813) );
  NAND2_X1 U13377 ( .A1(n11018), .A2(n11019), .ZN(n11017) );
  INV_X1 U13378 ( .A(n10813), .ZN(n10814) );
  NAND2_X1 U13379 ( .A1(n11017), .A2(n10815), .ZN(n10820) );
  XNOR2_X1 U13380 ( .A(n10809), .B(n15138), .ZN(n10992) );
  XNOR2_X1 U13381 ( .A(n10992), .B(n12636), .ZN(n10821) );
  INV_X1 U13382 ( .A(n10816), .ZN(n11072) );
  NAND2_X1 U13383 ( .A1(n11069), .A2(n11072), .ZN(n10818) );
  NAND3_X1 U13384 ( .A1(n11074), .A2(n11070), .A3(n15172), .ZN(n10817) );
  NAND2_X1 U13385 ( .A1(n10818), .A2(n10817), .ZN(n10819) );
  AOI21_X1 U13386 ( .B1(n10820), .B2(n10821), .A(n15043), .ZN(n10824) );
  INV_X1 U13387 ( .A(n10820), .ZN(n10823) );
  NAND2_X1 U13388 ( .A1(n10824), .A2(n10994), .ZN(n10825) );
  OAI211_X1 U13389 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11826), .A(n10826), .B(
        n10825), .ZN(P3_U3158) );
  NAND2_X1 U13390 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n13405) );
  NAND2_X1 U13391 ( .A1(n13376), .A2(n13316), .ZN(n10828) );
  NAND2_X1 U13392 ( .A1(n13374), .A2(n13315), .ZN(n10827) );
  AND2_X1 U13393 ( .A1(n10828), .A2(n10827), .ZN(n14994) );
  INV_X1 U13394 ( .A(n14994), .ZN(n10829) );
  NAND2_X1 U13395 ( .A1(n14576), .A2(n10829), .ZN(n10830) );
  OAI211_X1 U13396 ( .C1(n14581), .C2(n15199), .A(n13405), .B(n10830), .ZN(
        n10838) );
  NAND3_X1 U13397 ( .A1(n10831), .A2(n13334), .A3(n13376), .ZN(n10836) );
  OAI21_X1 U13398 ( .B1(n10833), .B2(n10832), .A(n14574), .ZN(n10835) );
  AOI21_X1 U13399 ( .B1(n10836), .B2(n10835), .A(n10834), .ZN(n10837) );
  AOI211_X1 U13400 ( .C1(n10839), .C2(n14578), .A(n10838), .B(n10837), .ZN(
        n10840) );
  INV_X1 U13401 ( .A(n10840), .ZN(P2_U3185) );
  INV_X1 U13402 ( .A(n11770), .ZN(n14874) );
  INV_X1 U13403 ( .A(n10841), .ZN(n10843) );
  OAI222_X1 U13404 ( .A1(n14874), .A2(P2_U3088), .B1(n13741), .B2(n10843), 
        .C1(n10842), .C2(n13739), .ZN(P2_U3312) );
  INV_X1 U13405 ( .A(n11316), .ZN(n14665) );
  OAI222_X1 U13406 ( .A1(n14410), .A2(n10844), .B1(n14403), .B2(n10843), .C1(
        P1_U3086), .C2(n14665), .ZN(P1_U3340) );
  OAI21_X1 U13407 ( .B1(n10847), .B2(n10846), .A(n10845), .ZN(n10850) );
  NAND2_X1 U13408 ( .A1(n13374), .A2(n13316), .ZN(n10849) );
  NAND2_X1 U13409 ( .A1(n13372), .A2(n13315), .ZN(n10848) );
  NAND2_X1 U13410 ( .A1(n10849), .A2(n10848), .ZN(n10876) );
  AOI21_X1 U13411 ( .B1(n10850), .B2(n14992), .A(n10876), .ZN(n10944) );
  INV_X1 U13412 ( .A(n10851), .ZN(n11009) );
  AOI211_X1 U13413 ( .C1(n10951), .C2(n10852), .A(n13202), .B(n11009), .ZN(
        n10946) );
  INV_X1 U13414 ( .A(n10951), .ZN(n10853) );
  NOR2_X1 U13415 ( .A1(n10853), .A2(n14951), .ZN(n10856) );
  OAI22_X1 U13416 ( .A1(n13512), .A2(n10854), .B1(n10879), .B2(n15200), .ZN(
        n10855) );
  AOI211_X1 U13417 ( .C1(n10946), .C2(n15195), .A(n10856), .B(n10855), .ZN(
        n10862) );
  OAI21_X1 U13418 ( .B1(n10859), .B2(n10858), .A(n10857), .ZN(n10860) );
  INV_X1 U13419 ( .A(n10860), .ZN(n10947) );
  NAND2_X1 U13420 ( .A1(n10947), .A2(n15196), .ZN(n10861) );
  OAI211_X1 U13421 ( .C1(n10944), .C2(n10410), .A(n10862), .B(n10861), .ZN(
        P2_U3256) );
  INV_X1 U13422 ( .A(n10863), .ZN(n10865) );
  AOI22_X1 U13423 ( .A1(n14703), .A2(n11036), .B1(n14241), .B2(n11044), .ZN(
        n10864) );
  OAI21_X1 U13424 ( .B1(n10865), .B2(n14706), .A(n10864), .ZN(n10868) );
  MUX2_X1 U13425 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10866), .S(n14225), .Z(
        n10867) );
  AOI211_X1 U13426 ( .C1(n14229), .C2(n10869), .A(n10868), .B(n10867), .ZN(
        n10870) );
  INV_X1 U13427 ( .A(n10870), .ZN(P1_U3287) );
  INV_X1 U13428 ( .A(n10880), .ZN(n10872) );
  NAND2_X1 U13429 ( .A1(n10872), .A2(n10871), .ZN(n10873) );
  NAND2_X1 U13430 ( .A1(n10874), .A2(n10873), .ZN(n10875) );
  XNOR2_X1 U13431 ( .A(n10951), .B(n13217), .ZN(n11180) );
  NAND2_X1 U13432 ( .A1(n13373), .A2(n13574), .ZN(n11181) );
  XNOR2_X1 U13433 ( .A(n11180), .B(n11181), .ZN(n10881) );
  NAND2_X1 U13434 ( .A1(n14576), .A2(n10876), .ZN(n10877) );
  OAI211_X1 U13435 ( .C1(n14581), .C2(n10879), .A(n10878), .B(n10877), .ZN(
        n10885) );
  AOI22_X1 U13436 ( .A1(n10880), .A2(n14574), .B1(n13334), .B2(n13374), .ZN(
        n10882) );
  NOR3_X1 U13437 ( .A1(n10883), .A2(n10882), .A3(n10881), .ZN(n10884) );
  AOI211_X1 U13438 ( .C1(n10951), .C2(n14578), .A(n10885), .B(n10884), .ZN(
        n10886) );
  OAI21_X1 U13439 ( .B1(n13350), .B2(n11184), .A(n10886), .ZN(P2_U3203) );
  INV_X1 U13440 ( .A(SI_21_), .ZN(n10889) );
  INV_X1 U13441 ( .A(n10887), .ZN(n10888) );
  OAI222_X1 U13442 ( .A1(n14525), .A2(n10889), .B1(n11389), .B2(n10888), .C1(
        P3_U3151), .C2(n10777), .ZN(P3_U3274) );
  NOR2_X1 U13443 ( .A1(n10891), .A2(n10890), .ZN(n12435) );
  NAND2_X1 U13444 ( .A1(n12423), .A2(n13914), .ZN(n10894) );
  NAND2_X1 U13445 ( .A1(n12417), .A2(n10892), .ZN(n10893) );
  NAND2_X1 U13446 ( .A1(n10894), .A2(n10893), .ZN(n10895) );
  XNOR2_X1 U13447 ( .A(n10895), .B(n12459), .ZN(n10902) );
  OAI22_X1 U13448 ( .A1(n12455), .A2(n10896), .B1(n14727), .B2(n10913), .ZN(
        n10901) );
  XNOR2_X1 U13449 ( .A(n10902), .B(n10901), .ZN(n12434) );
  AOI22_X1 U13450 ( .A1(n12422), .A2(n13913), .B1(n10929), .B2(n12423), .ZN(
        n10907) );
  OAI22_X1 U13451 ( .A1(n14736), .A2(n12458), .B1(n10905), .B2(n12456), .ZN(
        n10906) );
  XNOR2_X1 U13452 ( .A(n10906), .B(n12459), .ZN(n10927) );
  NAND2_X1 U13453 ( .A1(n10914), .A2(n12417), .ZN(n10911) );
  NAND2_X1 U13454 ( .A1(n13912), .A2(n12423), .ZN(n10910) );
  NAND2_X1 U13455 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  XNOR2_X1 U13456 ( .A(n10912), .B(n8097), .ZN(n10916) );
  AOI22_X1 U13457 ( .A1(n10914), .A2(n12418), .B1(n12422), .B2(n13912), .ZN(
        n10915) );
  OR2_X1 U13458 ( .A1(n10916), .A2(n10915), .ZN(n11032) );
  NAND2_X1 U13459 ( .A1(n6736), .A2(n11032), .ZN(n10917) );
  XNOR2_X1 U13460 ( .A(n11033), .B(n10917), .ZN(n10925) );
  INV_X1 U13461 ( .A(n14622), .ZN(n13865) );
  AOI22_X1 U13462 ( .A1(n14615), .A2(n10919), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10920) );
  OAI21_X1 U13463 ( .B1(n10921), .B2(n13868), .A(n10920), .ZN(n10922) );
  AOI21_X1 U13464 ( .B1(n10923), .B2(n13865), .A(n10922), .ZN(n10924) );
  OAI21_X1 U13465 ( .B1(n10925), .B2(n13889), .A(n10924), .ZN(P1_U3227) );
  XOR2_X1 U13466 ( .A(n10927), .B(n10926), .Z(n10933) );
  NOR2_X1 U13467 ( .A1(n14622), .A2(n10928), .ZN(n10932) );
  NAND2_X1 U13468 ( .A1(n14618), .A2(n10929), .ZN(n10930) );
  NAND2_X1 U13469 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13969) );
  OAI211_X1 U13470 ( .C1(n14733), .C2(n13831), .A(n10930), .B(n13969), .ZN(
        n10931) );
  AOI211_X1 U13471 ( .C1(n10933), .C2(n14613), .A(n10932), .B(n10931), .ZN(
        n10934) );
  INV_X1 U13472 ( .A(n10934), .ZN(P1_U3230) );
  NOR2_X1 U13473 ( .A1(n14525), .A2(SI_22_), .ZN(n10935) );
  AOI21_X1 U13474 ( .B1(n10936), .B2(P3_STATE_REG_SCAN_IN), .A(n10935), .ZN(
        n10937) );
  OAI21_X1 U13475 ( .B1(n10938), .B2(n11389), .A(n10937), .ZN(n10939) );
  INV_X1 U13476 ( .A(n10939), .ZN(P3_U3273) );
  INV_X1 U13477 ( .A(n10940), .ZN(n10942) );
  OAI222_X1 U13478 ( .A1(n14410), .A2(n10941), .B1(n14403), .B2(n10942), .C1(
        n14027), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13479 ( .A(n14893), .ZN(n10943) );
  OAI222_X1 U13480 ( .A1(P2_U3088), .A2(n10943), .B1(n13739), .B2(n15492), 
        .C1(n13741), .C2(n10942), .ZN(P2_U3311) );
  INV_X1 U13481 ( .A(n10944), .ZN(n10945) );
  AOI211_X1 U13482 ( .C1(n10947), .C2(n15024), .A(n10946), .B(n10945), .ZN(
        n10953) );
  INV_X1 U13483 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10948) );
  NOR2_X1 U13484 ( .A1(n15027), .A2(n10948), .ZN(n10949) );
  AOI21_X1 U13485 ( .B1(n10951), .B2(n9638), .A(n10949), .ZN(n10950) );
  OAI21_X1 U13486 ( .B1(n10953), .B2(n15025), .A(n10950), .ZN(P2_U3457) );
  AOI22_X1 U13487 ( .A1(n10951), .A2(n8743), .B1(n15035), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10952) );
  OAI21_X1 U13488 ( .B1(n10953), .B2(n15035), .A(n10952), .ZN(P2_U3508) );
  NOR3_X1 U13489 ( .A1(n12774), .A2(n15080), .A3(n15099), .ZN(n10963) );
  OR2_X1 U13490 ( .A1(n15071), .A2(n10954), .ZN(n10955) );
  MUX2_X1 U13491 ( .A(n10955), .B(n12765), .S(P3_IR_REG_0__SCAN_IN), .Z(n10962) );
  NAND2_X1 U13492 ( .A1(n15080), .A2(n10956), .ZN(n10958) );
  AOI22_X1 U13493 ( .A1(n15093), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10957) );
  NAND2_X1 U13494 ( .A1(n10958), .A2(n10957), .ZN(n10959) );
  AOI21_X1 U13495 ( .B1(n12774), .B2(n10960), .A(n10959), .ZN(n10961) );
  OAI211_X1 U13496 ( .C1(n10963), .C2(n10967), .A(n10962), .B(n10961), .ZN(
        P3_U3182) );
  INV_X1 U13497 ( .A(n10964), .ZN(n10966) );
  OAI21_X1 U13498 ( .B1(n10966), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10965), .ZN(
        n10977) );
  INV_X1 U13499 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10971) );
  XNOR2_X1 U13500 ( .A(n10968), .B(n10967), .ZN(n10969) );
  AOI22_X1 U13501 ( .A1(n15099), .A2(n10969), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10970) );
  OAI21_X1 U13502 ( .B1(n15088), .B2(n10971), .A(n10970), .ZN(n10976) );
  NAND2_X1 U13503 ( .A1(n10972), .A2(n9081), .ZN(n10973) );
  AOI21_X1 U13504 ( .B1(n10974), .B2(n10973), .A(n15103), .ZN(n10975) );
  AOI211_X1 U13505 ( .C1(n15080), .C2(n10977), .A(n10976), .B(n10975), .ZN(
        n10978) );
  OAI21_X1 U13506 ( .B1(n10979), .B2(n12765), .A(n10978), .ZN(P3_U3183) );
  OAI21_X1 U13507 ( .B1(n10981), .B2(n10983), .A(n10980), .ZN(n10982) );
  INV_X1 U13508 ( .A(n10982), .ZN(n14748) );
  XNOR2_X1 U13509 ( .A(n10984), .B(n10983), .ZN(n10985) );
  AOI222_X1 U13510 ( .A1(n14741), .A2(n10985), .B1(n13908), .B2(n14236), .C1(
        n13910), .C2(n14234), .ZN(n14747) );
  MUX2_X1 U13511 ( .A(n10986), .B(n14747), .S(n14225), .Z(n10990) );
  INV_X1 U13512 ( .A(n11346), .ZN(n10987) );
  AOI211_X1 U13513 ( .C1(n14745), .C2(n11055), .A(n14317), .B(n10987), .ZN(
        n14743) );
  OAI22_X1 U13514 ( .A1(n14244), .A2(n7069), .B1(n14698), .B2(n11574), .ZN(
        n10988) );
  AOI21_X1 U13515 ( .B1(n14743), .B2(n14251), .A(n10988), .ZN(n10989) );
  OAI211_X1 U13516 ( .C1(n14748), .C2(n14248), .A(n10990), .B(n10989), .ZN(
        P1_U3285) );
  INV_X1 U13517 ( .A(n10991), .ZN(n11328) );
  NAND2_X1 U13518 ( .A1(n10992), .A2(n12636), .ZN(n10993) );
  OAI21_X1 U13519 ( .B1(n10996), .B2(n10995), .A(n11137), .ZN(n10997) );
  NAND2_X1 U13520 ( .A1(n10997), .A2(n12613), .ZN(n11001) );
  AND2_X1 U13521 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11122) );
  OAI22_X1 U13522 ( .A1(n12609), .A2(n11492), .B1(n13015), .B2(n12618), .ZN(
        n10998) );
  AOI211_X1 U13523 ( .C1(n10999), .C2(n15040), .A(n11122), .B(n10998), .ZN(
        n11000) );
  OAI211_X1 U13524 ( .C1(n11328), .C2(n11826), .A(n11001), .B(n11000), .ZN(
        P3_U3170) );
  XOR2_X1 U13525 ( .A(n11002), .B(n11006), .Z(n11005) );
  OAI22_X1 U13526 ( .A1(n11004), .A2(n13340), .B1(n11003), .B2(n13342), .ZN(
        n11226) );
  AOI21_X1 U13527 ( .B1(n11005), .B2(n14992), .A(n11226), .ZN(n15012) );
  XOR2_X1 U13528 ( .A(n11007), .B(n11006), .Z(n15015) );
  INV_X1 U13529 ( .A(n11235), .ZN(n15013) );
  INV_X1 U13530 ( .A(n14942), .ZN(n11008) );
  OAI211_X1 U13531 ( .C1(n15013), .C2(n11009), .A(n11008), .B(n14997), .ZN(
        n15011) );
  OAI22_X1 U13532 ( .A1(n13512), .A2(n11010), .B1(n11228), .B2(n15200), .ZN(
        n11011) );
  AOI21_X1 U13533 ( .B1(n11235), .B2(n14937), .A(n11011), .ZN(n11012) );
  OAI21_X1 U13534 ( .B1(n15011), .B2(n13563), .A(n11012), .ZN(n11013) );
  AOI21_X1 U13535 ( .B1(n15015), .B2(n15196), .A(n11013), .ZN(n11014) );
  OAI21_X1 U13536 ( .B1(n14957), .B2(n15012), .A(n11014), .ZN(P2_U3255) );
  NOR2_X1 U13537 ( .A1(n12620), .A2(P3_U3151), .ZN(n15048) );
  INV_X1 U13538 ( .A(n12618), .ZN(n12606) );
  OAI22_X1 U13539 ( .A1(n12609), .A2(n13015), .B1(n12623), .B2(n11015), .ZN(
        n11016) );
  AOI21_X1 U13540 ( .B1(n12606), .B2(n9601), .A(n11016), .ZN(n11022) );
  OAI21_X1 U13541 ( .B1(n11019), .B2(n11018), .A(n11017), .ZN(n11020) );
  NAND2_X1 U13542 ( .A1(n11020), .A2(n12613), .ZN(n11021) );
  OAI211_X1 U13543 ( .C1(n10675), .C2(n15048), .A(n11022), .B(n11021), .ZN(
        P3_U3177) );
  INV_X1 U13544 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15403) );
  AOI21_X1 U13545 ( .B1(n12606), .B2(n15110), .A(n11023), .ZN(n11028) );
  INV_X1 U13546 ( .A(n12075), .ZN(n15109) );
  NAND3_X1 U13547 ( .A1(n10809), .A2(n15113), .A3(n15109), .ZN(n11024) );
  OAI211_X1 U13548 ( .C1(n6735), .C2(n15112), .A(n11025), .B(n11024), .ZN(
        n11026) );
  NAND2_X1 U13549 ( .A1(n11026), .A2(n12613), .ZN(n11027) );
  OAI211_X1 U13550 ( .C1(n15048), .C2(n15403), .A(n11028), .B(n11027), .ZN(
        P3_U3162) );
  INV_X1 U13551 ( .A(SI_23_), .ZN(n11031) );
  NAND2_X1 U13552 ( .A1(n11029), .A2(n13179), .ZN(n11030) );
  OAI211_X1 U13553 ( .C1(n11031), .C2(n14525), .A(n11030), .B(n12274), .ZN(
        P3_U3272) );
  NOR2_X1 U13554 ( .A1(n12455), .A2(n11034), .ZN(n11035) );
  AOI21_X1 U13555 ( .B1(n11036), .B2(n12423), .A(n11035), .ZN(n11248) );
  AOI22_X1 U13556 ( .A1(n11036), .A2(n12417), .B1(n12418), .B2(n13911), .ZN(
        n11037) );
  XNOR2_X1 U13557 ( .A(n11037), .B(n12459), .ZN(n11247) );
  XOR2_X1 U13558 ( .A(n11248), .B(n11247), .Z(n11038) );
  NAND2_X1 U13559 ( .A1(n11039), .A2(n11038), .ZN(n11246) );
  OAI211_X1 U13560 ( .C1(n11039), .C2(n11038), .A(n11246), .B(n14613), .ZN(
        n11046) );
  OAI21_X1 U13561 ( .B1(n13831), .B2(n11041), .A(n11040), .ZN(n11043) );
  NOR2_X1 U13562 ( .A1(n13868), .A2(n7070), .ZN(n11042) );
  AOI211_X1 U13563 ( .C1(n13865), .C2(n11044), .A(n11043), .B(n11042), .ZN(
        n11045) );
  NAND2_X1 U13564 ( .A1(n11046), .A2(n11045), .ZN(P1_U3239) );
  OAI21_X1 U13565 ( .B1(n11048), .B2(n11051), .A(n11047), .ZN(n14709) );
  INV_X1 U13566 ( .A(n14709), .ZN(n11056) );
  NAND2_X1 U13567 ( .A1(n13911), .A2(n14234), .ZN(n11050) );
  NAND2_X1 U13568 ( .A1(n13909), .A2(n14236), .ZN(n11049) );
  NAND2_X1 U13569 ( .A1(n11050), .A2(n11049), .ZN(n11254) );
  XNOR2_X1 U13570 ( .A(n11052), .B(n11051), .ZN(n11053) );
  NOR2_X1 U13571 ( .A1(n11053), .A2(n14329), .ZN(n11054) );
  AOI211_X1 U13572 ( .C1(n14730), .C2(n14709), .A(n11254), .B(n11054), .ZN(
        n14711) );
  OAI211_X1 U13573 ( .C1(n11249), .C2(n6733), .A(n14254), .B(n11055), .ZN(
        n14705) );
  OAI211_X1 U13574 ( .C1(n11056), .C2(n14723), .A(n14711), .B(n14705), .ZN(
        n11061) );
  OAI22_X1 U13575 ( .A1(n14304), .A2(n11249), .B1(n14759), .B2(n14005), .ZN(
        n11057) );
  AOI21_X1 U13576 ( .B1(n11061), .B2(n14759), .A(n11057), .ZN(n11058) );
  INV_X1 U13577 ( .A(n11058), .ZN(P1_U3535) );
  INV_X1 U13578 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11059) );
  OAI22_X1 U13579 ( .A1(n14381), .A2(n11249), .B1(n14752), .B2(n11059), .ZN(
        n11060) );
  AOI21_X1 U13580 ( .B1(n11061), .B2(n14752), .A(n11060), .ZN(n11062) );
  INV_X1 U13581 ( .A(n11062), .ZN(P1_U3480) );
  INV_X1 U13582 ( .A(n13068), .ZN(n13088) );
  NAND2_X1 U13583 ( .A1(n15110), .A2(n11078), .ZN(n12074) );
  INV_X1 U13584 ( .A(n12074), .ZN(n11063) );
  NOR2_X1 U13585 ( .A1(n12075), .A2(n11063), .ZN(n15044) );
  OR3_X1 U13586 ( .A1(n11064), .A2(n15155), .A3(n15044), .ZN(n11066) );
  NAND2_X1 U13587 ( .A1(n15117), .A2(n9601), .ZN(n11065) );
  AND2_X1 U13588 ( .A1(n11066), .A2(n11065), .ZN(n11130) );
  MUX2_X1 U13589 ( .A(n11067), .B(n11130), .S(n15192), .Z(n11068) );
  OAI21_X1 U13590 ( .B1(n13088), .B2(n11078), .A(n11068), .ZN(P3_U3459) );
  AND2_X1 U13591 ( .A1(n11069), .A2(n11073), .ZN(n11071) );
  NAND3_X1 U13592 ( .A1(n11074), .A2(n11073), .A3(n11072), .ZN(n11075) );
  MUX2_X1 U13593 ( .A(n9062), .B(n11130), .S(n15177), .Z(n11077) );
  OAI21_X1 U13594 ( .B1(n13169), .B2(n11078), .A(n11077), .ZN(P3_U3390) );
  INV_X1 U13595 ( .A(n14025), .ZN(n14678) );
  INV_X1 U13596 ( .A(n11079), .ZN(n11080) );
  OAI222_X1 U13597 ( .A1(P1_U3086), .A2(n14678), .B1(n14410), .B2(n15367), 
        .C1(n14403), .C2(n11080), .ZN(P1_U3338) );
  INV_X1 U13598 ( .A(n11773), .ZN(n14909) );
  OAI222_X1 U13599 ( .A1(P2_U3088), .A2(n14909), .B1(n11696), .B2(n11081), 
        .C1(n13729), .C2(n11080), .ZN(P2_U3310) );
  OAI22_X1 U13600 ( .A1(n11084), .A2(n11083), .B1(n11082), .B2(n11099), .ZN(
        n11112) );
  MUX2_X1 U13601 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12733), .Z(n11085) );
  XNOR2_X1 U13602 ( .A(n11085), .B(n11127), .ZN(n11113) );
  INV_X1 U13603 ( .A(n11085), .ZN(n11086) );
  AOI22_X1 U13604 ( .A1(n11112), .A2(n11113), .B1(n11127), .B2(n11086), .ZN(
        n11144) );
  INV_X1 U13605 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15182) );
  MUX2_X1 U13606 ( .A(n11087), .B(n15182), .S(n12725), .Z(n11089) );
  INV_X1 U13607 ( .A(n11089), .ZN(n11088) );
  NOR2_X1 U13608 ( .A1(n11088), .A2(n11159), .ZN(n15059) );
  NOR2_X1 U13609 ( .A1(n11089), .A2(n11164), .ZN(n11143) );
  NOR2_X1 U13610 ( .A1(n15059), .A2(n11143), .ZN(n11090) );
  XNOR2_X1 U13611 ( .A(n11144), .B(n11090), .ZN(n11111) );
  NAND2_X1 U13612 ( .A1(n11092), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13613 ( .A1(n11127), .A2(n11093), .ZN(n11094) );
  AND2_X1 U13614 ( .A1(n11095), .A2(n11094), .ZN(n11116) );
  NAND2_X1 U13615 ( .A1(n11115), .A2(n11116), .ZN(n11114) );
  NAND2_X1 U13616 ( .A1(n11114), .A2(n11095), .ZN(n11158) );
  XNOR2_X1 U13617 ( .A(n11158), .B(n11164), .ZN(n11096) );
  OAI21_X1 U13618 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11096), .A(n6734), .ZN(
        n11097) );
  NAND2_X1 U13619 ( .A1(n12774), .A2(n11097), .ZN(n11108) );
  INV_X1 U13620 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11103) );
  MUX2_X1 U13621 ( .A(n11103), .B(P3_REG1_REG_4__SCAN_IN), .S(n11127), .Z(
        n11119) );
  NAND2_X1 U13622 ( .A1(n11098), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U13623 ( .A1(n11100), .A2(n11099), .ZN(n11101) );
  NAND2_X1 U13624 ( .A1(n11102), .A2(n11101), .ZN(n11120) );
  NAND2_X1 U13625 ( .A1(n11119), .A2(n11120), .ZN(n11118) );
  XNOR2_X1 U13626 ( .A(n11162), .B(n11159), .ZN(n11165) );
  XNOR2_X1 U13627 ( .A(n11165), .B(n15182), .ZN(n11104) );
  NAND2_X1 U13628 ( .A1(n15080), .A2(n11104), .ZN(n11107) );
  NOR2_X1 U13629 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11105), .ZN(n11139) );
  AOI21_X1 U13630 ( .B1(n15093), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11139), .ZN(
        n11106) );
  NAND3_X1 U13631 ( .A1(n11108), .A2(n11107), .A3(n11106), .ZN(n11109) );
  AOI21_X1 U13632 ( .B1(n11164), .B2(n15097), .A(n11109), .ZN(n11110) );
  OAI21_X1 U13633 ( .B1(n15071), .B2(n11111), .A(n11110), .ZN(P3_U3187) );
  XOR2_X1 U13634 ( .A(n11113), .B(n11112), .Z(n11129) );
  OAI21_X1 U13635 ( .B1(n11116), .B2(n11115), .A(n11114), .ZN(n11117) );
  NAND2_X1 U13636 ( .A1(n12774), .A2(n11117), .ZN(n11125) );
  OAI21_X1 U13637 ( .B1(n11120), .B2(n11119), .A(n11118), .ZN(n11121) );
  NAND2_X1 U13638 ( .A1(n15080), .A2(n11121), .ZN(n11124) );
  AOI21_X1 U13639 ( .B1(n15093), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11122), .ZN(
        n11123) );
  NAND3_X1 U13640 ( .A1(n11125), .A2(n11124), .A3(n11123), .ZN(n11126) );
  AOI21_X1 U13641 ( .B1(n11127), .B2(n15097), .A(n11126), .ZN(n11128) );
  OAI21_X1 U13642 ( .B1(n11129), .B2(n15071), .A(n11128), .ZN(P3_U3186) );
  AOI22_X1 U13643 ( .A1(n12991), .A2(n15039), .B1(n12990), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11133) );
  MUX2_X1 U13644 ( .A(n11131), .B(n11130), .S(n6576), .Z(n11132) );
  NAND2_X1 U13645 ( .A1(n11133), .A2(n11132), .ZN(P3_U3233) );
  INV_X1 U13646 ( .A(n11134), .ZN(n11135) );
  NAND2_X1 U13647 ( .A1(n11135), .A2(n11266), .ZN(n11136) );
  XNOR2_X1 U13648 ( .A(n10809), .B(n15146), .ZN(n11491) );
  XNOR2_X1 U13649 ( .A(n11491), .B(n11492), .ZN(n11489) );
  XOR2_X1 U13650 ( .A(n11490), .B(n11489), .Z(n11142) );
  OAI22_X1 U13651 ( .A1(n12609), .A2(n11502), .B1(n11266), .B2(n12618), .ZN(
        n11138) );
  AOI211_X1 U13652 ( .C1(n11274), .C2(n15040), .A(n11139), .B(n11138), .ZN(
        n11141) );
  NAND2_X1 U13653 ( .A1(n12620), .A2(n11273), .ZN(n11140) );
  OAI211_X1 U13654 ( .C1(n11142), .C2(n15043), .A(n11141), .B(n11140), .ZN(
        P3_U3167) );
  NOR2_X1 U13655 ( .A1(n11144), .A2(n11143), .ZN(n15060) );
  INV_X1 U13656 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11145) );
  MUX2_X1 U13657 ( .A(n11146), .B(n11145), .S(n12733), .Z(n11147) );
  NAND2_X1 U13658 ( .A1(n11147), .A2(n15065), .ZN(n11156) );
  INV_X1 U13659 ( .A(n11147), .ZN(n11148) );
  NAND2_X1 U13660 ( .A1(n11148), .A2(n11161), .ZN(n11149) );
  AND2_X1 U13661 ( .A1(n11156), .A2(n11149), .ZN(n15058) );
  INV_X1 U13662 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11150) );
  MUX2_X1 U13663 ( .A(n11151), .B(n11150), .S(n12733), .Z(n11152) );
  INV_X1 U13664 ( .A(n11215), .ZN(n11198) );
  NAND2_X1 U13665 ( .A1(n11152), .A2(n11198), .ZN(n11202) );
  INV_X1 U13666 ( .A(n11152), .ZN(n11153) );
  NAND2_X1 U13667 ( .A1(n11153), .A2(n11215), .ZN(n11154) );
  NAND2_X1 U13668 ( .A1(n11202), .A2(n11154), .ZN(n11155) );
  NAND3_X1 U13669 ( .A1(n15062), .A2(n11156), .A3(n11155), .ZN(n11157) );
  AOI21_X1 U13670 ( .B1(n6729), .B2(n11157), .A(n15071), .ZN(n11175) );
  AOI22_X1 U13671 ( .A1(n15065), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11146), 
        .B2(n11161), .ZN(n15050) );
  NOR2_X1 U13672 ( .A1(n11151), .A2(n11160), .ZN(n11199) );
  AOI21_X1 U13673 ( .B1(n11151), .B2(n11160), .A(n11199), .ZN(n11173) );
  NAND2_X1 U13674 ( .A1(n15097), .A2(n11198), .ZN(n11172) );
  AOI22_X1 U13675 ( .A1(n15065), .A2(n11145), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n11161), .ZN(n15054) );
  INV_X1 U13676 ( .A(n11162), .ZN(n11163) );
  OAI22_X1 U13677 ( .A1(n11165), .A2(n15182), .B1(n11164), .B2(n11163), .ZN(
        n15053) );
  NAND2_X1 U13678 ( .A1(n15054), .A2(n15053), .ZN(n15052) );
  NAND2_X1 U13679 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n11166), .ZN(n11216) );
  OAI21_X1 U13680 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11166), .A(n11216), .ZN(
        n11167) );
  NAND2_X1 U13681 ( .A1(n15080), .A2(n11167), .ZN(n11170) );
  INV_X1 U13682 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11168) );
  NOR2_X1 U13683 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11168), .ZN(n11504) );
  AOI21_X1 U13684 ( .B1(n15093), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11504), .ZN(
        n11169) );
  AND2_X1 U13685 ( .A1(n11170), .A2(n11169), .ZN(n11171) );
  OAI211_X1 U13686 ( .C1(n11173), .C2(n15103), .A(n11172), .B(n11171), .ZN(
        n11174) );
  OR2_X1 U13687 ( .A1(n11175), .A2(n11174), .ZN(P3_U3189) );
  XNOR2_X1 U13688 ( .A(n14938), .B(n13255), .ZN(n11176) );
  NAND2_X1 U13689 ( .A1(n13371), .A2(n13574), .ZN(n11177) );
  NAND2_X1 U13690 ( .A1(n11176), .A2(n11177), .ZN(n11419) );
  INV_X1 U13691 ( .A(n11176), .ZN(n11179) );
  INV_X1 U13692 ( .A(n11177), .ZN(n11178) );
  NAND2_X1 U13693 ( .A1(n11179), .A2(n11178), .ZN(n11421) );
  NAND2_X1 U13694 ( .A1(n11419), .A2(n11421), .ZN(n11190) );
  INV_X1 U13695 ( .A(n11180), .ZN(n11182) );
  NAND2_X1 U13696 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  XNOR2_X1 U13697 ( .A(n11235), .B(n13255), .ZN(n11185) );
  NAND2_X1 U13698 ( .A1(n13372), .A2(n13574), .ZN(n11186) );
  XNOR2_X1 U13699 ( .A(n11185), .B(n11186), .ZN(n11232) );
  INV_X1 U13700 ( .A(n11185), .ZN(n11188) );
  INV_X1 U13701 ( .A(n11186), .ZN(n11187) );
  NAND2_X1 U13702 ( .A1(n11188), .A2(n11187), .ZN(n11189) );
  XOR2_X1 U13703 ( .A(n11190), .B(n11420), .Z(n11196) );
  OAI22_X1 U13704 ( .A1(n11192), .A2(n13340), .B1(n11191), .B2(n13342), .ZN(
        n14933) );
  AOI22_X1 U13705 ( .A1(n14576), .A2(n14933), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11193) );
  OAI21_X1 U13706 ( .B1(n14935), .B2(n14581), .A(n11193), .ZN(n11194) );
  AOI21_X1 U13707 ( .B1(n14938), .B2(n14578), .A(n11194), .ZN(n11195) );
  OAI21_X1 U13708 ( .B1(n11196), .B2(n13350), .A(n11195), .ZN(P2_U3208) );
  NOR2_X1 U13709 ( .A1(n11198), .A2(n11197), .ZN(n11200) );
  NOR2_X1 U13710 ( .A1(n11200), .A2(n11199), .ZN(n15075) );
  AOI22_X1 U13711 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15081), .B1(n11213), 
        .B2(n9196), .ZN(n15074) );
  NOR2_X1 U13712 ( .A1(n15075), .A2(n15074), .ZN(n15073) );
  AOI21_X1 U13713 ( .B1(n11207), .B2(n11201), .A(n11465), .ZN(n11225) );
  MUX2_X1 U13714 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12725), .Z(n11204) );
  INV_X1 U13715 ( .A(n11204), .ZN(n11205) );
  INV_X1 U13716 ( .A(n11202), .ZN(n11203) );
  XNOR2_X1 U13717 ( .A(n11204), .B(n11213), .ZN(n15070) );
  AOI21_X1 U13718 ( .B1(n15081), .B2(n11205), .A(n15069), .ZN(n11209) );
  INV_X1 U13719 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11206) );
  MUX2_X1 U13720 ( .A(n11207), .B(n11206), .S(n12725), .Z(n11208) );
  NOR2_X1 U13721 ( .A1(n11208), .A2(n11464), .ZN(n11210) );
  AND2_X1 U13722 ( .A1(n11208), .A2(n11464), .ZN(n11469) );
  OAI21_X1 U13723 ( .B1(n11210), .B2(n11469), .A(n11209), .ZN(n11211) );
  OAI21_X1 U13724 ( .B1(n6898), .B2(n11469), .A(n11211), .ZN(n11212) );
  NAND2_X1 U13725 ( .A1(n11212), .A2(n15099), .ZN(n11224) );
  INV_X1 U13726 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U13727 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11213), .B1(n15081), 
        .B2(n15186), .ZN(n15078) );
  NAND2_X1 U13728 ( .A1(n11215), .A2(n11214), .ZN(n11217) );
  NAND2_X1 U13729 ( .A1(n11217), .A2(n11216), .ZN(n15077) );
  NAND2_X1 U13730 ( .A1(n15078), .A2(n15077), .ZN(n15076) );
  OAI21_X1 U13731 ( .B1(n15081), .B2(n15186), .A(n15076), .ZN(n11472) );
  OAI21_X1 U13732 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n11218), .A(n11474), .ZN(
        n11222) );
  NOR2_X1 U13733 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11219), .ZN(n11737) );
  AOI21_X1 U13734 ( .B1(n15093), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11737), .ZN(
        n11220) );
  OAI21_X1 U13735 ( .B1(n12765), .B2(n11473), .A(n11220), .ZN(n11221) );
  AOI21_X1 U13736 ( .B1(n11222), .B2(n15080), .A(n11221), .ZN(n11223) );
  OAI211_X1 U13737 ( .C1(n11225), .C2(n15103), .A(n11224), .B(n11223), .ZN(
        P3_U3191) );
  NAND2_X1 U13738 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14826)
         );
  NAND2_X1 U13739 ( .A1(n14576), .A2(n11226), .ZN(n11227) );
  OAI211_X1 U13740 ( .C1(n14581), .C2(n11228), .A(n14826), .B(n11227), .ZN(
        n11234) );
  INV_X1 U13741 ( .A(n11229), .ZN(n11230) );
  AOI211_X1 U13742 ( .C1(n11232), .C2(n11231), .A(n13350), .B(n11230), .ZN(
        n11233) );
  AOI211_X1 U13743 ( .C1(n11235), .C2(n14578), .A(n11234), .B(n11233), .ZN(
        n11236) );
  INV_X1 U13744 ( .A(n11236), .ZN(P2_U3189) );
  XNOR2_X1 U13745 ( .A(n11237), .B(n11241), .ZN(n11238) );
  AOI22_X1 U13746 ( .A1(n13316), .A2(n13371), .B1(n13369), .B2(n13315), .ZN(
        n11428) );
  OAI21_X1 U13747 ( .B1(n11238), .B2(n13530), .A(n11428), .ZN(n11352) );
  INV_X1 U13748 ( .A(n11352), .ZN(n11245) );
  AOI211_X1 U13749 ( .C1(n11431), .C2(n14941), .A(n13202), .B(n7213), .ZN(
        n11353) );
  NOR2_X1 U13750 ( .A1(n11356), .A2(n14951), .ZN(n11240) );
  OAI22_X1 U13751 ( .A1(n13512), .A2(n11742), .B1(n11426), .B2(n15200), .ZN(
        n11239) );
  AOI211_X1 U13752 ( .C1(n11353), .C2(n15195), .A(n11240), .B(n11239), .ZN(
        n11244) );
  XNOR2_X1 U13753 ( .A(n11242), .B(n11241), .ZN(n11354) );
  NAND2_X1 U13754 ( .A1(n11354), .A2(n15196), .ZN(n11243) );
  OAI211_X1 U13755 ( .C1(n11245), .C2(n10410), .A(n11244), .B(n11243), .ZN(
        P2_U3253) );
  OAI21_X1 U13756 ( .B1(n11248), .B2(n11247), .A(n11246), .ZN(n11253) );
  OAI22_X1 U13757 ( .A1(n11249), .A2(n12458), .B1(n11575), .B2(n12456), .ZN(
        n11250) );
  XNOR2_X1 U13758 ( .A(n11250), .B(n12459), .ZN(n11564) );
  NOR2_X1 U13759 ( .A1(n12455), .A2(n11575), .ZN(n11251) );
  AOI21_X1 U13760 ( .B1(n14702), .B2(n12423), .A(n11251), .ZN(n11565) );
  XNOR2_X1 U13761 ( .A(n11564), .B(n11565), .ZN(n11252) );
  OAI211_X1 U13762 ( .C1(n11253), .C2(n11252), .A(n11568), .B(n14613), .ZN(
        n11258) );
  NAND2_X1 U13763 ( .A1(n14615), .A2(n11254), .ZN(n11255) );
  NAND2_X1 U13764 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13999) );
  OAI211_X1 U13765 ( .C1(n14622), .C2(n14699), .A(n11255), .B(n13999), .ZN(
        n11256) );
  AOI21_X1 U13766 ( .B1(n14702), .B2(n14618), .A(n11256), .ZN(n11257) );
  NAND2_X1 U13767 ( .A1(n11258), .A2(n11257), .ZN(P1_U3213) );
  OR2_X1 U13768 ( .A1(n11259), .A2(n12237), .ZN(n11260) );
  NAND2_X1 U13769 ( .A1(n11261), .A2(n11260), .ZN(n11269) );
  INV_X1 U13770 ( .A(n11269), .ZN(n15147) );
  INV_X1 U13771 ( .A(n11262), .ZN(n13027) );
  NAND2_X1 U13772 ( .A1(n6576), .A2(n13027), .ZN(n12875) );
  NAND2_X1 U13773 ( .A1(n11263), .A2(n12237), .ZN(n11264) );
  NAND2_X1 U13774 ( .A1(n11362), .A2(n11264), .ZN(n11268) );
  NAND2_X1 U13775 ( .A1(n15117), .A2(n12633), .ZN(n11265) );
  OAI21_X1 U13776 ( .B1(n11266), .B2(n15120), .A(n11265), .ZN(n11267) );
  AOI21_X1 U13777 ( .B1(n11268), .B2(n15114), .A(n11267), .ZN(n11271) );
  INV_X1 U13778 ( .A(n12867), .ZN(n13024) );
  NAND2_X1 U13779 ( .A1(n11269), .A2(n13024), .ZN(n11270) );
  NAND2_X1 U13780 ( .A1(n11271), .A2(n11270), .ZN(n15148) );
  MUX2_X1 U13781 ( .A(n15148), .B(P3_REG2_REG_5__SCAN_IN), .S(n15129), .Z(
        n11272) );
  INV_X1 U13782 ( .A(n11272), .ZN(n11276) );
  AOI22_X1 U13783 ( .A1(n12991), .A2(n11274), .B1(n12990), .B2(n11273), .ZN(
        n11275) );
  OAI211_X1 U13784 ( .C1(n15147), .C2(n12875), .A(n11276), .B(n11275), .ZN(
        P3_U3228) );
  INV_X1 U13785 ( .A(n11277), .ZN(n11280) );
  OAI211_X1 U13786 ( .C1(n11280), .C2(n11279), .A(n14741), .B(n11278), .ZN(
        n11281) );
  OAI21_X1 U13787 ( .B1(n11860), .B2(n14140), .A(n11281), .ZN(n11390) );
  INV_X1 U13788 ( .A(n11390), .ZN(n11293) );
  INV_X1 U13789 ( .A(n11863), .ZN(n11285) );
  INV_X1 U13790 ( .A(n11282), .ZN(n11345) );
  OAI211_X1 U13791 ( .C1(n11285), .C2(n11345), .A(n14254), .B(n11440), .ZN(
        n11283) );
  OAI21_X1 U13792 ( .B1(n11998), .B2(n14142), .A(n11283), .ZN(n11391) );
  OAI22_X1 U13793 ( .A1(n14225), .A2(n11284), .B1(n11859), .B2(n14698), .ZN(
        n11287) );
  NOR2_X1 U13794 ( .A1(n11285), .A2(n14244), .ZN(n11286) );
  AOI211_X1 U13795 ( .C1(n11391), .C2(n14251), .A(n11287), .B(n11286), .ZN(
        n11292) );
  OAI21_X1 U13796 ( .B1(n11290), .B2(n11289), .A(n11288), .ZN(n11392) );
  NAND2_X1 U13797 ( .A1(n11392), .A2(n14229), .ZN(n11291) );
  OAI211_X1 U13798 ( .C1(n11293), .C2(n14712), .A(n11292), .B(n11291), .ZN(
        P1_U3283) );
  INV_X1 U13799 ( .A(n11295), .ZN(n12232) );
  XNOR2_X1 U13800 ( .A(n11294), .B(n12232), .ZN(n15139) );
  AOI22_X1 U13801 ( .A1(n12985), .A2(n15116), .B1(n15117), .B2(n12635), .ZN(
        n11301) );
  INV_X1 U13802 ( .A(n13021), .ZN(n11297) );
  OAI21_X1 U13803 ( .B1(n11297), .B2(n11296), .A(n11295), .ZN(n11299) );
  NAND3_X1 U13804 ( .A1(n11299), .A2(n15114), .A3(n11298), .ZN(n11300) );
  OAI211_X1 U13805 ( .C1(n15139), .C2(n12867), .A(n11301), .B(n11300), .ZN(
        n15141) );
  INV_X1 U13806 ( .A(n15141), .ZN(n11307) );
  INV_X1 U13807 ( .A(n12875), .ZN(n11383) );
  INV_X1 U13808 ( .A(n15139), .ZN(n11305) );
  AOI22_X1 U13809 ( .A1(n12991), .A2(n11302), .B1(n12990), .B2(n9109), .ZN(
        n11303) );
  OAI21_X1 U13810 ( .B1(n9111), .B2(n6576), .A(n11303), .ZN(n11304) );
  AOI21_X1 U13811 ( .B1(n11383), .B2(n11305), .A(n11304), .ZN(n11306) );
  OAI21_X1 U13812 ( .B1(n15129), .B2(n11307), .A(n11306), .ZN(P3_U3230) );
  OAI21_X1 U13813 ( .B1(n11315), .B2(n10487), .A(n11308), .ZN(n11309) );
  INV_X1 U13814 ( .A(n11309), .ZN(n11310) );
  XNOR2_X1 U13815 ( .A(n11309), .B(n11316), .ZN(n14662) );
  NOR2_X1 U13816 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14662), .ZN(n14661) );
  AOI21_X1 U13817 ( .B1(n11310), .B2(n14665), .A(n14661), .ZN(n11313) );
  INV_X1 U13818 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11311) );
  MUX2_X1 U13819 ( .A(n11311), .B(P1_REG2_REG_16__SCAN_IN), .S(n14027), .Z(
        n11312) );
  NAND2_X1 U13820 ( .A1(n11312), .A2(n11313), .ZN(n14020) );
  OAI211_X1 U13821 ( .C1(n11313), .C2(n11312), .A(n14038), .B(n14020), .ZN(
        n11324) );
  NAND2_X1 U13822 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13798)
         );
  AOI21_X1 U13823 ( .B1(n7887), .B2(n11315), .A(n11314), .ZN(n11317) );
  INV_X1 U13824 ( .A(n11317), .ZN(n11318) );
  XNOR2_X1 U13825 ( .A(n11317), .B(n11316), .ZN(n14660) );
  NOR2_X1 U13826 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14660), .ZN(n14659) );
  AOI21_X1 U13827 ( .B1(n14665), .B2(n11318), .A(n14659), .ZN(n11320) );
  XNOR2_X1 U13828 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14027), .ZN(n11319) );
  NAND2_X1 U13829 ( .A1(n11319), .A2(n11320), .ZN(n14026) );
  OAI211_X1 U13830 ( .C1(n11320), .C2(n11319), .A(n14037), .B(n14026), .ZN(
        n11321) );
  NAND2_X1 U13831 ( .A1(n13798), .A2(n11321), .ZN(n11322) );
  AOI21_X1 U13832 ( .B1(n14655), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11322), 
        .ZN(n11323) );
  OAI211_X1 U13833 ( .C1(n14691), .C2(n14027), .A(n11324), .B(n11323), .ZN(
        P1_U3259) );
  OR2_X1 U13834 ( .A1(n11325), .A2(n9605), .ZN(n11327) );
  NAND2_X1 U13835 ( .A1(n11327), .A2(n11326), .ZN(n15145) );
  OAI22_X1 U13836 ( .A1(n13004), .A2(n15142), .B1(n11328), .B2(n15123), .ZN(
        n11334) );
  XNOR2_X1 U13837 ( .A(n11329), .B(n12096), .ZN(n11332) );
  NAND2_X1 U13838 ( .A1(n15145), .A2(n13024), .ZN(n11331) );
  AOI22_X1 U13839 ( .A1(n12985), .A2(n12636), .B1(n15117), .B2(n12634), .ZN(
        n11330) );
  OAI211_X1 U13840 ( .C1(n13019), .C2(n11332), .A(n11331), .B(n11330), .ZN(
        n15143) );
  MUX2_X1 U13841 ( .A(n15143), .B(P3_REG2_REG_4__SCAN_IN), .S(n15129), .Z(
        n11333) );
  AOI211_X1 U13842 ( .C1(n11383), .C2(n15145), .A(n11334), .B(n11333), .ZN(
        n11335) );
  INV_X1 U13843 ( .A(n11335), .ZN(P3_U3229) );
  OAI21_X1 U13844 ( .B1(n11337), .B2(n11341), .A(n11336), .ZN(n11457) );
  INV_X1 U13845 ( .A(n11457), .ZN(n11351) );
  INV_X1 U13846 ( .A(n11338), .ZN(n11339) );
  AOI21_X1 U13847 ( .B1(n11341), .B2(n11340), .A(n11339), .ZN(n11344) );
  AOI22_X1 U13848 ( .A1(n14234), .A2(n13909), .B1(n13907), .B2(n14236), .ZN(
        n11343) );
  NAND2_X1 U13849 ( .A1(n11457), .A2(n14730), .ZN(n11342) );
  OAI211_X1 U13850 ( .C1(n11344), .C2(n14329), .A(n11343), .B(n11342), .ZN(
        n11455) );
  NAND2_X1 U13851 ( .A1(n11455), .A2(n14225), .ZN(n11350) );
  AOI211_X1 U13852 ( .C1(n11716), .C2(n11346), .A(n14317), .B(n11345), .ZN(
        n11456) );
  INV_X1 U13853 ( .A(n11716), .ZN(n11726) );
  NOR2_X1 U13854 ( .A1(n11726), .A2(n14244), .ZN(n11348) );
  OAI22_X1 U13855 ( .A1(n14225), .A2(n10160), .B1(n11720), .B2(n14698), .ZN(
        n11347) );
  AOI211_X1 U13856 ( .C1(n11456), .C2(n14251), .A(n11348), .B(n11347), .ZN(
        n11349) );
  OAI211_X1 U13857 ( .C1(n11351), .C2(n14697), .A(n11350), .B(n11349), .ZN(
        P1_U3284) );
  AOI211_X1 U13858 ( .C1(n11354), .C2(n15024), .A(n11353), .B(n11352), .ZN(
        n11360) );
  INV_X1 U13859 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11355) );
  OAI22_X1 U13860 ( .A1(n11356), .A2(n13718), .B1(n15027), .B2(n11355), .ZN(
        n11357) );
  INV_X1 U13861 ( .A(n11357), .ZN(n11358) );
  OAI21_X1 U13862 ( .B1(n11360), .B2(n15025), .A(n11358), .ZN(P2_U3466) );
  AOI22_X1 U13863 ( .A1(n11431), .A2(n8743), .B1(n15035), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11359) );
  OAI21_X1 U13864 ( .B1(n11360), .B2(n15035), .A(n11359), .ZN(P2_U3511) );
  XOR2_X1 U13865 ( .A(n11361), .B(n12233), .Z(n15151) );
  AOI22_X1 U13866 ( .A1(n12985), .A2(n12634), .B1(n15117), .B2(n12632), .ZN(
        n11368) );
  INV_X1 U13867 ( .A(n11362), .ZN(n11364) );
  OAI21_X1 U13868 ( .B1(n11364), .B2(n11363), .A(n12233), .ZN(n11366) );
  NAND3_X1 U13869 ( .A1(n11366), .A2(n15114), .A3(n11365), .ZN(n11367) );
  OAI211_X1 U13870 ( .C1(n15151), .C2(n12867), .A(n11368), .B(n11367), .ZN(
        n15153) );
  INV_X1 U13871 ( .A(n15153), .ZN(n11373) );
  INV_X1 U13872 ( .A(n15151), .ZN(n11371) );
  AOI22_X1 U13873 ( .A1(n12991), .A2(n11496), .B1(n12990), .B2(n11515), .ZN(
        n11369) );
  OAI21_X1 U13874 ( .B1(n11146), .B2(n6576), .A(n11369), .ZN(n11370) );
  AOI21_X1 U13875 ( .B1(n11371), .B2(n11383), .A(n11370), .ZN(n11372) );
  OAI21_X1 U13876 ( .B1(n11373), .B2(n15129), .A(n11372), .ZN(P3_U3227) );
  XNOR2_X1 U13877 ( .A(n11374), .B(n12235), .ZN(n15157) );
  NAND2_X1 U13878 ( .A1(n15157), .A2(n13024), .ZN(n11380) );
  XNOR2_X1 U13879 ( .A(n11375), .B(n12235), .ZN(n11378) );
  NAND2_X1 U13880 ( .A1(n15117), .A2(n11728), .ZN(n11376) );
  OAI21_X1 U13881 ( .B1(n11502), .B2(n15120), .A(n11376), .ZN(n11377) );
  AOI21_X1 U13882 ( .B1(n11378), .B2(n15114), .A(n11377), .ZN(n11379) );
  AOI22_X1 U13883 ( .A1(n12991), .A2(n15154), .B1(n12990), .B2(n11488), .ZN(
        n11381) );
  OAI21_X1 U13884 ( .B1(n11151), .B2(n6576), .A(n11381), .ZN(n11382) );
  AOI21_X1 U13885 ( .B1(n15157), .B2(n11383), .A(n11382), .ZN(n11384) );
  OAI21_X1 U13886 ( .B1(n15159), .B2(n15129), .A(n11384), .ZN(P3_U3226) );
  INV_X1 U13887 ( .A(n11385), .ZN(n11388) );
  INV_X1 U13888 ( .A(SI_24_), .ZN(n11386) );
  OAI222_X1 U13889 ( .A1(n11389), .A2(n11388), .B1(P3_U3151), .B2(n11387), 
        .C1(n11386), .C2(n14525), .ZN(P3_U3271) );
  AOI211_X1 U13890 ( .C1(n14626), .C2(n11392), .A(n11391), .B(n11390), .ZN(
        n11395) );
  AOI22_X1 U13891 ( .A1(n11863), .A2(n8207), .B1(n14757), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11393) );
  OAI21_X1 U13892 ( .B1(n11395), .B2(n14757), .A(n11393), .ZN(P1_U3538) );
  AOI22_X1 U13893 ( .A1(n11863), .A2(n8212), .B1(n14751), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n11394) );
  OAI21_X1 U13894 ( .B1(n11395), .B2(n14751), .A(n11394), .ZN(P1_U3489) );
  XNOR2_X1 U13895 ( .A(n11396), .B(n8458), .ZN(n14603) );
  INV_X1 U13896 ( .A(n14603), .ZN(n11413) );
  INV_X1 U13897 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11397) );
  OAI22_X1 U13898 ( .A1(n13512), .A2(n11397), .B1(n11449), .B2(n15200), .ZN(
        n11398) );
  AOI21_X1 U13899 ( .B1(n14598), .B2(n14937), .A(n11398), .ZN(n11412) );
  NAND2_X1 U13900 ( .A1(n11400), .A2(n11399), .ZN(n11401) );
  NAND2_X1 U13901 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  NAND2_X1 U13902 ( .A1(n11403), .A2(n14992), .ZN(n11406) );
  NAND2_X1 U13903 ( .A1(n13368), .A2(n13315), .ZN(n11405) );
  NAND2_X1 U13904 ( .A1(n13370), .A2(n13316), .ZN(n11404) );
  AND2_X1 U13905 ( .A1(n11405), .A2(n11404), .ZN(n11450) );
  NAND2_X1 U13906 ( .A1(n11406), .A2(n11450), .ZN(n14602) );
  NAND2_X1 U13907 ( .A1(n14598), .A2(n11407), .ZN(n11408) );
  NAND3_X1 U13908 ( .A1(n11585), .A2(n14997), .A3(n11408), .ZN(n14600) );
  NOR2_X1 U13909 ( .A1(n14600), .A2(n11409), .ZN(n11410) );
  OAI21_X1 U13910 ( .B1(n14602), .B2(n11410), .A(n13512), .ZN(n11411) );
  OAI211_X1 U13911 ( .C1(n11413), .C2(n13604), .A(n11412), .B(n11411), .ZN(
        P2_U3252) );
  XNOR2_X1 U13912 ( .A(n11431), .B(n13255), .ZN(n11414) );
  NAND2_X1 U13913 ( .A1(n13370), .A2(n13574), .ZN(n11415) );
  NAND2_X1 U13914 ( .A1(n11414), .A2(n11415), .ZN(n11447) );
  INV_X1 U13915 ( .A(n11414), .ZN(n11417) );
  INV_X1 U13916 ( .A(n11415), .ZN(n11416) );
  NAND2_X1 U13917 ( .A1(n11417), .A2(n11416), .ZN(n11418) );
  NAND2_X1 U13918 ( .A1(n11447), .A2(n11418), .ZN(n11425) );
  NAND2_X1 U13919 ( .A1(n11422), .A2(n11421), .ZN(n11424) );
  INV_X1 U13920 ( .A(n11448), .ZN(n11423) );
  AOI21_X1 U13921 ( .B1(n11425), .B2(n11424), .A(n11423), .ZN(n11433) );
  NOR2_X1 U13922 ( .A1(n14581), .A2(n11426), .ZN(n11430) );
  OAI21_X1 U13923 ( .B1(n13318), .B2(n11428), .A(n11427), .ZN(n11429) );
  AOI211_X1 U13924 ( .C1(n11431), .C2(n14578), .A(n11430), .B(n11429), .ZN(
        n11432) );
  OAI21_X1 U13925 ( .B1(n11433), .B2(n13350), .A(n11432), .ZN(P2_U3196) );
  XNOR2_X1 U13926 ( .A(n11435), .B(n11434), .ZN(n11436) );
  OAI222_X1 U13927 ( .A1(n14142), .A2(n13840), .B1(n14140), .B2(n12010), .C1(
        n11436), .C2(n14329), .ZN(n11521) );
  INV_X1 U13928 ( .A(n11521), .ZN(n11446) );
  OAI21_X1 U13929 ( .B1(n11439), .B2(n11438), .A(n11437), .ZN(n11523) );
  AOI211_X1 U13930 ( .C1(n11525), .C2(n11440), .A(n14317), .B(n11655), .ZN(
        n11522) );
  NAND2_X1 U13931 ( .A1(n11522), .A2(n14251), .ZN(n11443) );
  INV_X1 U13932 ( .A(n11441), .ZN(n12013) );
  AOI22_X1 U13933 ( .A1(n14712), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12013), 
        .B2(n14241), .ZN(n11442) );
  OAI211_X1 U13934 ( .C1(n12016), .C2(n14244), .A(n11443), .B(n11442), .ZN(
        n11444) );
  AOI21_X1 U13935 ( .B1(n11523), .B2(n14229), .A(n11444), .ZN(n11445) );
  OAI21_X1 U13936 ( .B1(n11446), .B2(n14712), .A(n11445), .ZN(P1_U3282) );
  NAND2_X1 U13937 ( .A1(n13369), .A2(n13574), .ZN(n11869) );
  XNOR2_X1 U13938 ( .A(n11868), .B(n11869), .ZN(n11866) );
  XNOR2_X1 U13939 ( .A(n11867), .B(n11866), .ZN(n11454) );
  NOR2_X1 U13940 ( .A1(n14581), .A2(n11449), .ZN(n11452) );
  OAI22_X1 U13941 ( .A1(n13318), .A2(n11450), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8447), .ZN(n11451) );
  AOI211_X1 U13942 ( .C1(n14598), .C2(n14578), .A(n11452), .B(n11451), .ZN(
        n11453) );
  OAI21_X1 U13943 ( .B1(n11454), .B2(n13350), .A(n11453), .ZN(P2_U3206) );
  INV_X1 U13944 ( .A(n14723), .ZN(n14721) );
  AOI211_X1 U13945 ( .C1(n14721), .C2(n11457), .A(n11456), .B(n11455), .ZN(
        n11460) );
  AOI22_X1 U13946 ( .A1(n11716), .A2(n8212), .B1(n14751), .B2(
        P1_REG0_REG_9__SCAN_IN), .ZN(n11458) );
  OAI21_X1 U13947 ( .B1(n11460), .B2(n14751), .A(n11458), .ZN(P1_U3486) );
  AOI22_X1 U13948 ( .A1(n11716), .A2(n8207), .B1(n14757), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11459) );
  OAI21_X1 U13949 ( .B1(n11460), .B2(n14757), .A(n11459), .ZN(P1_U3537) );
  INV_X1 U13950 ( .A(n11461), .ZN(n11486) );
  OAI222_X1 U13951 ( .A1(n13739), .A2(n11462), .B1(n13741), .B2(n11486), .C1(
        n14925), .C2(P2_U3088), .ZN(P2_U3309) );
  NOR2_X1 U13952 ( .A1(n11464), .A2(n11463), .ZN(n11466) );
  NAND2_X1 U13953 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11471), .ZN(n11467) );
  OAI21_X1 U13954 ( .B1(n11471), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11467), 
        .ZN(n15102) );
  AOI21_X1 U13955 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11471), .A(n15101), 
        .ZN(n11533) );
  AOI21_X1 U13956 ( .B1(n11670), .B2(n11468), .A(n11534), .ZN(n11485) );
  MUX2_X1 U13957 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12725), .Z(n11470) );
  XNOR2_X1 U13958 ( .A(n11470), .B(n11471), .ZN(n15095) );
  MUX2_X1 U13959 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12725), .Z(n11537) );
  XNOR2_X1 U13960 ( .A(n11537), .B(n11539), .ZN(n11540) );
  XNOR2_X1 U13961 ( .A(n11541), .B(n11540), .ZN(n11483) );
  NAND2_X1 U13962 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11471), .ZN(n11476) );
  INV_X1 U13963 ( .A(n11471), .ZN(n15098) );
  INV_X1 U13964 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U13965 ( .A1(n15098), .A2(n15190), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11471), .ZN(n15092) );
  NAND2_X1 U13966 ( .A1(n11473), .A2(n11472), .ZN(n11475) );
  NAND2_X1 U13967 ( .A1(n11475), .A2(n11474), .ZN(n15091) );
  NAND2_X1 U13968 ( .A1(n15092), .A2(n15091), .ZN(n15090) );
  NAND2_X1 U13969 ( .A1(n11476), .A2(n15090), .ZN(n11544) );
  XOR2_X1 U13970 ( .A(n11545), .B(n11544), .Z(n11477) );
  OAI21_X1 U13971 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11477), .A(n11546), 
        .ZN(n11478) );
  NAND2_X1 U13972 ( .A1(n11478), .A2(n15080), .ZN(n11481) );
  NOR2_X1 U13973 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11479), .ZN(n12585) );
  AOI21_X1 U13974 ( .B1(n15093), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12585), 
        .ZN(n11480) );
  OAI211_X1 U13975 ( .C1(n12765), .C2(n11545), .A(n11481), .B(n11480), .ZN(
        n11482) );
  AOI21_X1 U13976 ( .B1(n11483), .B2(n15099), .A(n11482), .ZN(n11484) );
  OAI21_X1 U13977 ( .B1(n11485), .B2(n15103), .A(n11484), .ZN(P3_U3193) );
  INV_X1 U13978 ( .A(n14030), .ZN(n14690) );
  INV_X1 U13979 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11487) );
  OAI222_X1 U13980 ( .A1(P1_U3086), .A2(n14690), .B1(n14410), .B2(n11487), 
        .C1(n14413), .C2(n11486), .ZN(P1_U3337) );
  INV_X1 U13981 ( .A(n11488), .ZN(n11507) );
  NAND2_X1 U13982 ( .A1(n11490), .A2(n11489), .ZN(n11495) );
  INV_X1 U13983 ( .A(n11491), .ZN(n11493) );
  NAND2_X1 U13984 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  NAND2_X1 U13985 ( .A1(n11495), .A2(n11494), .ZN(n11511) );
  XNOR2_X1 U13986 ( .A(n10809), .B(n11496), .ZN(n11498) );
  XNOR2_X1 U13987 ( .A(n11498), .B(n11502), .ZN(n11512) );
  INV_X1 U13988 ( .A(n11498), .ZN(n11499) );
  NAND2_X1 U13989 ( .A1(n11499), .A2(n12633), .ZN(n11500) );
  XNOR2_X1 U13990 ( .A(n12235), .B(n10809), .ZN(n11594) );
  OAI211_X1 U13991 ( .C1(n11501), .C2(n11594), .A(n11597), .B(n12613), .ZN(
        n11506) );
  OAI22_X1 U13992 ( .A1(n12609), .A2(n11735), .B1(n11502), .B2(n12618), .ZN(
        n11503) );
  AOI211_X1 U13993 ( .C1(n15154), .C2(n15040), .A(n11504), .B(n11503), .ZN(
        n11505) );
  OAI211_X1 U13994 ( .C1(n11507), .C2(n11826), .A(n11506), .B(n11505), .ZN(
        P3_U3153) );
  AOI22_X1 U13995 ( .A1(n12606), .A2(n12634), .B1(n15038), .B2(n12632), .ZN(
        n11508) );
  NAND2_X1 U13996 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15066) );
  OAI211_X1 U13997 ( .C1(n15150), .C2(n12623), .A(n11508), .B(n15066), .ZN(
        n11514) );
  INV_X1 U13998 ( .A(n11509), .ZN(n11510) );
  AOI211_X1 U13999 ( .C1(n11512), .C2(n11511), .A(n15043), .B(n11510), .ZN(
        n11513) );
  AOI211_X1 U14000 ( .C1(n11515), .C2(n12620), .A(n11514), .B(n11513), .ZN(
        n11516) );
  INV_X1 U14001 ( .A(n11516), .ZN(P3_U3179) );
  INV_X1 U14002 ( .A(n11517), .ZN(n11519) );
  INV_X1 U14003 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11518) );
  OAI222_X1 U14004 ( .A1(n14040), .A2(P1_U3086), .B1(n14403), .B2(n11519), 
        .C1(n11518), .C2(n14410), .ZN(P1_U3336) );
  OAI222_X1 U14005 ( .A1(n13739), .A2(n11520), .B1(n13741), .B2(n11519), .C1(
        n13581), .C2(P2_U3088), .ZN(P2_U3308) );
  AOI211_X1 U14006 ( .C1(n14626), .C2(n11523), .A(n11522), .B(n11521), .ZN(
        n11527) );
  AOI22_X1 U14007 ( .A1(n11525), .A2(n8207), .B1(n14757), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11524) );
  OAI21_X1 U14008 ( .B1(n11527), .B2(n14757), .A(n11524), .ZN(P1_U3539) );
  AOI22_X1 U14009 ( .A1(n11525), .A2(n8212), .B1(n14751), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n11526) );
  OAI21_X1 U14010 ( .B1(n11527), .B2(n14751), .A(n11526), .ZN(P1_U3492) );
  OAI222_X1 U14011 ( .A1(n13739), .A2(n11529), .B1(P2_U3088), .B2(n11528), 
        .C1(n13729), .C2(n11530), .ZN(P2_U3307) );
  OAI222_X1 U14012 ( .A1(P1_U3086), .A2(n11532), .B1(n14410), .B2(n11531), 
        .C1(n14413), .C2(n11530), .ZN(P1_U3335) );
  AOI22_X1 U14013 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11897), .B1(n11887), 
        .B2(n11926), .ZN(n11535) );
  AOI21_X1 U14014 ( .B1(n11536), .B2(n11535), .A(n11886), .ZN(n11556) );
  INV_X1 U14015 ( .A(n11537), .ZN(n11538) );
  MUX2_X1 U14016 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12725), .Z(n11894) );
  XNOR2_X1 U14017 ( .A(n11894), .B(n11897), .ZN(n11542) );
  NAND2_X1 U14018 ( .A1(n11543), .A2(n11542), .ZN(n11895) );
  OAI211_X1 U14019 ( .C1(n11543), .C2(n11542), .A(n11895), .B(n15099), .ZN(
        n11555) );
  NAND2_X1 U14020 ( .A1(n11545), .A2(n11544), .ZN(n11547) );
  XNOR2_X1 U14021 ( .A(n11897), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U14022 ( .A1(n11548), .A2(n11549), .ZN(n11889) );
  OAI21_X1 U14023 ( .B1(n11549), .B2(n11548), .A(n11889), .ZN(n11553) );
  NOR2_X1 U14024 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11550), .ZN(n12529) );
  AOI21_X1 U14025 ( .B1(n15093), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12529), 
        .ZN(n11551) );
  OAI21_X1 U14026 ( .B1(n12765), .B2(n11887), .A(n11551), .ZN(n11552) );
  AOI21_X1 U14027 ( .B1(n11553), .B2(n15080), .A(n11552), .ZN(n11554) );
  OAI211_X1 U14028 ( .C1(n11556), .C2(n15103), .A(n11555), .B(n11554), .ZN(
        P3_U3194) );
  OAI222_X1 U14029 ( .A1(n13739), .A2(n11558), .B1(P2_U3088), .B2(n11557), 
        .C1(n13729), .C2(n11642), .ZN(P2_U3306) );
  INV_X1 U14030 ( .A(n11559), .ZN(n11561) );
  OAI222_X1 U14031 ( .A1(n14525), .A2(n11562), .B1(n11389), .B2(n11561), .C1(
        n11560), .C2(P3_U3151), .ZN(P3_U3270) );
  AOI22_X1 U14032 ( .A1(n14745), .A2(n12417), .B1(n12418), .B2(n13909), .ZN(
        n11563) );
  XNOR2_X1 U14033 ( .A(n11563), .B(n12459), .ZN(n11709) );
  AOI22_X1 U14034 ( .A1(n14745), .A2(n12423), .B1(n12422), .B2(n13909), .ZN(
        n11710) );
  XNOR2_X1 U14035 ( .A(n11709), .B(n11710), .ZN(n11572) );
  INV_X1 U14036 ( .A(n11565), .ZN(n11566) );
  NAND2_X1 U14037 ( .A1(n11564), .A2(n11566), .ZN(n11567) );
  INV_X1 U14038 ( .A(n11572), .ZN(n11569) );
  INV_X1 U14039 ( .A(n11713), .ZN(n11570) );
  AOI21_X1 U14040 ( .B1(n11572), .B2(n11571), .A(n11570), .ZN(n11579) );
  OAI21_X1 U14041 ( .B1(n14622), .B2(n11574), .A(n11573), .ZN(n11577) );
  OAI22_X1 U14042 ( .A1(n11575), .A2(n13884), .B1(n13883), .B2(n11860), .ZN(
        n11576) );
  AOI211_X1 U14043 ( .C1(n14745), .C2(n14618), .A(n11577), .B(n11576), .ZN(
        n11578) );
  OAI21_X1 U14044 ( .B1(n11579), .B2(n13889), .A(n11578), .ZN(P1_U3221) );
  XNOR2_X1 U14045 ( .A(n11580), .B(n11589), .ZN(n11583) );
  NAND2_X1 U14046 ( .A1(n13367), .A2(n13315), .ZN(n11582) );
  NAND2_X1 U14047 ( .A1(n13369), .A2(n13316), .ZN(n11581) );
  NAND2_X1 U14048 ( .A1(n11582), .A2(n11581), .ZN(n14577) );
  AOI21_X1 U14049 ( .B1(n11583), .B2(n14992), .A(n14577), .ZN(n14594) );
  INV_X1 U14050 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11584) );
  OAI22_X1 U14051 ( .A1(n13512), .A2(n11584), .B1(n14580), .B2(n15200), .ZN(
        n11588) );
  AOI21_X1 U14052 ( .B1(n14589), .B2(n11585), .A(n13202), .ZN(n11586) );
  NAND2_X1 U14053 ( .A1(n11586), .A2(n11680), .ZN(n14591) );
  NOR2_X1 U14054 ( .A1(n14591), .A2(n13563), .ZN(n11587) );
  AOI211_X1 U14055 ( .C1(n14937), .C2(n14589), .A(n11588), .B(n11587), .ZN(
        n11592) );
  NAND2_X1 U14056 ( .A1(n11590), .A2(n11589), .ZN(n14587) );
  NAND3_X1 U14057 ( .A1(n14588), .A2(n14587), .A3(n15196), .ZN(n11591) );
  OAI211_X1 U14058 ( .C1(n14594), .C2(n10410), .A(n11592), .B(n11591), .ZN(
        P2_U3251) );
  INV_X1 U14059 ( .A(n11593), .ZN(n11612) );
  INV_X1 U14060 ( .A(n11594), .ZN(n11595) );
  NAND2_X1 U14061 ( .A1(n11595), .A2(n12632), .ZN(n11596) );
  NAND2_X1 U14062 ( .A1(n11597), .A2(n11596), .ZN(n11599) );
  XNOR2_X1 U14063 ( .A(n10809), .B(n11603), .ZN(n11727) );
  XNOR2_X1 U14064 ( .A(n11727), .B(n11728), .ZN(n11598) );
  OAI211_X1 U14065 ( .C1(n11599), .C2(n11598), .A(n11731), .B(n12613), .ZN(
        n11605) );
  NAND2_X1 U14066 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15086) );
  INV_X1 U14067 ( .A(n15086), .ZN(n11602) );
  OAI22_X1 U14068 ( .A1(n12609), .A2(n11820), .B1(n11600), .B2(n12618), .ZN(
        n11601) );
  AOI211_X1 U14069 ( .C1(n11603), .C2(n15040), .A(n11602), .B(n11601), .ZN(
        n11604) );
  OAI211_X1 U14070 ( .C1(n11612), .C2(n11826), .A(n11605), .B(n11604), .ZN(
        P3_U3161) );
  XOR2_X1 U14071 ( .A(n11606), .B(n12234), .Z(n15161) );
  AOI21_X1 U14072 ( .B1(n12234), .B2(n11607), .A(n6725), .ZN(n11611) );
  AOI22_X1 U14073 ( .A1(n12985), .A2(n12632), .B1(n15117), .B2(n12631), .ZN(
        n11610) );
  INV_X1 U14074 ( .A(n15161), .ZN(n11608) );
  NAND2_X1 U14075 ( .A1(n11608), .A2(n13024), .ZN(n11609) );
  OAI211_X1 U14076 ( .C1(n11611), .C2(n13019), .A(n11610), .B(n11609), .ZN(
        n15162) );
  NAND2_X1 U14077 ( .A1(n15162), .A2(n6576), .ZN(n11615) );
  OAI22_X1 U14078 ( .A1(n13004), .A2(n15160), .B1(n11612), .B2(n15123), .ZN(
        n11613) );
  AOI21_X1 U14079 ( .B1(n15129), .B2(P3_REG2_REG_8__SCAN_IN), .A(n11613), .ZN(
        n11614) );
  OAI211_X1 U14080 ( .C1(n15161), .C2(n12875), .A(n11615), .B(n11614), .ZN(
        P3_U3225) );
  OAI222_X1 U14081 ( .A1(n13739), .A2(n11617), .B1(P2_U3088), .B2(n6585), .C1(
        n13729), .C2(n11616), .ZN(P2_U3305) );
  XOR2_X1 U14082 ( .A(n11618), .B(n12238), .Z(n15167) );
  AOI22_X1 U14083 ( .A1(n12985), .A2(n11728), .B1(n15117), .B2(n12630), .ZN(
        n11623) );
  OAI21_X1 U14084 ( .B1(n6725), .B2(n11619), .A(n12238), .ZN(n11621) );
  NAND3_X1 U14085 ( .A1(n11621), .A2(n15114), .A3(n11620), .ZN(n11622) );
  OAI211_X1 U14086 ( .C1(n15167), .C2(n12867), .A(n11623), .B(n11622), .ZN(
        n15169) );
  NAND2_X1 U14087 ( .A1(n15169), .A2(n6576), .ZN(n11627) );
  INV_X1 U14088 ( .A(n11738), .ZN(n11624) );
  OAI22_X1 U14089 ( .A1(n13004), .A2(n15165), .B1(n11624), .B2(n15123), .ZN(
        n11625) );
  AOI21_X1 U14090 ( .B1(n15129), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11625), .ZN(
        n11626) );
  OAI211_X1 U14091 ( .C1(n15167), .C2(n12875), .A(n11627), .B(n11626), .ZN(
        P3_U3224) );
  XNOR2_X1 U14092 ( .A(n11628), .B(n11630), .ZN(n11703) );
  INV_X1 U14093 ( .A(n11703), .ZN(n11641) );
  OAI21_X1 U14094 ( .B1(n11631), .B2(n11630), .A(n11629), .ZN(n11698) );
  NAND2_X1 U14095 ( .A1(n13843), .A2(n11654), .ZN(n11632) );
  NAND3_X1 U14096 ( .A1(n11841), .A2(n14254), .A3(n11632), .ZN(n11699) );
  NOR2_X1 U14097 ( .A1(n14225), .A2(n11633), .ZN(n11637) );
  NAND2_X1 U14098 ( .A1(n13905), .A2(n14234), .ZN(n11635) );
  NAND2_X1 U14099 ( .A1(n13903), .A2(n14236), .ZN(n11634) );
  AND2_X1 U14100 ( .A1(n11635), .A2(n11634), .ZN(n11700) );
  OAI22_X1 U14101 ( .A1(n14712), .A2(n11700), .B1(n13839), .B2(n14698), .ZN(
        n11636) );
  AOI211_X1 U14102 ( .C1(n13843), .C2(n14703), .A(n11637), .B(n11636), .ZN(
        n11638) );
  OAI21_X1 U14103 ( .B1(n11699), .B2(n14706), .A(n11638), .ZN(n11639) );
  AOI21_X1 U14104 ( .B1(n11698), .B2(n14229), .A(n11639), .ZN(n11640) );
  OAI21_X1 U14105 ( .B1(n14232), .B2(n11641), .A(n11640), .ZN(P1_U3280) );
  OAI222_X1 U14106 ( .A1(P1_U3086), .A2(n11644), .B1(n14410), .B2(n11643), 
        .C1(n14413), .C2(n11642), .ZN(P1_U3334) );
  OAI21_X1 U14107 ( .B1(n11647), .B2(n11646), .A(n11645), .ZN(n14539) );
  INV_X1 U14108 ( .A(n14539), .ZN(n11660) );
  XNOR2_X1 U14109 ( .A(n11649), .B(n11648), .ZN(n11652) );
  NAND2_X1 U14110 ( .A1(n14539), .A2(n14730), .ZN(n11651) );
  AOI22_X1 U14111 ( .A1(n14234), .A2(n13906), .B1(n13904), .B2(n14236), .ZN(
        n11650) );
  OAI211_X1 U14112 ( .C1(n14329), .C2(n11652), .A(n11651), .B(n11650), .ZN(
        n14537) );
  NAND2_X1 U14113 ( .A1(n14537), .A2(n14225), .ZN(n11659) );
  OAI22_X1 U14114 ( .A1(n14225), .A2(n11653), .B1(n11997), .B2(n14698), .ZN(
        n11657) );
  OAI211_X1 U14115 ( .C1(n14536), .C2(n11655), .A(n14254), .B(n11654), .ZN(
        n14535) );
  NOR2_X1 U14116 ( .A1(n14535), .A2(n14706), .ZN(n11656) );
  AOI211_X1 U14117 ( .C1(n14703), .C2(n12001), .A(n11657), .B(n11656), .ZN(
        n11658) );
  OAI211_X1 U14118 ( .C1(n11660), .C2(n14697), .A(n11659), .B(n11658), .ZN(
        P1_U3281) );
  INV_X1 U14119 ( .A(n11661), .ZN(n11663) );
  OAI222_X1 U14120 ( .A1(n14525), .A2(n15326), .B1(n11389), .B2(n11663), .C1(
        n11662), .C2(P3_U3151), .ZN(P3_U3269) );
  XNOR2_X1 U14121 ( .A(n11664), .B(n12243), .ZN(n11665) );
  NAND2_X1 U14122 ( .A1(n11665), .A2(n15114), .ZN(n11667) );
  AOI22_X1 U14123 ( .A1(n12985), .A2(n12630), .B1(n15117), .B2(n12628), .ZN(
        n11666) );
  NAND2_X1 U14124 ( .A1(n11667), .A2(n11666), .ZN(n14564) );
  INV_X1 U14125 ( .A(n14564), .ZN(n11675) );
  OAI21_X1 U14126 ( .B1(n11668), .B2(n12243), .A(n11669), .ZN(n14566) );
  INV_X1 U14127 ( .A(n13011), .ZN(n12961) );
  NOR2_X1 U14128 ( .A1(n6576), .A2(n11670), .ZN(n11673) );
  INV_X1 U14129 ( .A(n12586), .ZN(n11671) );
  OAI22_X1 U14130 ( .A1(n13004), .A2(n14563), .B1(n11671), .B2(n15123), .ZN(
        n11672) );
  AOI211_X1 U14131 ( .C1(n14566), .C2(n12961), .A(n11673), .B(n11672), .ZN(
        n11674) );
  OAI21_X1 U14132 ( .B1(n15129), .B2(n11675), .A(n11674), .ZN(P3_U3222) );
  XNOR2_X1 U14133 ( .A(n11676), .B(n11679), .ZN(n11677) );
  AOI22_X1 U14134 ( .A1(n13316), .A2(n13368), .B1(n13366), .B2(n13315), .ZN(
        n11881) );
  OAI21_X1 U14135 ( .B1(n11677), .B2(n13530), .A(n11881), .ZN(n14583) );
  INV_X1 U14136 ( .A(n14583), .ZN(n11686) );
  OAI21_X1 U14137 ( .B1(n6713), .B2(n11679), .A(n11678), .ZN(n14585) );
  OAI211_X1 U14138 ( .C1(n7210), .C2(n7211), .A(n14997), .B(n11803), .ZN(
        n14582) );
  INV_X1 U14139 ( .A(n11681), .ZN(n11883) );
  AOI22_X1 U14140 ( .A1(n14957), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11883), 
        .B2(n14948), .ZN(n11683) );
  NAND2_X1 U14141 ( .A1(n11878), .A2(n14937), .ZN(n11682) );
  OAI211_X1 U14142 ( .C1(n14582), .C2(n13563), .A(n11683), .B(n11682), .ZN(
        n11684) );
  AOI21_X1 U14143 ( .B1(n14585), .B2(n15196), .A(n11684), .ZN(n11685) );
  OAI21_X1 U14144 ( .B1(n14957), .B2(n11686), .A(n11685), .ZN(P2_U3250) );
  INV_X1 U14145 ( .A(n11687), .ZN(n11688) );
  OAI222_X1 U14146 ( .A1(n14525), .A2(n15275), .B1(n11389), .B2(n11688), .C1(
        P3_U3151), .C2(n12733), .ZN(P3_U3268) );
  NAND2_X1 U14147 ( .A1(n11693), .A2(n14405), .ZN(n11690) );
  OAI211_X1 U14148 ( .C1(n11691), .C2(n14410), .A(n11690), .B(n11689), .ZN(
        P1_U3332) );
  NAND2_X1 U14149 ( .A1(n11693), .A2(n11692), .ZN(n11695) );
  OAI211_X1 U14150 ( .C1(n11697), .C2(n11696), .A(n11695), .B(n11694), .ZN(
        P2_U3304) );
  INV_X1 U14151 ( .A(n11698), .ZN(n11701) );
  OAI211_X1 U14152 ( .C1(n11701), .C2(n14749), .A(n11700), .B(n11699), .ZN(
        n11702) );
  AOI21_X1 U14153 ( .B1(n11703), .B2(n14741), .A(n11702), .ZN(n11708) );
  INV_X1 U14154 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11704) );
  NOR2_X1 U14155 ( .A1(n14752), .A2(n11704), .ZN(n11705) );
  AOI21_X1 U14156 ( .B1(n13843), .B2(n8212), .A(n11705), .ZN(n11706) );
  OAI21_X1 U14157 ( .B1(n11708), .B2(n14751), .A(n11706), .ZN(P1_U3498) );
  AOI22_X1 U14158 ( .A1(n13843), .A2(n8207), .B1(n14757), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n11707) );
  OAI21_X1 U14159 ( .B1(n11708), .B2(n14757), .A(n11707), .ZN(P1_U3541) );
  INV_X1 U14160 ( .A(n11709), .ZN(n11712) );
  INV_X1 U14161 ( .A(n11710), .ZN(n11711) );
  NAND2_X1 U14162 ( .A1(n11716), .A2(n12423), .ZN(n11715) );
  NAND2_X1 U14163 ( .A1(n12422), .A2(n13908), .ZN(n11714) );
  NAND2_X1 U14164 ( .A1(n11715), .A2(n11714), .ZN(n11849) );
  XNOR2_X2 U14165 ( .A(n11848), .B(n11849), .ZN(n11719) );
  AOI22_X1 U14166 ( .A1(n11716), .A2(n12417), .B1(n12418), .B2(n13908), .ZN(
        n11717) );
  XOR2_X1 U14167 ( .A(n12459), .B(n11717), .Z(n11718) );
  OAI211_X1 U14168 ( .C1(n11719), .C2(n11718), .A(n11852), .B(n14613), .ZN(
        n11725) );
  NOR2_X1 U14169 ( .A1(n14622), .A2(n11720), .ZN(n11723) );
  OAI22_X1 U14170 ( .A1(n11721), .A2(n13884), .B1(n13883), .B2(n12010), .ZN(
        n11722) );
  AOI211_X1 U14171 ( .C1(P1_REG3_REG_9__SCAN_IN), .C2(P1_U3086), .A(n11723), 
        .B(n11722), .ZN(n11724) );
  OAI211_X1 U14172 ( .C1(n11726), .C2(n13868), .A(n11725), .B(n11724), .ZN(
        P1_U3231) );
  XNOR2_X1 U14173 ( .A(n10809), .B(n15165), .ZN(n11815) );
  XNOR2_X1 U14174 ( .A(n11815), .B(n12631), .ZN(n11734) );
  INV_X1 U14175 ( .A(n11727), .ZN(n11729) );
  NAND2_X1 U14176 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  INV_X1 U14177 ( .A(n11818), .ZN(n11732) );
  AOI21_X1 U14178 ( .B1(n11734), .B2(n11733), .A(n11732), .ZN(n11741) );
  OAI22_X1 U14179 ( .A1(n12609), .A2(n12588), .B1(n11735), .B2(n12618), .ZN(
        n11736) );
  AOI211_X1 U14180 ( .C1(n12119), .C2(n15040), .A(n11737), .B(n11736), .ZN(
        n11740) );
  NAND2_X1 U14181 ( .A1(n12620), .A2(n11738), .ZN(n11739) );
  OAI211_X1 U14182 ( .C1(n11741), .C2(n15043), .A(n11740), .B(n11739), .ZN(
        P3_U3171) );
  INV_X1 U14183 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n15271) );
  NAND2_X1 U14184 ( .A1(n11761), .A2(n11742), .ZN(n11743) );
  NAND2_X1 U14185 ( .A1(n11744), .A2(n11743), .ZN(n14844) );
  MUX2_X1 U14186 ( .A(n11397), .B(P2_REG2_REG_13__SCAN_IN), .S(n11765), .Z(
        n14843) );
  NAND2_X1 U14187 ( .A1(n11765), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11745) );
  NAND2_X1 U14188 ( .A1(n14845), .A2(n11745), .ZN(n11746) );
  XNOR2_X1 U14189 ( .A(n11746), .B(n14865), .ZN(n14859) );
  NAND2_X1 U14190 ( .A1(n14859), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14858) );
  NAND2_X1 U14191 ( .A1(n11746), .A2(n11767), .ZN(n11747) );
  NAND2_X1 U14192 ( .A1(n14858), .A2(n11747), .ZN(n11748) );
  XNOR2_X1 U14193 ( .A(n11748), .B(n14874), .ZN(n14870) );
  AOI21_X1 U14194 ( .B1(n11770), .B2(n11748), .A(n14872), .ZN(n14890) );
  INV_X1 U14195 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n15274) );
  NOR2_X1 U14196 ( .A1(n14893), .A2(n15274), .ZN(n11749) );
  AOI21_X1 U14197 ( .B1(n14893), .B2(n15274), .A(n11749), .ZN(n14889) );
  NOR2_X1 U14198 ( .A1(n14890), .A2(n14889), .ZN(n14888) );
  AOI21_X1 U14199 ( .B1(n14893), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14888), 
        .ZN(n14898) );
  INV_X1 U14200 ( .A(n14898), .ZN(n11754) );
  INV_X1 U14201 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11750) );
  OR2_X1 U14202 ( .A1(n11773), .A2(n11750), .ZN(n11752) );
  NAND2_X1 U14203 ( .A1(n11773), .A2(n11750), .ZN(n11751) );
  AND2_X1 U14204 ( .A1(n11752), .A2(n11751), .ZN(n14897) );
  INV_X1 U14205 ( .A(n14897), .ZN(n11753) );
  NAND2_X1 U14206 ( .A1(n11754), .A2(n11753), .ZN(n14900) );
  NAND2_X1 U14207 ( .A1(n11773), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11755) );
  XNOR2_X1 U14208 ( .A(n11757), .B(n11756), .ZN(n14914) );
  NAND2_X1 U14209 ( .A1(n14914), .A2(n8265), .ZN(n14913) );
  NAND2_X1 U14210 ( .A1(n11757), .A2(n14925), .ZN(n11758) );
  NAND2_X1 U14211 ( .A1(n14913), .A2(n11758), .ZN(n11759) );
  XNOR2_X1 U14212 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n11759), .ZN(n11781) );
  INV_X1 U14213 ( .A(n11781), .ZN(n11779) );
  XNOR2_X1 U14214 ( .A(n11773), .B(n15357), .ZN(n14901) );
  NAND2_X1 U14215 ( .A1(n14893), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11772) );
  NAND2_X1 U14216 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  NAND2_X1 U14217 ( .A1(n11763), .A2(n11762), .ZN(n14848) );
  INV_X1 U14218 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11764) );
  MUX2_X1 U14219 ( .A(n11764), .B(P2_REG1_REG_13__SCAN_IN), .S(n11765), .Z(
        n14847) );
  NAND2_X1 U14220 ( .A1(n11765), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U14221 ( .A1(n14849), .A2(n11766), .ZN(n14862) );
  INV_X1 U14222 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14596) );
  MUX2_X1 U14223 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14596), .S(n11767), .Z(
        n14861) );
  NAND2_X1 U14224 ( .A1(n14862), .A2(n14861), .ZN(n14860) );
  NAND2_X1 U14225 ( .A1(n11767), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U14226 ( .A1(n14860), .A2(n11768), .ZN(n11769) );
  XNOR2_X1 U14227 ( .A(n11769), .B(n14874), .ZN(n14873) );
  AOI21_X1 U14228 ( .B1(n11770), .B2(n11769), .A(n14875), .ZN(n14886) );
  XNOR2_X1 U14229 ( .A(n14893), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14885) );
  NOR2_X1 U14230 ( .A1(n14886), .A2(n14885), .ZN(n14884) );
  INV_X1 U14231 ( .A(n14884), .ZN(n11771) );
  NAND2_X1 U14232 ( .A1(n11772), .A2(n11771), .ZN(n14902) );
  NAND2_X1 U14233 ( .A1(n14901), .A2(n14902), .ZN(n14906) );
  NAND2_X1 U14234 ( .A1(n11773), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11774) );
  AND2_X1 U14235 ( .A1(n14906), .A2(n11774), .ZN(n11775) );
  XNOR2_X1 U14236 ( .A(n11775), .B(n14925), .ZN(n14918) );
  NOR2_X1 U14237 ( .A1(n14917), .A2(n14918), .ZN(n14919) );
  NOR2_X1 U14238 ( .A1(n11775), .A2(n14925), .ZN(n11776) );
  NOR2_X1 U14239 ( .A1(n14919), .A2(n11776), .ZN(n11777) );
  XNOR2_X1 U14240 ( .A(n11777), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n11780) );
  OAI21_X1 U14241 ( .B1(n11780), .B2(n14883), .A(n14926), .ZN(n11778) );
  AOI21_X1 U14242 ( .B1(n11779), .B2(n14915), .A(n11778), .ZN(n11783) );
  AOI22_X1 U14243 ( .A1(n11781), .A2(n14915), .B1(n14922), .B2(n11780), .ZN(
        n11782) );
  MUX2_X1 U14244 ( .A(n11783), .B(n11782), .S(n13581), .Z(n11784) );
  NAND2_X1 U14245 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13248)
         );
  OAI211_X1 U14246 ( .C1(n15271), .C2(n14930), .A(n11784), .B(n13248), .ZN(
        P2_U3233) );
  XNOR2_X1 U14247 ( .A(n11785), .B(n11791), .ZN(n14355) );
  AOI211_X1 U14248 ( .C1(n14351), .C2(n11842), .A(n14317), .B(n11971), .ZN(
        n14349) );
  INV_X1 U14249 ( .A(n14351), .ZN(n12337) );
  NAND2_X1 U14250 ( .A1(n13901), .A2(n14236), .ZN(n11786) );
  OAI21_X1 U14251 ( .B1(n13885), .B2(n14140), .A(n11786), .ZN(n14350) );
  INV_X1 U14252 ( .A(n13881), .ZN(n11787) );
  AOI22_X1 U14253 ( .A1(n14225), .A2(n14350), .B1(n11787), .B2(n14241), .ZN(
        n11789) );
  NAND2_X1 U14254 ( .A1(n14712), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11788) );
  OAI211_X1 U14255 ( .C1(n12337), .C2(n14244), .A(n11789), .B(n11788), .ZN(
        n11790) );
  AOI21_X1 U14256 ( .B1(n14349), .B2(n14251), .A(n11790), .ZN(n11794) );
  XNOR2_X1 U14257 ( .A(n11792), .B(n11791), .ZN(n14352) );
  NAND2_X1 U14258 ( .A1(n14352), .A2(n14121), .ZN(n11793) );
  OAI211_X1 U14259 ( .C1(n14355), .C2(n14248), .A(n11794), .B(n11793), .ZN(
        P1_U3278) );
  OAI222_X1 U14260 ( .A1(P2_U3088), .A2(n11796), .B1(n13741), .B2(n11827), 
        .C1(n11795), .C2(n13739), .ZN(P2_U3303) );
  INV_X1 U14261 ( .A(n11797), .ZN(n11800) );
  INV_X1 U14262 ( .A(n11810), .ZN(n11799) );
  OAI21_X1 U14263 ( .B1(n11800), .B2(n11799), .A(n11798), .ZN(n11802) );
  OAI22_X1 U14264 ( .A1(n13328), .A2(n13342), .B1(n11801), .B2(n13340), .ZN(
        n11945) );
  AOI21_X1 U14265 ( .B1(n11802), .B2(n14992), .A(n11945), .ZN(n13689) );
  NAND2_X1 U14266 ( .A1(n13687), .A2(n11803), .ZN(n11804) );
  NAND2_X1 U14267 ( .A1(n11804), .A2(n14997), .ZN(n11805) );
  NOR2_X1 U14268 ( .A1(n11957), .A2(n11805), .ZN(n13686) );
  NAND2_X1 U14269 ( .A1(n13687), .A2(n14937), .ZN(n11808) );
  INV_X1 U14270 ( .A(n11947), .ZN(n11806) );
  AOI22_X1 U14271 ( .A1(n14957), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n11806), 
        .B2(n14948), .ZN(n11807) );
  NAND2_X1 U14272 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  AOI21_X1 U14273 ( .B1(n13686), .B2(n15195), .A(n11809), .ZN(n11813) );
  OR2_X1 U14274 ( .A1(n11811), .A2(n11810), .ZN(n13685) );
  NAND3_X1 U14275 ( .A1(n13685), .A2(n15196), .A3(n13684), .ZN(n11812) );
  OAI211_X1 U14276 ( .C1(n13689), .C2(n10410), .A(n11813), .B(n11812), .ZN(
        P2_U3249) );
  INV_X1 U14277 ( .A(n11814), .ZN(n11918) );
  INV_X1 U14278 ( .A(n11815), .ZN(n11816) );
  NAND2_X1 U14279 ( .A1(n11816), .A2(n11820), .ZN(n11817) );
  XNOR2_X1 U14280 ( .A(n10809), .B(n15171), .ZN(n12279) );
  XNOR2_X1 U14281 ( .A(n12279), .B(n12588), .ZN(n11819) );
  OAI211_X1 U14282 ( .C1(n6732), .C2(n11819), .A(n12281), .B(n12613), .ZN(
        n11825) );
  NAND2_X1 U14283 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15106)
         );
  INV_X1 U14284 ( .A(n15106), .ZN(n11822) );
  OAI22_X1 U14285 ( .A1(n12609), .A2(n12583), .B1(n11820), .B2(n12618), .ZN(
        n11821) );
  AOI211_X1 U14286 ( .C1(n11823), .C2(n15040), .A(n11822), .B(n11821), .ZN(
        n11824) );
  OAI211_X1 U14287 ( .C1(n11918), .C2(n11826), .A(n11825), .B(n11824), .ZN(
        P3_U3157) );
  OAI222_X1 U14288 ( .A1(P1_U3086), .A2(n11829), .B1(n14410), .B2(n11828), 
        .C1(n14413), .C2(n11827), .ZN(P1_U3331) );
  XNOR2_X1 U14289 ( .A(n11831), .B(n11830), .ZN(n11832) );
  NAND2_X1 U14290 ( .A1(n11832), .A2(n14741), .ZN(n11836) );
  OR2_X1 U14291 ( .A1(n13799), .A2(n14142), .ZN(n11834) );
  NAND2_X1 U14292 ( .A1(n13904), .A2(n14234), .ZN(n11833) );
  NAND2_X1 U14293 ( .A1(n11834), .A2(n11833), .ZN(n14616) );
  INV_X1 U14294 ( .A(n14616), .ZN(n11835) );
  NAND2_X1 U14295 ( .A1(n11836), .A2(n11835), .ZN(n14625) );
  INV_X1 U14296 ( .A(n14625), .ZN(n11847) );
  INV_X1 U14297 ( .A(n11837), .ZN(n11838) );
  AOI21_X1 U14298 ( .B1(n11840), .B2(n11839), .A(n11838), .ZN(n14627) );
  OAI211_X1 U14299 ( .C1(n7071), .C2(n7072), .A(n14254), .B(n11842), .ZN(
        n14623) );
  OAI22_X1 U14300 ( .A1(n14225), .A2(n10487), .B1(n14621), .B2(n14698), .ZN(
        n11843) );
  AOI21_X1 U14301 ( .B1(n14617), .B2(n14703), .A(n11843), .ZN(n11844) );
  OAI21_X1 U14302 ( .B1(n14623), .B2(n14070), .A(n11844), .ZN(n11845) );
  AOI21_X1 U14303 ( .B1(n14627), .B2(n14229), .A(n11845), .ZN(n11846) );
  OAI21_X1 U14304 ( .B1(n14712), .B2(n11847), .A(n11846), .ZN(P1_U3279) );
  NAND2_X1 U14305 ( .A1(n11863), .A2(n12417), .ZN(n11854) );
  NAND2_X1 U14306 ( .A1(n12423), .A2(n13907), .ZN(n11853) );
  NAND2_X1 U14307 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  XNOR2_X1 U14308 ( .A(n11855), .B(n8097), .ZN(n11981) );
  NOR2_X1 U14309 ( .A1(n12455), .A2(n12010), .ZN(n11856) );
  AOI21_X1 U14310 ( .B1(n11863), .B2(n12418), .A(n11856), .ZN(n11980) );
  INV_X1 U14311 ( .A(n11980), .ZN(n11982) );
  XNOR2_X1 U14312 ( .A(n11981), .B(n11982), .ZN(n11857) );
  XNOR2_X1 U14313 ( .A(n11985), .B(n11857), .ZN(n11865) );
  OAI21_X1 U14314 ( .B1(n14622), .B2(n11859), .A(n11858), .ZN(n11862) );
  OAI22_X1 U14315 ( .A1(n11860), .A2(n13884), .B1(n13883), .B2(n11998), .ZN(
        n11861) );
  AOI211_X1 U14316 ( .C1(n11863), .C2(n14618), .A(n11862), .B(n11861), .ZN(
        n11864) );
  OAI21_X1 U14317 ( .B1(n11865), .B2(n13889), .A(n11864), .ZN(P1_U3217) );
  NAND2_X1 U14318 ( .A1(n13367), .A2(n13574), .ZN(n11941) );
  NAND2_X1 U14319 ( .A1(n14574), .A2(n11941), .ZN(n11880) );
  NAND2_X1 U14320 ( .A1(n13334), .A2(n13367), .ZN(n11879) );
  INV_X1 U14321 ( .A(n11868), .ZN(n11871) );
  INV_X1 U14322 ( .A(n11869), .ZN(n11870) );
  XNOR2_X1 U14323 ( .A(n14589), .B(n13255), .ZN(n11872) );
  NAND2_X1 U14324 ( .A1(n13368), .A2(n13574), .ZN(n11873) );
  NAND2_X1 U14325 ( .A1(n11872), .A2(n11873), .ZN(n11877) );
  INV_X1 U14326 ( .A(n11872), .ZN(n11875) );
  INV_X1 U14327 ( .A(n11873), .ZN(n11874) );
  NAND2_X1 U14328 ( .A1(n11875), .A2(n11874), .ZN(n11876) );
  AND2_X1 U14329 ( .A1(n11877), .A2(n11876), .ZN(n14573) );
  NAND2_X1 U14330 ( .A1(n14572), .A2(n14573), .ZN(n14571) );
  XOR2_X1 U14331 ( .A(n13217), .B(n11878), .Z(n11940) );
  MUX2_X1 U14332 ( .A(n11880), .B(n11879), .S(n11942), .Z(n11885) );
  OAI22_X1 U14333 ( .A1(n13318), .A2(n11881), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8481), .ZN(n11882) );
  AOI21_X1 U14334 ( .B1(n11883), .B2(n13322), .A(n11882), .ZN(n11884) );
  OAI211_X1 U14335 ( .C1(n7210), .C2(n13319), .A(n11885), .B(n11884), .ZN(
        P2_U3213) );
  INV_X1 U14336 ( .A(n12655), .ZN(n12647) );
  AOI21_X1 U14337 ( .B1(n13007), .B2(n11888), .A(n12639), .ZN(n11904) );
  INV_X1 U14338 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14492) );
  INV_X1 U14339 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11914) );
  XNOR2_X1 U14340 ( .A(n12647), .B(n12654), .ZN(n11890) );
  NAND2_X1 U14341 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11890), .ZN(n12656) );
  OAI21_X1 U14342 ( .B1(n11890), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12656), 
        .ZN(n11891) );
  NAND2_X1 U14343 ( .A1(n15080), .A2(n11891), .ZN(n11893) );
  AND2_X1 U14344 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12571) );
  INV_X1 U14345 ( .A(n12571), .ZN(n11892) );
  OAI211_X1 U14346 ( .C1(n14492), .C2(n15088), .A(n11893), .B(n11892), .ZN(
        n11902) );
  MUX2_X1 U14347 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12725), .Z(n12644) );
  XNOR2_X1 U14348 ( .A(n12644), .B(n12655), .ZN(n11899) );
  INV_X1 U14349 ( .A(n11894), .ZN(n11896) );
  OAI21_X1 U14350 ( .B1(n11897), .B2(n11896), .A(n11895), .ZN(n11898) );
  NOR2_X1 U14351 ( .A1(n11898), .A2(n11899), .ZN(n12645) );
  AOI21_X1 U14352 ( .B1(n11899), .B2(n11898), .A(n12645), .ZN(n11900) );
  NOR2_X1 U14353 ( .A1(n11900), .A2(n15071), .ZN(n11901) );
  AOI211_X1 U14354 ( .C1(n15097), .C2(n12647), .A(n11902), .B(n11901), .ZN(
        n11903) );
  OAI21_X1 U14355 ( .B1(n11904), .B2(n15103), .A(n11903), .ZN(P3_U3195) );
  OAI211_X1 U14356 ( .C1(n11907), .C2(n11906), .A(n11905), .B(n15114), .ZN(
        n11909) );
  AOI22_X1 U14357 ( .A1(n12985), .A2(n12629), .B1(n15117), .B2(n12984), .ZN(
        n11908) );
  AND2_X1 U14358 ( .A1(n11909), .A2(n11908), .ZN(n11927) );
  MUX2_X1 U14359 ( .A(n11927), .B(n11910), .S(n15176), .Z(n11913) );
  XNOR2_X1 U14360 ( .A(n11911), .B(n12244), .ZN(n11925) );
  INV_X1 U14361 ( .A(n13177), .ZN(n13161) );
  AOI22_X1 U14362 ( .A1(n11925), .A2(n13161), .B1(n13148), .B2(n12531), .ZN(
        n11912) );
  NAND2_X1 U14363 ( .A1(n11913), .A2(n11912), .ZN(P3_U3426) );
  MUX2_X1 U14364 ( .A(n11914), .B(n11927), .S(n15192), .Z(n11916) );
  INV_X1 U14365 ( .A(n13095), .ZN(n13083) );
  AOI22_X1 U14366 ( .A1(n11925), .A2(n13083), .B1(n13068), .B2(n12531), .ZN(
        n11915) );
  NAND2_X1 U14367 ( .A1(n11916), .A2(n11915), .ZN(P3_U3471) );
  XOR2_X1 U14368 ( .A(n11917), .B(n12239), .Z(n15175) );
  INV_X1 U14369 ( .A(n15175), .ZN(n11924) );
  OAI22_X1 U14370 ( .A1(n13004), .A2(n15171), .B1(n11918), .B2(n15123), .ZN(
        n11922) );
  XOR2_X1 U14371 ( .A(n11919), .B(n12239), .Z(n11920) );
  AOI222_X1 U14372 ( .A1(n15114), .A2(n11920), .B1(n12629), .B2(n15117), .C1(
        n12631), .C2(n12985), .ZN(n15170) );
  NOR2_X1 U14373 ( .A1(n15170), .A2(n15129), .ZN(n11921) );
  AOI211_X1 U14374 ( .C1(n15129), .C2(P3_REG2_REG_10__SCAN_IN), .A(n11922), 
        .B(n11921), .ZN(n11923) );
  OAI21_X1 U14375 ( .B1(n13011), .B2(n11924), .A(n11923), .ZN(P3_U3223) );
  INV_X1 U14376 ( .A(n11925), .ZN(n11930) );
  MUX2_X1 U14377 ( .A(n11927), .B(n11926), .S(n15129), .Z(n11929) );
  AOI22_X1 U14378 ( .A1(n12991), .A2(n12531), .B1(n12990), .B2(n12530), .ZN(
        n11928) );
  OAI211_X1 U14379 ( .C1(n11930), .C2(n13011), .A(n11929), .B(n11928), .ZN(
        P3_U3221) );
  INV_X1 U14380 ( .A(n11931), .ZN(n11935) );
  OAI222_X1 U14381 ( .A1(n14410), .A2(n11933), .B1(n14413), .B2(n11935), .C1(
        P1_U3086), .C2(n11932), .ZN(P1_U3330) );
  OAI222_X1 U14382 ( .A1(n13739), .A2(n11936), .B1(n13741), .B2(n11935), .C1(
        P2_U3088), .C2(n11934), .ZN(P2_U3302) );
  XNOR2_X1 U14383 ( .A(n13687), .B(n13255), .ZN(n11938) );
  NAND2_X1 U14384 ( .A1(n13366), .A2(n13574), .ZN(n11937) );
  NAND2_X1 U14385 ( .A1(n11938), .A2(n11937), .ZN(n12031) );
  OAI21_X1 U14386 ( .B1(n11938), .B2(n11937), .A(n12031), .ZN(n11944) );
  AOI21_X1 U14387 ( .B1(n11944), .B2(n11943), .A(n6721), .ZN(n11950) );
  NAND2_X1 U14388 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14895)
         );
  NAND2_X1 U14389 ( .A1(n14576), .A2(n11945), .ZN(n11946) );
  OAI211_X1 U14390 ( .C1(n14581), .C2(n11947), .A(n14895), .B(n11946), .ZN(
        n11948) );
  AOI21_X1 U14391 ( .B1(n13687), .B2(n14578), .A(n11948), .ZN(n11949) );
  OAI21_X1 U14392 ( .B1(n11950), .B2(n13350), .A(n11949), .ZN(P2_U3198) );
  XOR2_X1 U14393 ( .A(n11951), .B(n11955), .Z(n11953) );
  OAI22_X1 U14394 ( .A1(n13247), .A2(n13342), .B1(n11952), .B2(n13340), .ZN(
        n12037) );
  AOI21_X1 U14395 ( .B1(n11953), .B2(n14992), .A(n12037), .ZN(n13681) );
  OAI21_X1 U14396 ( .B1(n11956), .B2(n11955), .A(n11954), .ZN(n13683) );
  INV_X1 U14397 ( .A(n13683), .ZN(n11964) );
  OR2_X1 U14398 ( .A1(n11962), .A2(n11957), .ZN(n11958) );
  AND3_X1 U14399 ( .A1(n13595), .A2(n11958), .A3(n14997), .ZN(n13678) );
  NAND2_X1 U14400 ( .A1(n13678), .A2(n15195), .ZN(n11961) );
  INV_X1 U14401 ( .A(n12039), .ZN(n11959) );
  AOI22_X1 U14402 ( .A1(n14957), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n11959), 
        .B2(n14948), .ZN(n11960) );
  OAI211_X1 U14403 ( .C1(n11962), .C2(n14951), .A(n11961), .B(n11960), .ZN(
        n11963) );
  AOI21_X1 U14404 ( .B1(n11964), .B2(n15196), .A(n11963), .ZN(n11965) );
  OAI21_X1 U14405 ( .B1(n14957), .B2(n13681), .A(n11965), .ZN(P2_U3248) );
  XNOR2_X1 U14406 ( .A(n11966), .B(n11969), .ZN(n11967) );
  OAI222_X1 U14407 ( .A1(n14142), .A2(n13862), .B1(n14140), .B2(n13799), .C1(
        n11967), .C2(n14329), .ZN(n14345) );
  INV_X1 U14408 ( .A(n14345), .ZN(n11979) );
  OAI21_X1 U14409 ( .B1(n11970), .B2(n11969), .A(n11968), .ZN(n14347) );
  NOR2_X1 U14410 ( .A1(n14344), .A2(n11971), .ZN(n11972) );
  OR3_X1 U14411 ( .A1(n12023), .A2(n11972), .A3(n14317), .ZN(n14343) );
  NAND2_X1 U14412 ( .A1(n14712), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11973) );
  OAI21_X1 U14413 ( .B1(n14698), .B2(n13797), .A(n11973), .ZN(n11974) );
  AOI21_X1 U14414 ( .B1(n11975), .B2(n14703), .A(n11974), .ZN(n11976) );
  OAI21_X1 U14415 ( .B1(n14343), .B2(n14706), .A(n11976), .ZN(n11977) );
  AOI21_X1 U14416 ( .B1(n14347), .B2(n14229), .A(n11977), .ZN(n11978) );
  OAI21_X1 U14417 ( .B1(n11979), .B2(n14712), .A(n11978), .ZN(P1_U3277) );
  NAND2_X1 U14418 ( .A1(n11981), .A2(n11980), .ZN(n11984) );
  INV_X1 U14419 ( .A(n11981), .ZN(n11983) );
  OAI22_X1 U14420 ( .A1(n12016), .A2(n12456), .B1(n11998), .B2(n12455), .ZN(
        n11991) );
  OAI22_X1 U14421 ( .A1(n12016), .A2(n12458), .B1(n11998), .B2(n12456), .ZN(
        n11986) );
  XNOR2_X1 U14422 ( .A(n11986), .B(n12459), .ZN(n11990) );
  XOR2_X1 U14423 ( .A(n11991), .B(n11990), .Z(n12007) );
  OAI22_X1 U14424 ( .A1(n14536), .A2(n12458), .B1(n13840), .B2(n12456), .ZN(
        n11987) );
  XNOR2_X1 U14425 ( .A(n11987), .B(n8097), .ZN(n12327) );
  OR2_X1 U14426 ( .A1(n14536), .A2(n12456), .ZN(n11989) );
  NAND2_X1 U14427 ( .A1(n13905), .A2(n12422), .ZN(n11988) );
  NAND2_X1 U14428 ( .A1(n11989), .A2(n11988), .ZN(n12325) );
  XNOR2_X1 U14429 ( .A(n12327), .B(n12325), .ZN(n11994) );
  INV_X1 U14430 ( .A(n11990), .ZN(n11993) );
  INV_X1 U14431 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14432 ( .A1(n11993), .A2(n11992), .ZN(n11995) );
  NAND2_X1 U14433 ( .A1(n12326), .A2(n14613), .ZN(n12004) );
  AOI21_X1 U14434 ( .B1(n12005), .B2(n11995), .A(n11994), .ZN(n12003) );
  OAI22_X1 U14435 ( .A1(n14622), .A2(n11997), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11996), .ZN(n12000) );
  OAI22_X1 U14436 ( .A1(n11998), .A2(n13884), .B1(n13883), .B2(n12328), .ZN(
        n11999) );
  AOI211_X1 U14437 ( .C1(n12001), .C2(n14618), .A(n12000), .B(n11999), .ZN(
        n12002) );
  OAI21_X1 U14438 ( .B1(n12004), .B2(n12003), .A(n12002), .ZN(P1_U3224) );
  OAI21_X1 U14439 ( .B1(n12007), .B2(n12006), .A(n12005), .ZN(n12008) );
  NAND2_X1 U14440 ( .A1(n12008), .A2(n14613), .ZN(n12015) );
  INV_X1 U14441 ( .A(n12009), .ZN(n12012) );
  OAI22_X1 U14442 ( .A1(n12010), .A2(n13884), .B1(n13883), .B2(n13840), .ZN(
        n12011) );
  AOI211_X1 U14443 ( .C1(n12013), .C2(n13865), .A(n12012), .B(n12011), .ZN(
        n12014) );
  OAI211_X1 U14444 ( .C1(n12016), .C2(n13868), .A(n12015), .B(n12014), .ZN(
        P1_U3236) );
  XNOR2_X1 U14445 ( .A(n12018), .B(n12017), .ZN(n14342) );
  INV_X1 U14446 ( .A(n12019), .ZN(n12020) );
  AOI21_X1 U14447 ( .B1(n12022), .B2(n12021), .A(n12020), .ZN(n14340) );
  OAI211_X1 U14448 ( .C1(n14338), .C2(n12023), .A(n14254), .B(n14240), .ZN(
        n14337) );
  AND2_X1 U14449 ( .A1(n13901), .A2(n14234), .ZN(n12024) );
  AOI21_X1 U14450 ( .B1(n13900), .B2(n14236), .A(n12024), .ZN(n14336) );
  INV_X1 U14451 ( .A(n12025), .ZN(n13811) );
  OAI22_X1 U14452 ( .A1(n14712), .A2(n14336), .B1(n13811), .B2(n14698), .ZN(
        n12027) );
  NOR2_X1 U14453 ( .A1(n14338), .A2(n14244), .ZN(n12026) );
  AOI211_X1 U14454 ( .C1(n14712), .C2(P1_REG2_REG_17__SCAN_IN), .A(n12027), 
        .B(n12026), .ZN(n12028) );
  OAI21_X1 U14455 ( .B1(n14706), .B2(n14337), .A(n12028), .ZN(n12029) );
  AOI21_X1 U14456 ( .B1(n14340), .B2(n14121), .A(n12029), .ZN(n12030) );
  OAI21_X1 U14457 ( .B1(n14248), .B2(n14342), .A(n12030), .ZN(P1_U3276) );
  INV_X1 U14458 ( .A(n12031), .ZN(n12032) );
  XNOR2_X1 U14459 ( .A(n13679), .B(n13255), .ZN(n12034) );
  NAND2_X1 U14460 ( .A1(n13365), .A2(n13202), .ZN(n12033) );
  NAND2_X1 U14461 ( .A1(n12034), .A2(n12033), .ZN(n13189) );
  OAI21_X1 U14462 ( .B1(n12034), .B2(n12033), .A(n13189), .ZN(n12035) );
  AOI21_X1 U14463 ( .B1(n12036), .B2(n12035), .A(n13191), .ZN(n12042) );
  NAND2_X1 U14464 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14911)
         );
  NAND2_X1 U14465 ( .A1(n14576), .A2(n12037), .ZN(n12038) );
  OAI211_X1 U14466 ( .C1(n14581), .C2(n12039), .A(n14911), .B(n12038), .ZN(
        n12040) );
  AOI21_X1 U14467 ( .B1(n13679), .B2(n14578), .A(n12040), .ZN(n12041) );
  OAI21_X1 U14468 ( .B1(n12042), .B2(n13350), .A(n12041), .ZN(P2_U3200) );
  NAND2_X1 U14469 ( .A1(n13732), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U14470 ( .A1(n12044), .A2(n12043), .ZN(n12046) );
  NAND2_X1 U14471 ( .A1(n14398), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12045) );
  NAND2_X1 U14472 ( .A1(n12046), .A2(n12045), .ZN(n12052) );
  AOI22_X1 U14473 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12278), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n12444), .ZN(n12047) );
  INV_X1 U14474 ( .A(n12047), .ZN(n12048) );
  XNOR2_X1 U14475 ( .A(n12052), .B(n12048), .ZN(n12446) );
  NAND2_X1 U14476 ( .A1(n12446), .A2(n12055), .ZN(n12050) );
  OR2_X1 U14477 ( .A1(n12056), .A2(n12449), .ZN(n12049) );
  NAND2_X1 U14478 ( .A1(n12050), .A2(n12049), .ZN(n12069) );
  NOR2_X1 U14479 ( .A1(n12069), .A2(n12067), .ZN(n12223) );
  NOR2_X1 U14480 ( .A1(n12278), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12051) );
  OAI22_X1 U14481 ( .A1(n12052), .A2(n12051), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12444), .ZN(n12054) );
  XNOR2_X1 U14482 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12053) );
  XNOR2_X1 U14483 ( .A(n12054), .B(n12053), .ZN(n13180) );
  NAND2_X1 U14484 ( .A1(n13180), .A2(n12055), .ZN(n12058) );
  INV_X1 U14485 ( .A(SI_31_), .ZN(n13184) );
  OR2_X1 U14486 ( .A1(n12056), .A2(n13184), .ZN(n12057) );
  NAND2_X1 U14487 ( .A1(n6574), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12065) );
  INV_X1 U14488 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12060) );
  OR2_X1 U14489 ( .A1(n12061), .A2(n12060), .ZN(n12064) );
  INV_X1 U14490 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n15299) );
  OR2_X1 U14491 ( .A1(n12062), .A2(n15299), .ZN(n12063) );
  NAND2_X1 U14492 ( .A1(n12069), .A2(n12067), .ZN(n12068) );
  INV_X1 U14493 ( .A(n12069), .ZN(n14561) );
  INV_X1 U14494 ( .A(n12780), .ZN(n12624) );
  OAI21_X1 U14495 ( .B1(n14561), .B2(n12624), .A(n12254), .ZN(n12070) );
  XNOR2_X1 U14496 ( .A(n12072), .B(n12764), .ZN(n12268) );
  INV_X1 U14497 ( .A(n12256), .ZN(n12228) );
  NAND2_X1 U14498 ( .A1(n12077), .A2(n12074), .ZN(n12073) );
  NAND2_X1 U14499 ( .A1(n6565), .A2(n12073), .ZN(n12080) );
  OAI21_X1 U14500 ( .B1(n12075), .B2(n10803), .A(n12074), .ZN(n12076) );
  NAND2_X1 U14501 ( .A1(n12076), .A2(n6565), .ZN(n12078) );
  NAND2_X1 U14502 ( .A1(n12078), .A2(n12077), .ZN(n12079) );
  MUX2_X1 U14503 ( .A(n12080), .B(n12079), .S(n12213), .Z(n12084) );
  AND2_X1 U14504 ( .A1(n12081), .A2(n12094), .ZN(n12082) );
  NAND2_X1 U14505 ( .A1(n12085), .A2(n12087), .ZN(n12090) );
  NAND2_X1 U14506 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  NAND2_X1 U14507 ( .A1(n12211), .A2(n12088), .ZN(n12089) );
  NAND2_X1 U14508 ( .A1(n12090), .A2(n12089), .ZN(n12099) );
  MUX2_X1 U14509 ( .A(n12092), .B(n12091), .S(n12213), .Z(n12093) );
  NAND2_X1 U14510 ( .A1(n12093), .A2(n12237), .ZN(n12097) );
  AOI21_X1 U14511 ( .B1(n12099), .B2(n9605), .A(n12097), .ZN(n12103) );
  INV_X1 U14512 ( .A(n12094), .ZN(n12095) );
  NOR2_X1 U14513 ( .A1(n12096), .A2(n12095), .ZN(n12098) );
  AOI21_X1 U14514 ( .B1(n12099), .B2(n12098), .A(n12097), .ZN(n12101) );
  OR3_X1 U14515 ( .A1(n12101), .A2(n7167), .A3(n7169), .ZN(n12102) );
  OAI211_X1 U14516 ( .C1(n12103), .C2(n12211), .A(n12102), .B(n12105), .ZN(
        n12108) );
  NAND2_X1 U14517 ( .A1(n12105), .A2(n12104), .ZN(n12106) );
  NAND2_X1 U14518 ( .A1(n12213), .A2(n12106), .ZN(n12107) );
  NAND2_X1 U14519 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  OAI211_X1 U14520 ( .C1(n12211), .C2(n12110), .A(n12109), .B(n12235), .ZN(
        n12114) );
  MUX2_X1 U14521 ( .A(n12112), .B(n12111), .S(n12213), .Z(n12113) );
  NAND3_X1 U14522 ( .A1(n12114), .A2(n12234), .A3(n12113), .ZN(n12118) );
  MUX2_X1 U14523 ( .A(n12116), .B(n12115), .S(n12213), .Z(n12117) );
  NAND3_X1 U14524 ( .A1(n12118), .A2(n12238), .A3(n12117), .ZN(n12123) );
  MUX2_X1 U14525 ( .A(n12119), .B(n12631), .S(n12213), .Z(n12121) );
  AOI21_X1 U14526 ( .B1(n12121), .B2(n12120), .A(n12239), .ZN(n12122) );
  NAND2_X1 U14527 ( .A1(n12123), .A2(n12122), .ZN(n12124) );
  OAI21_X1 U14528 ( .B1(n12125), .B2(n12213), .A(n12124), .ZN(n12131) );
  INV_X1 U14529 ( .A(n12126), .ZN(n12127) );
  NAND2_X1 U14530 ( .A1(n12243), .A2(n12127), .ZN(n12129) );
  NAND3_X1 U14531 ( .A1(n12129), .A2(n12137), .A3(n12128), .ZN(n12130) );
  AOI22_X1 U14532 ( .A1(n12131), .A2(n12243), .B1(n12213), .B2(n12130), .ZN(
        n12136) );
  INV_X1 U14533 ( .A(n12132), .ZN(n12135) );
  OAI21_X1 U14534 ( .B1(n12583), .B2(n12587), .A(n12132), .ZN(n12133) );
  NAND2_X1 U14535 ( .A1(n12133), .A2(n12211), .ZN(n12134) );
  OAI21_X1 U14536 ( .B1(n12136), .B2(n12135), .A(n12134), .ZN(n12140) );
  INV_X1 U14537 ( .A(n12137), .ZN(n12138) );
  NAND2_X1 U14538 ( .A1(n12211), .A2(n12138), .ZN(n12139) );
  NAND3_X1 U14539 ( .A1(n12140), .A2(n12999), .A3(n12139), .ZN(n12144) );
  MUX2_X1 U14540 ( .A(n12142), .B(n12141), .S(n12213), .Z(n12143) );
  NAND4_X1 U14541 ( .A1(n12144), .A2(n12965), .A3(n9309), .A4(n12143), .ZN(
        n12150) );
  INV_X1 U14542 ( .A(n12965), .ZN(n12963) );
  OR2_X1 U14543 ( .A1(n13079), .A2(n12940), .ZN(n12145) );
  OAI211_X1 U14544 ( .C1(n12963), .C2(n12147), .A(n12146), .B(n12145), .ZN(
        n12148) );
  NAND2_X1 U14545 ( .A1(n12148), .A2(n12213), .ZN(n12149) );
  NAND2_X1 U14546 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  NAND2_X1 U14547 ( .A1(n12151), .A2(n12152), .ZN(n12157) );
  OAI211_X1 U14548 ( .C1(n12963), .C2(n12154), .A(n12153), .B(n12152), .ZN(
        n12155) );
  NAND2_X1 U14549 ( .A1(n12155), .A2(n12211), .ZN(n12156) );
  NAND2_X1 U14550 ( .A1(n12157), .A2(n12156), .ZN(n12159) );
  OR3_X1 U14551 ( .A1(n13079), .A2(n12940), .A3(n12213), .ZN(n12158) );
  NAND2_X1 U14552 ( .A1(n12159), .A2(n12158), .ZN(n12161) );
  NAND2_X1 U14553 ( .A1(n12161), .A2(n12160), .ZN(n12170) );
  INV_X1 U14554 ( .A(n12162), .ZN(n12173) );
  INV_X1 U14555 ( .A(n12163), .ZN(n12164) );
  NAND2_X1 U14556 ( .A1(n12171), .A2(n12164), .ZN(n12165) );
  AND3_X1 U14557 ( .A1(n12173), .A2(n12166), .A3(n12165), .ZN(n12167) );
  OAI21_X1 U14558 ( .B1(n12170), .B2(n12928), .A(n12167), .ZN(n12168) );
  NAND2_X1 U14559 ( .A1(n12168), .A2(n12172), .ZN(n12177) );
  AOI21_X1 U14560 ( .B1(n12170), .B2(n12169), .A(n12928), .ZN(n12175) );
  NAND2_X1 U14561 ( .A1(n12172), .A2(n12171), .ZN(n12174) );
  OAI21_X1 U14562 ( .B1(n12175), .B2(n12174), .A(n12173), .ZN(n12176) );
  MUX2_X1 U14563 ( .A(n12177), .B(n12176), .S(n12213), .Z(n12181) );
  NAND2_X1 U14564 ( .A1(n12182), .A2(n12183), .ZN(n12888) );
  INV_X1 U14565 ( .A(n12888), .ZN(n12886) );
  NAND2_X1 U14566 ( .A1(n12211), .A2(n12913), .ZN(n12179) );
  NAND2_X1 U14567 ( .A1(n12213), .A2(n12522), .ZN(n12178) );
  MUX2_X1 U14568 ( .A(n12179), .B(n12178), .S(n13142), .Z(n12180) );
  OAI211_X1 U14569 ( .C1(n12181), .C2(n12896), .A(n12886), .B(n12180), .ZN(
        n12186) );
  NAND2_X1 U14570 ( .A1(n12187), .A2(n12188), .ZN(n12877) );
  INV_X1 U14571 ( .A(n12877), .ZN(n12185) );
  MUX2_X1 U14572 ( .A(n12183), .B(n12182), .S(n12213), .Z(n12184) );
  NAND3_X1 U14573 ( .A1(n12186), .A2(n12185), .A3(n12184), .ZN(n12191) );
  MUX2_X1 U14574 ( .A(n12188), .B(n12187), .S(n12211), .Z(n12189) );
  AND2_X1 U14575 ( .A1(n12860), .A2(n12189), .ZN(n12190) );
  NAND4_X1 U14576 ( .A1(n12191), .A2(n12842), .A3(n12190), .A4(n12823), .ZN(
        n12204) );
  OR2_X1 U14577 ( .A1(n12837), .A2(n12847), .ZN(n12195) );
  INV_X1 U14578 ( .A(n12872), .ZN(n13127) );
  AND2_X1 U14579 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  MUX2_X1 U14580 ( .A(n12195), .B(n12194), .S(n12211), .Z(n12203) );
  NAND2_X1 U14581 ( .A1(n12200), .A2(n12196), .ZN(n12198) );
  AND2_X1 U14582 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  MUX2_X1 U14583 ( .A(n12200), .B(n12199), .S(n12213), .Z(n12201) );
  OR2_X1 U14584 ( .A1(n12201), .A2(n12829), .ZN(n12202) );
  NAND4_X1 U14585 ( .A1(n12204), .A2(n12813), .A3(n12203), .A4(n12202), .ZN(
        n12210) );
  MUX2_X1 U14586 ( .A(n12206), .B(n12205), .S(n12211), .Z(n12207) );
  INV_X1 U14587 ( .A(n12207), .ZN(n12208) );
  NOR2_X1 U14588 ( .A1(n12799), .A2(n12208), .ZN(n12209) );
  NAND3_X1 U14589 ( .A1(n12212), .A2(n12211), .A3(n12786), .ZN(n12222) );
  INV_X1 U14590 ( .A(n12212), .ZN(n12219) );
  NAND2_X1 U14591 ( .A1(n12214), .A2(n12213), .ZN(n12216) );
  NAND2_X1 U14592 ( .A1(n12216), .A2(n12215), .ZN(n12217) );
  NAND3_X1 U14593 ( .A1(n12219), .A2(n12218), .A3(n12217), .ZN(n12220) );
  NAND4_X1 U14594 ( .A1(n12222), .A2(n12221), .A3(n12254), .A4(n12220), .ZN(
        n12226) );
  INV_X1 U14595 ( .A(n12223), .ZN(n12225) );
  NAND2_X1 U14596 ( .A1(n12226), .A2(n6606), .ZN(n12227) );
  INV_X1 U14597 ( .A(n12262), .ZN(n12230) );
  NOR2_X1 U14598 ( .A1(n12230), .A2(n12229), .ZN(n12266) );
  NOR2_X1 U14599 ( .A1(n12829), .A2(n12845), .ZN(n12251) );
  NOR2_X1 U14600 ( .A1(n12232), .A2(n15113), .ZN(n12236) );
  NAND4_X1 U14601 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12242) );
  NAND4_X1 U14602 ( .A1(n13018), .A2(n9605), .A3(n12237), .A4(n15044), .ZN(
        n12241) );
  INV_X1 U14603 ( .A(n12238), .ZN(n12240) );
  NOR4_X1 U14604 ( .A1(n12242), .A2(n12241), .A3(n12240), .A4(n12239), .ZN(
        n12245) );
  NAND4_X1 U14605 ( .A1(n12245), .A2(n12999), .A3(n12244), .A4(n12243), .ZN(
        n12246) );
  NOR4_X1 U14606 ( .A1(n12937), .A2(n12247), .A3(n12963), .A4(n12246), .ZN(
        n12248) );
  NAND3_X1 U14607 ( .A1(n12909), .A2(n12248), .A3(n12956), .ZN(n12249) );
  NOR4_X1 U14608 ( .A1(n12888), .A2(n12877), .A3(n12928), .A4(n12249), .ZN(
        n12250) );
  NAND4_X1 U14609 ( .A1(n12898), .A2(n12813), .A3(n12251), .A4(n12250), .ZN(
        n12253) );
  NOR2_X1 U14610 ( .A1(n12253), .A2(n12252), .ZN(n12255) );
  INV_X1 U14611 ( .A(n12799), .ZN(n12801) );
  NAND4_X1 U14612 ( .A1(n12255), .A2(n12801), .A3(n12786), .A4(n12254), .ZN(
        n12258) );
  XNOR2_X1 U14613 ( .A(n12260), .B(n12259), .ZN(n12264) );
  OAI22_X1 U14614 ( .A1(n12264), .A2(n12263), .B1(n12262), .B2(n12261), .ZN(
        n12265) );
  AOI211_X1 U14615 ( .C1(n12268), .C2(n12267), .A(n12266), .B(n12265), .ZN(
        n12275) );
  NAND3_X1 U14616 ( .A1(n12270), .A2(n12269), .A3(n12733), .ZN(n12271) );
  OAI211_X1 U14617 ( .C1(n12272), .C2(n12274), .A(n12271), .B(P3_B_REG_SCAN_IN), .ZN(n12273) );
  OAI21_X1 U14618 ( .B1(n12275), .B2(n12274), .A(n12273), .ZN(P3_U3296) );
  INV_X1 U14619 ( .A(n12276), .ZN(n12445) );
  OAI222_X1 U14620 ( .A1(n13729), .A2(n12445), .B1(P2_U3088), .B2(n12277), 
        .C1(n12278), .C2(n13739), .ZN(P2_U3297) );
  NAND2_X1 U14621 ( .A1(n12279), .A2(n12630), .ZN(n12280) );
  XNOR2_X1 U14622 ( .A(n10809), .B(n12587), .ZN(n12283) );
  XNOR2_X2 U14623 ( .A(n12282), .B(n12283), .ZN(n12584) );
  INV_X1 U14624 ( .A(n12282), .ZN(n12284) );
  NAND2_X1 U14625 ( .A1(n12284), .A2(n12283), .ZN(n12285) );
  XNOR2_X1 U14626 ( .A(n10809), .B(n12531), .ZN(n12526) );
  INV_X1 U14627 ( .A(n12526), .ZN(n12286) );
  NAND2_X1 U14628 ( .A1(n12286), .A2(n12628), .ZN(n12287) );
  XNOR2_X1 U14629 ( .A(n13003), .B(n10809), .ZN(n12289) );
  INV_X1 U14630 ( .A(n12289), .ZN(n12288) );
  AND2_X1 U14631 ( .A1(n12289), .A2(n12984), .ZN(n12568) );
  XNOR2_X1 U14632 ( .A(n13087), .B(n10809), .ZN(n12290) );
  XNOR2_X1 U14633 ( .A(n12290), .B(n12969), .ZN(n12489) );
  XNOR2_X1 U14634 ( .A(n12974), .B(n10809), .ZN(n12291) );
  XNOR2_X1 U14635 ( .A(n12291), .B(n12983), .ZN(n12615) );
  NAND2_X1 U14636 ( .A1(n12616), .A2(n12615), .ZN(n12614) );
  INV_X1 U14637 ( .A(n12291), .ZN(n12292) );
  NAND2_X1 U14638 ( .A1(n12292), .A2(n12983), .ZN(n12293) );
  NAND2_X1 U14639 ( .A1(n12614), .A2(n12293), .ZN(n12548) );
  XNOR2_X1 U14640 ( .A(n13079), .B(n10809), .ZN(n12294) );
  XNOR2_X1 U14641 ( .A(n12294), .B(n12968), .ZN(n12547) );
  NAND2_X1 U14642 ( .A1(n12548), .A2(n12547), .ZN(n12546) );
  INV_X1 U14643 ( .A(n12294), .ZN(n12295) );
  NAND2_X1 U14644 ( .A1(n12295), .A2(n12968), .ZN(n12296) );
  NAND2_X1 U14645 ( .A1(n12546), .A2(n12296), .ZN(n12555) );
  XNOR2_X1 U14646 ( .A(n13076), .B(n10809), .ZN(n12297) );
  XNOR2_X1 U14647 ( .A(n12297), .B(n12949), .ZN(n12554) );
  NAND2_X1 U14648 ( .A1(n12555), .A2(n12554), .ZN(n12553) );
  INV_X1 U14649 ( .A(n12297), .ZN(n12298) );
  NAND2_X1 U14650 ( .A1(n12298), .A2(n12949), .ZN(n12299) );
  NAND2_X1 U14651 ( .A1(n12553), .A2(n12299), .ZN(n12599) );
  XNOR2_X1 U14652 ( .A(n12596), .B(n10809), .ZN(n12300) );
  XNOR2_X1 U14653 ( .A(n12300), .B(n12914), .ZN(n12598) );
  INV_X1 U14654 ( .A(n12300), .ZN(n12301) );
  NAND2_X1 U14655 ( .A1(n12301), .A2(n12914), .ZN(n12302) );
  NAND2_X1 U14656 ( .A1(n12597), .A2(n12302), .ZN(n12503) );
  XNOR2_X1 U14657 ( .A(n13066), .B(n7398), .ZN(n12303) );
  XNOR2_X1 U14658 ( .A(n12303), .B(n12900), .ZN(n12502) );
  NAND2_X1 U14659 ( .A1(n12503), .A2(n12502), .ZN(n12501) );
  INV_X1 U14660 ( .A(n12303), .ZN(n12304) );
  NAND2_X1 U14661 ( .A1(n12304), .A2(n12900), .ZN(n12305) );
  XNOR2_X1 U14662 ( .A(n13142), .B(n10809), .ZN(n12306) );
  XNOR2_X1 U14663 ( .A(n12306), .B(n12913), .ZN(n12561) );
  INV_X1 U14664 ( .A(n12306), .ZN(n12307) );
  NAND2_X1 U14665 ( .A1(n12307), .A2(n12913), .ZN(n12308) );
  XNOR2_X1 U14666 ( .A(n13136), .B(n7398), .ZN(n12309) );
  XNOR2_X1 U14667 ( .A(n12309), .B(n12901), .ZN(n12519) );
  INV_X1 U14668 ( .A(n12309), .ZN(n12310) );
  XNOR2_X1 U14669 ( .A(n13130), .B(n7398), .ZN(n12470) );
  XNOR2_X1 U14670 ( .A(n12480), .B(n12470), .ZN(n12577) );
  INV_X1 U14671 ( .A(n12470), .ZN(n12311) );
  AND2_X1 U14672 ( .A1(n12480), .A2(n12311), .ZN(n12312) );
  XNOR2_X1 U14673 ( .A(n12872), .B(n10809), .ZN(n12473) );
  XNOR2_X1 U14674 ( .A(n12855), .B(n10809), .ZN(n12472) );
  XOR2_X1 U14675 ( .A(n12826), .B(n12472), .Z(n12315) );
  XNOR2_X1 U14676 ( .A(n12316), .B(n12315), .ZN(n12321) );
  AOI22_X1 U14677 ( .A1(n15038), .A2(n12626), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12318) );
  NAND2_X1 U14678 ( .A1(n12620), .A2(n12851), .ZN(n12317) );
  OAI211_X1 U14679 ( .C1(n12881), .C2(n12618), .A(n12318), .B(n12317), .ZN(
        n12319) );
  AOI21_X1 U14680 ( .B1(n12855), .B2(n15040), .A(n12319), .ZN(n12320) );
  OAI21_X1 U14681 ( .B1(n12321), .B2(n15043), .A(n12320), .ZN(P3_U3169) );
  INV_X1 U14682 ( .A(n12322), .ZN(n12323) );
  OAI222_X1 U14683 ( .A1(n14525), .A2(n12324), .B1(n11389), .B2(n12323), .C1(
        P3_U3151), .C2(n10802), .ZN(P3_U3275) );
  NOR2_X1 U14684 ( .A1(n12455), .A2(n12328), .ZN(n12329) );
  AOI21_X1 U14685 ( .B1(n13843), .B2(n12423), .A(n12329), .ZN(n12331) );
  AOI22_X1 U14686 ( .A1(n13843), .A2(n12417), .B1(n12418), .B2(n13904), .ZN(
        n12330) );
  XNOR2_X1 U14687 ( .A(n12330), .B(n12459), .ZN(n12332) );
  XOR2_X1 U14688 ( .A(n12331), .B(n12332), .Z(n13836) );
  AOI22_X1 U14689 ( .A1(n14617), .A2(n12418), .B1(n12422), .B2(n13903), .ZN(
        n12334) );
  AOI22_X1 U14690 ( .A1(n14617), .A2(n12417), .B1(n12418), .B2(n13903), .ZN(
        n12333) );
  XNOR2_X1 U14691 ( .A(n12333), .B(n12459), .ZN(n12335) );
  XOR2_X1 U14692 ( .A(n12334), .B(n12335), .Z(n14611) );
  AOI22_X1 U14693 ( .A1(n14351), .A2(n12417), .B1(n12418), .B2(n13902), .ZN(
        n12336) );
  XNOR2_X1 U14694 ( .A(n12336), .B(n12459), .ZN(n12339) );
  OAI22_X1 U14695 ( .A1(n12337), .A2(n12456), .B1(n13799), .B2(n12455), .ZN(
        n13880) );
  INV_X1 U14696 ( .A(n12339), .ZN(n12340) );
  OAI22_X1 U14697 ( .A1(n14344), .A2(n12458), .B1(n13882), .B2(n12456), .ZN(
        n12341) );
  XNOR2_X1 U14698 ( .A(n12341), .B(n8097), .ZN(n12346) );
  OR2_X1 U14699 ( .A1(n14344), .A2(n12456), .ZN(n12343) );
  NAND2_X1 U14700 ( .A1(n12422), .A2(n13901), .ZN(n12342) );
  NAND2_X1 U14701 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  XNOR2_X1 U14702 ( .A(n12346), .B(n12344), .ZN(n13793) );
  INV_X1 U14703 ( .A(n12344), .ZN(n12345) );
  OAI22_X1 U14704 ( .A1(n14338), .A2(n12458), .B1(n13862), .B2(n12456), .ZN(
        n12347) );
  XNOR2_X1 U14705 ( .A(n12347), .B(n12459), .ZN(n12350) );
  OR2_X1 U14706 ( .A1(n14338), .A2(n12456), .ZN(n12349) );
  NAND2_X1 U14707 ( .A1(n14235), .A2(n12422), .ZN(n12348) );
  NAND2_X1 U14708 ( .A1(n12349), .A2(n12348), .ZN(n12351) );
  NAND2_X1 U14709 ( .A1(n12350), .A2(n12351), .ZN(n13807) );
  NAND2_X1 U14710 ( .A1(n13806), .A2(n13807), .ZN(n13805) );
  INV_X1 U14711 ( .A(n12350), .ZN(n12353) );
  INV_X1 U14712 ( .A(n12351), .ZN(n12352) );
  NAND2_X1 U14713 ( .A1(n12353), .A2(n12352), .ZN(n13809) );
  NAND2_X1 U14714 ( .A1(n13805), .A2(n13809), .ZN(n13857) );
  NAND2_X1 U14715 ( .A1(n14332), .A2(n12417), .ZN(n12355) );
  NAND2_X1 U14716 ( .A1(n13900), .A2(n12423), .ZN(n12354) );
  NAND2_X1 U14717 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  XNOR2_X1 U14718 ( .A(n12356), .B(n12459), .ZN(n12357) );
  AOI22_X1 U14719 ( .A1(n14332), .A2(n12418), .B1(n12422), .B2(n13900), .ZN(
        n12358) );
  XNOR2_X1 U14720 ( .A(n12357), .B(n12358), .ZN(n13858) );
  INV_X1 U14721 ( .A(n12357), .ZN(n12359) );
  NAND2_X1 U14722 ( .A1(n12359), .A2(n12358), .ZN(n12360) );
  AND2_X1 U14723 ( .A1(n14237), .A2(n12422), .ZN(n12361) );
  AOI21_X1 U14724 ( .B1(n14325), .B2(n12418), .A(n12361), .ZN(n12365) );
  NAND2_X1 U14725 ( .A1(n14325), .A2(n12417), .ZN(n12363) );
  NAND2_X1 U14726 ( .A1(n14237), .A2(n12423), .ZN(n12362) );
  NAND2_X1 U14727 ( .A1(n12363), .A2(n12362), .ZN(n12364) );
  XNOR2_X1 U14728 ( .A(n12364), .B(n12459), .ZN(n12367) );
  XOR2_X1 U14729 ( .A(n12365), .B(n12367), .Z(n13753) );
  INV_X1 U14730 ( .A(n12365), .ZN(n12366) );
  NAND2_X1 U14731 ( .A1(n12367), .A2(n12366), .ZN(n12368) );
  AND2_X1 U14732 ( .A1(n13899), .A2(n12422), .ZN(n12369) );
  AOI21_X1 U14733 ( .B1(n14315), .B2(n12418), .A(n12369), .ZN(n12372) );
  AOI22_X1 U14734 ( .A1(n14315), .A2(n12417), .B1(n12418), .B2(n13899), .ZN(
        n12370) );
  XNOR2_X1 U14735 ( .A(n12370), .B(n12459), .ZN(n12371) );
  XOR2_X1 U14736 ( .A(n12372), .B(n12371), .Z(n13826) );
  INV_X1 U14737 ( .A(n12371), .ZN(n12374) );
  INV_X1 U14738 ( .A(n12372), .ZN(n12373) );
  NAND2_X1 U14739 ( .A1(n12374), .A2(n12373), .ZN(n12375) );
  AOI22_X1 U14740 ( .A1(n14384), .A2(n12417), .B1(n12418), .B2(n13898), .ZN(
        n12376) );
  XNOR2_X1 U14741 ( .A(n12376), .B(n12459), .ZN(n12379) );
  AOI22_X1 U14742 ( .A1(n14384), .A2(n12418), .B1(n12422), .B2(n13898), .ZN(
        n12378) );
  XNOR2_X1 U14743 ( .A(n12379), .B(n12378), .ZN(n13777) );
  INV_X1 U14744 ( .A(n13777), .ZN(n12377) );
  NAND2_X1 U14745 ( .A1(n12379), .A2(n12378), .ZN(n12380) );
  OAI22_X1 U14746 ( .A1(n14380), .A2(n12458), .B1(n12381), .B2(n12456), .ZN(
        n12382) );
  XNOR2_X1 U14747 ( .A(n12382), .B(n12459), .ZN(n12384) );
  AND2_X1 U14748 ( .A1(n13897), .A2(n12422), .ZN(n12383) );
  AOI21_X1 U14749 ( .B1(n14186), .B2(n12418), .A(n12383), .ZN(n12385) );
  XNOR2_X1 U14750 ( .A(n12384), .B(n12385), .ZN(n13848) );
  INV_X1 U14751 ( .A(n12384), .ZN(n12386) );
  NAND2_X1 U14752 ( .A1(n12386), .A2(n12385), .ZN(n12387) );
  OAI22_X1 U14753 ( .A1(n14376), .A2(n12456), .B1(n14141), .B2(n12455), .ZN(
        n12392) );
  NAND2_X1 U14754 ( .A1(n6770), .A2(n12417), .ZN(n12389) );
  NAND2_X1 U14755 ( .A1(n12423), .A2(n13896), .ZN(n12388) );
  NAND2_X1 U14756 ( .A1(n12389), .A2(n12388), .ZN(n12390) );
  XNOR2_X1 U14757 ( .A(n12390), .B(n12459), .ZN(n12391) );
  XOR2_X1 U14758 ( .A(n12392), .B(n12391), .Z(n13746) );
  INV_X1 U14759 ( .A(n12391), .ZN(n12394) );
  INV_X1 U14760 ( .A(n12392), .ZN(n12393) );
  NAND2_X1 U14761 ( .A1(n14286), .A2(n12417), .ZN(n12396) );
  NAND2_X1 U14762 ( .A1(n12423), .A2(n13895), .ZN(n12395) );
  NAND2_X1 U14763 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  XNOR2_X1 U14764 ( .A(n12397), .B(n12459), .ZN(n12398) );
  AOI22_X1 U14765 ( .A1(n14286), .A2(n12418), .B1(n12422), .B2(n13895), .ZN(
        n12399) );
  XNOR2_X1 U14766 ( .A(n12398), .B(n12399), .ZN(n13819) );
  NAND2_X1 U14767 ( .A1(n13818), .A2(n13819), .ZN(n12402) );
  INV_X1 U14768 ( .A(n12398), .ZN(n12400) );
  NAND2_X1 U14769 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  OAI22_X1 U14770 ( .A1(n14371), .A2(n12456), .B1(n14143), .B2(n12455), .ZN(
        n12407) );
  NAND2_X1 U14771 ( .A1(n14135), .A2(n12417), .ZN(n12404) );
  NAND2_X1 U14772 ( .A1(n12423), .A2(n13894), .ZN(n12403) );
  NAND2_X1 U14773 ( .A1(n12404), .A2(n12403), .ZN(n12405) );
  XNOR2_X1 U14774 ( .A(n12405), .B(n12459), .ZN(n12406) );
  XOR2_X1 U14775 ( .A(n12407), .B(n12406), .Z(n13785) );
  INV_X1 U14776 ( .A(n12406), .ZN(n12409) );
  INV_X1 U14777 ( .A(n12407), .ZN(n12408) );
  NAND2_X1 U14778 ( .A1(n12409), .A2(n12408), .ZN(n12410) );
  NAND2_X1 U14779 ( .A1(n14270), .A2(n12417), .ZN(n12412) );
  NAND2_X1 U14780 ( .A1(n12418), .A2(n14093), .ZN(n12411) );
  NAND2_X1 U14781 ( .A1(n12412), .A2(n12411), .ZN(n12413) );
  XNOR2_X1 U14782 ( .A(n12413), .B(n12459), .ZN(n12414) );
  AOI22_X1 U14783 ( .A1(n14270), .A2(n12423), .B1(n12422), .B2(n14093), .ZN(
        n12415) );
  XNOR2_X1 U14784 ( .A(n12414), .B(n12415), .ZN(n13870) );
  INV_X1 U14785 ( .A(n12414), .ZN(n12416) );
  NAND2_X1 U14786 ( .A1(n14101), .A2(n12417), .ZN(n12420) );
  NAND2_X1 U14787 ( .A1(n12418), .A2(n13893), .ZN(n12419) );
  NAND2_X1 U14788 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  XNOR2_X1 U14789 ( .A(n12421), .B(n12459), .ZN(n12450) );
  AOI22_X1 U14790 ( .A1(n14101), .A2(n12423), .B1(n12422), .B2(n13893), .ZN(
        n12451) );
  XNOR2_X1 U14791 ( .A(n12450), .B(n12451), .ZN(n12453) );
  XNOR2_X1 U14792 ( .A(n12454), .B(n12453), .ZN(n12424) );
  NAND2_X1 U14793 ( .A1(n12424), .A2(n14613), .ZN(n12429) );
  NOR2_X1 U14794 ( .A1(n14622), .A2(n14102), .ZN(n12427) );
  OAI22_X1 U14795 ( .A1(n12425), .A2(n13884), .B1(n13883), .B2(n12457), .ZN(
        n12426) );
  AOI211_X1 U14796 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n12427), 
        .B(n12426), .ZN(n12428) );
  OAI211_X1 U14797 ( .C1(n14366), .C2(n13868), .A(n12429), .B(n12428), .ZN(
        P1_U3214) );
  INV_X1 U14798 ( .A(n12430), .ZN(n12432) );
  OAI222_X1 U14799 ( .A1(n14525), .A2(n12433), .B1(n11389), .B2(n12432), .C1(
        P3_U3151), .C2(n12431), .ZN(P3_U3267) );
  OAI21_X1 U14800 ( .B1(n12436), .B2(n12435), .A(n12434), .ZN(n12437) );
  NAND2_X1 U14801 ( .A1(n12437), .A2(n14613), .ZN(n12442) );
  AOI22_X1 U14802 ( .A1(n14615), .A2(n12438), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12439) );
  OAI21_X1 U14803 ( .B1(n14727), .B2(n13868), .A(n12439), .ZN(n12440) );
  AOI21_X1 U14804 ( .B1(n13865), .B2(n13948), .A(n12440), .ZN(n12441) );
  OAI21_X1 U14805 ( .B1(n12443), .B2(n12442), .A(n12441), .ZN(P1_U3218) );
  OAI222_X1 U14806 ( .A1(n14413), .A2(n12445), .B1(P1_U3086), .B2(n7649), .C1(
        n12444), .C2(n14410), .ZN(P1_U3325) );
  INV_X1 U14807 ( .A(n12446), .ZN(n12448) );
  OAI222_X1 U14808 ( .A1(n14525), .A2(n12449), .B1(n11389), .B2(n12448), .C1(
        P3_U3151), .C2(n12447), .ZN(P3_U3265) );
  INV_X1 U14809 ( .A(n12450), .ZN(n12452) );
  AOI22_X1 U14810 ( .A1(n12454), .A2(n12453), .B1(n12452), .B2(n12451), .ZN(
        n12464) );
  OAI22_X1 U14811 ( .A1(n14081), .A2(n10913), .B1(n12457), .B2(n12455), .ZN(
        n12462) );
  OAI22_X1 U14812 ( .A1(n14081), .A2(n12458), .B1(n12457), .B2(n12456), .ZN(
        n12460) );
  XNOR2_X1 U14813 ( .A(n12460), .B(n12459), .ZN(n12461) );
  XOR2_X1 U14814 ( .A(n12462), .B(n12461), .Z(n12463) );
  XNOR2_X1 U14815 ( .A(n12464), .B(n12463), .ZN(n12469) );
  INV_X1 U14816 ( .A(n14078), .ZN(n12465) );
  AOI22_X1 U14817 ( .A1(n14615), .A2(n12465), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12466) );
  OAI21_X1 U14818 ( .B1(n14077), .B2(n14622), .A(n12466), .ZN(n12467) );
  AOI21_X1 U14819 ( .B1(n7066), .B2(n14618), .A(n12467), .ZN(n12468) );
  OAI21_X1 U14820 ( .B1(n12469), .B2(n13889), .A(n12468), .ZN(P1_U3220) );
  XNOR2_X1 U14821 ( .A(n13037), .B(n7398), .ZN(n12508) );
  XNOR2_X1 U14822 ( .A(n12508), .B(n12790), .ZN(n12509) );
  OAI22_X1 U14823 ( .A1(n12472), .A2(n12863), .B1(n12881), .B2(n12473), .ZN(
        n12471) );
  AOI21_X1 U14824 ( .B1(n12470), .B2(n12890), .A(n12471), .ZN(n12479) );
  NOR3_X1 U14825 ( .A1(n12471), .A2(n12470), .A3(n12890), .ZN(n12478) );
  INV_X1 U14826 ( .A(n12472), .ZN(n12476) );
  AOI21_X1 U14827 ( .B1(n12473), .B2(n12881), .A(n12863), .ZN(n12475) );
  NAND3_X1 U14828 ( .A1(n12473), .A2(n12881), .A3(n12863), .ZN(n12474) );
  OAI21_X1 U14829 ( .B1(n12476), .B2(n12475), .A(n12474), .ZN(n12477) );
  XNOR2_X1 U14830 ( .A(n12837), .B(n7398), .ZN(n12481) );
  XNOR2_X1 U14831 ( .A(n12481), .B(n12626), .ZN(n12540) );
  XNOR2_X1 U14832 ( .A(n12816), .B(n10809), .ZN(n12482) );
  XNOR2_X1 U14833 ( .A(n12482), .B(n12825), .ZN(n12605) );
  XOR2_X1 U14834 ( .A(n12509), .B(n12510), .Z(n12487) );
  AOI22_X1 U14835 ( .A1(n12606), .A2(n12825), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12484) );
  NAND2_X1 U14836 ( .A1(n12620), .A2(n12806), .ZN(n12483) );
  OAI211_X1 U14837 ( .C1(n12804), .C2(n12609), .A(n12484), .B(n12483), .ZN(
        n12485) );
  AOI21_X1 U14838 ( .B1(n13037), .B2(n15040), .A(n12485), .ZN(n12486) );
  OAI21_X1 U14839 ( .B1(n12487), .B2(n15043), .A(n12486), .ZN(P3_U3154) );
  XOR2_X1 U14840 ( .A(n12489), .B(n12488), .Z(n12495) );
  NAND2_X1 U14841 ( .A1(n15038), .A2(n12983), .ZN(n12490) );
  NAND2_X1 U14842 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12661)
         );
  OAI211_X1 U14843 ( .C1(n12491), .C2(n12618), .A(n12490), .B(n12661), .ZN(
        n12492) );
  AOI21_X1 U14844 ( .B1(n12989), .B2(n12620), .A(n12492), .ZN(n12494) );
  NAND2_X1 U14845 ( .A1(n13087), .A2(n15040), .ZN(n12493) );
  OAI211_X1 U14846 ( .C1(n12495), .C2(n15043), .A(n12494), .B(n12493), .ZN(
        P3_U3155) );
  AOI22_X1 U14847 ( .A1(n12606), .A2(n12890), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12497) );
  NAND2_X1 U14848 ( .A1(n12620), .A2(n12868), .ZN(n12496) );
  OAI211_X1 U14849 ( .C1(n12863), .C2(n12609), .A(n12497), .B(n12496), .ZN(
        n12498) );
  AOI21_X1 U14850 ( .B1(n12872), .B2(n15040), .A(n12498), .ZN(n12499) );
  OAI21_X1 U14851 ( .B1(n12500), .B2(n15043), .A(n12499), .ZN(P3_U3156) );
  OAI211_X1 U14852 ( .C1(n12503), .C2(n12502), .A(n12501), .B(n12613), .ZN(
        n12507) );
  NAND2_X1 U14853 ( .A1(n15038), .A2(n12913), .ZN(n12504) );
  NAND2_X1 U14854 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12763)
         );
  OAI211_X1 U14855 ( .C1(n12941), .C2(n12618), .A(n12504), .B(n12763), .ZN(
        n12505) );
  AOI21_X1 U14856 ( .B1(n12919), .B2(n12620), .A(n12505), .ZN(n12506) );
  OAI211_X1 U14857 ( .C1(n12623), .C2(n13066), .A(n12507), .B(n12506), .ZN(
        P3_U3159) );
  OAI22_X1 U14858 ( .A1(n12510), .A2(n12509), .B1(n12508), .B2(n12790), .ZN(
        n12512) );
  XNOR2_X1 U14859 ( .A(n12789), .B(n10809), .ZN(n12511) );
  XNOR2_X1 U14860 ( .A(n12512), .B(n12511), .ZN(n12517) );
  AOI22_X1 U14861 ( .A1(n12606), .A2(n12790), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12513) );
  OAI21_X1 U14862 ( .B1(n12792), .B2(n12609), .A(n12513), .ZN(n12515) );
  NOR2_X1 U14863 ( .A1(n12795), .A2(n12623), .ZN(n12514) );
  AOI211_X1 U14864 ( .C1(n12620), .C2(n12793), .A(n12515), .B(n12514), .ZN(
        n12516) );
  OAI21_X1 U14865 ( .B1(n12517), .B2(n15043), .A(n12516), .ZN(P3_U3160) );
  AOI21_X1 U14866 ( .B1(n12519), .B2(n12518), .A(n6654), .ZN(n12525) );
  AOI22_X1 U14867 ( .A1(n15038), .A2(n12890), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12521) );
  NAND2_X1 U14868 ( .A1(n12620), .A2(n12893), .ZN(n12520) );
  OAI211_X1 U14869 ( .C1(n12522), .C2(n12618), .A(n12521), .B(n12520), .ZN(
        n12523) );
  AOI21_X1 U14870 ( .B1(n13136), .B2(n15040), .A(n12523), .ZN(n12524) );
  OAI21_X1 U14871 ( .B1(n12525), .B2(n15043), .A(n12524), .ZN(P3_U3163) );
  XNOR2_X1 U14872 ( .A(n12526), .B(n12628), .ZN(n12527) );
  XNOR2_X1 U14873 ( .A(n12528), .B(n12527), .ZN(n12537) );
  AOI21_X1 U14874 ( .B1(n15038), .B2(n12984), .A(n12529), .ZN(n12535) );
  NAND2_X1 U14875 ( .A1(n12620), .A2(n12530), .ZN(n12534) );
  NAND2_X1 U14876 ( .A1(n15040), .A2(n12531), .ZN(n12533) );
  OR2_X1 U14877 ( .A1(n12618), .A2(n12583), .ZN(n12532) );
  NAND4_X1 U14878 ( .A1(n12535), .A2(n12534), .A3(n12533), .A4(n12532), .ZN(
        n12536) );
  AOI21_X1 U14879 ( .B1(n12537), .B2(n12613), .A(n12536), .ZN(n12538) );
  INV_X1 U14880 ( .A(n12538), .ZN(P3_U3164) );
  XOR2_X1 U14881 ( .A(n12540), .B(n12539), .Z(n12545) );
  AOI22_X1 U14882 ( .A1(n15038), .A2(n12825), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12542) );
  NAND2_X1 U14883 ( .A1(n12620), .A2(n12833), .ZN(n12541) );
  OAI211_X1 U14884 ( .C1(n12863), .C2(n12618), .A(n12542), .B(n12541), .ZN(
        n12543) );
  AOI21_X1 U14885 ( .B1(n12837), .B2(n15040), .A(n12543), .ZN(n12544) );
  OAI21_X1 U14886 ( .B1(n12545), .B2(n15043), .A(n12544), .ZN(P3_U3165) );
  OAI211_X1 U14887 ( .C1(n12548), .C2(n12547), .A(n12546), .B(n12613), .ZN(
        n12552) );
  NAND2_X1 U14888 ( .A1(n15038), .A2(n12949), .ZN(n12549) );
  NAND2_X1 U14889 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12698)
         );
  OAI211_X1 U14890 ( .C1(n12951), .C2(n12618), .A(n12549), .B(n12698), .ZN(
        n12550) );
  AOI21_X1 U14891 ( .B1(n12957), .B2(n12620), .A(n12550), .ZN(n12551) );
  OAI211_X1 U14892 ( .C1(n12959), .C2(n12623), .A(n12552), .B(n12551), .ZN(
        P3_U3166) );
  INV_X1 U14893 ( .A(n13076), .ZN(n12944) );
  OAI211_X1 U14894 ( .C1(n12555), .C2(n12554), .A(n12553), .B(n12613), .ZN(
        n12559) );
  NAND2_X1 U14895 ( .A1(n15038), .A2(n12914), .ZN(n12556) );
  NAND2_X1 U14896 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12720)
         );
  OAI211_X1 U14897 ( .C1(n12940), .C2(n12618), .A(n12556), .B(n12720), .ZN(
        n12557) );
  AOI21_X1 U14898 ( .B1(n12942), .B2(n12620), .A(n12557), .ZN(n12558) );
  OAI211_X1 U14899 ( .C1(n12944), .C2(n12623), .A(n12559), .B(n12558), .ZN(
        P3_U3168) );
  OAI211_X1 U14900 ( .C1(n12562), .C2(n12561), .A(n12560), .B(n12613), .ZN(
        n12567) );
  AOI22_X1 U14901 ( .A1(n15038), .A2(n12901), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12564) );
  NAND2_X1 U14902 ( .A1(n12620), .A2(n12904), .ZN(n12563) );
  OAI211_X1 U14903 ( .C1(n12926), .C2(n12618), .A(n12564), .B(n12563), .ZN(
        n12565) );
  AOI21_X1 U14904 ( .B1(n13142), .B2(n15040), .A(n12565), .ZN(n12566) );
  NAND2_X1 U14905 ( .A1(n12567), .A2(n12566), .ZN(P3_U3173) );
  NOR2_X1 U14906 ( .A1(n6726), .A2(n12568), .ZN(n12569) );
  XNOR2_X1 U14907 ( .A(n12570), .B(n12569), .ZN(n12576) );
  INV_X1 U14908 ( .A(n13003), .ZN(n13092) );
  AOI21_X1 U14909 ( .B1(n15038), .B2(n12969), .A(n12571), .ZN(n12573) );
  NAND2_X1 U14910 ( .A1(n12620), .A2(n13005), .ZN(n12572) );
  OAI211_X1 U14911 ( .C1(n13001), .C2(n12618), .A(n12573), .B(n12572), .ZN(
        n12574) );
  AOI21_X1 U14912 ( .B1(n13092), .B2(n15040), .A(n12574), .ZN(n12575) );
  OAI21_X1 U14913 ( .B1(n12576), .B2(n15043), .A(n12575), .ZN(P3_U3174) );
  XNOR2_X1 U14914 ( .A(n12577), .B(n12890), .ZN(n12582) );
  AOI22_X1 U14915 ( .A1(n12606), .A2(n12901), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12579) );
  NAND2_X1 U14916 ( .A1(n12620), .A2(n12883), .ZN(n12578) );
  OAI211_X1 U14917 ( .C1(n12881), .C2(n12609), .A(n12579), .B(n12578), .ZN(
        n12580) );
  AOI21_X1 U14918 ( .B1(n13130), .B2(n15040), .A(n12580), .ZN(n12581) );
  OAI21_X1 U14919 ( .B1(n12582), .B2(n15043), .A(n12581), .ZN(P3_U3175) );
  XNOR2_X1 U14920 ( .A(n12584), .B(n12583), .ZN(n12594) );
  AOI21_X1 U14921 ( .B1(n15038), .B2(n12628), .A(n12585), .ZN(n12592) );
  NAND2_X1 U14922 ( .A1(n12620), .A2(n12586), .ZN(n12591) );
  NAND2_X1 U14923 ( .A1(n15040), .A2(n12587), .ZN(n12590) );
  OR2_X1 U14924 ( .A1(n12618), .A2(n12588), .ZN(n12589) );
  NAND4_X1 U14925 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12593) );
  AOI21_X1 U14926 ( .B1(n12594), .B2(n12613), .A(n12593), .ZN(n12595) );
  INV_X1 U14927 ( .A(n12595), .ZN(P3_U3176) );
  INV_X1 U14928 ( .A(n12596), .ZN(n13154) );
  OAI211_X1 U14929 ( .C1(n12599), .C2(n12598), .A(n12597), .B(n12613), .ZN(
        n12603) );
  NAND2_X1 U14930 ( .A1(n15038), .A2(n12900), .ZN(n12600) );
  NAND2_X1 U14931 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12742)
         );
  OAI211_X1 U14932 ( .C1(n12925), .C2(n12618), .A(n12600), .B(n12742), .ZN(
        n12601) );
  AOI21_X1 U14933 ( .B1(n12931), .B2(n12620), .A(n12601), .ZN(n12602) );
  OAI211_X1 U14934 ( .C1(n13154), .C2(n12623), .A(n12603), .B(n12602), .ZN(
        P3_U3178) );
  XOR2_X1 U14935 ( .A(n12605), .B(n12604), .Z(n12612) );
  AOI22_X1 U14936 ( .A1(n12606), .A2(n12626), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12608) );
  NAND2_X1 U14937 ( .A1(n12620), .A2(n12817), .ZN(n12607) );
  OAI211_X1 U14938 ( .C1(n12815), .C2(n12609), .A(n12608), .B(n12607), .ZN(
        n12610) );
  AOI21_X1 U14939 ( .B1(n12816), .B2(n15040), .A(n12610), .ZN(n12611) );
  OAI21_X1 U14940 ( .B1(n12612), .B2(n15043), .A(n12611), .ZN(P3_U3180) );
  INV_X1 U14941 ( .A(n12974), .ZN(n13164) );
  OAI211_X1 U14942 ( .C1(n12616), .C2(n12615), .A(n12614), .B(n12613), .ZN(
        n12622) );
  NAND2_X1 U14943 ( .A1(n15038), .A2(n12968), .ZN(n12617) );
  NAND2_X1 U14944 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12673)
         );
  OAI211_X1 U14945 ( .C1(n13002), .C2(n12618), .A(n12617), .B(n12673), .ZN(
        n12619) );
  AOI21_X1 U14946 ( .B1(n12973), .B2(n12620), .A(n12619), .ZN(n12621) );
  OAI211_X1 U14947 ( .C1(n13164), .C2(n12623), .A(n12622), .B(n12621), .ZN(
        P3_U3181) );
  MUX2_X1 U14948 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12624), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14949 ( .A(n12625), .B(P3_DATAO_REG_28__SCAN_IN), .S(n12637), .Z(
        P3_U3519) );
  MUX2_X1 U14950 ( .A(n12790), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12637), .Z(
        P3_U3518) );
  MUX2_X1 U14951 ( .A(n12825), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12637), .Z(
        P3_U3517) );
  MUX2_X1 U14952 ( .A(n12626), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12637), .Z(
        P3_U3516) );
  MUX2_X1 U14953 ( .A(n12826), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12637), .Z(
        P3_U3515) );
  MUX2_X1 U14954 ( .A(n12627), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12637), .Z(
        P3_U3514) );
  MUX2_X1 U14955 ( .A(n12901), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12637), .Z(
        P3_U3512) );
  MUX2_X1 U14956 ( .A(n12913), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12637), .Z(
        P3_U3511) );
  MUX2_X1 U14957 ( .A(n12914), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12637), .Z(
        P3_U3509) );
  MUX2_X1 U14958 ( .A(n12949), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12637), .Z(
        P3_U3508) );
  MUX2_X1 U14959 ( .A(n12968), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12637), .Z(
        P3_U3507) );
  MUX2_X1 U14960 ( .A(n12983), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12637), .Z(
        P3_U3506) );
  MUX2_X1 U14961 ( .A(n12969), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12637), .Z(
        P3_U3505) );
  MUX2_X1 U14962 ( .A(n12984), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12637), .Z(
        P3_U3504) );
  MUX2_X1 U14963 ( .A(n12628), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12637), .Z(
        P3_U3503) );
  MUX2_X1 U14964 ( .A(n12629), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12637), .Z(
        P3_U3502) );
  MUX2_X1 U14965 ( .A(n12630), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12637), .Z(
        P3_U3501) );
  MUX2_X1 U14966 ( .A(n12631), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12637), .Z(
        P3_U3500) );
  MUX2_X1 U14967 ( .A(n12632), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12637), .Z(
        P3_U3498) );
  MUX2_X1 U14968 ( .A(n12633), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12637), .Z(
        P3_U3497) );
  MUX2_X1 U14969 ( .A(n12634), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12637), .Z(
        P3_U3496) );
  MUX2_X1 U14970 ( .A(n12635), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12637), .Z(
        P3_U3495) );
  MUX2_X1 U14971 ( .A(n12636), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12637), .Z(
        P3_U3494) );
  MUX2_X1 U14972 ( .A(n9601), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12637), .Z(
        P3_U3492) );
  MUX2_X1 U14973 ( .A(n15110), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12637), .Z(
        P3_U3491) );
  NOR2_X1 U14974 ( .A1(n12647), .A2(n12638), .ZN(n12640) );
  OR2_X1 U14975 ( .A1(n12660), .A2(n12641), .ZN(n12676) );
  OAI21_X1 U14976 ( .B1(n12642), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12676), 
        .ZN(n12650) );
  AOI21_X1 U14977 ( .B1(n12643), .B2(n12650), .A(n12668), .ZN(n12667) );
  INV_X1 U14978 ( .A(n12644), .ZN(n12646) );
  INV_X1 U14979 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12648) );
  OR2_X1 U14980 ( .A1(n12660), .A2(n12648), .ZN(n12675) );
  NAND2_X1 U14981 ( .A1(n12660), .A2(n12648), .ZN(n12649) );
  AND2_X1 U14982 ( .A1(n12675), .A2(n12649), .ZN(n12659) );
  INV_X1 U14983 ( .A(n12650), .ZN(n12651) );
  MUX2_X1 U14984 ( .A(n12659), .B(n12651), .S(n12754), .Z(n12652) );
  OAI211_X1 U14985 ( .C1(n12653), .C2(n12652), .A(n12678), .B(n15099), .ZN(
        n12666) );
  NAND2_X1 U14986 ( .A1(n12655), .A2(n12654), .ZN(n12657) );
  NAND2_X1 U14987 ( .A1(n12657), .A2(n12656), .ZN(n12658) );
  NAND2_X1 U14988 ( .A1(n12658), .A2(n12659), .ZN(n12670) );
  OAI21_X1 U14989 ( .B1(n12659), .B2(n12658), .A(n12670), .ZN(n12664) );
  INV_X1 U14990 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14495) );
  NAND2_X1 U14991 ( .A1(n15097), .A2(n12660), .ZN(n12662) );
  OAI211_X1 U14992 ( .C1(n14495), .C2(n15088), .A(n12662), .B(n12661), .ZN(
        n12663) );
  AOI21_X1 U14993 ( .B1(n12664), .B2(n15080), .A(n12663), .ZN(n12665) );
  OAI211_X1 U14994 ( .C1(n12667), .C2(n15103), .A(n12666), .B(n12665), .ZN(
        P3_U3196) );
  INV_X1 U14995 ( .A(n12688), .ZN(n14528) );
  NOR2_X1 U14996 ( .A1(n12680), .A2(n12669), .ZN(n12689) );
  AOI21_X1 U14997 ( .B1(n12680), .B2(n12669), .A(n12689), .ZN(n12686) );
  INV_X1 U14998 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14502) );
  NAND2_X1 U14999 ( .A1(n12675), .A2(n12670), .ZN(n12693) );
  XNOR2_X1 U15000 ( .A(n12688), .B(n12693), .ZN(n12671) );
  NAND2_X1 U15001 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12671), .ZN(n12694) );
  OAI21_X1 U15002 ( .B1(n12671), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12694), 
        .ZN(n12672) );
  NAND2_X1 U15003 ( .A1(n15080), .A2(n12672), .ZN(n12674) );
  OAI211_X1 U15004 ( .C1(n14502), .C2(n15088), .A(n12674), .B(n12673), .ZN(
        n12684) );
  MUX2_X1 U15005 ( .A(n12676), .B(n12675), .S(n12725), .Z(n12677) );
  INV_X1 U15006 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12679) );
  MUX2_X1 U15007 ( .A(n12680), .B(n12679), .S(n12725), .Z(n12681) );
  NOR2_X1 U15008 ( .A1(n12682), .A2(n12681), .ZN(n12700) );
  AOI211_X1 U15009 ( .C1(n12682), .C2(n12681), .A(n15071), .B(n12700), .ZN(
        n12683) );
  AOI211_X1 U15010 ( .C1(n15097), .C2(n12688), .A(n12684), .B(n12683), .ZN(
        n12685) );
  OAI21_X1 U15011 ( .B1(n12686), .B2(n15103), .A(n12685), .ZN(P3_U3197) );
  NOR2_X1 U15012 ( .A1(n12688), .A2(n12687), .ZN(n12690) );
  AOI22_X1 U15013 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12718), .B1(n12723), 
        .B2(n12709), .ZN(n12691) );
  AOI21_X1 U15014 ( .B1(n12692), .B2(n12691), .A(n12711), .ZN(n12708) );
  NAND2_X1 U15015 ( .A1(n14528), .A2(n12693), .ZN(n12695) );
  NAND2_X1 U15016 ( .A1(n12695), .A2(n12694), .ZN(n12697) );
  XNOR2_X1 U15017 ( .A(n12718), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12696) );
  NAND2_X1 U15018 ( .A1(n12696), .A2(n12697), .ZN(n12716) );
  OAI21_X1 U15019 ( .B1(n12697), .B2(n12696), .A(n12716), .ZN(n12706) );
  INV_X1 U15020 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14508) );
  NAND2_X1 U15021 ( .A1(n15097), .A2(n12718), .ZN(n12699) );
  OAI211_X1 U15022 ( .C1(n14508), .C2(n15088), .A(n12699), .B(n12698), .ZN(
        n12705) );
  AOI21_X1 U15023 ( .B1(n14528), .B2(n12701), .A(n12700), .ZN(n12703) );
  MUX2_X1 U15024 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12725), .Z(n12724) );
  XNOR2_X1 U15025 ( .A(n12724), .B(n12723), .ZN(n12702) );
  NOR2_X1 U15026 ( .A1(n12703), .A2(n12702), .ZN(n12722) );
  AOI211_X1 U15027 ( .C1(n12703), .C2(n12702), .A(n15071), .B(n12722), .ZN(
        n12704) );
  AOI211_X1 U15028 ( .C1(n15080), .C2(n12706), .A(n12705), .B(n12704), .ZN(
        n12707) );
  OAI21_X1 U15029 ( .B1(n12708), .B2(n15103), .A(n12707), .ZN(P3_U3198) );
  NOR2_X1 U15030 ( .A1(n12718), .A2(n12709), .ZN(n12710) );
  INV_X1 U15031 ( .A(n12749), .ZN(n12713) );
  AOI21_X1 U15032 ( .B1(n12715), .B2(n12714), .A(n12713), .ZN(n12732) );
  INV_X1 U15033 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15331) );
  INV_X1 U15034 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12717) );
  OAI21_X1 U15035 ( .B1(n12718), .B2(n12717), .A(n12716), .ZN(n12738) );
  XNOR2_X1 U15036 ( .A(n12740), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U15037 ( .A1(n15080), .A2(n12719), .ZN(n12721) );
  OAI211_X1 U15038 ( .C1(n15088), .C2(n15331), .A(n12721), .B(n12720), .ZN(
        n12729) );
  AOI21_X1 U15039 ( .B1(n12724), .B2(n12723), .A(n12722), .ZN(n12727) );
  MUX2_X1 U15040 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12725), .Z(n12735) );
  XOR2_X1 U15041 ( .A(n12735), .B(n12730), .Z(n12726) );
  NOR2_X1 U15042 ( .A1(n12727), .A2(n12726), .ZN(n12734) );
  AOI211_X1 U15043 ( .C1(n12727), .C2(n12726), .A(n15071), .B(n12734), .ZN(
        n12728) );
  AOI211_X1 U15044 ( .C1(n15097), .C2(n12730), .A(n12729), .B(n12728), .ZN(
        n12731) );
  OAI21_X1 U15045 ( .B1(n12732), .B2(n15103), .A(n12731), .ZN(P3_U3199) );
  MUX2_X1 U15046 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12733), .Z(n12737) );
  AOI21_X1 U15047 ( .B1(n12737), .B2(n12736), .A(n12755), .ZN(n12753) );
  INV_X1 U15048 ( .A(n15080), .ZN(n12744) );
  XOR2_X1 U15049 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12758), .Z(n12759) );
  XOR2_X1 U15050 ( .A(n12759), .B(n12760), .Z(n12743) );
  NAND2_X1 U15051 ( .A1(n15093), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12741) );
  OAI211_X1 U15052 ( .C1(n12744), .C2(n12743), .A(n12742), .B(n12741), .ZN(
        n12745) );
  AOI21_X1 U15053 ( .B1(n12758), .B2(n15097), .A(n12745), .ZN(n12752) );
  OR2_X1 U15054 ( .A1(n12758), .A2(n15465), .ZN(n12769) );
  NAND2_X1 U15055 ( .A1(n12758), .A2(n15465), .ZN(n12746) );
  NAND2_X1 U15056 ( .A1(n12769), .A2(n12746), .ZN(n12747) );
  AND3_X1 U15057 ( .A1(n12749), .A2(n12748), .A3(n12747), .ZN(n12750) );
  OAI21_X1 U15058 ( .B1(n12771), .B2(n12750), .A(n12774), .ZN(n12751) );
  OAI211_X1 U15059 ( .C1(n12753), .C2(n15071), .A(n12752), .B(n12751), .ZN(
        P3_U3200) );
  XNOR2_X1 U15060 ( .A(n12764), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12762) );
  XNOR2_X1 U15061 ( .A(n12764), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12772) );
  MUX2_X1 U15062 ( .A(n12762), .B(n12772), .S(n12754), .Z(n12757) );
  XOR2_X1 U15063 ( .A(n12757), .B(n12756), .Z(n12778) );
  INV_X1 U15064 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n15330) );
  OAI22_X1 U15065 ( .A1(n12760), .A2(n12759), .B1(n12758), .B2(n15330), .ZN(
        n12761) );
  XOR2_X1 U15066 ( .A(n12762), .B(n12761), .Z(n12768) );
  OAI21_X1 U15067 ( .B1(n15088), .B2(n7545), .A(n12763), .ZN(n12767) );
  NOR2_X1 U15068 ( .A1(n12765), .A2(n12764), .ZN(n12766) );
  INV_X1 U15069 ( .A(n12769), .ZN(n12770) );
  XNOR2_X1 U15070 ( .A(n12773), .B(n12772), .ZN(n12775) );
  NAND2_X1 U15071 ( .A1(n12775), .A2(n12774), .ZN(n12776) );
  OAI211_X1 U15072 ( .C1(n12778), .C2(n15071), .A(n12777), .B(n12776), .ZN(
        P3_U3201) );
  OR2_X1 U15073 ( .A1(n12781), .A2(n12780), .ZN(n14560) );
  OAI21_X1 U15074 ( .B1(n15129), .B2(n14560), .A(n12782), .ZN(n12784) );
  AOI21_X1 U15075 ( .B1(n15129), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12784), 
        .ZN(n12783) );
  OAI21_X1 U15076 ( .B1(n13097), .B2(n13004), .A(n12783), .ZN(P3_U3202) );
  AOI21_X1 U15077 ( .B1(n15129), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12784), 
        .ZN(n12785) );
  OAI21_X1 U15078 ( .B1(n14561), .B2(n13004), .A(n12785), .ZN(P3_U3203) );
  XNOR2_X1 U15079 ( .A(n12787), .B(n12786), .ZN(n13107) );
  NAND2_X1 U15080 ( .A1(n12985), .A2(n12790), .ZN(n12791) );
  AOI22_X1 U15081 ( .A1(n15129), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n12990), 
        .B2(n12793), .ZN(n12794) );
  OAI21_X1 U15082 ( .B1(n12795), .B2(n13004), .A(n12794), .ZN(n12796) );
  AOI21_X1 U15083 ( .B1(n13032), .B2(n6576), .A(n12796), .ZN(n12797) );
  OAI21_X1 U15084 ( .B1(n13107), .B2(n13011), .A(n12797), .ZN(P3_U3205) );
  AOI21_X1 U15085 ( .B1(n12800), .B2(n12799), .A(n12798), .ZN(n13111) );
  XNOR2_X1 U15086 ( .A(n12802), .B(n12801), .ZN(n12803) );
  OAI222_X1 U15087 ( .A1(n15120), .A2(n12805), .B1(n13016), .B2(n12804), .C1(
        n13019), .C2(n12803), .ZN(n13036) );
  AOI22_X1 U15088 ( .A1(n15129), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n12990), 
        .B2(n12806), .ZN(n12807) );
  OAI21_X1 U15089 ( .B1(n12808), .B2(n13004), .A(n12807), .ZN(n12809) );
  AOI21_X1 U15090 ( .B1(n13036), .B2(n6576), .A(n12809), .ZN(n12810) );
  OAI21_X1 U15091 ( .B1(n13111), .B2(n13011), .A(n12810), .ZN(P3_U3206) );
  XNOR2_X1 U15092 ( .A(n12811), .B(n12813), .ZN(n13041) );
  INV_X1 U15093 ( .A(n13041), .ZN(n12821) );
  XOR2_X1 U15094 ( .A(n12813), .B(n12812), .Z(n12814) );
  OAI222_X1 U15095 ( .A1(n15120), .A2(n12847), .B1(n13016), .B2(n12815), .C1(
        n12814), .C2(n13019), .ZN(n13040) );
  INV_X1 U15096 ( .A(n12816), .ZN(n13115) );
  AOI22_X1 U15097 ( .A1(n15129), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n12990), 
        .B2(n12817), .ZN(n12818) );
  OAI21_X1 U15098 ( .B1(n13115), .B2(n13004), .A(n12818), .ZN(n12819) );
  AOI21_X1 U15099 ( .B1(n13040), .B2(n6576), .A(n12819), .ZN(n12820) );
  OAI21_X1 U15100 ( .B1(n13011), .B2(n12821), .A(n12820), .ZN(P3_U3207) );
  OAI21_X1 U15101 ( .B1(n12824), .B2(n12823), .A(n12822), .ZN(n13045) );
  INV_X1 U15102 ( .A(n13045), .ZN(n12840) );
  AOI22_X1 U15103 ( .A1(n12985), .A2(n12826), .B1(n15117), .B2(n12825), .ZN(
        n12832) );
  AND2_X1 U15104 ( .A1(n12844), .A2(n12827), .ZN(n12830) );
  OAI211_X1 U15105 ( .C1(n12830), .C2(n12829), .A(n12828), .B(n15114), .ZN(
        n12831) );
  OAI211_X1 U15106 ( .C1(n12840), .C2(n12867), .A(n12832), .B(n12831), .ZN(
        n13044) );
  NAND2_X1 U15107 ( .A1(n13044), .A2(n6576), .ZN(n12839) );
  INV_X1 U15108 ( .A(n12833), .ZN(n12834) );
  OAI22_X1 U15109 ( .A1(n6576), .A2(n12835), .B1(n12834), .B2(n15123), .ZN(
        n12836) );
  AOI21_X1 U15110 ( .B1(n12837), .B2(n12991), .A(n12836), .ZN(n12838) );
  OAI211_X1 U15111 ( .C1(n12840), .C2(n12875), .A(n12839), .B(n12838), .ZN(
        P3_U3208) );
  OAI21_X1 U15112 ( .B1(n12843), .B2(n12842), .A(n12841), .ZN(n13048) );
  INV_X1 U15113 ( .A(n13048), .ZN(n12858) );
  OAI21_X1 U15114 ( .B1(n12846), .B2(n12845), .A(n12844), .ZN(n12849) );
  OAI22_X1 U15115 ( .A1(n13016), .A2(n12847), .B1(n12881), .B2(n15120), .ZN(
        n12848) );
  AOI21_X1 U15116 ( .B1(n12849), .B2(n15114), .A(n12848), .ZN(n12850) );
  OAI21_X1 U15117 ( .B1(n12858), .B2(n12867), .A(n12850), .ZN(n13047) );
  NAND2_X1 U15118 ( .A1(n13047), .A2(n6576), .ZN(n12857) );
  INV_X1 U15119 ( .A(n12851), .ZN(n12852) );
  OAI22_X1 U15120 ( .A1(n6576), .A2(n12853), .B1(n12852), .B2(n15123), .ZN(
        n12854) );
  AOI21_X1 U15121 ( .B1(n12855), .B2(n12991), .A(n12854), .ZN(n12856) );
  OAI211_X1 U15122 ( .C1(n12858), .C2(n12875), .A(n12857), .B(n12856), .ZN(
        P3_U3209) );
  XNOR2_X1 U15123 ( .A(n12859), .B(n12860), .ZN(n13051) );
  XNOR2_X1 U15124 ( .A(n12861), .B(n12860), .ZN(n12865) );
  OAI22_X1 U15125 ( .A1(n13016), .A2(n12863), .B1(n12862), .B2(n15120), .ZN(
        n12864) );
  AOI21_X1 U15126 ( .B1(n12865), .B2(n15114), .A(n12864), .ZN(n12866) );
  OAI21_X1 U15127 ( .B1(n13051), .B2(n12867), .A(n12866), .ZN(n13052) );
  NAND2_X1 U15128 ( .A1(n13052), .A2(n6576), .ZN(n12874) );
  INV_X1 U15129 ( .A(n12868), .ZN(n12869) );
  OAI22_X1 U15130 ( .A1(n6576), .A2(n12870), .B1(n12869), .B2(n15123), .ZN(
        n12871) );
  AOI21_X1 U15131 ( .B1(n12872), .B2(n12991), .A(n12871), .ZN(n12873) );
  OAI211_X1 U15132 ( .C1(n12875), .C2(n13051), .A(n12874), .B(n12873), .ZN(
        P3_U3210) );
  XNOR2_X1 U15133 ( .A(n12876), .B(n12877), .ZN(n13133) );
  XNOR2_X1 U15134 ( .A(n12878), .B(n12877), .ZN(n12879) );
  OAI222_X1 U15135 ( .A1(n13016), .A2(n12881), .B1(n15120), .B2(n12880), .C1(
        n13019), .C2(n12879), .ZN(n13056) );
  INV_X1 U15136 ( .A(n13056), .ZN(n13128) );
  MUX2_X1 U15137 ( .A(n12882), .B(n13128), .S(n6576), .Z(n12885) );
  AOI22_X1 U15138 ( .A1(n13130), .A2(n12991), .B1(n12990), .B2(n12883), .ZN(
        n12884) );
  OAI211_X1 U15139 ( .C1(n13133), .C2(n13011), .A(n12885), .B(n12884), .ZN(
        P3_U3211) );
  XNOR2_X1 U15140 ( .A(n12887), .B(n12886), .ZN(n13139) );
  XNOR2_X1 U15141 ( .A(n12889), .B(n12888), .ZN(n12891) );
  AOI222_X1 U15142 ( .A1(n15114), .A2(n12891), .B1(n12890), .B2(n15117), .C1(
        n12913), .C2(n12985), .ZN(n13134) );
  MUX2_X1 U15143 ( .A(n12892), .B(n13134), .S(n6576), .Z(n12895) );
  AOI22_X1 U15144 ( .A1(n13136), .A2(n12991), .B1(n12990), .B2(n12893), .ZN(
        n12894) );
  OAI211_X1 U15145 ( .C1(n13139), .C2(n13011), .A(n12895), .B(n12894), .ZN(
        P3_U3212) );
  XNOR2_X1 U15146 ( .A(n12897), .B(n12896), .ZN(n13145) );
  XNOR2_X1 U15147 ( .A(n12899), .B(n12898), .ZN(n12902) );
  AOI222_X1 U15148 ( .A1(n15114), .A2(n12902), .B1(n12901), .B2(n15117), .C1(
        n12900), .C2(n12985), .ZN(n13140) );
  MUX2_X1 U15149 ( .A(n12903), .B(n13140), .S(n6576), .Z(n12906) );
  AOI22_X1 U15150 ( .A1(n13142), .A2(n12991), .B1(n12990), .B2(n12904), .ZN(
        n12905) );
  OAI211_X1 U15151 ( .C1(n13145), .C2(n13011), .A(n12906), .B(n12905), .ZN(
        P3_U3213) );
  XNOR2_X1 U15152 ( .A(n12907), .B(n12909), .ZN(n13150) );
  NOR2_X1 U15153 ( .A1(n13066), .A2(n13004), .ZN(n12918) );
  NAND2_X1 U15154 ( .A1(n12921), .A2(n12908), .ZN(n12910) );
  NAND2_X1 U15155 ( .A1(n12910), .A2(n12909), .ZN(n12912) );
  NAND3_X1 U15156 ( .A1(n12912), .A2(n15114), .A3(n12911), .ZN(n12916) );
  AOI22_X1 U15157 ( .A1(n12985), .A2(n12914), .B1(n15117), .B2(n12913), .ZN(
        n12915) );
  NAND2_X1 U15158 ( .A1(n12916), .A2(n12915), .ZN(n13146) );
  MUX2_X1 U15159 ( .A(n13146), .B(P3_REG2_REG_19__SCAN_IN), .S(n15129), .Z(
        n12917) );
  AOI211_X1 U15160 ( .C1(n12990), .C2(n12919), .A(n12918), .B(n12917), .ZN(
        n12920) );
  OAI21_X1 U15161 ( .B1(n13150), .B2(n13011), .A(n12920), .ZN(P3_U3214) );
  INV_X1 U15162 ( .A(n12921), .ZN(n12922) );
  AOI21_X1 U15163 ( .B1(n9377), .B2(n12923), .A(n12922), .ZN(n12924) );
  OAI222_X1 U15164 ( .A1(n13016), .A2(n12926), .B1(n15120), .B2(n12925), .C1(
        n13019), .C2(n12924), .ZN(n13072) );
  INV_X1 U15165 ( .A(n12927), .ZN(n12930) );
  AND2_X1 U15166 ( .A1(n12929), .A2(n12928), .ZN(n13071) );
  NOR3_X1 U15167 ( .A1(n12930), .A2(n13071), .A3(n13011), .ZN(n12934) );
  AOI22_X1 U15168 ( .A1(n15129), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12990), 
        .B2(n12931), .ZN(n12932) );
  OAI21_X1 U15169 ( .B1(n13154), .B2(n13004), .A(n12932), .ZN(n12933) );
  AOI211_X1 U15170 ( .C1(n13072), .C2(n6576), .A(n12934), .B(n12933), .ZN(
        n12935) );
  INV_X1 U15171 ( .A(n12935), .ZN(P3_U3215) );
  XNOR2_X1 U15172 ( .A(n12936), .B(n12937), .ZN(n13157) );
  XNOR2_X1 U15173 ( .A(n12938), .B(n12937), .ZN(n12939) );
  OAI222_X1 U15174 ( .A1(n13016), .A2(n12941), .B1(n15120), .B2(n12940), .C1(
        n12939), .C2(n13019), .ZN(n13075) );
  AOI22_X1 U15175 ( .A1(n15129), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12990), 
        .B2(n12942), .ZN(n12943) );
  OAI21_X1 U15176 ( .B1(n12944), .B2(n13004), .A(n12943), .ZN(n12945) );
  AOI21_X1 U15177 ( .B1(n13075), .B2(n6576), .A(n12945), .ZN(n12946) );
  OAI21_X1 U15178 ( .B1(n13011), .B2(n13157), .A(n12946), .ZN(P3_U3216) );
  INV_X1 U15179 ( .A(n12956), .ZN(n12947) );
  XNOR2_X1 U15180 ( .A(n12948), .B(n12947), .ZN(n12953) );
  NAND2_X1 U15181 ( .A1(n15117), .A2(n12949), .ZN(n12950) );
  OAI21_X1 U15182 ( .B1(n12951), .B2(n15120), .A(n12950), .ZN(n12952) );
  AOI21_X1 U15183 ( .B1(n12953), .B2(n15114), .A(n12952), .ZN(n13081) );
  OAI21_X1 U15184 ( .B1(n12954), .B2(n12956), .A(n12955), .ZN(n13160) );
  AOI22_X1 U15185 ( .A1(n15129), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12990), 
        .B2(n12957), .ZN(n12958) );
  OAI21_X1 U15186 ( .B1(n12959), .B2(n13004), .A(n12958), .ZN(n12960) );
  AOI21_X1 U15187 ( .B1(n13160), .B2(n12961), .A(n12960), .ZN(n12962) );
  OAI21_X1 U15188 ( .B1(n13081), .B2(n15129), .A(n12962), .ZN(P3_U3217) );
  XNOR2_X1 U15189 ( .A(n12964), .B(n12963), .ZN(n13165) );
  XNOR2_X1 U15190 ( .A(n12966), .B(n12965), .ZN(n12967) );
  NAND2_X1 U15191 ( .A1(n12967), .A2(n15114), .ZN(n12971) );
  AOI22_X1 U15192 ( .A1(n12985), .A2(n12969), .B1(n15117), .B2(n12968), .ZN(
        n12970) );
  NAND2_X1 U15193 ( .A1(n12971), .A2(n12970), .ZN(n13163) );
  MUX2_X1 U15194 ( .A(P3_REG2_REG_15__SCAN_IN), .B(n13163), .S(n6576), .Z(
        n12972) );
  INV_X1 U15195 ( .A(n12972), .ZN(n12976) );
  AOI22_X1 U15196 ( .A1(n12991), .A2(n12974), .B1(n12990), .B2(n12973), .ZN(
        n12975) );
  OAI211_X1 U15197 ( .C1(n13165), .C2(n13011), .A(n12976), .B(n12975), .ZN(
        P3_U3218) );
  XNOR2_X1 U15198 ( .A(n12977), .B(n9309), .ZN(n13171) );
  NAND2_X1 U15199 ( .A1(n12978), .A2(n12979), .ZN(n12980) );
  NAND2_X1 U15200 ( .A1(n12980), .A2(n9309), .ZN(n12982) );
  NAND3_X1 U15201 ( .A1(n12982), .A2(n15114), .A3(n12981), .ZN(n12987) );
  AOI22_X1 U15202 ( .A1(n12985), .A2(n12984), .B1(n15117), .B2(n12983), .ZN(
        n12986) );
  NAND2_X1 U15203 ( .A1(n12987), .A2(n12986), .ZN(n13168) );
  MUX2_X1 U15204 ( .A(n13168), .B(P3_REG2_REG_14__SCAN_IN), .S(n15129), .Z(
        n12988) );
  INV_X1 U15205 ( .A(n12988), .ZN(n12993) );
  AOI22_X1 U15206 ( .A1(n12991), .A2(n13087), .B1(n12990), .B2(n12989), .ZN(
        n12992) );
  OAI211_X1 U15207 ( .C1(n13171), .C2(n13011), .A(n12993), .B(n12992), .ZN(
        P3_U3219) );
  XNOR2_X1 U15208 ( .A(n12995), .B(n12994), .ZN(n13178) );
  INV_X1 U15209 ( .A(n12996), .ZN(n12998) );
  INV_X1 U15210 ( .A(n12978), .ZN(n12997) );
  AOI21_X1 U15211 ( .B1(n12999), .B2(n12998), .A(n12997), .ZN(n13000) );
  OAI222_X1 U15212 ( .A1(n13016), .A2(n13002), .B1(n15120), .B2(n13001), .C1(
        n13019), .C2(n13000), .ZN(n13091) );
  NOR2_X1 U15213 ( .A1(n13004), .A2(n13003), .ZN(n13009) );
  INV_X1 U15214 ( .A(n13005), .ZN(n13006) );
  OAI22_X1 U15215 ( .A1(n6576), .A2(n13007), .B1(n13006), .B2(n15123), .ZN(
        n13008) );
  AOI211_X1 U15216 ( .C1(n13091), .C2(n6576), .A(n13009), .B(n13008), .ZN(
        n13010) );
  OAI21_X1 U15217 ( .B1(n13011), .B2(n13178), .A(n13010), .ZN(P3_U3220) );
  OAI21_X1 U15218 ( .B1(n13013), .B2(n13018), .A(n13012), .ZN(n15137) );
  OAI22_X1 U15219 ( .A1(n13016), .A2(n13015), .B1(n13014), .B2(n15120), .ZN(
        n13023) );
  NAND3_X1 U15220 ( .A1(n15111), .A2(n13018), .A3(n13017), .ZN(n13020) );
  AOI21_X1 U15221 ( .B1(n13021), .B2(n13020), .A(n13019), .ZN(n13022) );
  AOI211_X1 U15222 ( .C1(n13024), .C2(n15137), .A(n13023), .B(n13022), .ZN(
        n15134) );
  NAND2_X1 U15223 ( .A1(n15155), .A2(n13025), .ZN(n15133) );
  OAI22_X1 U15224 ( .A1(n15124), .A2(n15133), .B1(n15123), .B2(n10675), .ZN(
        n13026) );
  AOI21_X1 U15225 ( .B1(n15137), .B2(n13027), .A(n13026), .ZN(n13028) );
  NAND2_X1 U15226 ( .A1(n15134), .A2(n13028), .ZN(n13029) );
  MUX2_X1 U15227 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n13029), .S(n6576), .Z(
        P3_U3231) );
  INV_X1 U15228 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13030) );
  MUX2_X1 U15229 ( .A(n13030), .B(n14560), .S(n15192), .Z(n13031) );
  OAI21_X1 U15230 ( .B1(n13097), .B2(n13088), .A(n13031), .ZN(P3_U3490) );
  INV_X1 U15231 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13034) );
  OAI21_X1 U15232 ( .B1(n13107), .B2(n13095), .A(n13035), .ZN(P3_U3487) );
  INV_X1 U15233 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13038) );
  AOI21_X1 U15234 ( .B1(n15155), .B2(n13037), .A(n13036), .ZN(n13108) );
  OAI21_X1 U15235 ( .B1(n13111), .B2(n13095), .A(n13039), .ZN(P3_U3486) );
  INV_X1 U15236 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13042) );
  AOI21_X1 U15237 ( .B1(n13041), .B2(n15174), .A(n13040), .ZN(n13112) );
  MUX2_X1 U15238 ( .A(n13042), .B(n13112), .S(n15192), .Z(n13043) );
  OAI21_X1 U15239 ( .B1(n13115), .B2(n13088), .A(n13043), .ZN(P3_U3485) );
  INV_X1 U15240 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n15493) );
  INV_X1 U15241 ( .A(n15166), .ZN(n15156) );
  AOI21_X1 U15242 ( .B1(n15156), .B2(n13045), .A(n13044), .ZN(n13116) );
  MUX2_X1 U15243 ( .A(n15493), .B(n13116), .S(n15192), .Z(n13046) );
  OAI21_X1 U15244 ( .B1(n13119), .B2(n13088), .A(n13046), .ZN(P3_U3484) );
  INV_X1 U15245 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13049) );
  AOI21_X1 U15246 ( .B1(n15156), .B2(n13048), .A(n13047), .ZN(n13120) );
  MUX2_X1 U15247 ( .A(n13049), .B(n13120), .S(n15192), .Z(n13050) );
  OAI21_X1 U15248 ( .B1(n13123), .B2(n13088), .A(n13050), .ZN(P3_U3483) );
  INV_X1 U15249 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13054) );
  INV_X1 U15250 ( .A(n13051), .ZN(n13053) );
  AOI21_X1 U15251 ( .B1(n15156), .B2(n13053), .A(n13052), .ZN(n13124) );
  MUX2_X1 U15252 ( .A(n13054), .B(n13124), .S(n15192), .Z(n13055) );
  OAI21_X1 U15253 ( .B1(n13127), .B2(n13088), .A(n13055), .ZN(P3_U3482) );
  MUX2_X1 U15254 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n13056), .S(n15192), .Z(
        n13059) );
  OAI22_X1 U15255 ( .A1(n13133), .A2(n13095), .B1(n13057), .B2(n13088), .ZN(
        n13058) );
  OR2_X1 U15256 ( .A1(n13059), .A2(n13058), .ZN(P3_U3481) );
  INV_X1 U15257 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13060) );
  MUX2_X1 U15258 ( .A(n13060), .B(n13134), .S(n15192), .Z(n13062) );
  NAND2_X1 U15259 ( .A1(n13136), .A2(n13068), .ZN(n13061) );
  OAI211_X1 U15260 ( .C1(n13139), .C2(n13095), .A(n13062), .B(n13061), .ZN(
        P3_U3480) );
  INV_X1 U15261 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13063) );
  MUX2_X1 U15262 ( .A(n13063), .B(n13140), .S(n15192), .Z(n13065) );
  NAND2_X1 U15263 ( .A1(n13142), .A2(n13068), .ZN(n13064) );
  OAI211_X1 U15264 ( .C1(n13145), .C2(n13095), .A(n13065), .B(n13064), .ZN(
        P3_U3479) );
  MUX2_X1 U15265 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13146), .S(n15192), .Z(
        n13067) );
  AOI21_X1 U15266 ( .B1(n13068), .B2(n6854), .A(n13067), .ZN(n13069) );
  OAI21_X1 U15267 ( .B1(n13150), .B2(n13095), .A(n13069), .ZN(P3_U3478) );
  INV_X1 U15268 ( .A(n15174), .ZN(n13070) );
  NOR2_X1 U15269 ( .A1(n13071), .A2(n13070), .ZN(n13073) );
  AOI21_X1 U15270 ( .B1(n13073), .B2(n12927), .A(n13072), .ZN(n13151) );
  MUX2_X1 U15271 ( .A(n15330), .B(n13151), .S(n15192), .Z(n13074) );
  OAI21_X1 U15272 ( .B1(n13154), .B2(n13088), .A(n13074), .ZN(P3_U3477) );
  INV_X1 U15273 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13077) );
  AOI21_X1 U15274 ( .B1(n15155), .B2(n13076), .A(n13075), .ZN(n13155) );
  MUX2_X1 U15275 ( .A(n13077), .B(n13155), .S(n15192), .Z(n13078) );
  OAI21_X1 U15276 ( .B1(n13095), .B2(n13157), .A(n13078), .ZN(P3_U3476) );
  NAND2_X1 U15277 ( .A1(n13079), .A2(n15155), .ZN(n13080) );
  NAND2_X1 U15278 ( .A1(n13081), .A2(n13080), .ZN(n13158) );
  MUX2_X1 U15279 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13158), .S(n15192), .Z(
        n13082) );
  AOI21_X1 U15280 ( .B1(n13083), .B2(n13160), .A(n13082), .ZN(n13084) );
  INV_X1 U15281 ( .A(n13084), .ZN(P3_U3475) );
  MUX2_X1 U15282 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13163), .S(n15192), .Z(
        n13086) );
  OAI22_X1 U15283 ( .A1(n13165), .A2(n13095), .B1(n13164), .B2(n13088), .ZN(
        n13085) );
  OR2_X1 U15284 ( .A1(n13086), .A2(n13085), .ZN(P3_U3474) );
  MUX2_X1 U15285 ( .A(n13168), .B(P3_REG1_REG_14__SCAN_IN), .S(n15189), .Z(
        n13090) );
  INV_X1 U15286 ( .A(n13087), .ZN(n13170) );
  OAI22_X1 U15287 ( .A1(n13171), .A2(n13095), .B1(n13170), .B2(n13088), .ZN(
        n13089) );
  OR2_X1 U15288 ( .A1(n13090), .A2(n13089), .ZN(P3_U3473) );
  INV_X1 U15289 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13093) );
  AOI21_X1 U15290 ( .B1(n15155), .B2(n13092), .A(n13091), .ZN(n13174) );
  MUX2_X1 U15291 ( .A(n13093), .B(n13174), .S(n15192), .Z(n13094) );
  OAI21_X1 U15292 ( .B1(n13095), .B2(n13178), .A(n13094), .ZN(P3_U3472) );
  MUX2_X1 U15293 ( .A(n12060), .B(n14560), .S(n15177), .Z(n13096) );
  OAI21_X1 U15294 ( .B1(n13097), .B2(n13169), .A(n13096), .ZN(P3_U3458) );
  OAI21_X1 U15295 ( .B1(n13103), .B2(n13177), .A(n13102), .ZN(P3_U3456) );
  OAI21_X1 U15296 ( .B1(n13107), .B2(n13177), .A(n13106), .ZN(P3_U3455) );
  OAI21_X1 U15297 ( .B1(n13111), .B2(n13177), .A(n13110), .ZN(P3_U3454) );
  MUX2_X1 U15298 ( .A(n13113), .B(n13112), .S(n15177), .Z(n13114) );
  OAI21_X1 U15299 ( .B1(n13115), .B2(n13169), .A(n13114), .ZN(P3_U3453) );
  MUX2_X1 U15300 ( .A(n13117), .B(n13116), .S(n15177), .Z(n13118) );
  OAI21_X1 U15301 ( .B1(n13119), .B2(n13169), .A(n13118), .ZN(P3_U3452) );
  MUX2_X1 U15302 ( .A(n13121), .B(n13120), .S(n15177), .Z(n13122) );
  OAI21_X1 U15303 ( .B1(n13123), .B2(n13169), .A(n13122), .ZN(P3_U3451) );
  MUX2_X1 U15304 ( .A(n13125), .B(n13124), .S(n15177), .Z(n13126) );
  OAI21_X1 U15305 ( .B1(n13127), .B2(n13169), .A(n13126), .ZN(P3_U3450) );
  MUX2_X1 U15306 ( .A(n13129), .B(n13128), .S(n15177), .Z(n13132) );
  NAND2_X1 U15307 ( .A1(n13130), .A2(n13148), .ZN(n13131) );
  OAI211_X1 U15308 ( .C1(n13133), .C2(n13177), .A(n13132), .B(n13131), .ZN(
        P3_U3449) );
  MUX2_X1 U15309 ( .A(n13135), .B(n13134), .S(n15177), .Z(n13138) );
  NAND2_X1 U15310 ( .A1(n13136), .A2(n13148), .ZN(n13137) );
  OAI211_X1 U15311 ( .C1(n13139), .C2(n13177), .A(n13138), .B(n13137), .ZN(
        P3_U3448) );
  MUX2_X1 U15312 ( .A(n13141), .B(n13140), .S(n15177), .Z(n13144) );
  NAND2_X1 U15313 ( .A1(n13142), .A2(n13148), .ZN(n13143) );
  OAI211_X1 U15314 ( .C1(n13145), .C2(n13177), .A(n13144), .B(n13143), .ZN(
        P3_U3447) );
  MUX2_X1 U15315 ( .A(n13146), .B(P3_REG0_REG_19__SCAN_IN), .S(n15176), .Z(
        n13147) );
  AOI21_X1 U15316 ( .B1(n13148), .B2(n6854), .A(n13147), .ZN(n13149) );
  OAI21_X1 U15317 ( .B1(n13150), .B2(n13177), .A(n13149), .ZN(P3_U3446) );
  MUX2_X1 U15318 ( .A(n13152), .B(n13151), .S(n15177), .Z(n13153) );
  OAI21_X1 U15319 ( .B1(n13154), .B2(n13169), .A(n13153), .ZN(P3_U3444) );
  MUX2_X1 U15320 ( .A(n15298), .B(n13155), .S(n15177), .Z(n13156) );
  OAI21_X1 U15321 ( .B1(n13157), .B2(n13177), .A(n13156), .ZN(P3_U3441) );
  MUX2_X1 U15322 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13158), .S(n15177), .Z(
        n13159) );
  AOI21_X1 U15323 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n13162) );
  INV_X1 U15324 ( .A(n13162), .ZN(P3_U3438) );
  MUX2_X1 U15325 ( .A(n13163), .B(P3_REG0_REG_15__SCAN_IN), .S(n15176), .Z(
        n13167) );
  OAI22_X1 U15326 ( .A1(n13165), .A2(n13177), .B1(n13164), .B2(n13169), .ZN(
        n13166) );
  OR2_X1 U15327 ( .A1(n13167), .A2(n13166), .ZN(P3_U3435) );
  MUX2_X1 U15328 ( .A(n13168), .B(P3_REG0_REG_14__SCAN_IN), .S(n15176), .Z(
        n13173) );
  OAI22_X1 U15329 ( .A1(n13171), .A2(n13177), .B1(n13170), .B2(n13169), .ZN(
        n13172) );
  OR2_X1 U15330 ( .A1(n13173), .A2(n13172), .ZN(P3_U3432) );
  MUX2_X1 U15331 ( .A(n13175), .B(n13174), .S(n15177), .Z(n13176) );
  OAI21_X1 U15332 ( .B1(n13178), .B2(n13177), .A(n13176), .ZN(P3_U3429) );
  NAND2_X1 U15333 ( .A1(n13180), .A2(n13179), .ZN(n13183) );
  OR4_X1 U15334 ( .A1(n13181), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n9056), .ZN(n13182) );
  OAI211_X1 U15335 ( .C1(n13184), .C2(n14525), .A(n13183), .B(n13182), .ZN(
        P3_U3264) );
  INV_X1 U15336 ( .A(n13185), .ZN(n13187) );
  OAI222_X1 U15337 ( .A1(n14525), .A2(n13188), .B1(n11389), .B2(n13187), .C1(
        P3_U3151), .C2(n13186), .ZN(P3_U3266) );
  XNOR2_X1 U15338 ( .A(n13657), .B(n13217), .ZN(n13198) );
  INV_X1 U15339 ( .A(n13198), .ZN(n13200) );
  NAND2_X1 U15340 ( .A1(n13361), .A2(n13574), .ZN(n13199) );
  XNOR2_X1 U15341 ( .A(n13713), .B(n13255), .ZN(n13197) );
  NAND2_X1 U15342 ( .A1(n13362), .A2(n13574), .ZN(n13196) );
  NOR2_X1 U15343 ( .A1(n13329), .A2(n14997), .ZN(n13245) );
  INV_X1 U15344 ( .A(n13189), .ZN(n13190) );
  NAND2_X1 U15345 ( .A1(n13364), .A2(n13202), .ZN(n13192) );
  XNOR2_X1 U15346 ( .A(n13193), .B(n13192), .ZN(n13326) );
  INV_X1 U15347 ( .A(n13192), .ZN(n13194) );
  XNOR2_X1 U15348 ( .A(n13197), .B(n13196), .ZN(n13303) );
  XOR2_X1 U15349 ( .A(n13217), .B(n13583), .Z(n13195) );
  NAND2_X1 U15350 ( .A1(n7511), .A2(n13245), .ZN(n13244) );
  XNOR2_X1 U15351 ( .A(n13198), .B(n13199), .ZN(n13271) );
  NAND2_X1 U15352 ( .A1(n13272), .A2(n13271), .ZN(n13270) );
  XNOR2_X1 U15353 ( .A(n13537), .B(n13217), .ZN(n13203) );
  INV_X1 U15354 ( .A(n13203), .ZN(n13201) );
  XNOR2_X1 U15355 ( .A(n13204), .B(n13201), .ZN(n13314) );
  NAND2_X1 U15356 ( .A1(n13314), .A2(n7529), .ZN(n13313) );
  XNOR2_X1 U15357 ( .A(n13647), .B(n13217), .ZN(n13206) );
  NAND2_X1 U15358 ( .A1(n13359), .A2(n13202), .ZN(n13234) );
  INV_X1 U15359 ( .A(n13206), .ZN(n13207) );
  XNOR2_X1 U15360 ( .A(n13705), .B(n13217), .ZN(n13283) );
  NAND2_X1 U15361 ( .A1(n13358), .A2(n13202), .ZN(n13209) );
  NOR2_X1 U15362 ( .A1(n13283), .A2(n13209), .ZN(n13210) );
  AOI21_X1 U15363 ( .B1(n13283), .B2(n13209), .A(n13210), .ZN(n13292) );
  INV_X1 U15364 ( .A(n13210), .ZN(n13211) );
  XNOR2_X1 U15365 ( .A(n13487), .B(n13255), .ZN(n13335) );
  NOR2_X1 U15366 ( .A1(n13341), .A2(n14997), .ZN(n13212) );
  NAND2_X1 U15367 ( .A1(n13335), .A2(n13212), .ZN(n13218) );
  INV_X1 U15368 ( .A(n13335), .ZN(n13214) );
  INV_X1 U15369 ( .A(n13212), .ZN(n13213) );
  NAND2_X1 U15370 ( .A1(n13214), .A2(n13213), .ZN(n13215) );
  AND2_X1 U15371 ( .A1(n13218), .A2(n13215), .ZN(n13280) );
  NAND2_X1 U15372 ( .A1(n13216), .A2(n13280), .ZN(n13284) );
  XNOR2_X1 U15373 ( .A(n13630), .B(n13217), .ZN(n13220) );
  NAND2_X1 U15374 ( .A1(n13356), .A2(n13202), .ZN(n13221) );
  XNOR2_X1 U15375 ( .A(n13220), .B(n13221), .ZN(n13337) );
  INV_X1 U15376 ( .A(n13220), .ZN(n13222) );
  NAND2_X1 U15377 ( .A1(n13222), .A2(n13221), .ZN(n13223) );
  XNOR2_X1 U15378 ( .A(n13623), .B(n13255), .ZN(n13253) );
  NOR2_X1 U15379 ( .A1(n13343), .A2(n14997), .ZN(n13224) );
  NAND2_X1 U15380 ( .A1(n13253), .A2(n13224), .ZN(n13259) );
  OAI21_X1 U15381 ( .B1(n13253), .B2(n13224), .A(n13259), .ZN(n13226) );
  INV_X1 U15382 ( .A(n13226), .ZN(n13227) );
  NAND2_X1 U15383 ( .A1(n13228), .A2(n14578), .ZN(n13232) );
  NAND2_X1 U15384 ( .A1(n13354), .A2(n13315), .ZN(n13230) );
  NAND2_X1 U15385 ( .A1(n13356), .A2(n13316), .ZN(n13229) );
  NAND2_X1 U15386 ( .A1(n13230), .A2(n13229), .ZN(n13457) );
  AOI22_X1 U15387 ( .A1(n14576), .A2(n13457), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13231) );
  OAI211_X1 U15388 ( .C1(n14581), .C2(n13460), .A(n13232), .B(n13231), .ZN(
        n13233) );
  INV_X1 U15389 ( .A(n13647), .ZN(n13243) );
  NAND2_X1 U15390 ( .A1(n13334), .A2(n13359), .ZN(n13237) );
  NAND2_X1 U15391 ( .A1(n14574), .A2(n13234), .ZN(n13236) );
  MUX2_X1 U15392 ( .A(n13237), .B(n13236), .S(n13235), .Z(n13242) );
  INV_X1 U15393 ( .A(n13238), .ZN(n13522) );
  AOI22_X1 U15394 ( .A1(n13360), .A2(n13316), .B1(n13315), .B2(n13358), .ZN(
        n13517) );
  INV_X1 U15395 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13239) );
  OAI22_X1 U15396 ( .A1(n13517), .A2(n13318), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13239), .ZN(n13240) );
  AOI21_X1 U15397 ( .B1(n13522), .B2(n13322), .A(n13240), .ZN(n13241) );
  OAI211_X1 U15398 ( .C1(n13243), .C2(n13319), .A(n13242), .B(n13241), .ZN(
        P2_U3188) );
  OAI21_X1 U15399 ( .B1(n7511), .B2(n13245), .A(n13244), .ZN(n13246) );
  XNOR2_X1 U15400 ( .A(n13300), .B(n13246), .ZN(n13252) );
  OAI22_X1 U15401 ( .A1(n13273), .A2(n13342), .B1(n13247), .B2(n13340), .ZN(
        n13578) );
  NAND2_X1 U15402 ( .A1(n13578), .A2(n14576), .ZN(n13249) );
  OAI211_X1 U15403 ( .C1(n14581), .C2(n13584), .A(n13249), .B(n13248), .ZN(
        n13250) );
  AOI21_X1 U15404 ( .B1(n13583), .B2(n14578), .A(n13250), .ZN(n13251) );
  OAI21_X1 U15405 ( .B1(n13252), .B2(n13350), .A(n13251), .ZN(P2_U3191) );
  NAND3_X1 U15406 ( .A1(n13253), .A2(n13334), .A3(n13355), .ZN(n13254) );
  NAND2_X1 U15407 ( .A1(n13354), .A2(n13202), .ZN(n13256) );
  XNOR2_X1 U15408 ( .A(n13256), .B(n13255), .ZN(n13257) );
  XNOR2_X1 U15409 ( .A(n13617), .B(n13257), .ZN(n13260) );
  NAND2_X1 U15410 ( .A1(n13258), .A2(n13260), .ZN(n13269) );
  INV_X1 U15411 ( .A(n13259), .ZN(n13261) );
  NOR3_X1 U15412 ( .A1(n13261), .A2(n13260), .A3(n13350), .ZN(n13266) );
  NAND2_X1 U15413 ( .A1(n13617), .A2(n14578), .ZN(n13264) );
  NAND2_X1 U15414 ( .A1(n13353), .A2(n13315), .ZN(n13262) );
  OAI21_X1 U15415 ( .B1(n13343), .B2(n13340), .A(n13262), .ZN(n13441) );
  AOI22_X1 U15416 ( .A1(n14576), .A2(n13441), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13263) );
  OAI211_X1 U15417 ( .C1(n13449), .C2(n14581), .A(n13264), .B(n13263), .ZN(
        n13265) );
  AOI21_X1 U15418 ( .B1(n13267), .B2(n13266), .A(n13265), .ZN(n13268) );
  NAND2_X1 U15419 ( .A1(n13269), .A2(n13268), .ZN(P2_U3192) );
  INV_X1 U15420 ( .A(n13657), .ZN(n13550) );
  OAI211_X1 U15421 ( .C1(n13272), .C2(n13271), .A(n13270), .B(n14574), .ZN(
        n13278) );
  OAI22_X1 U15422 ( .A1(n13274), .A2(n13342), .B1(n13273), .B2(n13340), .ZN(
        n13545) );
  INV_X1 U15423 ( .A(n13545), .ZN(n13275) );
  OAI22_X1 U15424 ( .A1(n13275), .A2(n13318), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15325), .ZN(n13276) );
  AOI21_X1 U15425 ( .B1(n13548), .B2(n13322), .A(n13276), .ZN(n13277) );
  OAI211_X1 U15426 ( .C1(n13550), .C2(n13319), .A(n13278), .B(n13277), .ZN(
        P2_U3195) );
  INV_X1 U15427 ( .A(n13280), .ZN(n13281) );
  AOI21_X1 U15428 ( .B1(n13279), .B2(n13281), .A(n13350), .ZN(n13286) );
  NOR3_X1 U15429 ( .A1(n13283), .A2(n13282), .A3(n13299), .ZN(n13285) );
  OAI21_X1 U15430 ( .B1(n13286), .B2(n13285), .A(n13284), .ZN(n13291) );
  INV_X1 U15431 ( .A(n13287), .ZN(n13485) );
  AOI22_X1 U15432 ( .A1(n13358), .A2(n13316), .B1(n13315), .B2(n13356), .ZN(
        n13491) );
  INV_X1 U15433 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13288) );
  OAI22_X1 U15434 ( .A1(n13318), .A2(n13491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13288), .ZN(n13289) );
  AOI21_X1 U15435 ( .B1(n13485), .B2(n13322), .A(n13289), .ZN(n13290) );
  OAI211_X1 U15436 ( .C1(n13487), .C2(n13319), .A(n13291), .B(n13290), .ZN(
        P2_U3197) );
  OAI211_X1 U15437 ( .C1(n13293), .C2(n13292), .A(n13279), .B(n14574), .ZN(
        n13298) );
  INV_X1 U15438 ( .A(n13294), .ZN(n13508) );
  AOI22_X1 U15439 ( .A1(n13357), .A2(n13315), .B1(n13316), .B2(n13359), .ZN(
        n13504) );
  OAI22_X1 U15440 ( .A1(n13318), .A2(n13504), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13295), .ZN(n13296) );
  AOI21_X1 U15441 ( .B1(n13508), .B2(n13322), .A(n13296), .ZN(n13297) );
  OAI211_X1 U15442 ( .C1(n13705), .C2(n13319), .A(n13298), .B(n13297), .ZN(
        P2_U3201) );
  NOR3_X1 U15443 ( .A1(n13300), .A2(n13329), .A3(n13299), .ZN(n13301) );
  AOI21_X1 U15444 ( .B1(n14574), .B2(n13302), .A(n13301), .ZN(n13312) );
  INV_X1 U15445 ( .A(n13303), .ZN(n13311) );
  NAND2_X1 U15446 ( .A1(n13713), .A2(n14578), .ZN(n13307) );
  NAND2_X1 U15447 ( .A1(n13361), .A2(n13315), .ZN(n13305) );
  NAND2_X1 U15448 ( .A1(n13363), .A2(n13316), .ZN(n13304) );
  NAND2_X1 U15449 ( .A1(n13305), .A2(n13304), .ZN(n13568) );
  AOI22_X1 U15450 ( .A1(n13568), .A2(n14576), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13306) );
  OAI211_X1 U15451 ( .C1(n14581), .C2(n13560), .A(n13307), .B(n13306), .ZN(
        n13308) );
  AOI21_X1 U15452 ( .B1(n13309), .B2(n14574), .A(n13308), .ZN(n13310) );
  OAI21_X1 U15453 ( .B1(n13312), .B2(n13311), .A(n13310), .ZN(P2_U3205) );
  AOI22_X1 U15454 ( .A1(n13314), .A2(n14574), .B1(n13334), .B2(n13360), .ZN(
        n13324) );
  AOI22_X1 U15455 ( .A1(n13361), .A2(n13316), .B1(n13315), .B2(n13359), .ZN(
        n13529) );
  OAI22_X1 U15456 ( .A1(n13529), .A2(n13318), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13317), .ZN(n13321) );
  NOR2_X1 U15457 ( .A1(n13709), .A2(n13319), .ZN(n13320) );
  AOI211_X1 U15458 ( .C1(n13322), .C2(n13538), .A(n13321), .B(n13320), .ZN(
        n13323) );
  OAI21_X1 U15459 ( .B1(n13325), .B2(n13324), .A(n13323), .ZN(P2_U3207) );
  XNOR2_X1 U15460 ( .A(n13327), .B(n13326), .ZN(n13333) );
  OAI22_X1 U15461 ( .A1(n13329), .A2(n13342), .B1(n13328), .B2(n13340), .ZN(
        n13592) );
  NAND2_X1 U15462 ( .A1(n13592), .A2(n14576), .ZN(n13330) );
  NAND2_X1 U15463 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14928)
         );
  OAI211_X1 U15464 ( .C1(n14581), .C2(n13596), .A(n13330), .B(n14928), .ZN(
        n13331) );
  AOI21_X1 U15465 ( .B1(n13674), .B2(n14578), .A(n13331), .ZN(n13332) );
  OAI21_X1 U15466 ( .B1(n13333), .B2(n13350), .A(n13332), .ZN(P2_U3210) );
  NAND3_X1 U15467 ( .A1(n13335), .A2(n13334), .A3(n13357), .ZN(n13336) );
  OAI21_X1 U15468 ( .B1(n13284), .B2(n13350), .A(n13336), .ZN(n13339) );
  INV_X1 U15469 ( .A(n13337), .ZN(n13338) );
  NAND2_X1 U15470 ( .A1(n13339), .A2(n13338), .ZN(n13349) );
  NOR2_X1 U15471 ( .A1(n13341), .A2(n13340), .ZN(n13345) );
  NOR2_X1 U15472 ( .A1(n13343), .A2(n13342), .ZN(n13344) );
  OR2_X1 U15473 ( .A1(n13345), .A2(n13344), .ZN(n13470) );
  AOI22_X1 U15474 ( .A1(n14576), .A2(n13470), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13346) );
  OAI21_X1 U15475 ( .B1(n13473), .B2(n14581), .A(n13346), .ZN(n13347) );
  AOI21_X1 U15476 ( .B1(n13630), .B2(n14578), .A(n13347), .ZN(n13348) );
  OAI211_X1 U15477 ( .C1(n13351), .C2(n13350), .A(n13349), .B(n13348), .ZN(
        P2_U3212) );
  MUX2_X1 U15478 ( .A(n13421), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13379), .Z(
        P2_U3562) );
  MUX2_X1 U15479 ( .A(n13352), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13379), .Z(
        P2_U3561) );
  MUX2_X1 U15480 ( .A(n13353), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13379), .Z(
        P2_U3560) );
  MUX2_X1 U15481 ( .A(n13354), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13379), .Z(
        P2_U3559) );
  MUX2_X1 U15482 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13355), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15483 ( .A(n13356), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13379), .Z(
        P2_U3557) );
  MUX2_X1 U15484 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13357), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15485 ( .A(n13358), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13379), .Z(
        P2_U3555) );
  MUX2_X1 U15486 ( .A(n13359), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13379), .Z(
        P2_U3554) );
  MUX2_X1 U15487 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13360), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15488 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13361), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15489 ( .A(n13362), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13379), .Z(
        P2_U3551) );
  MUX2_X1 U15490 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13363), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15491 ( .A(n13364), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13379), .Z(
        P2_U3549) );
  MUX2_X1 U15492 ( .A(n13365), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13379), .Z(
        P2_U3548) );
  MUX2_X1 U15493 ( .A(n13366), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13379), .Z(
        P2_U3547) );
  MUX2_X1 U15494 ( .A(n13367), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13379), .Z(
        P2_U3546) );
  MUX2_X1 U15495 ( .A(n13368), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13379), .Z(
        P2_U3545) );
  MUX2_X1 U15496 ( .A(n13369), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13379), .Z(
        P2_U3544) );
  MUX2_X1 U15497 ( .A(n13370), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13379), .Z(
        P2_U3543) );
  MUX2_X1 U15498 ( .A(n13371), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13379), .Z(
        P2_U3542) );
  MUX2_X1 U15499 ( .A(n13372), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13379), .Z(
        P2_U3541) );
  MUX2_X1 U15500 ( .A(n13373), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13379), .Z(
        P2_U3540) );
  MUX2_X1 U15501 ( .A(n13374), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13379), .Z(
        P2_U3539) );
  MUX2_X1 U15502 ( .A(n13375), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13379), .Z(
        P2_U3538) );
  MUX2_X1 U15503 ( .A(n13376), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13379), .Z(
        P2_U3537) );
  MUX2_X1 U15504 ( .A(n13377), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13379), .Z(
        P2_U3536) );
  MUX2_X1 U15505 ( .A(n13378), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13379), .Z(
        P2_U3535) );
  MUX2_X1 U15506 ( .A(n13380), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13379), .Z(
        P2_U3534) );
  MUX2_X1 U15507 ( .A(n13381), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13379), .Z(
        P2_U3533) );
  MUX2_X1 U15508 ( .A(n9903), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13379), .Z(
        P2_U3532) );
  MUX2_X1 U15509 ( .A(n8750), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13379), .Z(
        P2_U3531) );
  INV_X1 U15510 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n15386) );
  OAI22_X1 U15511 ( .A1(n14926), .A2(n13382), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15386), .ZN(n13383) );
  AOI21_X1 U15512 ( .B1(n14760), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n13383), .ZN(
        n13392) );
  OAI211_X1 U15513 ( .C1(n13386), .C2(n13385), .A(n14915), .B(n13384), .ZN(
        n13391) );
  OAI211_X1 U15514 ( .C1(n13389), .C2(n13388), .A(n14922), .B(n13387), .ZN(
        n13390) );
  NAND3_X1 U15515 ( .A1(n13392), .A2(n13391), .A3(n13390), .ZN(P2_U3216) );
  NAND2_X1 U15516 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n13393) );
  OAI21_X1 U15517 ( .B1(n14926), .B2(n13394), .A(n13393), .ZN(n13395) );
  AOI21_X1 U15518 ( .B1(n14760), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13395), .ZN(
        n13404) );
  OAI211_X1 U15519 ( .C1(n13398), .C2(n13397), .A(n14922), .B(n13396), .ZN(
        n13403) );
  OAI211_X1 U15520 ( .C1(n13401), .C2(n13400), .A(n14915), .B(n13399), .ZN(
        n13402) );
  NAND3_X1 U15521 ( .A1(n13404), .A2(n13403), .A3(n13402), .ZN(P2_U3217) );
  OAI21_X1 U15522 ( .B1(n14926), .B2(n13406), .A(n13405), .ZN(n13407) );
  AOI21_X1 U15523 ( .B1(n14760), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n13407), .ZN(
        n13416) );
  OAI211_X1 U15524 ( .C1(n13410), .C2(n13409), .A(n14915), .B(n13408), .ZN(
        n13415) );
  OAI211_X1 U15525 ( .C1(n13413), .C2(n13412), .A(n14922), .B(n13411), .ZN(
        n13414) );
  NAND3_X1 U15526 ( .A1(n13416), .A2(n13415), .A3(n13414), .ZN(P2_U3221) );
  NAND2_X1 U15527 ( .A1(n7203), .A2(n13424), .ZN(n13417) );
  XNOR2_X1 U15528 ( .A(n13417), .B(n13694), .ZN(n13609) );
  NAND2_X1 U15529 ( .A1(n13609), .A2(n13418), .ZN(n13423) );
  INV_X1 U15530 ( .A(n13419), .ZN(n13420) );
  AND2_X1 U15531 ( .A1(n13421), .A2(n13420), .ZN(n13608) );
  INV_X1 U15532 ( .A(n13608), .ZN(n13612) );
  NOR2_X1 U15533 ( .A1(n13612), .A2(n10410), .ZN(n13428) );
  AOI21_X1 U15534 ( .B1(n14957), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13428), 
        .ZN(n13422) );
  OAI211_X1 U15535 ( .C1(n13694), .C2(n14951), .A(n13423), .B(n13422), .ZN(
        P2_U3234) );
  NAND2_X1 U15536 ( .A1(n13426), .A2(n14997), .ZN(n13613) );
  NOR2_X1 U15537 ( .A1(n7203), .A2(n14951), .ZN(n13427) );
  AOI211_X1 U15538 ( .C1(n14957), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13428), 
        .B(n13427), .ZN(n13429) );
  OAI21_X1 U15539 ( .B1(n13613), .B2(n13563), .A(n13429), .ZN(P2_U3235) );
  INV_X1 U15540 ( .A(n13430), .ZN(n13438) );
  NOR2_X1 U15541 ( .A1(n6921), .A2(n14951), .ZN(n13435) );
  INV_X1 U15542 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13433) );
  OAI22_X1 U15543 ( .A1(n13512), .A2(n13433), .B1(n13432), .B2(n15200), .ZN(
        n13434) );
  AOI211_X1 U15544 ( .C1(n13436), .C2(n15195), .A(n13435), .B(n13434), .ZN(
        n13437) );
  INV_X1 U15545 ( .A(n13439), .ZN(n13440) );
  AOI21_X1 U15546 ( .B1(n13440), .B2(n13446), .A(n13530), .ZN(n13443) );
  AOI21_X1 U15547 ( .B1(n13443), .B2(n13442), .A(n13441), .ZN(n13619) );
  OAI21_X1 U15548 ( .B1(n13446), .B2(n13445), .A(n13444), .ZN(n13620) );
  INV_X1 U15549 ( .A(n13620), .ZN(n13454) );
  AOI21_X1 U15550 ( .B1(n13617), .B2(n13459), .A(n13202), .ZN(n13448) );
  AND2_X1 U15551 ( .A1(n13448), .A2(n13447), .ZN(n13616) );
  NAND2_X1 U15552 ( .A1(n13616), .A2(n15195), .ZN(n13452) );
  INV_X1 U15553 ( .A(n13449), .ZN(n13450) );
  AOI22_X1 U15554 ( .A1(n14957), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n13450), 
        .B2(n14948), .ZN(n13451) );
  OAI211_X1 U15555 ( .C1(n7202), .C2(n14951), .A(n13452), .B(n13451), .ZN(
        n13453) );
  AOI21_X1 U15556 ( .B1(n13454), .B2(n15196), .A(n13453), .ZN(n13455) );
  OAI21_X1 U15557 ( .B1(n13619), .B2(n10410), .A(n13455), .ZN(P2_U3237) );
  XNOR2_X1 U15558 ( .A(n13456), .B(n13466), .ZN(n13458) );
  AOI21_X1 U15559 ( .B1(n13458), .B2(n14992), .A(n13457), .ZN(n13628) );
  OAI211_X1 U15560 ( .C1(n13623), .C2(n13472), .A(n14997), .B(n13459), .ZN(
        n13622) );
  INV_X1 U15561 ( .A(n13622), .ZN(n13464) );
  INV_X1 U15562 ( .A(n13460), .ZN(n13461) );
  AOI22_X1 U15563 ( .A1(n14957), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13461), 
        .B2(n14948), .ZN(n13462) );
  OAI21_X1 U15564 ( .B1(n13623), .B2(n14951), .A(n13462), .ZN(n13463) );
  AOI21_X1 U15565 ( .B1(n13464), .B2(n15195), .A(n13463), .ZN(n13468) );
  NAND2_X1 U15566 ( .A1(n13466), .A2(n13465), .ZN(n13621) );
  NAND3_X1 U15567 ( .A1(n13625), .A2(n13621), .A3(n15196), .ZN(n13467) );
  OAI211_X1 U15568 ( .C1(n13628), .C2(n10410), .A(n13468), .B(n13467), .ZN(
        P2_U3238) );
  XOR2_X1 U15569 ( .A(n13469), .B(n13477), .Z(n13471) );
  AOI21_X1 U15570 ( .B1(n13471), .B2(n14992), .A(n13470), .ZN(n13632) );
  AOI211_X1 U15571 ( .C1(n13630), .C2(n13484), .A(n13202), .B(n13472), .ZN(
        n13629) );
  INV_X1 U15572 ( .A(n13630), .ZN(n13476) );
  INV_X1 U15573 ( .A(n13473), .ZN(n13474) );
  AOI22_X1 U15574 ( .A1(n14957), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13474), 
        .B2(n14948), .ZN(n13475) );
  OAI21_X1 U15575 ( .B1(n13476), .B2(n14951), .A(n13475), .ZN(n13480) );
  XNOR2_X1 U15576 ( .A(n13478), .B(n13477), .ZN(n13633) );
  NOR2_X1 U15577 ( .A1(n13633), .A2(n13604), .ZN(n13479) );
  AOI211_X1 U15578 ( .C1(n13629), .C2(n15195), .A(n13480), .B(n13479), .ZN(
        n13481) );
  OAI21_X1 U15579 ( .B1(n14957), .B2(n13632), .A(n13481), .ZN(P2_U3239) );
  XOR2_X1 U15580 ( .A(n13482), .B(n13489), .Z(n13638) );
  OR2_X1 U15581 ( .A1(n13487), .A2(n13506), .ZN(n13483) );
  AND3_X1 U15582 ( .A1(n13484), .A2(n13483), .A3(n14997), .ZN(n13634) );
  AOI22_X1 U15583 ( .A1(n14957), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13485), 
        .B2(n14948), .ZN(n13486) );
  OAI21_X1 U15584 ( .B1(n13487), .B2(n14951), .A(n13486), .ZN(n13495) );
  OAI21_X1 U15585 ( .B1(n13490), .B2(n13489), .A(n13488), .ZN(n13493) );
  INV_X1 U15586 ( .A(n13491), .ZN(n13492) );
  AOI21_X1 U15587 ( .B1(n13493), .B2(n14992), .A(n13492), .ZN(n13637) );
  NOR2_X1 U15588 ( .A1(n13637), .A2(n10410), .ZN(n13494) );
  AOI211_X1 U15589 ( .C1(n13634), .C2(n15195), .A(n13495), .B(n13494), .ZN(
        n13496) );
  OAI21_X1 U15590 ( .B1(n13638), .B2(n13604), .A(n13496), .ZN(P2_U3240) );
  XOR2_X1 U15591 ( .A(n13497), .B(n13499), .Z(n13642) );
  INV_X1 U15592 ( .A(n13642), .ZN(n13514) );
  INV_X1 U15593 ( .A(n13499), .ZN(n13501) );
  NAND3_X1 U15594 ( .A1(n13498), .A2(n13501), .A3(n13500), .ZN(n13502) );
  AND2_X1 U15595 ( .A1(n13503), .A2(n13502), .ZN(n13505) );
  OAI21_X1 U15596 ( .B1(n13505), .B2(n13530), .A(n13504), .ZN(n13640) );
  NOR2_X1 U15597 ( .A1(n13521), .A2(n13705), .ZN(n13507) );
  NOR2_X1 U15598 ( .A1(n13639), .A2(n13563), .ZN(n13511) );
  AOI22_X1 U15599 ( .A1(n14957), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13508), 
        .B2(n14948), .ZN(n13509) );
  OAI21_X1 U15600 ( .B1(n13705), .B2(n14951), .A(n13509), .ZN(n13510) );
  AOI211_X1 U15601 ( .C1(n13640), .C2(n13512), .A(n13511), .B(n13510), .ZN(
        n13513) );
  OAI21_X1 U15602 ( .B1(n13604), .B2(n13514), .A(n13513), .ZN(P2_U3241) );
  XOR2_X1 U15603 ( .A(n13515), .B(n13516), .Z(n13650) );
  OAI21_X1 U15604 ( .B1(n13516), .B2(n6706), .A(n13498), .ZN(n13519) );
  INV_X1 U15605 ( .A(n13517), .ZN(n13518) );
  AOI21_X1 U15606 ( .B1(n13519), .B2(n14992), .A(n13518), .ZN(n13649) );
  INV_X1 U15607 ( .A(n13649), .ZN(n13526) );
  AND2_X1 U15608 ( .A1(n13647), .A2(n13534), .ZN(n13520) );
  OR3_X1 U15609 ( .A1(n13521), .A2(n13520), .A3(n13202), .ZN(n13645) );
  AOI22_X1 U15610 ( .A1(n14957), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13522), 
        .B2(n14948), .ZN(n13524) );
  NAND2_X1 U15611 ( .A1(n13647), .A2(n14937), .ZN(n13523) );
  OAI211_X1 U15612 ( .C1(n13645), .C2(n13563), .A(n13524), .B(n13523), .ZN(
        n13525) );
  AOI21_X1 U15613 ( .B1(n13526), .B2(n13512), .A(n13525), .ZN(n13527) );
  OAI21_X1 U15614 ( .B1(n13604), .B2(n13650), .A(n13527), .ZN(P2_U3242) );
  XNOR2_X1 U15615 ( .A(n13528), .B(n13532), .ZN(n13531) );
  OAI21_X1 U15616 ( .B1(n13531), .B2(n13530), .A(n13529), .ZN(n13651) );
  INV_X1 U15617 ( .A(n13651), .ZN(n13543) );
  XOR2_X1 U15618 ( .A(n13533), .B(n13532), .Z(n13653) );
  INV_X1 U15619 ( .A(n13547), .ZN(n13536) );
  INV_X1 U15620 ( .A(n13534), .ZN(n13535) );
  AOI211_X1 U15621 ( .C1(n13537), .C2(n13536), .A(n13574), .B(n13535), .ZN(
        n13652) );
  NAND2_X1 U15622 ( .A1(n13652), .A2(n15195), .ZN(n13540) );
  AOI22_X1 U15623 ( .A1(n13538), .A2(n14948), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n10410), .ZN(n13539) );
  OAI211_X1 U15624 ( .C1(n13709), .C2(n14951), .A(n13540), .B(n13539), .ZN(
        n13541) );
  AOI21_X1 U15625 ( .B1(n15196), .B2(n13653), .A(n13541), .ZN(n13542) );
  OAI21_X1 U15626 ( .B1(n14957), .B2(n13543), .A(n13542), .ZN(P2_U3243) );
  XNOR2_X1 U15627 ( .A(n13544), .B(n13551), .ZN(n13546) );
  AOI21_X1 U15628 ( .B1(n13546), .B2(n14992), .A(n13545), .ZN(n13658) );
  AOI211_X1 U15629 ( .C1(n13657), .C2(n13557), .A(n13202), .B(n13547), .ZN(
        n13656) );
  AOI22_X1 U15630 ( .A1(n13548), .A2(n14948), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14957), .ZN(n13549) );
  OAI21_X1 U15631 ( .B1(n13550), .B2(n14951), .A(n13549), .ZN(n13554) );
  XNOR2_X1 U15632 ( .A(n13552), .B(n13551), .ZN(n13660) );
  NOR2_X1 U15633 ( .A1(n13660), .A2(n13604), .ZN(n13553) );
  AOI211_X1 U15634 ( .C1(n13656), .C2(n15195), .A(n13554), .B(n13553), .ZN(
        n13555) );
  OAI21_X1 U15635 ( .B1(n14957), .B2(n13658), .A(n13555), .ZN(P2_U3244) );
  XNOR2_X1 U15636 ( .A(n13556), .B(n13564), .ZN(n13661) );
  AOI21_X1 U15637 ( .B1(n13573), .B2(n13713), .A(n13202), .ZN(n13558) );
  NAND2_X1 U15638 ( .A1(n13558), .A2(n13557), .ZN(n13662) );
  NAND2_X1 U15639 ( .A1(n14957), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13559) );
  OAI21_X1 U15640 ( .B1(n13560), .B2(n15200), .A(n13559), .ZN(n13561) );
  AOI21_X1 U15641 ( .B1(n13713), .B2(n14937), .A(n13561), .ZN(n13562) );
  OAI21_X1 U15642 ( .B1(n13662), .B2(n13563), .A(n13562), .ZN(n13571) );
  NAND2_X1 U15643 ( .A1(n13565), .A2(n13564), .ZN(n13566) );
  NAND2_X1 U15644 ( .A1(n13567), .A2(n13566), .ZN(n13569) );
  AOI21_X1 U15645 ( .B1(n13569), .B2(n14992), .A(n13568), .ZN(n13663) );
  NOR2_X1 U15646 ( .A1(n13663), .A2(n10410), .ZN(n13570) );
  AOI211_X1 U15647 ( .C1(n15196), .C2(n13661), .A(n13571), .B(n13570), .ZN(
        n13572) );
  INV_X1 U15648 ( .A(n13572), .ZN(P2_U3245) );
  AOI211_X1 U15649 ( .C1(n13583), .C2(n13594), .A(n13574), .B(n6914), .ZN(
        n13668) );
  XNOR2_X1 U15650 ( .A(n13575), .B(n13576), .ZN(n13582) );
  XNOR2_X1 U15651 ( .A(n13577), .B(n13576), .ZN(n13579) );
  AOI21_X1 U15652 ( .B1(n13579), .B2(n14992), .A(n13578), .ZN(n13580) );
  OAI21_X1 U15653 ( .B1(n13582), .B2(n14974), .A(n13580), .ZN(n13667) );
  AOI21_X1 U15654 ( .B1(n13668), .B2(n13581), .A(n13667), .ZN(n13590) );
  INV_X1 U15655 ( .A(n13582), .ZN(n13669) );
  INV_X1 U15656 ( .A(n13584), .ZN(n13585) );
  AOI22_X1 U15657 ( .A1(n14957), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13585), 
        .B2(n14948), .ZN(n13586) );
  OAI21_X1 U15658 ( .B1(n7205), .B2(n14951), .A(n13586), .ZN(n13587) );
  AOI21_X1 U15659 ( .B1(n13669), .B2(n13588), .A(n13587), .ZN(n13589) );
  OAI21_X1 U15660 ( .B1(n13590), .B2(n10410), .A(n13589), .ZN(P2_U3246) );
  XNOR2_X1 U15661 ( .A(n13591), .B(n13603), .ZN(n13593) );
  AOI21_X1 U15662 ( .B1(n13593), .B2(n14992), .A(n13592), .ZN(n13675) );
  AOI211_X1 U15663 ( .C1(n13674), .C2(n13595), .A(n13202), .B(n7206), .ZN(
        n13673) );
  INV_X1 U15664 ( .A(n13674), .ZN(n13599) );
  INV_X1 U15665 ( .A(n13596), .ZN(n13597) );
  AOI22_X1 U15666 ( .A1(n14957), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13597), 
        .B2(n14948), .ZN(n13598) );
  OAI21_X1 U15667 ( .B1(n13599), .B2(n14951), .A(n13598), .ZN(n13606) );
  INV_X1 U15668 ( .A(n13600), .ZN(n13601) );
  AOI21_X1 U15669 ( .B1(n13603), .B2(n13602), .A(n13601), .ZN(n13677) );
  NOR2_X1 U15670 ( .A1(n13677), .A2(n13604), .ZN(n13605) );
  AOI211_X1 U15671 ( .C1(n13673), .C2(n15195), .A(n13606), .B(n13605), .ZN(
        n13607) );
  OAI21_X1 U15672 ( .B1(n14957), .B2(n13675), .A(n13607), .ZN(P2_U3247) );
  INV_X1 U15673 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13610) );
  AOI21_X1 U15674 ( .B1(n13609), .B2(n14997), .A(n13608), .ZN(n13691) );
  MUX2_X1 U15675 ( .A(n13610), .B(n13691), .S(n15037), .Z(n13611) );
  OAI21_X1 U15676 ( .B1(n13694), .B2(n13672), .A(n13611), .ZN(P2_U3530) );
  INV_X1 U15677 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13614) );
  MUX2_X1 U15678 ( .A(n13614), .B(n13695), .S(n15037), .Z(n13615) );
  OAI21_X1 U15679 ( .B1(n7203), .B2(n13672), .A(n13615), .ZN(P2_U3529) );
  AOI21_X1 U15680 ( .B1(n14597), .B2(n13617), .A(n13616), .ZN(n13618) );
  MUX2_X1 U15681 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13698), .S(n15037), .Z(
        P2_U3527) );
  AND2_X1 U15682 ( .A1(n13621), .A2(n15024), .ZN(n13626) );
  OAI21_X1 U15683 ( .B1(n13623), .B2(n15018), .A(n13622), .ZN(n13624) );
  AOI21_X1 U15684 ( .B1(n13626), .B2(n13625), .A(n13624), .ZN(n13627) );
  NAND2_X1 U15685 ( .A1(n13628), .A2(n13627), .ZN(n13699) );
  MUX2_X1 U15686 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13699), .S(n15037), .Z(
        P2_U3526) );
  AOI21_X1 U15687 ( .B1(n14597), .B2(n13630), .A(n13629), .ZN(n13631) );
  OAI211_X1 U15688 ( .C1(n13682), .C2(n13633), .A(n13632), .B(n13631), .ZN(
        n13700) );
  MUX2_X1 U15689 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13700), .S(n15037), .Z(
        P2_U3525) );
  AOI21_X1 U15690 ( .B1(n14597), .B2(n13635), .A(n13634), .ZN(n13636) );
  OAI211_X1 U15691 ( .C1(n13638), .C2(n13682), .A(n13637), .B(n13636), .ZN(
        n13701) );
  MUX2_X1 U15692 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13701), .S(n15037), .Z(
        P2_U3524) );
  INV_X1 U15693 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13643) );
  INV_X1 U15694 ( .A(n13639), .ZN(n13641) );
  AOI211_X1 U15695 ( .C1(n13642), .C2(n15024), .A(n13641), .B(n13640), .ZN(
        n13702) );
  MUX2_X1 U15696 ( .A(n13643), .B(n13702), .S(n15037), .Z(n13644) );
  OAI21_X1 U15697 ( .B1(n13705), .B2(n13672), .A(n13644), .ZN(P2_U3523) );
  INV_X1 U15698 ( .A(n13645), .ZN(n13646) );
  AOI21_X1 U15699 ( .B1(n14597), .B2(n13647), .A(n13646), .ZN(n13648) );
  OAI211_X1 U15700 ( .C1(n13650), .C2(n13682), .A(n13649), .B(n13648), .ZN(
        n13706) );
  MUX2_X1 U15701 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13706), .S(n15037), .Z(
        P2_U3522) );
  INV_X1 U15702 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13654) );
  AOI211_X1 U15703 ( .C1(n15024), .C2(n13653), .A(n13652), .B(n13651), .ZN(
        n13707) );
  MUX2_X1 U15704 ( .A(n13654), .B(n13707), .S(n15037), .Z(n13655) );
  OAI21_X1 U15705 ( .B1(n13709), .B2(n13672), .A(n13655), .ZN(P2_U3521) );
  AOI21_X1 U15706 ( .B1(n14597), .B2(n13657), .A(n13656), .ZN(n13659) );
  OAI211_X1 U15707 ( .C1(n13682), .C2(n13660), .A(n13659), .B(n13658), .ZN(
        n13710) );
  MUX2_X1 U15708 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13710), .S(n15037), .Z(
        P2_U3520) );
  NAND2_X1 U15709 ( .A1(n13661), .A2(n15024), .ZN(n13664) );
  NAND3_X1 U15710 ( .A1(n13664), .A2(n13663), .A3(n13662), .ZN(n13711) );
  MUX2_X1 U15711 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13711), .S(n15037), .Z(
        n13665) );
  AOI21_X1 U15712 ( .B1(n8743), .B2(n13713), .A(n13665), .ZN(n13666) );
  INV_X1 U15713 ( .A(n13666), .ZN(P2_U3519) );
  INV_X1 U15714 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13670) );
  INV_X1 U15715 ( .A(n14970), .ZN(n15006) );
  AOI211_X1 U15716 ( .C1(n13669), .C2(n15006), .A(n13668), .B(n13667), .ZN(
        n13715) );
  MUX2_X1 U15717 ( .A(n13670), .B(n13715), .S(n15037), .Z(n13671) );
  OAI21_X1 U15718 ( .B1(n7205), .B2(n13672), .A(n13671), .ZN(P2_U3518) );
  AOI21_X1 U15719 ( .B1(n14597), .B2(n13674), .A(n13673), .ZN(n13676) );
  OAI211_X1 U15720 ( .C1(n13682), .C2(n13677), .A(n13676), .B(n13675), .ZN(
        n13719) );
  MUX2_X1 U15721 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13719), .S(n15037), .Z(
        P2_U3517) );
  AOI21_X1 U15722 ( .B1(n14597), .B2(n13679), .A(n13678), .ZN(n13680) );
  OAI211_X1 U15723 ( .C1(n13683), .C2(n13682), .A(n13681), .B(n13680), .ZN(
        n13720) );
  MUX2_X1 U15724 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13720), .S(n15037), .Z(
        P2_U3516) );
  NAND3_X1 U15725 ( .A1(n13685), .A2(n15024), .A3(n13684), .ZN(n13690) );
  AOI21_X1 U15726 ( .B1(n14597), .B2(n13687), .A(n13686), .ZN(n13688) );
  NAND3_X1 U15727 ( .A1(n13690), .A2(n13689), .A3(n13688), .ZN(n13721) );
  MUX2_X1 U15728 ( .A(n13721), .B(P2_REG1_REG_16__SCAN_IN), .S(n15035), .Z(
        P2_U3515) );
  INV_X1 U15729 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13692) );
  MUX2_X1 U15730 ( .A(n13692), .B(n13691), .S(n15027), .Z(n13693) );
  OAI21_X1 U15731 ( .B1(n13694), .B2(n13718), .A(n13693), .ZN(P2_U3498) );
  MUX2_X1 U15732 ( .A(n13696), .B(n13695), .S(n15027), .Z(n13697) );
  OAI21_X1 U15733 ( .B1(n7203), .B2(n13718), .A(n13697), .ZN(P2_U3497) );
  MUX2_X1 U15734 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13698), .S(n15027), .Z(
        P2_U3495) );
  MUX2_X1 U15735 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13699), .S(n15027), .Z(
        P2_U3494) );
  MUX2_X1 U15736 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13700), .S(n15027), .Z(
        P2_U3493) );
  MUX2_X1 U15737 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13701), .S(n15027), .Z(
        P2_U3492) );
  MUX2_X1 U15738 ( .A(n13703), .B(n13702), .S(n15027), .Z(n13704) );
  OAI21_X1 U15739 ( .B1(n13705), .B2(n13718), .A(n13704), .ZN(P2_U3491) );
  MUX2_X1 U15740 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13706), .S(n15027), .Z(
        P2_U3490) );
  MUX2_X1 U15741 ( .A(n15354), .B(n13707), .S(n15027), .Z(n13708) );
  OAI21_X1 U15742 ( .B1(n13709), .B2(n13718), .A(n13708), .ZN(P2_U3489) );
  MUX2_X1 U15743 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13710), .S(n15027), .Z(
        P2_U3488) );
  MUX2_X1 U15744 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13711), .S(n15027), .Z(
        n13712) );
  AOI21_X1 U15745 ( .B1(n9638), .B2(n13713), .A(n13712), .ZN(n13714) );
  INV_X1 U15746 ( .A(n13714), .ZN(P2_U3487) );
  INV_X1 U15747 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13716) );
  MUX2_X1 U15748 ( .A(n13716), .B(n13715), .S(n15027), .Z(n13717) );
  OAI21_X1 U15749 ( .B1(n7205), .B2(n13718), .A(n13717), .ZN(P2_U3486) );
  MUX2_X1 U15750 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13719), .S(n15027), .Z(
        P2_U3484) );
  MUX2_X1 U15751 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13720), .S(n15027), .Z(
        P2_U3481) );
  MUX2_X1 U15752 ( .A(n13721), .B(P2_REG0_REG_16__SCAN_IN), .S(n15025), .Z(
        P2_U3478) );
  INV_X1 U15753 ( .A(n13722), .ZN(n14397) );
  INV_X1 U15754 ( .A(n13723), .ZN(n13725) );
  NOR4_X1 U15755 ( .A1(n13725), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13724), .A4(
        P2_U3088), .ZN(n13726) );
  AOI21_X1 U15756 ( .B1(n13735), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13726), 
        .ZN(n13727) );
  OAI21_X1 U15757 ( .B1(n14397), .B2(n13741), .A(n13727), .ZN(P2_U3296) );
  INV_X1 U15758 ( .A(n13728), .ZN(n14399) );
  OAI222_X1 U15759 ( .A1(n13739), .A2(n13732), .B1(P2_U3088), .B2(n13730), 
        .C1(n13729), .C2(n14399), .ZN(P2_U3298) );
  INV_X1 U15760 ( .A(n13733), .ZN(n14402) );
  AOI21_X1 U15761 ( .B1(n13735), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13734), 
        .ZN(n13736) );
  OAI21_X1 U15762 ( .B1(n14402), .B2(n13741), .A(n13736), .ZN(P2_U3299) );
  INV_X1 U15763 ( .A(n14406), .ZN(n13737) );
  OAI222_X1 U15764 ( .A1(n13739), .A2(n13738), .B1(n13741), .B2(n13737), .C1(
        n8659), .C2(P2_U3088), .ZN(P2_U3300) );
  OAI222_X1 U15765 ( .A1(P2_U3088), .A2(n13742), .B1(n13741), .B2(n14412), 
        .C1(n13740), .C2(n13739), .ZN(P2_U3301) );
  INV_X1 U15766 ( .A(n13743), .ZN(n13744) );
  MUX2_X1 U15767 ( .A(n13744), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15768 ( .A(n13746), .B(n13745), .Z(n13752) );
  NAND2_X1 U15769 ( .A1(n13897), .A2(n14234), .ZN(n13748) );
  NAND2_X1 U15770 ( .A1(n13895), .A2(n14236), .ZN(n13747) );
  NAND2_X1 U15771 ( .A1(n13748), .A2(n13747), .ZN(n14164) );
  AOI22_X1 U15772 ( .A1(n14164), .A2(n14615), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13749) );
  OAI21_X1 U15773 ( .B1(n14165), .B2(n14622), .A(n13749), .ZN(n13750) );
  AOI21_X1 U15774 ( .B1(n6770), .B2(n14618), .A(n13750), .ZN(n13751) );
  OAI21_X1 U15775 ( .B1(n13752), .B2(n13889), .A(n13751), .ZN(P1_U3216) );
  AOI21_X1 U15776 ( .B1(n13754), .B2(n13753), .A(n13889), .ZN(n13756) );
  NAND2_X1 U15777 ( .A1(n13756), .A2(n13755), .ZN(n13762) );
  NAND2_X1 U15778 ( .A1(n13899), .A2(n14236), .ZN(n13758) );
  NAND2_X1 U15779 ( .A1(n13900), .A2(n14234), .ZN(n13757) );
  NAND2_X1 U15780 ( .A1(n13758), .A2(n13757), .ZN(n14324) );
  NOR2_X1 U15781 ( .A1(n13759), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14043) );
  NOR2_X1 U15782 ( .A1(n14622), .A2(n14220), .ZN(n13760) );
  AOI211_X1 U15783 ( .C1(n14615), .C2(n14324), .A(n14043), .B(n13760), .ZN(
        n13761) );
  OAI211_X1 U15784 ( .C1(n7067), .C2(n13868), .A(n13762), .B(n13761), .ZN(
        P1_U3219) );
  NOR2_X1 U15785 ( .A1(n13764), .A2(n13763), .ZN(n13766) );
  OAI21_X1 U15786 ( .B1(n13766), .B2(n13765), .A(n14613), .ZN(n13773) );
  INV_X1 U15787 ( .A(n13884), .ZN(n13768) );
  AOI22_X1 U15788 ( .A1(n13768), .A2(n6758), .B1(n13767), .B2(n13915), .ZN(
        n13772) );
  AOI22_X1 U15789 ( .A1(n13770), .A2(n14618), .B1(n13769), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n13771) );
  NAND3_X1 U15790 ( .A1(n13773), .A2(n13772), .A3(n13771), .ZN(P1_U3222) );
  INV_X1 U15791 ( .A(n13774), .ZN(n13775) );
  AOI21_X1 U15792 ( .B1(n13777), .B2(n13776), .A(n13775), .ZN(n13783) );
  NAND2_X1 U15793 ( .A1(n13897), .A2(n14236), .ZN(n13779) );
  NAND2_X1 U15794 ( .A1(n13899), .A2(n14234), .ZN(n13778) );
  NAND2_X1 U15795 ( .A1(n13779), .A2(n13778), .ZN(n14196) );
  AOI22_X1 U15796 ( .A1(n14196), .A2(n14615), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13780) );
  OAI21_X1 U15797 ( .B1(n14197), .B2(n14622), .A(n13780), .ZN(n13781) );
  AOI21_X1 U15798 ( .B1(n14384), .B2(n14618), .A(n13781), .ZN(n13782) );
  OAI21_X1 U15799 ( .B1(n13783), .B2(n13889), .A(n13782), .ZN(P1_U3223) );
  XOR2_X1 U15800 ( .A(n13785), .B(n13784), .Z(n13791) );
  NAND2_X1 U15801 ( .A1(n13895), .A2(n14234), .ZN(n13787) );
  NAND2_X1 U15802 ( .A1(n14093), .A2(n14236), .ZN(n13786) );
  NAND2_X1 U15803 ( .A1(n13787), .A2(n13786), .ZN(n14129) );
  AOI22_X1 U15804 ( .A1(n14615), .A2(n14129), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13788) );
  OAI21_X1 U15805 ( .B1(n14130), .B2(n14622), .A(n13788), .ZN(n13789) );
  AOI21_X1 U15806 ( .B1(n14135), .B2(n14618), .A(n13789), .ZN(n13790) );
  OAI21_X1 U15807 ( .B1(n13791), .B2(n13889), .A(n13790), .ZN(P1_U3225) );
  INV_X1 U15808 ( .A(n13792), .ZN(n13796) );
  AOI21_X1 U15809 ( .B1(n13794), .B2(n13878), .A(n13793), .ZN(n13795) );
  OAI21_X1 U15810 ( .B1(n13796), .B2(n13795), .A(n14613), .ZN(n13804) );
  INV_X1 U15811 ( .A(n13797), .ZN(n13802) );
  INV_X1 U15812 ( .A(n13798), .ZN(n13801) );
  OAI22_X1 U15813 ( .A1(n13799), .A2(n13884), .B1(n13883), .B2(n13862), .ZN(
        n13800) );
  AOI211_X1 U15814 ( .C1(n13865), .C2(n13802), .A(n13801), .B(n13800), .ZN(
        n13803) );
  OAI211_X1 U15815 ( .C1(n14344), .C2(n13868), .A(n13804), .B(n13803), .ZN(
        P1_U3226) );
  INV_X1 U15816 ( .A(n13805), .ZN(n13810) );
  AOI21_X1 U15817 ( .B1(n13807), .B2(n13809), .A(n13806), .ZN(n13808) );
  AOI21_X1 U15818 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n13817) );
  NAND2_X1 U15819 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14680)
         );
  OAI21_X1 U15820 ( .B1(n14622), .B2(n13811), .A(n14680), .ZN(n13814) );
  OAI22_X1 U15821 ( .A1(n13812), .A2(n13883), .B1(n13884), .B2(n13882), .ZN(
        n13813) );
  AOI211_X1 U15822 ( .C1(n13815), .C2(n14618), .A(n13814), .B(n13813), .ZN(
        n13816) );
  OAI21_X1 U15823 ( .B1(n13817), .B2(n13889), .A(n13816), .ZN(P1_U3228) );
  XOR2_X1 U15824 ( .A(n13819), .B(n13818), .Z(n13824) );
  INV_X1 U15825 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13820) );
  OAI22_X1 U15826 ( .A1(n14622), .A2(n14152), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13820), .ZN(n13822) );
  OAI22_X1 U15827 ( .A1(n14141), .A2(n13884), .B1(n13883), .B2(n14143), .ZN(
        n13821) );
  AOI211_X1 U15828 ( .C1(n14286), .C2(n14618), .A(n13822), .B(n13821), .ZN(
        n13823) );
  OAI21_X1 U15829 ( .B1(n13824), .B2(n13889), .A(n13823), .ZN(P1_U3229) );
  INV_X1 U15830 ( .A(n14315), .ZN(n13835) );
  OAI211_X1 U15831 ( .C1(n13827), .C2(n13826), .A(n13825), .B(n14613), .ZN(
        n13834) );
  INV_X1 U15832 ( .A(n13828), .ZN(n14210) );
  AND2_X1 U15833 ( .A1(n14237), .A2(n14234), .ZN(n13829) );
  AOI21_X1 U15834 ( .B1(n13898), .B2(n14236), .A(n13829), .ZN(n14313) );
  INV_X1 U15835 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13830) );
  OAI22_X1 U15836 ( .A1(n14313), .A2(n13831), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13830), .ZN(n13832) );
  AOI21_X1 U15837 ( .B1(n14210), .B2(n13865), .A(n13832), .ZN(n13833) );
  OAI211_X1 U15838 ( .C1(n13835), .C2(n13868), .A(n13834), .B(n13833), .ZN(
        P1_U3233) );
  XNOR2_X1 U15839 ( .A(n13837), .B(n13836), .ZN(n13845) );
  OAI21_X1 U15840 ( .B1(n14622), .B2(n13839), .A(n13838), .ZN(n13842) );
  OAI22_X1 U15841 ( .A1(n13840), .A2(n13884), .B1(n13883), .B2(n13885), .ZN(
        n13841) );
  AOI211_X1 U15842 ( .C1(n13843), .C2(n14618), .A(n13842), .B(n13841), .ZN(
        n13844) );
  OAI21_X1 U15843 ( .B1(n13845), .B2(n13889), .A(n13844), .ZN(P1_U3234) );
  OAI21_X1 U15844 ( .B1(n13848), .B2(n13847), .A(n13846), .ZN(n13849) );
  NAND2_X1 U15845 ( .A1(n13849), .A2(n14613), .ZN(n13855) );
  NAND2_X1 U15846 ( .A1(n13898), .A2(n14234), .ZN(n13851) );
  NAND2_X1 U15847 ( .A1(n13896), .A2(n14236), .ZN(n13850) );
  NAND2_X1 U15848 ( .A1(n13851), .A2(n13850), .ZN(n14182) );
  AOI22_X1 U15849 ( .A1(n14182), .A2(n14615), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13854) );
  NAND2_X1 U15850 ( .A1(n14186), .A2(n14618), .ZN(n13853) );
  NAND2_X1 U15851 ( .A1(n13865), .A2(n14183), .ZN(n13852) );
  NAND4_X1 U15852 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        P1_U3235) );
  INV_X1 U15853 ( .A(n14332), .ZN(n14245) );
  OAI21_X1 U15854 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n13859) );
  NAND2_X1 U15855 ( .A1(n13859), .A2(n14613), .ZN(n13867) );
  INV_X1 U15856 ( .A(n13860), .ZN(n14242) );
  NAND2_X1 U15857 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14693)
         );
  INV_X1 U15858 ( .A(n14693), .ZN(n13864) );
  OAI22_X1 U15859 ( .A1(n13862), .A2(n13884), .B1(n13883), .B2(n13861), .ZN(
        n13863) );
  AOI211_X1 U15860 ( .C1(n13865), .C2(n14242), .A(n13864), .B(n13863), .ZN(
        n13866) );
  OAI211_X1 U15861 ( .C1(n14245), .C2(n13868), .A(n13867), .B(n13866), .ZN(
        P1_U3238) );
  XOR2_X1 U15862 ( .A(n13870), .B(n13869), .Z(n13876) );
  NAND2_X1 U15863 ( .A1(n13894), .A2(n14234), .ZN(n13872) );
  NAND2_X1 U15864 ( .A1(n13893), .A2(n14236), .ZN(n13871) );
  NAND2_X1 U15865 ( .A1(n13872), .A2(n13871), .ZN(n14269) );
  AOI22_X1 U15866 ( .A1(n14615), .A2(n14269), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13873) );
  OAI21_X1 U15867 ( .B1(n14115), .B2(n14622), .A(n13873), .ZN(n13874) );
  AOI21_X1 U15868 ( .B1(n14270), .B2(n14618), .A(n13874), .ZN(n13875) );
  OAI21_X1 U15869 ( .B1(n13876), .B2(n13889), .A(n13875), .ZN(P1_U3240) );
  NAND2_X1 U15870 ( .A1(n13878), .A2(n13877), .ZN(n13879) );
  XOR2_X1 U15871 ( .A(n13880), .B(n13879), .Z(n13890) );
  NAND2_X1 U15872 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14667)
         );
  OAI21_X1 U15873 ( .B1(n14622), .B2(n13881), .A(n14667), .ZN(n13887) );
  OAI22_X1 U15874 ( .A1(n13885), .A2(n13884), .B1(n13883), .B2(n13882), .ZN(
        n13886) );
  AOI211_X1 U15875 ( .C1(n14351), .C2(n14618), .A(n13887), .B(n13886), .ZN(
        n13888) );
  OAI21_X1 U15876 ( .B1(n13890), .B2(n13889), .A(n13888), .ZN(P1_U3241) );
  MUX2_X1 U15877 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14050), .S(P1_U4016), .Z(
        P1_U3591) );
  CLKBUF_X2 U15878 ( .A(P1_U4016), .Z(n13916) );
  MUX2_X1 U15879 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13891), .S(n13916), .Z(
        P1_U3590) );
  MUX2_X1 U15880 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13892), .S(n13916), .Z(
        P1_U3589) );
  MUX2_X1 U15881 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14092), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15882 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13893), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15883 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14093), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15884 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13894), .S(n13916), .Z(
        P1_U3585) );
  MUX2_X1 U15885 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13895), .S(n13916), .Z(
        P1_U3584) );
  MUX2_X1 U15886 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13896), .S(n13916), .Z(
        P1_U3583) );
  MUX2_X1 U15887 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13897), .S(n13916), .Z(
        P1_U3582) );
  MUX2_X1 U15888 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13898), .S(n13916), .Z(
        P1_U3581) );
  MUX2_X1 U15889 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13899), .S(n13916), .Z(
        P1_U3580) );
  MUX2_X1 U15890 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14237), .S(n13916), .Z(
        P1_U3579) );
  MUX2_X1 U15891 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13900), .S(n13916), .Z(
        P1_U3578) );
  MUX2_X1 U15892 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14235), .S(n13916), .Z(
        P1_U3577) );
  MUX2_X1 U15893 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13901), .S(n13916), .Z(
        P1_U3576) );
  MUX2_X1 U15894 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13902), .S(n13916), .Z(
        P1_U3575) );
  MUX2_X1 U15895 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13903), .S(n13916), .Z(
        P1_U3574) );
  MUX2_X1 U15896 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13904), .S(n13916), .Z(
        P1_U3573) );
  MUX2_X1 U15897 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13905), .S(n13916), .Z(
        P1_U3572) );
  MUX2_X1 U15898 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13906), .S(n13916), .Z(
        P1_U3571) );
  MUX2_X1 U15899 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13907), .S(n13916), .Z(
        P1_U3570) );
  MUX2_X1 U15900 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13908), .S(n13916), .Z(
        P1_U3569) );
  MUX2_X1 U15901 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13909), .S(n13916), .Z(
        P1_U3568) );
  MUX2_X1 U15902 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13910), .S(n13916), .Z(
        P1_U3567) );
  MUX2_X1 U15903 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13911), .S(n13916), .Z(
        P1_U3566) );
  MUX2_X1 U15904 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13912), .S(n13916), .Z(
        P1_U3565) );
  MUX2_X1 U15905 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13913), .S(n13916), .Z(
        P1_U3564) );
  MUX2_X1 U15906 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13914), .S(n13916), .Z(
        P1_U3563) );
  MUX2_X1 U15907 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13915), .S(n13916), .Z(
        P1_U3562) );
  MUX2_X1 U15908 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13917), .S(n13916), .Z(
        P1_U3561) );
  MUX2_X1 U15909 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6758), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15910 ( .C1(n13931), .C2(n13920), .A(n14038), .B(n13919), .ZN(
        n13930) );
  MUX2_X1 U15911 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n13922), .S(n13921), .Z(
        n13923) );
  OAI21_X1 U15912 ( .B1(n14652), .B2(n13935), .A(n13923), .ZN(n13924) );
  NAND3_X1 U15913 ( .A1(n14037), .A2(n13925), .A3(n13924), .ZN(n13929) );
  NAND2_X1 U15914 ( .A1(n14002), .A2(n13926), .ZN(n13928) );
  AOI22_X1 U15915 ( .A1(n14655), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13927) );
  NAND4_X1 U15916 ( .A1(n13930), .A2(n13929), .A3(n13928), .A4(n13927), .ZN(
        P1_U3244) );
  INV_X1 U15917 ( .A(n13931), .ZN(n13933) );
  MUX2_X1 U15918 ( .A(n13933), .B(n13932), .S(n6586), .Z(n13937) );
  OAI21_X1 U15919 ( .B1(n6586), .B2(P1_REG2_REG_0__SCAN_IN), .A(n13934), .ZN(
        n14651) );
  NAND2_X1 U15920 ( .A1(n14651), .A2(n13935), .ZN(n13936) );
  OAI211_X1 U15921 ( .C1(n13937), .C2(n14401), .A(P1_U4016), .B(n13936), .ZN(
        n13982) );
  AOI22_X1 U15922 ( .A1(n14655), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13947) );
  OAI211_X1 U15923 ( .C1(n13939), .C2(n13938), .A(n14037), .B(n13953), .ZN(
        n13943) );
  OAI211_X1 U15924 ( .C1(n13941), .C2(n13940), .A(n14038), .B(n13957), .ZN(
        n13942) );
  OAI211_X1 U15925 ( .C1(n14691), .C2(n13944), .A(n13943), .B(n13942), .ZN(
        n13945) );
  INV_X1 U15926 ( .A(n13945), .ZN(n13946) );
  NAND3_X1 U15927 ( .A1(n13982), .A2(n13947), .A3(n13946), .ZN(P1_U3245) );
  OAI22_X1 U15928 ( .A1(n14695), .A2(n14461), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13948), .ZN(n13949) );
  AOI21_X1 U15929 ( .B1(n13950), .B2(n14002), .A(n13949), .ZN(n13962) );
  MUX2_X1 U15930 ( .A(n10049), .B(P1_REG1_REG_3__SCAN_IN), .S(n13950), .Z(
        n13951) );
  NAND3_X1 U15931 ( .A1(n13953), .A2(n13952), .A3(n13951), .ZN(n13954) );
  NAND3_X1 U15932 ( .A1(n14037), .A2(n13976), .A3(n13954), .ZN(n13961) );
  INV_X1 U15933 ( .A(n13968), .ZN(n13959) );
  NAND3_X1 U15934 ( .A1(n13957), .A2(n13956), .A3(n13955), .ZN(n13958) );
  NAND3_X1 U15935 ( .A1(n14038), .A2(n13959), .A3(n13958), .ZN(n13960) );
  NAND3_X1 U15936 ( .A1(n13962), .A2(n13961), .A3(n13960), .ZN(P1_U3246) );
  INV_X1 U15937 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14423) );
  MUX2_X1 U15938 ( .A(n13963), .B(P1_REG2_REG_4__SCAN_IN), .S(n13972), .Z(
        n13966) );
  INV_X1 U15939 ( .A(n13964), .ZN(n13965) );
  NAND2_X1 U15940 ( .A1(n13966), .A2(n13965), .ZN(n13967) );
  OAI211_X1 U15941 ( .C1(n13968), .C2(n13967), .A(n14038), .B(n13993), .ZN(
        n13970) );
  OAI211_X1 U15942 ( .C1(n14423), .C2(n14695), .A(n13970), .B(n13969), .ZN(
        n13971) );
  INV_X1 U15943 ( .A(n13971), .ZN(n13981) );
  NAND2_X1 U15944 ( .A1(n14002), .A2(n13972), .ZN(n13980) );
  INV_X1 U15945 ( .A(n13973), .ZN(n13978) );
  NAND3_X1 U15946 ( .A1(n13976), .A2(n13975), .A3(n13974), .ZN(n13977) );
  NAND3_X1 U15947 ( .A1(n14037), .A2(n13978), .A3(n13977), .ZN(n13979) );
  NAND4_X1 U15948 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        P1_U3247) );
  INV_X1 U15949 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14466) );
  NAND2_X1 U15950 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13983) );
  OAI21_X1 U15951 ( .B1(n14695), .B2(n14466), .A(n13983), .ZN(n13984) );
  AOI21_X1 U15952 ( .B1(n13985), .B2(n14002), .A(n13984), .ZN(n13998) );
  OAI21_X1 U15953 ( .B1(n13988), .B2(n13987), .A(n13986), .ZN(n13989) );
  NAND2_X1 U15954 ( .A1(n14037), .A2(n13989), .ZN(n13997) );
  INV_X1 U15955 ( .A(n13990), .ZN(n13995) );
  NAND3_X1 U15956 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(n13994) );
  NAND3_X1 U15957 ( .A1(n14038), .A2(n13995), .A3(n13994), .ZN(n13996) );
  NAND3_X1 U15958 ( .A1(n13998), .A2(n13997), .A3(n13996), .ZN(P1_U3248) );
  INV_X1 U15959 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14000) );
  OAI21_X1 U15960 ( .B1(n14695), .B2(n14000), .A(n13999), .ZN(n14001) );
  AOI21_X1 U15961 ( .B1(n14004), .B2(n14002), .A(n14001), .ZN(n14019) );
  INV_X1 U15962 ( .A(n14003), .ZN(n14007) );
  MUX2_X1 U15963 ( .A(n14005), .B(P1_REG1_REG_7__SCAN_IN), .S(n14004), .Z(
        n14006) );
  NAND2_X1 U15964 ( .A1(n14007), .A2(n14006), .ZN(n14009) );
  OAI211_X1 U15965 ( .C1(n14010), .C2(n14009), .A(n14037), .B(n14008), .ZN(
        n14018) );
  INV_X1 U15966 ( .A(n14011), .ZN(n14016) );
  NAND3_X1 U15967 ( .A1(n14014), .A2(n14013), .A3(n14012), .ZN(n14015) );
  NAND3_X1 U15968 ( .A1(n14038), .A2(n14016), .A3(n14015), .ZN(n14017) );
  NAND3_X1 U15969 ( .A1(n14019), .A2(n14018), .A3(n14017), .ZN(P1_U3250) );
  INV_X1 U15970 ( .A(n14554), .ZN(n14046) );
  INV_X1 U15971 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14021) );
  AOI22_X1 U15972 ( .A1(n14025), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14021), 
        .B2(n14678), .ZN(n14675) );
  OAI21_X1 U15973 ( .B1(n11311), .B2(n14027), .A(n14020), .ZN(n14674) );
  NAND2_X1 U15974 ( .A1(n14675), .A2(n14674), .ZN(n14673) );
  OAI21_X1 U15975 ( .B1(n14021), .B2(n14678), .A(n14673), .ZN(n14022) );
  XOR2_X1 U15976 ( .A(n14030), .B(n14022), .Z(n14685) );
  NAND2_X1 U15977 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14685), .ZN(n14684) );
  NAND2_X1 U15978 ( .A1(n14030), .A2(n14022), .ZN(n14023) );
  NAND2_X1 U15979 ( .A1(n14684), .A2(n14023), .ZN(n14024) );
  XOR2_X1 U15980 ( .A(n14024), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14039) );
  INV_X1 U15981 ( .A(n14039), .ZN(n14035) );
  INV_X1 U15982 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14028) );
  AOI22_X1 U15983 ( .A1(n14025), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n14028), 
        .B2(n14678), .ZN(n14672) );
  INV_X1 U15984 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n15430) );
  OAI21_X1 U15985 ( .B1(n15430), .B2(n14027), .A(n14026), .ZN(n14671) );
  NAND2_X1 U15986 ( .A1(n14672), .A2(n14671), .ZN(n14670) );
  OAI21_X1 U15987 ( .B1(n14028), .B2(n14678), .A(n14670), .ZN(n14029) );
  XOR2_X1 U15988 ( .A(n14030), .B(n14029), .Z(n14683) );
  NAND2_X1 U15989 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14683), .ZN(n14682) );
  NAND2_X1 U15990 ( .A1(n14030), .A2(n14029), .ZN(n14031) );
  NAND2_X1 U15991 ( .A1(n14682), .A2(n14031), .ZN(n14033) );
  XNOR2_X1 U15992 ( .A(n14033), .B(n14032), .ZN(n14036) );
  OAI21_X1 U15993 ( .B1(n14036), .B2(n14689), .A(n14691), .ZN(n14034) );
  AOI21_X1 U15994 ( .B1(n14038), .B2(n14035), .A(n14034), .ZN(n14042) );
  AOI22_X1 U15995 ( .A1(n14039), .A2(n14038), .B1(n14037), .B2(n14036), .ZN(
        n14041) );
  MUX2_X1 U15996 ( .A(n14042), .B(n14041), .S(n14040), .Z(n14045) );
  INV_X1 U15997 ( .A(n14043), .ZN(n14044) );
  OAI211_X1 U15998 ( .C1(n14046), .C2(n14695), .A(n14045), .B(n14044), .ZN(
        P1_U3262) );
  NAND2_X1 U15999 ( .A1(n14360), .A2(n14054), .ZN(n14053) );
  XOR2_X1 U16000 ( .A(n14047), .B(n14053), .Z(n14255) );
  NAND2_X1 U16001 ( .A1(n14255), .A2(n14048), .ZN(n14052) );
  AND2_X1 U16002 ( .A1(n14050), .A2(n14049), .ZN(n14253) );
  INV_X1 U16003 ( .A(n14253), .ZN(n14259) );
  NOR2_X1 U16004 ( .A1(n14712), .A2(n14259), .ZN(n14055) );
  AOI21_X1 U16005 ( .B1(n14712), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14055), 
        .ZN(n14051) );
  OAI211_X1 U16006 ( .C1(n14358), .C2(n14244), .A(n14052), .B(n14051), .ZN(
        P1_U3263) );
  OAI21_X1 U16007 ( .B1(n14360), .B2(n14054), .A(n14053), .ZN(n14258) );
  NAND2_X1 U16008 ( .A1(n14712), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14057) );
  INV_X1 U16009 ( .A(n14055), .ZN(n14056) );
  OAI211_X1 U16010 ( .C1(n14360), .C2(n14244), .A(n14057), .B(n14056), .ZN(
        n14058) );
  INV_X1 U16011 ( .A(n14058), .ZN(n14059) );
  OAI21_X1 U16012 ( .B1(n14258), .B2(n14214), .A(n14059), .ZN(P1_U3264) );
  INV_X1 U16013 ( .A(n14060), .ZN(n14075) );
  OAI22_X1 U16014 ( .A1(n14063), .A2(n14062), .B1(n14061), .B2(n14698), .ZN(
        n14066) );
  NOR2_X1 U16015 ( .A1(n14712), .A2(n14064), .ZN(n14065) );
  AOI211_X1 U16016 ( .C1(n14712), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14066), 
        .B(n14065), .ZN(n14069) );
  NAND2_X1 U16017 ( .A1(n14067), .A2(n14703), .ZN(n14068) );
  OAI211_X1 U16018 ( .C1(n14071), .C2(n14070), .A(n14069), .B(n14068), .ZN(
        n14072) );
  AOI21_X1 U16019 ( .B1(n14073), .B2(n14121), .A(n14072), .ZN(n14074) );
  OAI21_X1 U16020 ( .B1(n14075), .B2(n14248), .A(n14074), .ZN(P1_U3356) );
  INV_X1 U16021 ( .A(n14076), .ZN(n14083) );
  OAI22_X1 U16022 ( .A1(n14712), .A2(n14078), .B1(n14077), .B2(n14698), .ZN(
        n14079) );
  AOI21_X1 U16023 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(n14712), .A(n14079), 
        .ZN(n14080) );
  OAI21_X1 U16024 ( .B1(n14081), .B2(n14244), .A(n14080), .ZN(n14082) );
  AOI21_X1 U16025 ( .B1(n14083), .B2(n14251), .A(n14082), .ZN(n14086) );
  NAND2_X1 U16026 ( .A1(n14084), .A2(n14121), .ZN(n14085) );
  OAI211_X1 U16027 ( .C1(n14087), .C2(n14248), .A(n14086), .B(n14085), .ZN(
        P1_U3265) );
  INV_X1 U16028 ( .A(n14088), .ZN(n14089) );
  NAND2_X1 U16029 ( .A1(n14091), .A2(n14090), .ZN(n14097) );
  NAND2_X1 U16030 ( .A1(n14092), .A2(n14236), .ZN(n14095) );
  OAI21_X1 U16031 ( .B1(n14100), .B2(n14099), .A(n14098), .ZN(n14264) );
  AOI211_X1 U16032 ( .C1(n14101), .C2(n14114), .A(n14317), .B(n6617), .ZN(
        n14265) );
  NAND2_X1 U16033 ( .A1(n14265), .A2(n14251), .ZN(n14105) );
  INV_X1 U16034 ( .A(n14102), .ZN(n14103) );
  AOI22_X1 U16035 ( .A1(n14712), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14103), 
        .B2(n14241), .ZN(n14104) );
  OAI211_X1 U16036 ( .C1(n14366), .C2(n14244), .A(n14105), .B(n14104), .ZN(
        n14106) );
  AOI21_X1 U16037 ( .B1(n14264), .B2(n14229), .A(n14106), .ZN(n14107) );
  OAI21_X1 U16038 ( .B1(n14712), .B2(n14263), .A(n14107), .ZN(P1_U3266) );
  XNOR2_X1 U16039 ( .A(n14109), .B(n14108), .ZN(n14276) );
  OAI21_X1 U16040 ( .B1(n14112), .B2(n14111), .A(n14110), .ZN(n14274) );
  OAI21_X1 U16041 ( .B1(n8142), .B2(n14113), .A(n14114), .ZN(n14272) );
  INV_X1 U16042 ( .A(n14269), .ZN(n14116) );
  OAI22_X1 U16043 ( .A1(n14712), .A2(n14116), .B1(n14115), .B2(n14698), .ZN(
        n14118) );
  NOR2_X1 U16044 ( .A1(n8142), .A2(n14244), .ZN(n14117) );
  AOI211_X1 U16045 ( .C1(n14712), .C2(P1_REG2_REG_26__SCAN_IN), .A(n14118), 
        .B(n14117), .ZN(n14119) );
  OAI21_X1 U16046 ( .B1(n14214), .B2(n14272), .A(n14119), .ZN(n14120) );
  AOI21_X1 U16047 ( .B1(n14121), .B2(n14274), .A(n14120), .ZN(n14122) );
  OAI21_X1 U16048 ( .B1(n14248), .B2(n14276), .A(n14122), .ZN(P1_U3267) );
  XNOR2_X1 U16049 ( .A(n14124), .B(n14123), .ZN(n14282) );
  XNOR2_X1 U16050 ( .A(n14126), .B(n14125), .ZN(n14277) );
  AOI21_X1 U16051 ( .B1(n14135), .B2(n14150), .A(n14317), .ZN(n14128) );
  NAND2_X1 U16052 ( .A1(n14128), .A2(n14127), .ZN(n14279) );
  INV_X1 U16053 ( .A(n14129), .ZN(n14278) );
  NAND2_X1 U16054 ( .A1(n14712), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14133) );
  INV_X1 U16055 ( .A(n14130), .ZN(n14131) );
  NAND2_X1 U16056 ( .A1(n14241), .A2(n14131), .ZN(n14132) );
  OAI211_X1 U16057 ( .C1(n14712), .C2(n14278), .A(n14133), .B(n14132), .ZN(
        n14134) );
  AOI21_X1 U16058 ( .B1(n14135), .B2(n14703), .A(n14134), .ZN(n14136) );
  OAI21_X1 U16059 ( .B1(n14279), .B2(n14706), .A(n14136), .ZN(n14137) );
  AOI21_X1 U16060 ( .B1(n14277), .B2(n14229), .A(n14137), .ZN(n14138) );
  OAI21_X1 U16061 ( .B1(n14232), .B2(n14282), .A(n14138), .ZN(P1_U3268) );
  OAI21_X1 U16062 ( .B1(n6640), .B2(n14147), .A(n14139), .ZN(n14156) );
  OAI22_X1 U16063 ( .A1(n14143), .A2(n14142), .B1(n14141), .B2(n14140), .ZN(
        n14149) );
  INV_X1 U16064 ( .A(n14144), .ZN(n14145) );
  AOI211_X1 U16065 ( .C1(n14147), .C2(n14146), .A(n14329), .B(n14145), .ZN(
        n14148) );
  AOI211_X1 U16066 ( .C1(n14730), .C2(n14156), .A(n14149), .B(n14148), .ZN(
        n14288) );
  INV_X1 U16067 ( .A(n14150), .ZN(n14151) );
  AOI211_X1 U16068 ( .C1(n14286), .C2(n14168), .A(n14317), .B(n14151), .ZN(
        n14285) );
  INV_X1 U16069 ( .A(n14286), .ZN(n14155) );
  INV_X1 U16070 ( .A(n14152), .ZN(n14153) );
  AOI22_X1 U16071 ( .A1(n14712), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14153), 
        .B2(n14241), .ZN(n14154) );
  OAI21_X1 U16072 ( .B1(n14155), .B2(n14244), .A(n14154), .ZN(n14158) );
  INV_X1 U16073 ( .A(n14156), .ZN(n14289) );
  NOR2_X1 U16074 ( .A1(n14289), .A2(n14697), .ZN(n14157) );
  AOI211_X1 U16075 ( .C1(n14285), .C2(n14251), .A(n14158), .B(n14157), .ZN(
        n14159) );
  OAI21_X1 U16076 ( .B1(n14288), .B2(n14712), .A(n14159), .ZN(P1_U3269) );
  OAI21_X1 U16077 ( .B1(n14162), .B2(n14161), .A(n14160), .ZN(n14163) );
  INV_X1 U16078 ( .A(n14163), .ZN(n14292) );
  INV_X1 U16079 ( .A(n14164), .ZN(n14291) );
  INV_X1 U16080 ( .A(n14165), .ZN(n14166) );
  AOI22_X1 U16081 ( .A1(n14712), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14166), 
        .B2(n14241), .ZN(n14167) );
  OAI21_X1 U16082 ( .B1(n14291), .B2(n14712), .A(n14167), .ZN(n14171) );
  INV_X1 U16083 ( .A(n14181), .ZN(n14169) );
  OAI211_X1 U16084 ( .C1(n14169), .C2(n14376), .A(n14254), .B(n14168), .ZN(
        n14290) );
  NOR2_X1 U16085 ( .A1(n14290), .A2(n14706), .ZN(n14170) );
  AOI211_X1 U16086 ( .C1(n14703), .C2(n6770), .A(n14171), .B(n14170), .ZN(
        n14176) );
  XNOR2_X1 U16087 ( .A(n14174), .B(n14173), .ZN(n14294) );
  NAND2_X1 U16088 ( .A1(n14294), .A2(n14229), .ZN(n14175) );
  OAI211_X1 U16089 ( .C1(n14292), .C2(n14232), .A(n14176), .B(n14175), .ZN(
        P1_U3270) );
  XNOR2_X1 U16090 ( .A(n14177), .B(n7121), .ZN(n14301) );
  OAI21_X1 U16091 ( .B1(n14180), .B2(n14179), .A(n14178), .ZN(n14296) );
  OAI211_X1 U16092 ( .C1(n14380), .C2(n14195), .A(n14254), .B(n14181), .ZN(
        n14298) );
  INV_X1 U16093 ( .A(n14182), .ZN(n14297) );
  AOI22_X1 U16094 ( .A1(n14183), .A2(n14241), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14712), .ZN(n14184) );
  OAI21_X1 U16095 ( .B1(n14297), .B2(n14712), .A(n14184), .ZN(n14185) );
  AOI21_X1 U16096 ( .B1(n14186), .B2(n14703), .A(n14185), .ZN(n14187) );
  OAI21_X1 U16097 ( .B1(n14298), .B2(n14706), .A(n14187), .ZN(n14188) );
  AOI21_X1 U16098 ( .B1(n14296), .B2(n14229), .A(n14188), .ZN(n14189) );
  OAI21_X1 U16099 ( .B1(n14301), .B2(n14232), .A(n14189), .ZN(P1_U3271) );
  XNOR2_X1 U16100 ( .A(n14190), .B(n14191), .ZN(n14310) );
  XNOR2_X1 U16101 ( .A(n14192), .B(n14191), .ZN(n14305) );
  NAND2_X1 U16102 ( .A1(n6612), .A2(n14384), .ZN(n14193) );
  NAND2_X1 U16103 ( .A1(n14193), .A2(n14254), .ZN(n14194) );
  OR2_X1 U16104 ( .A1(n14195), .A2(n14194), .ZN(n14307) );
  NOR2_X1 U16105 ( .A1(n14307), .A2(n14706), .ZN(n14202) );
  INV_X1 U16106 ( .A(n14196), .ZN(n14306) );
  NAND2_X1 U16107 ( .A1(n14384), .A2(n14703), .ZN(n14200) );
  INV_X1 U16108 ( .A(n14197), .ZN(n14198) );
  AOI22_X1 U16109 ( .A1(n14198), .A2(n14241), .B1(n14712), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14199) );
  OAI211_X1 U16110 ( .C1(n14712), .C2(n14306), .A(n14200), .B(n14199), .ZN(
        n14201) );
  AOI211_X1 U16111 ( .C1(n14305), .C2(n14229), .A(n14202), .B(n14201), .ZN(
        n14203) );
  OAI21_X1 U16112 ( .B1(n14232), .B2(n14310), .A(n14203), .ZN(P1_U3272) );
  OAI21_X1 U16113 ( .B1(n6724), .B2(n14208), .A(n14204), .ZN(n14322) );
  INV_X1 U16114 ( .A(n14205), .ZN(n14206) );
  AOI21_X1 U16115 ( .B1(n14208), .B2(n14207), .A(n14206), .ZN(n14320) );
  NAND2_X1 U16116 ( .A1(n14218), .A2(n14315), .ZN(n14209) );
  NAND2_X1 U16117 ( .A1(n6612), .A2(n14209), .ZN(n14318) );
  AOI22_X1 U16118 ( .A1(n14712), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14210), 
        .B2(n14241), .ZN(n14211) );
  OAI21_X1 U16119 ( .B1(n14313), .B2(n14712), .A(n14211), .ZN(n14212) );
  AOI21_X1 U16120 ( .B1(n14315), .B2(n14703), .A(n14212), .ZN(n14213) );
  OAI21_X1 U16121 ( .B1(n14318), .B2(n14214), .A(n14213), .ZN(n14215) );
  AOI21_X1 U16122 ( .B1(n14320), .B2(n14229), .A(n14215), .ZN(n14216) );
  OAI21_X1 U16123 ( .B1(n14232), .B2(n14322), .A(n14216), .ZN(P1_U3273) );
  XOR2_X1 U16124 ( .A(n14217), .B(n14227), .Z(n14330) );
  AOI21_X1 U16125 ( .B1(n14325), .B2(n14239), .A(n14317), .ZN(n14219) );
  AND2_X1 U16126 ( .A1(n14219), .A2(n14218), .ZN(n14323) );
  INV_X1 U16127 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U16128 ( .A1(n14325), .A2(n14703), .ZN(n14223) );
  NOR2_X1 U16129 ( .A1(n14220), .A2(n14698), .ZN(n14221) );
  AOI21_X1 U16130 ( .B1(n14324), .B2(n14225), .A(n14221), .ZN(n14222) );
  OAI211_X1 U16131 ( .C1(n14225), .C2(n14224), .A(n14223), .B(n14222), .ZN(
        n14226) );
  AOI21_X1 U16132 ( .B1(n14323), .B2(n14251), .A(n14226), .ZN(n14231) );
  XNOR2_X1 U16133 ( .A(n14228), .B(n14227), .ZN(n14326) );
  NAND2_X1 U16134 ( .A1(n14326), .A2(n14229), .ZN(n14230) );
  OAI211_X1 U16135 ( .C1(n14330), .C2(n14232), .A(n14231), .B(n14230), .ZN(
        P1_U3274) );
  XOR2_X1 U16136 ( .A(n14233), .B(n14246), .Z(n14238) );
  AOI222_X1 U16137 ( .A1(n14741), .A2(n14238), .B1(n14237), .B2(n14236), .C1(
        n14235), .C2(n14234), .ZN(n14334) );
  AOI211_X1 U16138 ( .C1(n14332), .C2(n14240), .A(n14317), .B(n7068), .ZN(
        n14331) );
  AOI22_X1 U16139 ( .A1(n14712), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14242), 
        .B2(n14241), .ZN(n14243) );
  OAI21_X1 U16140 ( .B1(n14245), .B2(n14244), .A(n14243), .ZN(n14250) );
  XOR2_X1 U16141 ( .A(n14247), .B(n14246), .Z(n14335) );
  NOR2_X1 U16142 ( .A1(n14335), .A2(n14248), .ZN(n14249) );
  AOI211_X1 U16143 ( .C1(n14331), .C2(n14251), .A(n14250), .B(n14249), .ZN(
        n14252) );
  OAI21_X1 U16144 ( .B1(n14712), .B2(n14334), .A(n14252), .ZN(P1_U3275) );
  AOI21_X1 U16145 ( .B1(n14255), .B2(n14254), .A(n14253), .ZN(n14356) );
  INV_X1 U16146 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14256) );
  MUX2_X1 U16147 ( .A(n14356), .B(n14256), .S(n14757), .Z(n14257) );
  OAI21_X1 U16148 ( .B1(n14358), .B2(n14304), .A(n14257), .ZN(P1_U3559) );
  OR2_X1 U16149 ( .A1(n14258), .A2(n14317), .ZN(n14260) );
  NAND2_X1 U16150 ( .A1(n14260), .A2(n14259), .ZN(n14359) );
  MUX2_X1 U16151 ( .A(n14359), .B(P1_REG1_REG_30__SCAN_IN), .S(n14757), .Z(
        n14262) );
  NOR2_X1 U16152 ( .A1(n14360), .A2(n14304), .ZN(n14261) );
  INV_X1 U16153 ( .A(n14263), .ZN(n14266) );
  OAI21_X1 U16154 ( .B1(n14366), .B2(n14304), .A(n14268), .ZN(P1_U3555) );
  AOI21_X1 U16155 ( .B1(n14270), .B2(n14744), .A(n14269), .ZN(n14271) );
  OAI21_X1 U16156 ( .B1(n14272), .B2(n14317), .A(n14271), .ZN(n14273) );
  AOI21_X1 U16157 ( .B1(n14274), .B2(n14741), .A(n14273), .ZN(n14275) );
  OAI21_X1 U16158 ( .B1(n14276), .B2(n14749), .A(n14275), .ZN(n14367) );
  MUX2_X1 U16159 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14367), .S(n14759), .Z(
        P1_U3554) );
  NAND2_X1 U16160 ( .A1(n14277), .A2(n14626), .ZN(n14281) );
  AND2_X1 U16161 ( .A1(n14279), .A2(n14278), .ZN(n14280) );
  OAI211_X1 U16162 ( .C1(n14329), .C2(n14282), .A(n14281), .B(n14280), .ZN(
        n14368) );
  MUX2_X1 U16163 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14368), .S(n14759), .Z(
        n14283) );
  INV_X1 U16164 ( .A(n14283), .ZN(n14284) );
  OAI21_X1 U16165 ( .B1(n14371), .B2(n14304), .A(n14284), .ZN(P1_U3553) );
  AOI21_X1 U16166 ( .B1(n14286), .B2(n14744), .A(n14285), .ZN(n14287) );
  OAI211_X1 U16167 ( .C1(n14289), .C2(n14723), .A(n14288), .B(n14287), .ZN(
        n14372) );
  MUX2_X1 U16168 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14372), .S(n14759), .Z(
        P1_U3552) );
  OAI211_X1 U16169 ( .C1(n14292), .C2(n14329), .A(n14291), .B(n14290), .ZN(
        n14293) );
  AOI21_X1 U16170 ( .B1(n14294), .B2(n14626), .A(n14293), .ZN(n14373) );
  MUX2_X1 U16171 ( .A(n15397), .B(n14373), .S(n14759), .Z(n14295) );
  OAI21_X1 U16172 ( .B1(n14376), .B2(n14304), .A(n14295), .ZN(P1_U3551) );
  NAND2_X1 U16173 ( .A1(n14296), .A2(n14626), .ZN(n14300) );
  AND2_X1 U16174 ( .A1(n14298), .A2(n14297), .ZN(n14299) );
  OAI211_X1 U16175 ( .C1(n14329), .C2(n14301), .A(n14300), .B(n14299), .ZN(
        n14377) );
  MUX2_X1 U16176 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14377), .S(n14759), .Z(
        n14302) );
  INV_X1 U16177 ( .A(n14302), .ZN(n14303) );
  OAI21_X1 U16178 ( .B1(n14304), .B2(n14380), .A(n14303), .ZN(P1_U3550) );
  NAND2_X1 U16179 ( .A1(n14305), .A2(n14626), .ZN(n14309) );
  AND2_X1 U16180 ( .A1(n14307), .A2(n14306), .ZN(n14308) );
  OAI211_X1 U16181 ( .C1(n14329), .C2(n14310), .A(n14309), .B(n14308), .ZN(
        n14382) );
  MUX2_X1 U16182 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14382), .S(n14759), .Z(
        n14311) );
  AOI21_X1 U16183 ( .B1(n8207), .B2(n14384), .A(n14311), .ZN(n14312) );
  INV_X1 U16184 ( .A(n14312), .ZN(P1_U3549) );
  INV_X1 U16185 ( .A(n14313), .ZN(n14314) );
  AOI21_X1 U16186 ( .B1(n14315), .B2(n14744), .A(n14314), .ZN(n14316) );
  OAI21_X1 U16187 ( .B1(n14318), .B2(n14317), .A(n14316), .ZN(n14319) );
  AOI21_X1 U16188 ( .B1(n14320), .B2(n14626), .A(n14319), .ZN(n14321) );
  OAI21_X1 U16189 ( .B1(n14329), .B2(n14322), .A(n14321), .ZN(n14386) );
  MUX2_X1 U16190 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14386), .S(n14759), .Z(
        P1_U3548) );
  AOI211_X1 U16191 ( .C1(n14325), .C2(n14744), .A(n14324), .B(n14323), .ZN(
        n14328) );
  NAND2_X1 U16192 ( .A1(n14326), .A2(n14626), .ZN(n14327) );
  OAI211_X1 U16193 ( .C1(n14330), .C2(n14329), .A(n14328), .B(n14327), .ZN(
        n14387) );
  MUX2_X1 U16194 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14387), .S(n14759), .Z(
        P1_U3547) );
  AOI21_X1 U16195 ( .B1(n14332), .B2(n14744), .A(n14331), .ZN(n14333) );
  OAI211_X1 U16196 ( .C1(n14749), .C2(n14335), .A(n14334), .B(n14333), .ZN(
        n14388) );
  MUX2_X1 U16197 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14388), .S(n14759), .Z(
        P1_U3546) );
  INV_X1 U16198 ( .A(n14744), .ZN(n14735) );
  OAI211_X1 U16199 ( .C1(n14338), .C2(n14735), .A(n14337), .B(n14336), .ZN(
        n14339) );
  AOI21_X1 U16200 ( .B1(n14340), .B2(n14741), .A(n14339), .ZN(n14341) );
  OAI21_X1 U16201 ( .B1(n14749), .B2(n14342), .A(n14341), .ZN(n14389) );
  MUX2_X1 U16202 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14389), .S(n14759), .Z(
        P1_U3545) );
  OAI21_X1 U16203 ( .B1(n14344), .B2(n14735), .A(n14343), .ZN(n14346) );
  AOI211_X1 U16204 ( .C1(n14626), .C2(n14347), .A(n14346), .B(n14345), .ZN(
        n14348) );
  INV_X1 U16205 ( .A(n14348), .ZN(n14390) );
  MUX2_X1 U16206 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14390), .S(n14759), .Z(
        P1_U3544) );
  AOI211_X1 U16207 ( .C1(n14351), .C2(n14744), .A(n14350), .B(n14349), .ZN(
        n14354) );
  NAND2_X1 U16208 ( .A1(n14352), .A2(n14741), .ZN(n14353) );
  OAI211_X1 U16209 ( .C1(n14749), .C2(n14355), .A(n14354), .B(n14353), .ZN(
        n14391) );
  MUX2_X1 U16210 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14391), .S(n14759), .Z(
        P1_U3543) );
  MUX2_X1 U16211 ( .A(n14356), .B(n15464), .S(n14751), .Z(n14357) );
  OAI21_X1 U16212 ( .B1(n14358), .B2(n14381), .A(n14357), .ZN(P1_U3527) );
  MUX2_X1 U16213 ( .A(n14359), .B(P1_REG0_REG_30__SCAN_IN), .S(n14751), .Z(
        n14362) );
  NOR2_X1 U16214 ( .A1(n14360), .A2(n14381), .ZN(n14361) );
  INV_X1 U16215 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14364) );
  MUX2_X1 U16216 ( .A(n14364), .B(n14363), .S(n14752), .Z(n14365) );
  OAI21_X1 U16217 ( .B1(n14366), .B2(n14381), .A(n14365), .ZN(P1_U3523) );
  MUX2_X1 U16218 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14367), .S(n14752), .Z(
        P1_U3522) );
  MUX2_X1 U16219 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14368), .S(n14752), .Z(
        n14369) );
  INV_X1 U16220 ( .A(n14369), .ZN(n14370) );
  OAI21_X1 U16221 ( .B1(n14371), .B2(n14381), .A(n14370), .ZN(P1_U3521) );
  MUX2_X1 U16222 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14372), .S(n14752), .Z(
        P1_U3520) );
  INV_X1 U16223 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14374) );
  MUX2_X1 U16224 ( .A(n14374), .B(n14373), .S(n14752), .Z(n14375) );
  OAI21_X1 U16225 ( .B1(n14376), .B2(n14381), .A(n14375), .ZN(P1_U3519) );
  MUX2_X1 U16226 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14377), .S(n14752), .Z(
        n14378) );
  INV_X1 U16227 ( .A(n14378), .ZN(n14379) );
  OAI21_X1 U16228 ( .B1(n14381), .B2(n14380), .A(n14379), .ZN(P1_U3518) );
  MUX2_X1 U16229 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14382), .S(n14752), .Z(
        n14383) );
  AOI21_X1 U16230 ( .B1(n8212), .B2(n14384), .A(n14383), .ZN(n14385) );
  INV_X1 U16231 ( .A(n14385), .ZN(P1_U3517) );
  MUX2_X1 U16232 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14386), .S(n14752), .Z(
        P1_U3516) );
  MUX2_X1 U16233 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14387), .S(n14752), .Z(
        P1_U3515) );
  MUX2_X1 U16234 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14388), .S(n14752), .Z(
        P1_U3513) );
  MUX2_X1 U16235 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14389), .S(n14752), .Z(
        P1_U3510) );
  MUX2_X1 U16236 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14390), .S(n14752), .Z(
        P1_U3507) );
  MUX2_X1 U16237 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14391), .S(n14752), .Z(
        P1_U3504) );
  NOR4_X1 U16238 ( .A1(n14393), .A2(P1_IR_REG_30__SCAN_IN), .A3(n7918), .A4(
        P1_U3086), .ZN(n14394) );
  AOI21_X1 U16239 ( .B1(n14395), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14394), 
        .ZN(n14396) );
  OAI21_X1 U16240 ( .B1(n14397), .B2(n14403), .A(n14396), .ZN(P1_U3324) );
  OAI222_X1 U16241 ( .A1(P1_U3086), .A2(n14400), .B1(n14413), .B2(n14399), 
        .C1(n14398), .C2(n14410), .ZN(P1_U3326) );
  OAI222_X1 U16242 ( .A1(n14410), .A2(n14404), .B1(n14403), .B2(n14402), .C1(
        P1_U3086), .C2(n14401), .ZN(P1_U3327) );
  NAND2_X1 U16243 ( .A1(n14406), .A2(n14405), .ZN(n14408) );
  OAI211_X1 U16244 ( .C1(n14409), .C2(n14410), .A(n14408), .B(n14407), .ZN(
        P1_U3328) );
  OAI222_X1 U16245 ( .A1(P1_U3086), .A2(n14414), .B1(n14413), .B2(n14412), 
        .C1(n14411), .C2(n14410), .ZN(P1_U3329) );
  MUX2_X1 U16246 ( .A(n8143), .B(n14415), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16247 ( .A(n14416), .ZN(n14417) );
  MUX2_X1 U16248 ( .A(n14417), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16249 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14869) );
  INV_X1 U16250 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14857) );
  INV_X1 U16251 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14441) );
  INV_X1 U16252 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14418) );
  XOR2_X1 U16253 ( .A(n14418), .B(n14441), .Z(n14487) );
  XNOR2_X1 U16254 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14443) );
  XOR2_X1 U16255 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n14481) );
  XNOR2_X1 U16256 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n14447) );
  NAND2_X1 U16257 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14420), .ZN(n14421) );
  NAND2_X1 U16258 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14422), .ZN(n14424) );
  NAND2_X1 U16259 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14425), .ZN(n14427) );
  NAND2_X1 U16260 ( .A1(n14465), .A2(n14466), .ZN(n14426) );
  INV_X1 U16261 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15068) );
  NAND2_X1 U16262 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15068), .ZN(n14428) );
  INV_X1 U16263 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U16264 ( .A1(n14431), .A2(n14430), .ZN(n14433) );
  XNOR2_X1 U16265 ( .A(n14431), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14475) );
  NAND2_X1 U16266 ( .A1(n14475), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14432) );
  NAND2_X1 U16267 ( .A1(n14433), .A2(n14432), .ZN(n14448) );
  NAND2_X1 U16268 ( .A1(n14447), .A2(n14448), .ZN(n14434) );
  XNOR2_X1 U16269 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .ZN(n14445) );
  NAND2_X1 U16270 ( .A1(n14446), .A2(n14445), .ZN(n14437) );
  NAND2_X1 U16271 ( .A1(n14443), .A2(n14444), .ZN(n14438) );
  XOR2_X1 U16272 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14442) );
  XNOR2_X1 U16273 ( .A(n14491), .B(n14442), .ZN(n14639) );
  INV_X1 U16274 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14842) );
  XOR2_X1 U16275 ( .A(n14444), .B(n14443), .Z(n14631) );
  XOR2_X1 U16276 ( .A(n14446), .B(n14445), .Z(n14532) );
  XOR2_X1 U16277 ( .A(n14448), .B(n14447), .Z(n14479) );
  NAND2_X1 U16278 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14450), .ZN(n14464) );
  INV_X1 U16279 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14787) );
  INV_X1 U16280 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14521) );
  XNOR2_X1 U16281 ( .A(n14452), .B(n14451), .ZN(n14519) );
  XNOR2_X1 U16282 ( .A(n14453), .B(n14454), .ZN(n14456) );
  NAND2_X1 U16283 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14456), .ZN(n14458) );
  AOI21_X1 U16284 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14455), .A(n14454), .ZN(
        n15517) );
  NOR2_X1 U16285 ( .A1(n15517), .A2(n15516), .ZN(n15525) );
  NAND2_X1 U16286 ( .A1(n14458), .A2(n14457), .ZN(n14520) );
  NAND2_X1 U16287 ( .A1(n14519), .A2(n14520), .ZN(n14459) );
  NOR2_X1 U16288 ( .A1(n14519), .A2(n14520), .ZN(n14518) );
  XNOR2_X1 U16289 ( .A(n14461), .B(n14460), .ZN(n15522) );
  NOR2_X1 U16290 ( .A1(n15521), .A2(n15522), .ZN(n14463) );
  INV_X1 U16291 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U16292 ( .A1(n15521), .A2(n15522), .ZN(n15520) );
  OAI21_X1 U16293 ( .B1(n14463), .B2(n14462), .A(n15520), .ZN(n15513) );
  NOR2_X1 U16294 ( .A1(n14468), .A2(n14467), .ZN(n14470) );
  NOR2_X1 U16295 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15515), .ZN(n14469) );
  NAND2_X1 U16296 ( .A1(n14471), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14474) );
  XOR2_X1 U16297 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n14472) );
  XOR2_X1 U16298 ( .A(n14473), .B(n14472), .Z(n14523) );
  NAND2_X1 U16299 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14476), .ZN(n14477) );
  XOR2_X1 U16300 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14475), .Z(n15519) );
  XNOR2_X1 U16301 ( .A(n14481), .B(n14480), .ZN(n14483) );
  NAND2_X1 U16302 ( .A1(n14482), .A2(n14483), .ZN(n14485) );
  INV_X1 U16303 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14828) );
  XNOR2_X1 U16304 ( .A(n14487), .B(n14486), .ZN(n14635) );
  INV_X1 U16305 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14488) );
  NAND2_X1 U16306 ( .A1(n14634), .A2(n14635), .ZN(n14633) );
  XNOR2_X1 U16307 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14493) );
  AND2_X1 U16308 ( .A1(n14492), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14490) );
  XNOR2_X1 U16309 ( .A(n14493), .B(n14497), .ZN(n14643) );
  XNOR2_X1 U16310 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14499) );
  NOR2_X1 U16311 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14495), .ZN(n14498) );
  INV_X1 U16312 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14496) );
  OAI22_X1 U16313 ( .A1(n14498), .A2(n14497), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14496), .ZN(n14503) );
  XOR2_X1 U16314 ( .A(n14499), .B(n14503), .Z(n14501) );
  NOR2_X1 U16315 ( .A1(n14500), .A2(n14501), .ZN(n14646) );
  NAND2_X1 U16316 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14508), .ZN(n14509) );
  OAI21_X1 U16317 ( .B1(n14508), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14509), 
        .ZN(n14505) );
  INV_X1 U16318 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14669) );
  NOR2_X1 U16319 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14669), .ZN(n14504) );
  OAI22_X1 U16320 ( .A1(n14504), .A2(n14503), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14502), .ZN(n14510) );
  XOR2_X1 U16321 ( .A(n14505), .B(n14510), .Z(n14506) );
  NOR2_X1 U16322 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14508), .ZN(n14511) );
  OAI21_X1 U16323 ( .B1(n14511), .B2(n14510), .A(n14509), .ZN(n14512) );
  XOR2_X1 U16324 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14512), .Z(n14513) );
  XNOR2_X1 U16325 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14513), .ZN(n14544) );
  INV_X1 U16326 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15424) );
  NAND2_X1 U16327 ( .A1(n14543), .A2(n14544), .ZN(n14542) );
  NOR2_X1 U16328 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14512), .ZN(n14515) );
  AND2_X1 U16329 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14513), .ZN(n14514) );
  NOR2_X1 U16330 ( .A1(n14515), .A2(n14514), .ZN(n14552) );
  XOR2_X1 U16331 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14551) );
  XNOR2_X1 U16332 ( .A(n14552), .B(n14551), .ZN(n14547) );
  XNOR2_X1 U16333 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14546), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16334 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14516) );
  OAI21_X1 U16335 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n14516), 
        .ZN(U28) );
  AOI21_X1 U16336 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14517) );
  OAI21_X1 U16337 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14517), 
        .ZN(U29) );
  AOI21_X1 U16338 ( .B1(n14520), .B2(n14519), .A(n14518), .ZN(n14522) );
  XNOR2_X1 U16339 ( .A(n14522), .B(n14521), .ZN(SUB_1596_U61) );
  XOR2_X1 U16340 ( .A(n14524), .B(n14523), .Z(SUB_1596_U57) );
  OAI22_X1 U16341 ( .A1(n14526), .A2(n11389), .B1(SI_15_), .B2(n14525), .ZN(
        n14527) );
  AOI21_X1 U16342 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n14528), .A(n14527), .ZN(
        P3_U3280) );
  XNOR2_X1 U16343 ( .A(n14529), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16344 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14530), .Z(SUB_1596_U54) );
  OAI21_X1 U16345 ( .B1(n14533), .B2(n14532), .A(n14531), .ZN(n14534) );
  XNOR2_X1 U16346 ( .A(n14534), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI21_X1 U16347 ( .B1(n14536), .B2(n14735), .A(n14535), .ZN(n14538) );
  AOI211_X1 U16348 ( .C1(n14721), .C2(n14539), .A(n14538), .B(n14537), .ZN(
        n14541) );
  INV_X1 U16349 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14540) );
  AOI22_X1 U16350 ( .A1(n14752), .A2(n14541), .B1(n14540), .B2(n14751), .ZN(
        P1_U3495) );
  AOI22_X1 U16351 ( .A1(n14759), .A2(n14541), .B1(n10200), .B2(n14757), .ZN(
        P1_U3540) );
  OAI21_X1 U16352 ( .B1(n14544), .B2(n14543), .A(n14542), .ZN(n14545) );
  XNOR2_X1 U16353 ( .A(n14545), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16354 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n14546), .ZN(n14550) );
  NOR2_X1 U16355 ( .A1(n14548), .A2(n14547), .ZN(n14549) );
  INV_X1 U16356 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14696) );
  NOR2_X1 U16357 ( .A1(n14552), .A2(n14551), .ZN(n14553) );
  AOI21_X1 U16358 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14696), .A(n14553), 
        .ZN(n14557) );
  XNOR2_X1 U16359 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(n14554), .ZN(n14555) );
  XNOR2_X1 U16360 ( .A(n7545), .B(n14555), .ZN(n14556) );
  XNOR2_X1 U16361 ( .A(n14557), .B(n14556), .ZN(n14558) );
  XNOR2_X1 U16362 ( .A(n14559), .B(n14558), .ZN(SUB_1596_U4) );
  OAI21_X1 U16363 ( .B1(n14561), .B2(n15172), .A(n14560), .ZN(n14568) );
  OAI22_X1 U16364 ( .A1(n15189), .A2(n14568), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15192), .ZN(n14562) );
  INV_X1 U16365 ( .A(n14562), .ZN(P3_U3489) );
  NOR2_X1 U16366 ( .A1(n15172), .A2(n14563), .ZN(n14565) );
  AOI211_X1 U16367 ( .C1(n15174), .C2(n14566), .A(n14565), .B(n14564), .ZN(
        n14570) );
  INV_X1 U16368 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U16369 ( .A1(n15192), .A2(n14570), .B1(n14567), .B2(n15189), .ZN(
        P3_U3470) );
  OAI22_X1 U16370 ( .A1(n15176), .A2(n14568), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n15177), .ZN(n14569) );
  INV_X1 U16371 ( .A(n14569), .ZN(P3_U3457) );
  AOI22_X1 U16372 ( .A1(n15177), .A2(n14570), .B1(n9256), .B2(n15176), .ZN(
        P3_U3423) );
  OAI21_X1 U16373 ( .B1(n14573), .B2(n14572), .A(n14571), .ZN(n14575) );
  AOI222_X1 U16374 ( .A1(n14578), .A2(n14589), .B1(n14577), .B2(n14576), .C1(
        n14575), .C2(n14574), .ZN(n14579) );
  NAND2_X1 U16375 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14867)
         );
  OAI211_X1 U16376 ( .C1(n14581), .C2(n14580), .A(n14579), .B(n14867), .ZN(
        P2_U3187) );
  OAI21_X1 U16377 ( .B1(n7210), .B2(n15018), .A(n14582), .ZN(n14584) );
  AOI211_X1 U16378 ( .C1(n15024), .C2(n14585), .A(n14584), .B(n14583), .ZN(
        n14607) );
  INV_X1 U16379 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14586) );
  AOI22_X1 U16380 ( .A1(n15037), .A2(n14607), .B1(n14586), .B2(n15035), .ZN(
        P2_U3514) );
  NAND3_X1 U16381 ( .A1(n14588), .A2(n14587), .A3(n15024), .ZN(n14593) );
  NAND2_X1 U16382 ( .A1(n14589), .A2(n14597), .ZN(n14590) );
  AND2_X1 U16383 ( .A1(n14591), .A2(n14590), .ZN(n14592) );
  AND2_X1 U16384 ( .A1(n14593), .A2(n14592), .ZN(n14595) );
  AOI22_X1 U16385 ( .A1(n15037), .A2(n14608), .B1(n14596), .B2(n15035), .ZN(
        P2_U3513) );
  NAND2_X1 U16386 ( .A1(n14598), .A2(n14597), .ZN(n14599) );
  NAND2_X1 U16387 ( .A1(n14600), .A2(n14599), .ZN(n14601) );
  NOR2_X1 U16388 ( .A1(n14602), .A2(n14601), .ZN(n14605) );
  NAND2_X1 U16389 ( .A1(n14603), .A2(n15024), .ZN(n14604) );
  AND2_X1 U16390 ( .A1(n14605), .A2(n14604), .ZN(n14610) );
  AOI22_X1 U16391 ( .A1(n15037), .A2(n14610), .B1(n11764), .B2(n15035), .ZN(
        P2_U3512) );
  INV_X1 U16392 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14606) );
  AOI22_X1 U16393 ( .A1(n15027), .A2(n14607), .B1(n14606), .B2(n15025), .ZN(
        P2_U3475) );
  INV_X1 U16394 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15475) );
  AOI22_X1 U16395 ( .A1(n15027), .A2(n14608), .B1(n15475), .B2(n15025), .ZN(
        P2_U3472) );
  INV_X1 U16396 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14609) );
  AOI22_X1 U16397 ( .A1(n15027), .A2(n14610), .B1(n14609), .B2(n15025), .ZN(
        P2_U3469) );
  XNOR2_X1 U16398 ( .A(n14612), .B(n14611), .ZN(n14614) );
  AOI222_X1 U16399 ( .A1(n14618), .A2(n14617), .B1(n14616), .B2(n14615), .C1(
        n14614), .C2(n14613), .ZN(n14620) );
  OAI211_X1 U16400 ( .C1(n14622), .C2(n14621), .A(n14620), .B(n14619), .ZN(
        P1_U3215) );
  OAI21_X1 U16401 ( .B1(n7071), .B2(n14735), .A(n14623), .ZN(n14624) );
  AOI211_X1 U16402 ( .C1(n14627), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        n14628) );
  AOI22_X1 U16403 ( .A1(n14759), .A2(n14628), .B1(n7887), .B2(n14757), .ZN(
        P1_U3542) );
  INV_X1 U16404 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15416) );
  AOI22_X1 U16405 ( .A1(n14752), .A2(n14628), .B1(n15416), .B2(n14751), .ZN(
        P1_U3501) );
  AOI21_X1 U16406 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14632) );
  XNOR2_X1 U16407 ( .A(n14632), .B(n14842), .ZN(SUB_1596_U69) );
  OAI21_X1 U16408 ( .B1(n14635), .B2(n14634), .A(n14633), .ZN(n14636) );
  XNOR2_X1 U16409 ( .A(n14636), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16410 ( .B1(n14639), .B2(n14638), .A(n14637), .ZN(n14640) );
  XNOR2_X1 U16411 ( .A(n14640), .B(n14857), .ZN(SUB_1596_U67) );
  AOI21_X1 U16412 ( .B1(n14643), .B2(n14642), .A(n14641), .ZN(n14644) );
  XNOR2_X1 U16413 ( .A(n14644), .B(n14869), .ZN(SUB_1596_U66) );
  NOR2_X1 U16414 ( .A1(n14646), .A2(n14645), .ZN(n14647) );
  XOR2_X1 U16415 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14647), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16416 ( .A1(n14649), .A2(n14648), .ZN(n14650) );
  XOR2_X1 U16417 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14650), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16418 ( .B1(n6586), .B2(n14652), .A(n14651), .ZN(n14654) );
  XNOR2_X1 U16419 ( .A(n14654), .B(P1_IR_REG_0__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16420 ( .A1(n14655), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14656) );
  OAI21_X1 U16421 ( .B1(n14658), .B2(n14657), .A(n14656), .ZN(P1_U3243) );
  AOI21_X1 U16422 ( .B1(n14660), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14659), 
        .ZN(n14664) );
  AOI21_X1 U16423 ( .B1(n14662), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14661), 
        .ZN(n14663) );
  OAI222_X1 U16424 ( .A1(n14691), .A2(n14665), .B1(n14689), .B2(n14664), .C1(
        n14687), .C2(n14663), .ZN(n14666) );
  INV_X1 U16425 ( .A(n14666), .ZN(n14668) );
  OAI211_X1 U16426 ( .C1(n14669), .C2(n14695), .A(n14668), .B(n14667), .ZN(
        P1_U3258) );
  INV_X1 U16427 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15428) );
  OAI21_X1 U16428 ( .B1(n14672), .B2(n14671), .A(n14670), .ZN(n14677) );
  OAI21_X1 U16429 ( .B1(n14675), .B2(n14674), .A(n14673), .ZN(n14676) );
  OAI222_X1 U16430 ( .A1(n14691), .A2(n14678), .B1(n14689), .B2(n14677), .C1(
        n14687), .C2(n14676), .ZN(n14679) );
  INV_X1 U16431 ( .A(n14679), .ZN(n14681) );
  OAI211_X1 U16432 ( .C1(n15428), .C2(n14695), .A(n14681), .B(n14680), .ZN(
        P1_U3260) );
  OAI21_X1 U16433 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n14683), .A(n14682), 
        .ZN(n14688) );
  OAI21_X1 U16434 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n14685), .A(n14684), 
        .ZN(n14686) );
  OAI222_X1 U16435 ( .A1(n14691), .A2(n14690), .B1(n14689), .B2(n14688), .C1(
        n14687), .C2(n14686), .ZN(n14692) );
  INV_X1 U16436 ( .A(n14692), .ZN(n14694) );
  OAI211_X1 U16437 ( .C1(n14696), .C2(n14695), .A(n14694), .B(n14693), .ZN(
        P1_U3261) );
  INV_X1 U16438 ( .A(n14697), .ZN(n14708) );
  INV_X1 U16439 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n14700) );
  OAI22_X1 U16440 ( .A1(n14225), .A2(n14700), .B1(n14699), .B2(n14698), .ZN(
        n14701) );
  AOI21_X1 U16441 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n14704) );
  OAI21_X1 U16442 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n14707) );
  AOI21_X1 U16443 ( .B1(n14709), .B2(n14708), .A(n14707), .ZN(n14710) );
  OAI21_X1 U16444 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(P1_U3286) );
  AND2_X1 U16445 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14714), .ZN(P1_U3294) );
  AND2_X1 U16446 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14714), .ZN(P1_U3295) );
  NOR2_X1 U16447 ( .A1(n14713), .A2(n15311), .ZN(P1_U3296) );
  AND2_X1 U16448 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14714), .ZN(P1_U3297) );
  AND2_X1 U16449 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14714), .ZN(P1_U3298) );
  NOR2_X1 U16450 ( .A1(n14713), .A2(n15459), .ZN(P1_U3299) );
  AND2_X1 U16451 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14714), .ZN(P1_U3300) );
  AND2_X1 U16452 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14714), .ZN(P1_U3301) );
  NOR2_X1 U16453 ( .A1(n14713), .A2(n15450), .ZN(P1_U3302) );
  AND2_X1 U16454 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14714), .ZN(P1_U3303) );
  AND2_X1 U16455 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14714), .ZN(P1_U3304) );
  AND2_X1 U16456 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14714), .ZN(P1_U3305) );
  AND2_X1 U16457 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14714), .ZN(P1_U3306) );
  AND2_X1 U16458 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14714), .ZN(P1_U3307) );
  AND2_X1 U16459 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14714), .ZN(P1_U3308) );
  AND2_X1 U16460 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14714), .ZN(P1_U3309) );
  AND2_X1 U16461 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14714), .ZN(P1_U3310) );
  AND2_X1 U16462 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14714), .ZN(P1_U3311) );
  AND2_X1 U16463 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14714), .ZN(P1_U3312) );
  AND2_X1 U16464 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14714), .ZN(P1_U3313) );
  NOR2_X1 U16465 ( .A1(n14713), .A2(n15270), .ZN(P1_U3314) );
  AND2_X1 U16466 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14714), .ZN(P1_U3315) );
  AND2_X1 U16467 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14714), .ZN(P1_U3316) );
  AND2_X1 U16468 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14714), .ZN(P1_U3317) );
  AND2_X1 U16469 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14714), .ZN(P1_U3318) );
  AND2_X1 U16470 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14714), .ZN(P1_U3319) );
  AND2_X1 U16471 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14714), .ZN(P1_U3320) );
  AND2_X1 U16472 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14714), .ZN(P1_U3321) );
  AND2_X1 U16473 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14714), .ZN(P1_U3322) );
  AND2_X1 U16474 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14714), .ZN(P1_U3323) );
  OAI21_X1 U16475 ( .B1(n14716), .B2(n14735), .A(n14715), .ZN(n14719) );
  INV_X1 U16476 ( .A(n14717), .ZN(n14718) );
  AOI211_X1 U16477 ( .C1(n14721), .C2(n14720), .A(n14719), .B(n14718), .ZN(
        n14753) );
  INV_X1 U16478 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14722) );
  AOI22_X1 U16479 ( .A1(n14752), .A2(n14753), .B1(n14722), .B2(n14751), .ZN(
        P1_U3465) );
  INV_X1 U16480 ( .A(n14724), .ZN(n14731) );
  NOR2_X1 U16481 ( .A1(n14724), .A2(n14723), .ZN(n14729) );
  OAI211_X1 U16482 ( .C1(n14727), .C2(n14735), .A(n14726), .B(n14725), .ZN(
        n14728) );
  AOI211_X1 U16483 ( .C1(n14731), .C2(n14730), .A(n14729), .B(n14728), .ZN(
        n14754) );
  INV_X1 U16484 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U16485 ( .A1(n14752), .A2(n14754), .B1(n14732), .B2(n14751), .ZN(
        P1_U3468) );
  OAI211_X1 U16486 ( .C1(n14736), .C2(n14735), .A(n14734), .B(n14733), .ZN(
        n14739) );
  NOR2_X1 U16487 ( .A1(n14737), .A2(n14749), .ZN(n14738) );
  AOI211_X1 U16488 ( .C1(n14741), .C2(n14740), .A(n14739), .B(n14738), .ZN(
        n14756) );
  INV_X1 U16489 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14742) );
  AOI22_X1 U16490 ( .A1(n14752), .A2(n14756), .B1(n14742), .B2(n14751), .ZN(
        P1_U3471) );
  AOI21_X1 U16491 ( .B1(n14745), .B2(n14744), .A(n14743), .ZN(n14746) );
  OAI211_X1 U16492 ( .C1(n14749), .C2(n14748), .A(n14747), .B(n14746), .ZN(
        n14750) );
  INV_X1 U16493 ( .A(n14750), .ZN(n14758) );
  INV_X1 U16494 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U16495 ( .A1(n14752), .A2(n14758), .B1(n15510), .B2(n14751), .ZN(
        P1_U3483) );
  AOI22_X1 U16496 ( .A1(n14759), .A2(n14753), .B1(n10046), .B2(n14757), .ZN(
        P1_U3530) );
  AOI22_X1 U16497 ( .A1(n14759), .A2(n14754), .B1(n10049), .B2(n14757), .ZN(
        P1_U3531) );
  AOI22_X1 U16498 ( .A1(n14759), .A2(n14756), .B1(n14755), .B2(n14757), .ZN(
        P1_U3532) );
  AOI22_X1 U16499 ( .A1(n14759), .A2(n14758), .B1(n10056), .B2(n14757), .ZN(
        P1_U3536) );
  NOR2_X1 U16500 ( .A1(n14760), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16501 ( .A1(n14760), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14774) );
  OAI211_X1 U16502 ( .C1(n14763), .C2(n14762), .A(n14922), .B(n14761), .ZN(
        n14770) );
  INV_X1 U16503 ( .A(n14764), .ZN(n14766) );
  NAND2_X1 U16504 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14765) );
  NAND2_X1 U16505 ( .A1(n14766), .A2(n14765), .ZN(n14767) );
  NAND3_X1 U16506 ( .A1(n14915), .A2(n14768), .A3(n14767), .ZN(n14769) );
  OAI211_X1 U16507 ( .C1(n14926), .C2(n14771), .A(n14770), .B(n14769), .ZN(
        n14772) );
  INV_X1 U16508 ( .A(n14772), .ZN(n14773) );
  NAND2_X1 U16509 ( .A1(n14774), .A2(n14773), .ZN(P2_U3215) );
  OAI211_X1 U16510 ( .C1(n14777), .C2(n14776), .A(n14915), .B(n14775), .ZN(
        n14782) );
  OAI211_X1 U16511 ( .C1(n14780), .C2(n14779), .A(n14922), .B(n14778), .ZN(
        n14781) );
  OAI211_X1 U16512 ( .C1(n14926), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        n14784) );
  INV_X1 U16513 ( .A(n14784), .ZN(n14786) );
  NAND2_X1 U16514 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14785) );
  OAI211_X1 U16515 ( .C1(n14930), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        P2_U3218) );
  INV_X1 U16516 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n14800) );
  OAI211_X1 U16517 ( .C1(n14790), .C2(n14789), .A(n14915), .B(n14788), .ZN(
        n14795) );
  OAI211_X1 U16518 ( .C1(n14793), .C2(n14792), .A(n14922), .B(n14791), .ZN(
        n14794) );
  OAI211_X1 U16519 ( .C1(n14926), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14797) );
  INV_X1 U16520 ( .A(n14797), .ZN(n14799) );
  NAND2_X1 U16521 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14798) );
  OAI211_X1 U16522 ( .C1(n14930), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        P2_U3219) );
  INV_X1 U16523 ( .A(n14801), .ZN(n14810) );
  OAI211_X1 U16524 ( .C1(n14804), .C2(n14803), .A(n14922), .B(n14802), .ZN(
        n14809) );
  OAI211_X1 U16525 ( .C1(n14807), .C2(n14806), .A(n14915), .B(n14805), .ZN(
        n14808) );
  OAI211_X1 U16526 ( .C1(n14926), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        n14811) );
  INV_X1 U16527 ( .A(n14811), .ZN(n14813) );
  OAI211_X1 U16528 ( .C1(n14930), .C2(n7057), .A(n14813), .B(n14812), .ZN(
        P2_U3220) );
  NAND2_X1 U16529 ( .A1(n14815), .A2(n14814), .ZN(n14816) );
  NAND3_X1 U16530 ( .A1(n14817), .A2(n14922), .A3(n14816), .ZN(n14823) );
  NAND2_X1 U16531 ( .A1(n14819), .A2(n14818), .ZN(n14820) );
  NAND3_X1 U16532 ( .A1(n14821), .A2(n14915), .A3(n14820), .ZN(n14822) );
  OAI211_X1 U16533 ( .C1(n14926), .C2(n14824), .A(n14823), .B(n14822), .ZN(
        n14825) );
  INV_X1 U16534 ( .A(n14825), .ZN(n14827) );
  OAI211_X1 U16535 ( .C1(n14828), .C2(n14930), .A(n14827), .B(n14826), .ZN(
        P2_U3224) );
  OAI211_X1 U16536 ( .C1(n14831), .C2(n14830), .A(n14829), .B(n14922), .ZN(
        n14832) );
  OAI21_X1 U16537 ( .B1(n14926), .B2(n14833), .A(n14832), .ZN(n14839) );
  NAND2_X1 U16538 ( .A1(n14835), .A2(n14834), .ZN(n14836) );
  AOI21_X1 U16539 ( .B1(n14837), .B2(n14836), .A(n14887), .ZN(n14838) );
  NOR2_X1 U16540 ( .A1(n14839), .A2(n14838), .ZN(n14841) );
  NAND2_X1 U16541 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14840)
         );
  OAI211_X1 U16542 ( .C1(n14842), .C2(n14930), .A(n14841), .B(n14840), .ZN(
        P2_U3225) );
  AOI21_X1 U16543 ( .B1(n14844), .B2(n14843), .A(n14887), .ZN(n14846) );
  NAND2_X1 U16544 ( .A1(n14846), .A2(n14845), .ZN(n14852) );
  AOI21_X1 U16545 ( .B1(n14848), .B2(n14847), .A(n14883), .ZN(n14850) );
  NAND2_X1 U16546 ( .A1(n14850), .A2(n14849), .ZN(n14851) );
  OAI211_X1 U16547 ( .C1(n14926), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        n14854) );
  INV_X1 U16548 ( .A(n14854), .ZN(n14856) );
  NAND2_X1 U16549 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14855)
         );
  OAI211_X1 U16550 ( .C1(n14857), .C2(n14930), .A(n14856), .B(n14855), .ZN(
        P2_U3227) );
  OAI211_X1 U16551 ( .C1(n14859), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14858), 
        .B(n14915), .ZN(n14864) );
  OAI211_X1 U16552 ( .C1(n14862), .C2(n14861), .A(n14860), .B(n14922), .ZN(
        n14863) );
  OAI211_X1 U16553 ( .C1(n14926), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        n14866) );
  INV_X1 U16554 ( .A(n14866), .ZN(n14868) );
  OAI211_X1 U16555 ( .C1(n14869), .C2(n14930), .A(n14868), .B(n14867), .ZN(
        P2_U3228) );
  INV_X1 U16556 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14882) );
  OAI21_X1 U16557 ( .B1(n14870), .B2(P2_REG2_REG_15__SCAN_IN), .A(n14915), 
        .ZN(n14871) );
  OR2_X1 U16558 ( .A1(n14872), .A2(n14871), .ZN(n14879) );
  OAI21_X1 U16559 ( .B1(n14873), .B2(P2_REG1_REG_15__SCAN_IN), .A(n14922), 
        .ZN(n14876) );
  OAI22_X1 U16560 ( .A1(n14876), .A2(n14875), .B1(n14874), .B2(n14926), .ZN(
        n14877) );
  INV_X1 U16561 ( .A(n14877), .ZN(n14878) );
  AND2_X1 U16562 ( .A1(n14879), .A2(n14878), .ZN(n14881) );
  NAND2_X1 U16563 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14880)
         );
  OAI211_X1 U16564 ( .C1(n14882), .C2(n14930), .A(n14881), .B(n14880), .ZN(
        P2_U3229) );
  INV_X1 U16565 ( .A(n14926), .ZN(n14894) );
  AOI211_X1 U16566 ( .C1(n14886), .C2(n14885), .A(n14884), .B(n14883), .ZN(
        n14892) );
  AOI211_X1 U16567 ( .C1(n14890), .C2(n14889), .A(n14888), .B(n14887), .ZN(
        n14891) );
  AOI211_X1 U16568 ( .C1(n14894), .C2(n14893), .A(n14892), .B(n14891), .ZN(
        n14896) );
  OAI211_X1 U16569 ( .C1(n6745), .C2(n14930), .A(n14896), .B(n14895), .ZN(
        P2_U3230) );
  NAND2_X1 U16570 ( .A1(n14898), .A2(n14897), .ZN(n14899) );
  NAND3_X1 U16571 ( .A1(n14915), .A2(n14900), .A3(n14899), .ZN(n14908) );
  INV_X1 U16572 ( .A(n14901), .ZN(n14904) );
  INV_X1 U16573 ( .A(n14902), .ZN(n14903) );
  NAND2_X1 U16574 ( .A1(n14904), .A2(n14903), .ZN(n14905) );
  NAND3_X1 U16575 ( .A1(n14922), .A2(n14906), .A3(n14905), .ZN(n14907) );
  OAI211_X1 U16576 ( .C1(n14926), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        n14910) );
  INV_X1 U16577 ( .A(n14910), .ZN(n14912) );
  OAI211_X1 U16578 ( .C1(n15424), .C2(n14930), .A(n14912), .B(n14911), .ZN(
        P2_U3231) );
  INV_X1 U16579 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14931) );
  OAI21_X1 U16580 ( .B1(n14914), .B2(n8265), .A(n14913), .ZN(n14916) );
  NAND2_X1 U16581 ( .A1(n14916), .A2(n14915), .ZN(n14924) );
  NAND2_X1 U16582 ( .A1(n14918), .A2(n14917), .ZN(n14921) );
  INV_X1 U16583 ( .A(n14919), .ZN(n14920) );
  NAND3_X1 U16584 ( .A1(n14922), .A2(n14921), .A3(n14920), .ZN(n14923) );
  OAI211_X1 U16585 ( .C1(n14926), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        n14927) );
  INV_X1 U16586 ( .A(n14927), .ZN(n14929) );
  OAI211_X1 U16587 ( .C1(n14931), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        P2_U3232) );
  XNOR2_X1 U16588 ( .A(n14932), .B(n14939), .ZN(n14934) );
  AOI21_X1 U16589 ( .B1(n14934), .B2(n14992), .A(n14933), .ZN(n15020) );
  INV_X1 U16590 ( .A(n14935), .ZN(n14936) );
  AOI222_X1 U16591 ( .A1(n14938), .A2(n14937), .B1(P2_REG2_REG_11__SCAN_IN), 
        .B2(n10410), .C1(n14948), .C2(n14936), .ZN(n14945) );
  XNOR2_X1 U16592 ( .A(n14940), .B(n14939), .ZN(n15023) );
  OAI211_X1 U16593 ( .C1(n15019), .C2(n14942), .A(n14997), .B(n14941), .ZN(
        n15017) );
  INV_X1 U16594 ( .A(n15017), .ZN(n14943) );
  AOI22_X1 U16595 ( .A1(n15023), .A2(n15196), .B1(n15195), .B2(n14943), .ZN(
        n14944) );
  OAI211_X1 U16596 ( .C1(n14957), .C2(n15020), .A(n14945), .B(n14944), .ZN(
        P2_U3254) );
  NAND2_X1 U16597 ( .A1(n14946), .A2(n15195), .ZN(n14950) );
  AOI22_X1 U16598 ( .A1(n14957), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14948), .ZN(n14949) );
  OAI211_X1 U16599 ( .C1(n14952), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14953) );
  AOI21_X1 U16600 ( .B1(n15196), .B2(n14954), .A(n14953), .ZN(n14955) );
  OAI21_X1 U16601 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(P2_U3263) );
  NOR2_X1 U16602 ( .A1(n14966), .A2(n14958), .ZN(n14959) );
  AND2_X1 U16603 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14960), .ZN(P2_U3266) );
  INV_X1 U16604 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15458) );
  NOR2_X1 U16605 ( .A1(n14959), .A2(n15458), .ZN(P2_U3267) );
  INV_X1 U16606 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15400) );
  NOR2_X1 U16607 ( .A1(n14959), .A2(n15400), .ZN(P2_U3268) );
  AND2_X1 U16608 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14960), .ZN(P2_U3269) );
  AND2_X1 U16609 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14960), .ZN(P2_U3270) );
  AND2_X1 U16610 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14960), .ZN(P2_U3271) );
  INV_X1 U16611 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15399) );
  NOR2_X1 U16612 ( .A1(n14959), .A2(n15399), .ZN(P2_U3272) );
  AND2_X1 U16613 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14960), .ZN(P2_U3273) );
  AND2_X1 U16614 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14960), .ZN(P2_U3274) );
  AND2_X1 U16615 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14960), .ZN(P2_U3275) );
  AND2_X1 U16616 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14960), .ZN(P2_U3276) );
  AND2_X1 U16617 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14960), .ZN(P2_U3277) );
  AND2_X1 U16618 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14960), .ZN(P2_U3278) );
  AND2_X1 U16619 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14960), .ZN(P2_U3279) );
  AND2_X1 U16620 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14960), .ZN(P2_U3280) );
  AND2_X1 U16621 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14960), .ZN(P2_U3281) );
  AND2_X1 U16622 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14960), .ZN(P2_U3282) );
  AND2_X1 U16623 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14960), .ZN(P2_U3283) );
  AND2_X1 U16624 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14960), .ZN(P2_U3284) );
  AND2_X1 U16625 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14960), .ZN(P2_U3285) );
  AND2_X1 U16626 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14960), .ZN(P2_U3286) );
  AND2_X1 U16627 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14960), .ZN(P2_U3287) );
  AND2_X1 U16628 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14960), .ZN(P2_U3288) );
  AND2_X1 U16629 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14960), .ZN(P2_U3289) );
  AND2_X1 U16630 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14960), .ZN(P2_U3290) );
  AND2_X1 U16631 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14960), .ZN(P2_U3291) );
  AND2_X1 U16632 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14960), .ZN(P2_U3292) );
  AND2_X1 U16633 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14960), .ZN(P2_U3293) );
  AND2_X1 U16634 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14960), .ZN(P2_U3294) );
  AND2_X1 U16635 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14960), .ZN(P2_U3295) );
  AOI22_X1 U16636 ( .A1(n14963), .A2(n14962), .B1(n14961), .B2(n14966), .ZN(
        P2_U3416) );
  INV_X1 U16637 ( .A(n14964), .ZN(n14965) );
  AOI21_X1 U16638 ( .B1(n14966), .B2(n15487), .A(n14965), .ZN(P2_U3417) );
  INV_X1 U16639 ( .A(n14967), .ZN(n14973) );
  OAI22_X1 U16640 ( .A1(n14971), .A2(n14970), .B1(n14969), .B2(n14968), .ZN(
        n14972) );
  NOR2_X1 U16641 ( .A1(n14973), .A2(n14972), .ZN(n15028) );
  AOI22_X1 U16642 ( .A1(n15027), .A2(n15028), .B1(n8281), .B2(n15025), .ZN(
        P2_U3430) );
  INV_X1 U16643 ( .A(n14981), .ZN(n14975) );
  NOR2_X1 U16644 ( .A1(n14975), .A2(n14974), .ZN(n14980) );
  OAI211_X1 U16645 ( .C1(n14978), .C2(n15018), .A(n14977), .B(n14976), .ZN(
        n14979) );
  AOI211_X1 U16646 ( .C1(n14981), .C2(n15006), .A(n14980), .B(n14979), .ZN(
        n15029) );
  INV_X1 U16647 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U16648 ( .A1(n15027), .A2(n15029), .B1(n14982), .B2(n15025), .ZN(
        P2_U3445) );
  OAI22_X1 U16649 ( .A1(n14984), .A2(n13202), .B1(n7208), .B2(n15018), .ZN(
        n14985) );
  AOI21_X1 U16650 ( .B1(n14986), .B2(n15006), .A(n14985), .ZN(n14987) );
  AND2_X1 U16651 ( .A1(n14988), .A2(n14987), .ZN(n15030) );
  INV_X1 U16652 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U16653 ( .A1(n15027), .A2(n15030), .B1(n14989), .B2(n15025), .ZN(
        P2_U3448) );
  XNOR2_X1 U16654 ( .A(n14991), .B(n14990), .ZN(n14993) );
  NAND2_X1 U16655 ( .A1(n14993), .A2(n14992), .ZN(n14995) );
  NAND2_X1 U16656 ( .A1(n14995), .A2(n14994), .ZN(n15198) );
  OAI211_X1 U16657 ( .C1(n15201), .C2(n7209), .A(n14997), .B(n14996), .ZN(
        n15193) );
  OAI21_X1 U16658 ( .B1(n15201), .B2(n15018), .A(n15193), .ZN(n14998) );
  NOR2_X1 U16659 ( .A1(n15198), .A2(n14998), .ZN(n15002) );
  XNOR2_X1 U16660 ( .A(n15000), .B(n14999), .ZN(n15197) );
  NAND2_X1 U16661 ( .A1(n15197), .A2(n15024), .ZN(n15001) );
  AND2_X1 U16662 ( .A1(n15002), .A2(n15001), .ZN(n15031) );
  INV_X1 U16663 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15479) );
  AOI22_X1 U16664 ( .A1(n15027), .A2(n15031), .B1(n15479), .B2(n15025), .ZN(
        P2_U3451) );
  OAI21_X1 U16665 ( .B1(n7207), .B2(n15018), .A(n15004), .ZN(n15005) );
  AOI21_X1 U16666 ( .B1(n15007), .B2(n15006), .A(n15005), .ZN(n15008) );
  AND2_X1 U16667 ( .A1(n15009), .A2(n15008), .ZN(n15033) );
  INV_X1 U16668 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15010) );
  AOI22_X1 U16669 ( .A1(n15027), .A2(n15033), .B1(n15010), .B2(n15025), .ZN(
        P2_U3454) );
  OAI211_X1 U16670 ( .C1(n15013), .C2(n15018), .A(n15012), .B(n15011), .ZN(
        n15014) );
  AOI21_X1 U16671 ( .B1(n15024), .B2(n15015), .A(n15014), .ZN(n15034) );
  INV_X1 U16672 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U16673 ( .A1(n15027), .A2(n15034), .B1(n15016), .B2(n15025), .ZN(
        P2_U3460) );
  OAI21_X1 U16674 ( .B1(n15019), .B2(n15018), .A(n15017), .ZN(n15022) );
  INV_X1 U16675 ( .A(n15020), .ZN(n15021) );
  AOI211_X1 U16676 ( .C1(n15024), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15036) );
  INV_X1 U16677 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U16678 ( .A1(n15027), .A2(n15036), .B1(n15026), .B2(n15025), .ZN(
        P2_U3463) );
  AOI22_X1 U16679 ( .A1(n15037), .A2(n15028), .B1(n8289), .B2(n15035), .ZN(
        P2_U3499) );
  AOI22_X1 U16680 ( .A1(n15037), .A2(n15029), .B1(n10091), .B2(n15035), .ZN(
        P2_U3504) );
  AOI22_X1 U16681 ( .A1(n15037), .A2(n15030), .B1(n15443), .B2(n15035), .ZN(
        P2_U3505) );
  AOI22_X1 U16682 ( .A1(n15037), .A2(n15031), .B1(n15444), .B2(n15035), .ZN(
        P2_U3506) );
  AOI22_X1 U16683 ( .A1(n15037), .A2(n15033), .B1(n15032), .B2(n15035), .ZN(
        P2_U3507) );
  AOI22_X1 U16684 ( .A1(n15037), .A2(n15034), .B1(n10280), .B2(n15035), .ZN(
        P2_U3509) );
  AOI22_X1 U16685 ( .A1(n15037), .A2(n15036), .B1(n15387), .B2(n15035), .ZN(
        P2_U3510) );
  NOR2_X1 U16686 ( .A1(P3_U3897), .A2(n15093), .ZN(P3_U3150) );
  INV_X1 U16687 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U16688 ( .A1(n15038), .A2(n9601), .ZN(n15042) );
  NAND2_X1 U16689 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  OAI211_X1 U16690 ( .C1(n15044), .C2(n15043), .A(n15042), .B(n15041), .ZN(
        n15045) );
  INV_X1 U16691 ( .A(n15045), .ZN(n15046) );
  OAI21_X1 U16692 ( .B1(n15048), .B2(n15047), .A(n15046), .ZN(P3_U3172) );
  AOI21_X1 U16693 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(n15057) );
  OAI21_X1 U16694 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15055) );
  NAND2_X1 U16695 ( .A1(n15080), .A2(n15055), .ZN(n15056) );
  OAI21_X1 U16696 ( .B1(n15103), .B2(n15057), .A(n15056), .ZN(n15064) );
  OR3_X1 U16697 ( .A1(n15060), .A2(n15059), .A3(n15058), .ZN(n15061) );
  AOI21_X1 U16698 ( .B1(n15062), .B2(n15061), .A(n15071), .ZN(n15063) );
  AOI211_X1 U16699 ( .C1(n15097), .C2(n15065), .A(n15064), .B(n15063), .ZN(
        n15067) );
  OAI211_X1 U16700 ( .C1(n15068), .C2(n15088), .A(n15067), .B(n15066), .ZN(
        P3_U3188) );
  INV_X1 U16701 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15089) );
  AOI21_X1 U16702 ( .B1(n6728), .B2(n15070), .A(n15069), .ZN(n15072) );
  NOR2_X1 U16703 ( .A1(n15072), .A2(n15071), .ZN(n15085) );
  AOI21_X1 U16704 ( .B1(n15075), .B2(n15074), .A(n15073), .ZN(n15083) );
  OAI21_X1 U16705 ( .B1(n15078), .B2(n15077), .A(n15076), .ZN(n15079) );
  AOI22_X1 U16706 ( .A1(n15097), .A2(n15081), .B1(n15080), .B2(n15079), .ZN(
        n15082) );
  OAI21_X1 U16707 ( .B1(n15083), .B2(n15103), .A(n15082), .ZN(n15084) );
  NOR2_X1 U16708 ( .A1(n15085), .A2(n15084), .ZN(n15087) );
  OAI211_X1 U16709 ( .C1(n15089), .C2(n15088), .A(n15087), .B(n15086), .ZN(
        P3_U3190) );
  OAI21_X1 U16710 ( .B1(n15092), .B2(n15091), .A(n15090), .ZN(n15094) );
  AOI22_X1 U16711 ( .A1(n15094), .A2(n15080), .B1(n15093), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n15108) );
  XNOR2_X1 U16712 ( .A(n15096), .B(n15095), .ZN(n15100) );
  AOI22_X1 U16713 ( .A1(n15100), .A2(n15099), .B1(n15098), .B2(n15097), .ZN(
        n15107) );
  AOI21_X1 U16714 ( .B1(n6727), .B2(n15102), .A(n15101), .ZN(n15104) );
  OR2_X1 U16715 ( .A1(n15104), .A2(n15103), .ZN(n15105) );
  NAND4_X1 U16716 ( .A1(n15108), .A2(n15107), .A3(n15106), .A4(n15105), .ZN(
        P3_U3192) );
  XNOR2_X1 U16717 ( .A(n15113), .B(n15109), .ZN(n15132) );
  INV_X1 U16718 ( .A(n15110), .ZN(n15121) );
  OAI21_X1 U16719 ( .B1(n15113), .B2(n15112), .A(n15111), .ZN(n15115) );
  NAND2_X1 U16720 ( .A1(n15115), .A2(n15114), .ZN(n15119) );
  NAND2_X1 U16721 ( .A1(n15117), .A2(n15116), .ZN(n15118) );
  OAI211_X1 U16722 ( .C1(n15121), .C2(n15120), .A(n15119), .B(n15118), .ZN(
        n15130) );
  NOR2_X1 U16723 ( .A1(n15172), .A2(n15122), .ZN(n15131) );
  INV_X1 U16724 ( .A(n15131), .ZN(n15125) );
  OAI22_X1 U16725 ( .A1(n15125), .A2(n15124), .B1(n15403), .B2(n15123), .ZN(
        n15126) );
  AOI211_X1 U16726 ( .C1(n15127), .C2(n15132), .A(n15130), .B(n15126), .ZN(
        n15128) );
  AOI22_X1 U16727 ( .A1(n15129), .A2(n9081), .B1(n15128), .B2(n6576), .ZN(
        P3_U3232) );
  AOI211_X1 U16728 ( .C1(n15174), .C2(n15132), .A(n15131), .B(n15130), .ZN(
        n15178) );
  AOI22_X1 U16729 ( .A1(n15177), .A2(n15178), .B1(n9080), .B2(n15176), .ZN(
        P3_U3393) );
  INV_X1 U16730 ( .A(n15133), .ZN(n15136) );
  INV_X1 U16731 ( .A(n15134), .ZN(n15135) );
  AOI211_X1 U16732 ( .C1(n15156), .C2(n15137), .A(n15136), .B(n15135), .ZN(
        n15179) );
  AOI22_X1 U16733 ( .A1(n15177), .A2(n15179), .B1(n9086), .B2(n15176), .ZN(
        P3_U3396) );
  OAI22_X1 U16734 ( .A1(n15139), .A2(n15166), .B1(n15172), .B2(n15138), .ZN(
        n15140) );
  NOR2_X1 U16735 ( .A1(n15141), .A2(n15140), .ZN(n15180) );
  AOI22_X1 U16736 ( .A1(n15177), .A2(n15180), .B1(n9110), .B2(n15176), .ZN(
        P3_U3399) );
  NOR2_X1 U16737 ( .A1(n15172), .A2(n15142), .ZN(n15144) );
  AOI211_X1 U16738 ( .C1(n15156), .C2(n15145), .A(n15144), .B(n15143), .ZN(
        n15181) );
  AOI22_X1 U16739 ( .A1(n15177), .A2(n15181), .B1(n9120), .B2(n15176), .ZN(
        P3_U3402) );
  OAI22_X1 U16740 ( .A1(n15147), .A2(n15166), .B1(n15172), .B2(n15146), .ZN(
        n15149) );
  NOR2_X1 U16741 ( .A1(n15149), .A2(n15148), .ZN(n15183) );
  AOI22_X1 U16742 ( .A1(n15177), .A2(n15183), .B1(n9144), .B2(n15176), .ZN(
        P3_U3405) );
  OAI22_X1 U16743 ( .A1(n15151), .A2(n15166), .B1(n15150), .B2(n15172), .ZN(
        n15152) );
  NOR2_X1 U16744 ( .A1(n15153), .A2(n15152), .ZN(n15184) );
  AOI22_X1 U16745 ( .A1(n15177), .A2(n15184), .B1(n9162), .B2(n15176), .ZN(
        P3_U3408) );
  AOI22_X1 U16746 ( .A1(n15157), .A2(n15156), .B1(n15155), .B2(n15154), .ZN(
        n15158) );
  AND2_X1 U16747 ( .A1(n15159), .A2(n15158), .ZN(n15185) );
  AOI22_X1 U16748 ( .A1(n15177), .A2(n15185), .B1(n9173), .B2(n15176), .ZN(
        P3_U3411) );
  OAI22_X1 U16749 ( .A1(n15161), .A2(n15166), .B1(n15160), .B2(n15172), .ZN(
        n15163) );
  NOR2_X1 U16750 ( .A1(n15163), .A2(n15162), .ZN(n15187) );
  INV_X1 U16751 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U16752 ( .A1(n15177), .A2(n15187), .B1(n15164), .B2(n15176), .ZN(
        P3_U3414) );
  OAI22_X1 U16753 ( .A1(n15167), .A2(n15166), .B1(n15172), .B2(n15165), .ZN(
        n15168) );
  NOR2_X1 U16754 ( .A1(n15169), .A2(n15168), .ZN(n15188) );
  AOI22_X1 U16755 ( .A1(n15177), .A2(n15188), .B1(n9213), .B2(n15176), .ZN(
        P3_U3417) );
  OAI21_X1 U16756 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(n15173) );
  AOI21_X1 U16757 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(n15191) );
  AOI22_X1 U16758 ( .A1(n15177), .A2(n15191), .B1(n9230), .B2(n15176), .ZN(
        P3_U3420) );
  AOI22_X1 U16759 ( .A1(n15192), .A2(n15178), .B1(n10669), .B2(n15189), .ZN(
        P3_U3460) );
  AOI22_X1 U16760 ( .A1(n15192), .A2(n15179), .B1(n10666), .B2(n15189), .ZN(
        P3_U3461) );
  INV_X1 U16761 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U16762 ( .A1(n15192), .A2(n15180), .B1(n15352), .B2(n15189), .ZN(
        P3_U3462) );
  AOI22_X1 U16763 ( .A1(n15192), .A2(n15181), .B1(n11103), .B2(n15189), .ZN(
        P3_U3463) );
  AOI22_X1 U16764 ( .A1(n15192), .A2(n15183), .B1(n15182), .B2(n15189), .ZN(
        P3_U3464) );
  AOI22_X1 U16765 ( .A1(n15192), .A2(n15184), .B1(n11145), .B2(n15189), .ZN(
        P3_U3465) );
  AOI22_X1 U16766 ( .A1(n15192), .A2(n15185), .B1(n11150), .B2(n15189), .ZN(
        P3_U3466) );
  AOI22_X1 U16767 ( .A1(n15192), .A2(n15187), .B1(n15186), .B2(n15189), .ZN(
        P3_U3467) );
  AOI22_X1 U16768 ( .A1(n15192), .A2(n15188), .B1(n11206), .B2(n15189), .ZN(
        P3_U3468) );
  AOI22_X1 U16769 ( .A1(n15192), .A2(n15191), .B1(n15190), .B2(n15189), .ZN(
        P3_U3469) );
  INV_X1 U16770 ( .A(n15193), .ZN(n15194) );
  AOI22_X1 U16771 ( .A1(n15197), .A2(n15196), .B1(n15195), .B2(n15194), .ZN(
        n15205) );
  MUX2_X1 U16772 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n15198), .S(n13512), .Z(
        n15203) );
  OAI22_X1 U16773 ( .A1(n15201), .A2(n14951), .B1(n15200), .B2(n15199), .ZN(
        n15202) );
  NOR2_X1 U16774 ( .A1(n15203), .A2(n15202), .ZN(n15204) );
  NAND2_X1 U16775 ( .A1(n15205), .A2(n15204), .ZN(n15512) );
  NAND2_X1 U16776 ( .A1(keyinput51), .A2(keyinput110), .ZN(n15206) );
  NOR3_X1 U16777 ( .A1(keyinput53), .A2(keyinput25), .A3(n15206), .ZN(n15207)
         );
  NAND4_X1 U16778 ( .A1(keyinput28), .A2(keyinput49), .A3(keyinput127), .A4(
        n15207), .ZN(n15219) );
  NOR2_X1 U16779 ( .A1(keyinput68), .A2(keyinput95), .ZN(n15208) );
  NAND3_X1 U16780 ( .A1(keyinput121), .A2(keyinput104), .A3(n15208), .ZN(
        n15218) );
  NAND4_X1 U16781 ( .A1(keyinput22), .A2(keyinput81), .A3(keyinput112), .A4(
        keyinput7), .ZN(n15217) );
  NAND2_X1 U16782 ( .A1(keyinput45), .A2(keyinput85), .ZN(n15209) );
  NOR3_X1 U16783 ( .A1(keyinput11), .A2(keyinput12), .A3(n15209), .ZN(n15215)
         );
  NOR4_X1 U16784 ( .A1(keyinput42), .A2(keyinput33), .A3(keyinput71), .A4(
        keyinput86), .ZN(n15214) );
  INV_X1 U16785 ( .A(keyinput107), .ZN(n15210) );
  NOR4_X1 U16786 ( .A1(keyinput2), .A2(keyinput103), .A3(keyinput9), .A4(
        n15210), .ZN(n15213) );
  NAND3_X1 U16787 ( .A1(keyinput37), .A2(keyinput66), .A3(keyinput69), .ZN(
        n15211) );
  NOR2_X1 U16788 ( .A1(keyinput118), .A2(n15211), .ZN(n15212) );
  NAND4_X1 U16789 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        n15216) );
  NOR4_X1 U16790 ( .A1(n15219), .A2(n15218), .A3(n15217), .A4(n15216), .ZN(
        n15268) );
  NAND2_X1 U16791 ( .A1(keyinput102), .A2(keyinput19), .ZN(n15220) );
  NOR3_X1 U16792 ( .A1(keyinput113), .A2(keyinput40), .A3(n15220), .ZN(n15221)
         );
  NAND3_X1 U16793 ( .A1(keyinput1), .A2(keyinput31), .A3(n15221), .ZN(n15235)
         );
  INV_X1 U16794 ( .A(keyinput47), .ZN(n15222) );
  NOR4_X1 U16795 ( .A1(keyinput65), .A2(keyinput92), .A3(keyinput38), .A4(
        n15222), .ZN(n15233) );
  NAND2_X1 U16796 ( .A1(keyinput82), .A2(keyinput79), .ZN(n15223) );
  NOR3_X1 U16797 ( .A1(keyinput16), .A2(keyinput57), .A3(n15223), .ZN(n15232)
         );
  NOR2_X1 U16798 ( .A1(keyinput119), .A2(keyinput41), .ZN(n15224) );
  NAND3_X1 U16799 ( .A1(keyinput123), .A2(keyinput56), .A3(n15224), .ZN(n15230) );
  INV_X1 U16800 ( .A(keyinput23), .ZN(n15225) );
  NAND4_X1 U16801 ( .A1(keyinput10), .A2(keyinput88), .A3(keyinput100), .A4(
        n15225), .ZN(n15229) );
  NAND4_X1 U16802 ( .A1(keyinput78), .A2(keyinput109), .A3(keyinput126), .A4(
        keyinput83), .ZN(n15228) );
  NOR2_X1 U16803 ( .A1(keyinput14), .A2(keyinput44), .ZN(n15226) );
  NAND3_X1 U16804 ( .A1(keyinput97), .A2(keyinput101), .A3(n15226), .ZN(n15227) );
  NOR4_X1 U16805 ( .A1(n15230), .A2(n15229), .A3(n15228), .A4(n15227), .ZN(
        n15231) );
  NAND3_X1 U16806 ( .A1(n15233), .A2(n15232), .A3(n15231), .ZN(n15234) );
  NOR4_X1 U16807 ( .A1(keyinput39), .A2(keyinput72), .A3(n15235), .A4(n15234), 
        .ZN(n15267) );
  NAND2_X1 U16808 ( .A1(keyinput76), .A2(keyinput35), .ZN(n15236) );
  NOR3_X1 U16809 ( .A1(keyinput94), .A2(keyinput61), .A3(n15236), .ZN(n15237)
         );
  NAND3_X1 U16810 ( .A1(keyinput27), .A2(keyinput73), .A3(n15237), .ZN(n15248)
         );
  NAND4_X1 U16811 ( .A1(keyinput90), .A2(keyinput29), .A3(keyinput6), .A4(
        keyinput32), .ZN(n15238) );
  NOR3_X1 U16812 ( .A1(keyinput26), .A2(keyinput17), .A3(n15238), .ZN(n15246)
         );
  INV_X1 U16813 ( .A(keyinput98), .ZN(n15239) );
  NAND4_X1 U16814 ( .A1(keyinput93), .A2(keyinput116), .A3(keyinput125), .A4(
        n15239), .ZN(n15244) );
  NAND4_X1 U16815 ( .A1(keyinput0), .A2(keyinput87), .A3(keyinput43), .A4(
        keyinput46), .ZN(n15243) );
  NOR2_X1 U16816 ( .A1(keyinput36), .A2(keyinput24), .ZN(n15240) );
  NAND3_X1 U16817 ( .A1(keyinput115), .A2(keyinput50), .A3(n15240), .ZN(n15242) );
  OR4_X1 U16818 ( .A1(keyinput84), .A2(keyinput114), .A3(keyinput62), .A4(
        keyinput120), .ZN(n15241) );
  NOR4_X1 U16819 ( .A1(n15244), .A2(n15243), .A3(n15242), .A4(n15241), .ZN(
        n15245) );
  NAND4_X1 U16820 ( .A1(keyinput75), .A2(keyinput5), .A3(n15246), .A4(n15245), 
        .ZN(n15247) );
  NOR4_X1 U16821 ( .A1(keyinput21), .A2(keyinput99), .A3(n15248), .A4(n15247), 
        .ZN(n15266) );
  NOR2_X1 U16822 ( .A1(keyinput96), .A2(keyinput4), .ZN(n15249) );
  NAND3_X1 U16823 ( .A1(keyinput70), .A2(keyinput34), .A3(n15249), .ZN(n15264)
         );
  INV_X1 U16824 ( .A(keyinput48), .ZN(n15250) );
  NAND4_X1 U16825 ( .A1(keyinput77), .A2(keyinput67), .A3(keyinput30), .A4(
        n15250), .ZN(n15263) );
  NOR2_X1 U16826 ( .A1(keyinput58), .A2(keyinput52), .ZN(n15251) );
  NAND3_X1 U16827 ( .A1(keyinput89), .A2(keyinput111), .A3(n15251), .ZN(n15252) );
  NOR3_X1 U16828 ( .A1(keyinput64), .A2(keyinput54), .A3(n15252), .ZN(n15253)
         );
  NAND3_X1 U16829 ( .A1(keyinput122), .A2(keyinput15), .A3(n15253), .ZN(n15262) );
  NOR4_X1 U16830 ( .A1(keyinput80), .A2(keyinput55), .A3(keyinput20), .A4(
        keyinput106), .ZN(n15260) );
  NAND3_X1 U16831 ( .A1(keyinput105), .A2(keyinput63), .A3(keyinput59), .ZN(
        n15254) );
  NOR2_X1 U16832 ( .A1(keyinput108), .A2(n15254), .ZN(n15259) );
  INV_X1 U16833 ( .A(keyinput124), .ZN(n15255) );
  NOR4_X1 U16834 ( .A1(keyinput117), .A2(keyinput8), .A3(keyinput60), .A4(
        n15255), .ZN(n15258) );
  NAND2_X1 U16835 ( .A1(keyinput3), .A2(keyinput91), .ZN(n15256) );
  NOR3_X1 U16836 ( .A1(keyinput18), .A2(keyinput74), .A3(n15256), .ZN(n15257)
         );
  NAND4_X1 U16837 ( .A1(n15260), .A2(n15259), .A3(n15258), .A4(n15257), .ZN(
        n15261) );
  NOR4_X1 U16838 ( .A1(n15264), .A2(n15263), .A3(n15262), .A4(n15261), .ZN(
        n15265) );
  NAND4_X1 U16839 ( .A1(n15268), .A2(n15267), .A3(n15266), .A4(n15265), .ZN(
        n15509) );
  AOI22_X1 U16840 ( .A1(n15271), .A2(keyinput29), .B1(keyinput6), .B2(n15270), 
        .ZN(n15269) );
  OAI221_X1 U16841 ( .B1(n15271), .B2(keyinput29), .C1(n15270), .C2(keyinput6), 
        .A(n15269), .ZN(n15282) );
  INV_X1 U16842 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U16843 ( .A1(n15274), .A2(keyinput32), .B1(n15273), .B2(keyinput0), 
        .ZN(n15272) );
  OAI221_X1 U16844 ( .B1(n15274), .B2(keyinput32), .C1(n15273), .C2(keyinput0), 
        .A(n15272), .ZN(n15281) );
  INV_X1 U16845 ( .A(SI_27_), .ZN(n15275) );
  XOR2_X1 U16846 ( .A(n15275), .B(keyinput5), .Z(n15279) );
  XNOR2_X1 U16847 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput26), .ZN(n15278) );
  XNOR2_X1 U16848 ( .A(P2_REG0_REG_26__SCAN_IN), .B(keyinput17), .ZN(n15277)
         );
  XNOR2_X1 U16849 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput90), .ZN(n15276) );
  NAND4_X1 U16850 ( .A1(n15279), .A2(n15278), .A3(n15277), .A4(n15276), .ZN(
        n15280) );
  NOR3_X1 U16851 ( .A1(n15282), .A2(n15281), .A3(n15280), .ZN(n15323) );
  INV_X1 U16852 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15284) );
  AOI22_X1 U16853 ( .A1(n15285), .A2(keyinput46), .B1(keyinput98), .B2(n15284), 
        .ZN(n15283) );
  OAI221_X1 U16854 ( .B1(n15285), .B2(keyinput46), .C1(n15284), .C2(keyinput98), .A(n15283), .ZN(n15294) );
  XNOR2_X1 U16855 ( .A(n15286), .B(keyinput84), .ZN(n15293) );
  XNOR2_X1 U16856 ( .A(keyinput125), .B(n10200), .ZN(n15292) );
  XNOR2_X1 U16857 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput43), .ZN(n15290)
         );
  XNOR2_X1 U16858 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput87), .ZN(n15289) );
  XNOR2_X1 U16859 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput93), .ZN(n15288) );
  XNOR2_X1 U16860 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput116), .ZN(n15287)
         );
  NAND4_X1 U16861 ( .A1(n15290), .A2(n15289), .A3(n15288), .A4(n15287), .ZN(
        n15291) );
  NOR4_X1 U16862 ( .A1(n15294), .A2(n15293), .A3(n15292), .A4(n15291), .ZN(
        n15322) );
  AOI22_X1 U16863 ( .A1(n15296), .A2(keyinput120), .B1(n12680), .B2(keyinput35), .ZN(n15295) );
  OAI221_X1 U16864 ( .B1(n15296), .B2(keyinput120), .C1(n12680), .C2(
        keyinput35), .A(n15295), .ZN(n15306) );
  AOI22_X1 U16865 ( .A1(n15299), .A2(keyinput50), .B1(keyinput62), .B2(n15298), 
        .ZN(n15297) );
  OAI221_X1 U16866 ( .B1(n15299), .B2(keyinput50), .C1(n15298), .C2(keyinput62), .A(n15297), .ZN(n15305) );
  XNOR2_X1 U16867 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput115), .ZN(n15303) );
  XNOR2_X1 U16868 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput114), .ZN(n15302) );
  XNOR2_X1 U16869 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput36), .ZN(n15301)
         );
  XNOR2_X1 U16870 ( .A(keyinput24), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n15300) );
  NAND4_X1 U16871 ( .A1(n15303), .A2(n15302), .A3(n15301), .A4(n15300), .ZN(
        n15304) );
  NOR3_X1 U16872 ( .A1(n15306), .A2(n15305), .A3(n15304), .ZN(n15321) );
  AOI22_X1 U16873 ( .A1(n15308), .A2(keyinput99), .B1(keyinput27), .B2(n11760), 
        .ZN(n15307) );
  OAI221_X1 U16874 ( .B1(n15308), .B2(keyinput99), .C1(n11760), .C2(keyinput27), .A(n15307), .ZN(n15319) );
  INV_X1 U16875 ( .A(keyinput67), .ZN(n15310) );
  AOI22_X1 U16876 ( .A1(n15311), .A2(keyinput73), .B1(P3_DATAO_REG_2__SCAN_IN), 
        .B2(n15310), .ZN(n15309) );
  OAI221_X1 U16877 ( .B1(n15311), .B2(keyinput73), .C1(n15310), .C2(
        P3_DATAO_REG_2__SCAN_IN), .A(n15309), .ZN(n15318) );
  INV_X1 U16878 ( .A(keyinput61), .ZN(n15312) );
  XOR2_X1 U16879 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n15312), .Z(n15316) );
  XNOR2_X1 U16880 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput94), .ZN(n15315)
         );
  XNOR2_X1 U16881 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput21), .ZN(n15314)
         );
  XNOR2_X1 U16882 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput76), .ZN(n15313) );
  NAND4_X1 U16883 ( .A1(n15316), .A2(n15315), .A3(n15314), .A4(n15313), .ZN(
        n15317) );
  NOR3_X1 U16884 ( .A1(n15319), .A2(n15318), .A3(n15317), .ZN(n15320) );
  NAND4_X1 U16885 ( .A1(n15323), .A2(n15322), .A3(n15321), .A4(n15320), .ZN(
        n15507) );
  AOI22_X1 U16886 ( .A1(n15326), .A2(keyinput70), .B1(keyinput34), .B2(n15325), 
        .ZN(n15324) );
  OAI221_X1 U16887 ( .B1(n15326), .B2(keyinput70), .C1(n15325), .C2(keyinput34), .A(n15324), .ZN(n15337) );
  AOI22_X1 U16888 ( .A1(n7692), .A2(keyinput30), .B1(n15328), .B2(keyinput96), 
        .ZN(n15327) );
  OAI221_X1 U16889 ( .B1(n7692), .B2(keyinput30), .C1(n15328), .C2(keyinput96), 
        .A(n15327), .ZN(n15336) );
  AOI22_X1 U16890 ( .A1(n15331), .A2(keyinput77), .B1(n15330), .B2(keyinput48), 
        .ZN(n15329) );
  OAI221_X1 U16891 ( .B1(n15331), .B2(keyinput77), .C1(n15330), .C2(keyinput48), .A(n15329), .ZN(n15335) );
  XNOR2_X1 U16892 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput64), .ZN(n15333) );
  XNOR2_X1 U16893 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput4), .ZN(n15332) );
  NAND2_X1 U16894 ( .A1(n15333), .A2(n15332), .ZN(n15334) );
  NOR4_X1 U16895 ( .A1(n15337), .A2(n15336), .A3(n15335), .A4(n15334), .ZN(
        n15383) );
  AOI22_X1 U16896 ( .A1(n15339), .A2(keyinput52), .B1(keyinput122), .B2(n11010), .ZN(n15338) );
  OAI221_X1 U16897 ( .B1(n15339), .B2(keyinput52), .C1(n11010), .C2(
        keyinput122), .A(n15338), .ZN(n15349) );
  AOI22_X1 U16898 ( .A1(n15341), .A2(keyinput58), .B1(keyinput111), .B2(n8265), 
        .ZN(n15340) );
  OAI221_X1 U16899 ( .B1(n15341), .B2(keyinput58), .C1(n8265), .C2(keyinput111), .A(n15340), .ZN(n15348) );
  INV_X1 U16900 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n15343) );
  AOI22_X1 U16901 ( .A1(n15343), .A2(keyinput54), .B1(keyinput89), .B2(n9120), 
        .ZN(n15342) );
  OAI221_X1 U16902 ( .B1(n15343), .B2(keyinput54), .C1(n9120), .C2(keyinput89), 
        .A(n15342), .ZN(n15347) );
  XOR2_X1 U16903 ( .A(n12853), .B(keyinput59), .Z(n15345) );
  XNOR2_X1 U16904 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput15), .ZN(n15344) );
  NAND2_X1 U16905 ( .A1(n15345), .A2(n15344), .ZN(n15346) );
  NOR4_X1 U16906 ( .A1(n15349), .A2(n15348), .A3(n15347), .A4(n15346), .ZN(
        n15382) );
  AOI22_X1 U16907 ( .A1(n15352), .A2(keyinput108), .B1(keyinput80), .B2(n15351), .ZN(n15350) );
  OAI221_X1 U16908 ( .B1(n15352), .B2(keyinput108), .C1(n15351), .C2(
        keyinput80), .A(n15350), .ZN(n15364) );
  AOI22_X1 U16909 ( .A1(n15354), .A2(keyinput55), .B1(n8407), .B2(keyinput20), 
        .ZN(n15353) );
  OAI221_X1 U16910 ( .B1(n15354), .B2(keyinput55), .C1(n8407), .C2(keyinput20), 
        .A(n15353), .ZN(n15363) );
  INV_X1 U16911 ( .A(keyinput63), .ZN(n15356) );
  AOI22_X1 U16912 ( .A1(n15357), .A2(keyinput106), .B1(P1_WR_REG_SCAN_IN), 
        .B2(n15356), .ZN(n15355) );
  OAI221_X1 U16913 ( .B1(n15357), .B2(keyinput106), .C1(n15356), .C2(
        P1_WR_REG_SCAN_IN), .A(n15355), .ZN(n15362) );
  AOI22_X1 U16914 ( .A1(n15360), .A2(keyinput105), .B1(keyinput91), .B2(n15359), .ZN(n15358) );
  OAI221_X1 U16915 ( .B1(n15360), .B2(keyinput105), .C1(n15359), .C2(
        keyinput91), .A(n15358), .ZN(n15361) );
  NOR4_X1 U16916 ( .A1(n15364), .A2(n15363), .A3(n15362), .A4(n15361), .ZN(
        n15381) );
  AOI22_X1 U16917 ( .A1(n15367), .A2(keyinput8), .B1(keyinput117), .B2(n15366), 
        .ZN(n15365) );
  OAI221_X1 U16918 ( .B1(n15367), .B2(keyinput8), .C1(n15366), .C2(keyinput117), .A(n15365), .ZN(n15379) );
  AOI22_X1 U16919 ( .A1(n15370), .A2(keyinput18), .B1(keyinput3), .B2(n15369), 
        .ZN(n15368) );
  OAI221_X1 U16920 ( .B1(n15370), .B2(keyinput18), .C1(n15369), .C2(keyinput3), 
        .A(n15368), .ZN(n15378) );
  INV_X1 U16921 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U16922 ( .A1(n15373), .A2(keyinput74), .B1(n15372), .B2(keyinput124), .ZN(n15371) );
  OAI221_X1 U16923 ( .B1(n15373), .B2(keyinput74), .C1(n15372), .C2(
        keyinput124), .A(n15371), .ZN(n15377) );
  XNOR2_X1 U16924 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput28), .ZN(n15375)
         );
  XNOR2_X1 U16925 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput60), .ZN(n15374) );
  NAND2_X1 U16926 ( .A1(n15375), .A2(n15374), .ZN(n15376) );
  NOR4_X1 U16927 ( .A1(n15379), .A2(n15378), .A3(n15377), .A4(n15376), .ZN(
        n15380) );
  NAND4_X1 U16928 ( .A1(n15383), .A2(n15382), .A3(n15381), .A4(n15380), .ZN(
        n15506) );
  AOI22_X1 U16929 ( .A1(n15385), .A2(keyinput82), .B1(keyinput65), .B2(n13433), 
        .ZN(n15384) );
  OAI221_X1 U16930 ( .B1(n15385), .B2(keyinput82), .C1(n13433), .C2(keyinput65), .A(n15384), .ZN(n15395) );
  XNOR2_X1 U16931 ( .A(keyinput79), .B(n15386), .ZN(n15394) );
  XNOR2_X1 U16932 ( .A(keyinput47), .B(n15387), .ZN(n15393) );
  XNOR2_X1 U16933 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput10), .ZN(n15391) );
  XNOR2_X1 U16934 ( .A(P3_IR_REG_26__SCAN_IN), .B(keyinput57), .ZN(n15390) );
  XNOR2_X1 U16935 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput38), .ZN(n15389) );
  XNOR2_X1 U16936 ( .A(keyinput92), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n15388) );
  NAND4_X1 U16937 ( .A1(n15391), .A2(n15390), .A3(n15389), .A4(n15388), .ZN(
        n15392) );
  NOR4_X1 U16938 ( .A1(n15395), .A2(n15394), .A3(n15393), .A4(n15392), .ZN(
        n15441) );
  AOI22_X1 U16939 ( .A1(n15397), .A2(keyinput72), .B1(n12060), .B2(keyinput113), .ZN(n15396) );
  OAI221_X1 U16940 ( .B1(n15397), .B2(keyinput72), .C1(n12060), .C2(
        keyinput113), .A(n15396), .ZN(n15409) );
  AOI22_X1 U16941 ( .A1(n15400), .A2(keyinput40), .B1(keyinput1), .B2(n15399), 
        .ZN(n15398) );
  OAI221_X1 U16942 ( .B1(n15400), .B2(keyinput40), .C1(n15399), .C2(keyinput1), 
        .A(n15398), .ZN(n15408) );
  AOI22_X1 U16943 ( .A1(n7660), .A2(keyinput102), .B1(keyinput16), .B2(n15402), 
        .ZN(n15401) );
  OAI221_X1 U16944 ( .B1(n7660), .B2(keyinput102), .C1(n15402), .C2(keyinput16), .A(n15401), .ZN(n15407) );
  XOR2_X1 U16945 ( .A(n15403), .B(keyinput31), .Z(n15405) );
  XNOR2_X1 U16946 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput39), .ZN(n15404)
         );
  NAND2_X1 U16947 ( .A1(n15405), .A2(n15404), .ZN(n15406) );
  NOR4_X1 U16948 ( .A1(n15409), .A2(n15408), .A3(n15407), .A4(n15406), .ZN(
        n15440) );
  AOI22_X1 U16949 ( .A1(n15411), .A2(keyinput83), .B1(keyinput75), .B2(n10669), 
        .ZN(n15410) );
  OAI221_X1 U16950 ( .B1(n15411), .B2(keyinput83), .C1(n10669), .C2(keyinput75), .A(n15410), .ZN(n15422) );
  AOI22_X1 U16951 ( .A1(n12870), .A2(keyinput44), .B1(keyinput78), .B2(n15413), 
        .ZN(n15412) );
  OAI221_X1 U16952 ( .B1(n12870), .B2(keyinput44), .C1(n15413), .C2(keyinput78), .A(n15412), .ZN(n15421) );
  INV_X1 U16953 ( .A(keyinput126), .ZN(n15415) );
  AOI22_X1 U16954 ( .A1(n7112), .A2(keyinput101), .B1(P3_DATAO_REG_19__SCAN_IN), .B2(n15415), .ZN(n15414) );
  OAI221_X1 U16955 ( .B1(n7112), .B2(keyinput101), .C1(n15415), .C2(
        P3_DATAO_REG_19__SCAN_IN), .A(n15414), .ZN(n15420) );
  XOR2_X1 U16956 ( .A(n15416), .B(keyinput109), .Z(n15418) );
  XNOR2_X1 U16957 ( .A(SI_7_), .B(keyinput14), .ZN(n15417) );
  NAND2_X1 U16958 ( .A1(n15418), .A2(n15417), .ZN(n15419) );
  NOR4_X1 U16959 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15439) );
  AOI22_X1 U16960 ( .A1(n15425), .A2(keyinput23), .B1(keyinput88), .B2(n15424), 
        .ZN(n15423) );
  OAI221_X1 U16961 ( .B1(n15425), .B2(keyinput23), .C1(n15424), .C2(keyinput88), .A(n15423), .ZN(n15437) );
  AOI22_X1 U16962 ( .A1(n15428), .A2(keyinput41), .B1(n15427), .B2(keyinput97), 
        .ZN(n15426) );
  OAI221_X1 U16963 ( .B1(n15428), .B2(keyinput41), .C1(n15427), .C2(keyinput97), .A(n15426), .ZN(n15436) );
  AOI22_X1 U16964 ( .A1(n15431), .A2(keyinput100), .B1(keyinput119), .B2(
        n15430), .ZN(n15429) );
  OAI221_X1 U16965 ( .B1(n15431), .B2(keyinput100), .C1(n15430), .C2(
        keyinput119), .A(n15429), .ZN(n15435) );
  XNOR2_X1 U16966 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput123), .ZN(n15433)
         );
  XNOR2_X1 U16967 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput56), .ZN(n15432)
         );
  NAND2_X1 U16968 ( .A1(n15433), .A2(n15432), .ZN(n15434) );
  NOR4_X1 U16969 ( .A1(n15437), .A2(n15436), .A3(n15435), .A4(n15434), .ZN(
        n15438) );
  NAND4_X1 U16970 ( .A1(n15441), .A2(n15440), .A3(n15439), .A4(n15438), .ZN(
        n15505) );
  AOI22_X1 U16971 ( .A1(n15444), .A2(keyinput45), .B1(n15443), .B2(keyinput71), 
        .ZN(n15442) );
  OAI221_X1 U16972 ( .B1(n15444), .B2(keyinput45), .C1(n15443), .C2(keyinput71), .A(n15442), .ZN(n15456) );
  INV_X1 U16973 ( .A(keyinput12), .ZN(n15446) );
  AOI22_X1 U16974 ( .A1(n15447), .A2(keyinput85), .B1(P3_DATAO_REG_28__SCAN_IN), .B2(n15446), .ZN(n15445) );
  OAI221_X1 U16975 ( .B1(n15447), .B2(keyinput85), .C1(n15446), .C2(
        P3_DATAO_REG_28__SCAN_IN), .A(n15445), .ZN(n15455) );
  AOI22_X1 U16976 ( .A1(n15450), .A2(keyinput86), .B1(keyinput22), .B2(n15449), 
        .ZN(n15448) );
  OAI221_X1 U16977 ( .B1(n15450), .B2(keyinput86), .C1(n15449), .C2(keyinput22), .A(n15448), .ZN(n15454) );
  XOR2_X1 U16978 ( .A(n7050), .B(keyinput11), .Z(n15452) );
  XNOR2_X1 U16979 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput33), .ZN(n15451) );
  NAND2_X1 U16980 ( .A1(n15452), .A2(n15451), .ZN(n15453) );
  NOR4_X1 U16981 ( .A1(n15456), .A2(n15455), .A3(n15454), .A4(n15453), .ZN(
        n15503) );
  AOI22_X1 U16982 ( .A1(n15459), .A2(keyinput53), .B1(keyinput110), .B2(n15458), .ZN(n15457) );
  OAI221_X1 U16983 ( .B1(n15459), .B2(keyinput53), .C1(n15458), .C2(
        keyinput110), .A(n15457), .ZN(n15471) );
  INV_X1 U16984 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n15462) );
  INV_X1 U16985 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U16986 ( .A1(n15462), .A2(keyinput25), .B1(n15461), .B2(keyinput42), 
        .ZN(n15460) );
  OAI221_X1 U16987 ( .B1(n15462), .B2(keyinput25), .C1(n15461), .C2(keyinput42), .A(n15460), .ZN(n15470) );
  AOI22_X1 U16988 ( .A1(n15465), .A2(keyinput127), .B1(keyinput51), .B2(n15464), .ZN(n15463) );
  OAI221_X1 U16989 ( .B1(n15465), .B2(keyinput127), .C1(n15464), .C2(
        keyinput51), .A(n15463), .ZN(n15469) );
  INV_X1 U16990 ( .A(keyinput13), .ZN(n15467) );
  XNOR2_X1 U16991 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput49), .ZN(n15466) );
  OAI21_X1 U16992 ( .B1(P1_REG0_REG_8__SCAN_IN), .B2(n15467), .A(n15466), .ZN(
        n15468) );
  NOR4_X1 U16993 ( .A1(n15471), .A2(n15470), .A3(n15469), .A4(n15468), .ZN(
        n15502) );
  AOI22_X1 U16994 ( .A1(n9046), .A2(keyinput103), .B1(keyinput107), .B2(n15473), .ZN(n15472) );
  OAI221_X1 U16995 ( .B1(n9046), .B2(keyinput103), .C1(n15473), .C2(
        keyinput107), .A(n15472), .ZN(n15485) );
  AOI22_X1 U16996 ( .A1(n15476), .A2(keyinput69), .B1(n15475), .B2(keyinput37), 
        .ZN(n15474) );
  OAI221_X1 U16997 ( .B1(n15476), .B2(keyinput69), .C1(n15475), .C2(keyinput37), .A(n15474), .ZN(n15484) );
  INV_X1 U16998 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U16999 ( .A1(n15478), .A2(keyinput9), .B1(n8008), .B2(keyinput19), 
        .ZN(n15477) );
  OAI221_X1 U17000 ( .B1(n15478), .B2(keyinput9), .C1(n8008), .C2(keyinput19), 
        .A(n15477), .ZN(n15483) );
  XOR2_X1 U17001 ( .A(n15479), .B(keyinput118), .Z(n15481) );
  XNOR2_X1 U17002 ( .A(P3_IR_REG_13__SCAN_IN), .B(keyinput2), .ZN(n15480) );
  NAND2_X1 U17003 ( .A1(n15481), .A2(n15480), .ZN(n15482) );
  NOR4_X1 U17004 ( .A1(n15485), .A2(n15484), .A3(n15483), .A4(n15482), .ZN(
        n15501) );
  AOI22_X1 U17005 ( .A1(n15488), .A2(keyinput95), .B1(keyinput68), .B2(n15487), 
        .ZN(n15486) );
  OAI221_X1 U17006 ( .B1(n15488), .B2(keyinput95), .C1(n15487), .C2(keyinput68), .A(n15486), .ZN(n15499) );
  INV_X1 U17007 ( .A(keyinput121), .ZN(n15490) );
  AOI22_X1 U17008 ( .A1(n9510), .A2(keyinput7), .B1(P3_DATAO_REG_22__SCAN_IN), 
        .B2(n15490), .ZN(n15489) );
  OAI221_X1 U17009 ( .B1(n9510), .B2(keyinput7), .C1(n15490), .C2(
        P3_DATAO_REG_22__SCAN_IN), .A(n15489), .ZN(n15498) );
  AOI22_X1 U17010 ( .A1(n15493), .A2(keyinput104), .B1(n15492), .B2(keyinput66), .ZN(n15491) );
  OAI221_X1 U17011 ( .B1(n15493), .B2(keyinput104), .C1(n15492), .C2(
        keyinput66), .A(n15491), .ZN(n15497) );
  XNOR2_X1 U17012 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput81), .ZN(n15495) );
  XNOR2_X1 U17013 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput112), .ZN(n15494)
         );
  NAND2_X1 U17014 ( .A1(n15495), .A2(n15494), .ZN(n15496) );
  NOR4_X1 U17015 ( .A1(n15499), .A2(n15498), .A3(n15497), .A4(n15496), .ZN(
        n15500) );
  NAND4_X1 U17016 ( .A1(n15503), .A2(n15502), .A3(n15501), .A4(n15500), .ZN(
        n15504) );
  NOR4_X1 U17017 ( .A1(n15507), .A2(n15506), .A3(n15505), .A4(n15504), .ZN(
        n15508) );
  OAI221_X1 U17018 ( .B1(n15510), .B2(keyinput13), .C1(n15510), .C2(n15509), 
        .A(n15508), .ZN(n15511) );
  XNOR2_X1 U17019 ( .A(n15512), .B(n15511), .ZN(P2_U3258) );
  XOR2_X1 U17020 ( .A(n15514), .B(n15513), .Z(SUB_1596_U59) );
  XNOR2_X1 U17021 ( .A(n15515), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17022 ( .B1(n15517), .B2(n15516), .A(n15525), .ZN(SUB_1596_U53) );
  XOR2_X1 U17023 ( .A(n15518), .B(n15519), .Z(SUB_1596_U56) );
  OAI21_X1 U17024 ( .B1(n15522), .B2(n15521), .A(n15520), .ZN(n15523) );
  XNOR2_X1 U17025 ( .A(n15523), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U17026 ( .A(n15525), .B(n15524), .Z(SUB_1596_U5) );
  AND2_X1 U7587 ( .A1(n12277), .A2(n13730), .ZN(n8928) );
  CLKBUF_X1 U7324 ( .A(n9117), .Z(n12059) );
  CLKBUF_X1 U7336 ( .A(n10375), .Z(n12455) );
  CLKBUF_X1 U7354 ( .A(n7928), .Z(n7988) );
  CLKBUF_X1 U7414 ( .A(n9945), .Z(n7046) );
  XNOR2_X1 U7575 ( .A(n9057), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9064) );
  INV_X2 U8000 ( .A(n13574), .ZN(n14997) );
  OR2_X2 U9023 ( .A1(n8309), .A2(n8308), .ZN(n10343) );
  CLKBUF_X1 U9241 ( .A(n8044), .Z(n8070) );
  AND2_X1 U10013 ( .A1(n7145), .A2(n7144), .ZN(n9642) );
endmodule

