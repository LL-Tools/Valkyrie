

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673;

  AND2_X1 U4972 ( .A1(n6082), .A2(n6081), .ZN(n9245) );
  INV_X2 U4973 ( .A(n4909), .ZN(n9170) );
  INV_X1 U4974 ( .A(n6378), .ZN(n8306) );
  CLKBUF_X2 U4975 ( .A(n6046), .Z(n4909) );
  INV_X1 U4976 ( .A(n8473), .ZN(n8477) );
  OR2_X1 U4977 ( .A1(n6527), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6343) );
  INV_X1 U4978 ( .A(n10022), .ZN(n5638) );
  INV_X1 U4979 ( .A(n8300), .ZN(n6677) );
  INV_X1 U4980 ( .A(n8688), .ZN(n8272) );
  INV_X1 U4982 ( .A(n9170), .ZN(n6214) );
  NAND2_X1 U4983 ( .A1(n6236), .A2(n9544), .ZN(n5654) );
  NOR2_X1 U4984 ( .A1(n9874), .A2(n9960), .ZN(n9858) );
  NOR2_X1 U4985 ( .A1(n8029), .A2(n9980), .ZN(n8102) );
  NAND2_X1 U4986 ( .A1(n7831), .A2(n9778), .ZN(n9383) );
  AND3_X1 U4987 ( .A1(n5466), .A2(n5590), .A3(n5477), .ZN(n5634) );
  OAI211_X1 U4988 ( .C1(n5703), .C2(n6792), .A(n5147), .B(n5146), .ZN(n7234)
         );
  NAND2_X1 U4989 ( .A1(n6071), .A2(n6070), .ZN(n9943) );
  INV_X1 U4990 ( .A(n6312), .ZN(n9146) );
  XNOR2_X2 U4992 ( .A(n5515), .B(SI_5_), .ZN(n5757) );
  NAND4_X2 U4993 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n8522)
         );
  OAI22_X2 U4994 ( .A1(n8731), .A2(n8737), .B1(n8744), .B2(n8835), .ZN(n8720)
         );
  XNOR2_X1 U4995 ( .A(n5596), .B(n5595), .ZN(n6245) );
  AOI21_X2 U4996 ( .B1(n7840), .B2(n7724), .A(n7723), .ZN(n7866) );
  NAND2_X2 U4997 ( .A1(n5378), .A2(n5375), .ZN(n6863) );
  OAI21_X2 U4998 ( .B1(n5971), .B2(n5555), .A(n5554), .ZN(n5990) );
  AND2_X4 U4999 ( .A1(n10021), .A2(n5638), .ZN(n4916) );
  INV_X1 U5000 ( .A(n5639), .ZN(n10021) );
  XNOR2_X2 U5001 ( .A(n8672), .B(n8326), .ZN(n8653) );
  NAND2_X4 U5002 ( .A1(n6313), .A2(n9146), .ZN(n6374) );
  NAND2_X2 U5003 ( .A1(n6366), .A2(n6365), .ZN(n6878) );
  OR2_X1 U5004 ( .A1(n6082), .A2(n6081), .ZN(n9244) );
  NAND2_X1 U5005 ( .A1(n8167), .A2(n4919), .ZN(n8169) );
  INV_X1 U5006 ( .A(n8522), .ZN(n8699) );
  INV_X1 U5007 ( .A(n9573), .ZN(n7535) );
  INV_X1 U5008 ( .A(n7073), .ZN(n7273) );
  INV_X1 U5009 ( .A(n5284), .ZN(n10446) );
  NAND4_X1 U5010 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n9573)
         );
  INV_X1 U5011 ( .A(n9383), .ZN(n9394) );
  NAND2_X1 U5012 ( .A1(n5290), .A2(n5291), .ZN(n5643) );
  NOR2_X1 U5013 ( .A1(n5295), .A2(n4930), .ZN(n9908) );
  NAND2_X1 U5014 ( .A1(n9208), .A2(n9209), .ZN(n6270) );
  AOI21_X1 U5015 ( .B1(n6765), .B2(n8793), .A(n6764), .ZN(n8682) );
  AND2_X1 U5016 ( .A1(n8653), .A2(n5255), .ZN(n5254) );
  AOI21_X1 U5017 ( .B1(n5318), .B2(n5320), .A(n5317), .ZN(n9796) );
  NAND2_X1 U5018 ( .A1(n6658), .A2(n6657), .ZN(n8672) );
  NAND2_X1 U5019 ( .A1(n9456), .A2(n9523), .ZN(n9695) );
  AND2_X1 U5020 ( .A1(n9835), .A2(n4915), .ZN(n9766) );
  OAI22_X1 U5021 ( .A1(n8122), .A2(n5197), .B1(n4955), .B2(n5196), .ZN(n6027)
         );
  NAND2_X1 U5022 ( .A1(n8111), .A2(n9353), .ZN(n9881) );
  NAND2_X1 U5023 ( .A1(n8068), .A2(n8067), .ZN(n8066) );
  AND2_X1 U5024 ( .A1(n5249), .A2(n4956), .ZN(n8068) );
  NAND2_X1 U5025 ( .A1(n5602), .A2(n5601), .ZN(n9950) );
  XNOR2_X1 U5026 ( .A(n6069), .B(n6084), .ZN(n7819) );
  NAND2_X1 U5027 ( .A1(n6305), .A2(n6304), .ZN(n8851) );
  NAND2_X1 U5028 ( .A1(n5220), .A2(n5219), .ZN(n5842) );
  NAND2_X1 U5029 ( .A1(n5052), .A2(n5256), .ZN(n7834) );
  AND2_X1 U5030 ( .A1(n5578), .A2(n5577), .ZN(n6089) );
  NAND2_X1 U5031 ( .A1(n5288), .A2(n5287), .ZN(n7807) );
  NAND2_X1 U5032 ( .A1(n8006), .A2(n8005), .ZN(n8029) );
  NAND2_X1 U5033 ( .A1(n6775), .A2(n5173), .ZN(n6777) );
  NAND2_X1 U5034 ( .A1(n7404), .A2(n10448), .ZN(n9868) );
  BUF_X1 U5035 ( .A(n6917), .Z(n6943) );
  NAND2_X2 U5036 ( .A1(n5674), .A2(n5673), .ZN(n9574) );
  NAND2_X1 U5037 ( .A1(n8335), .A2(n8343), .ZN(n7128) );
  AND3_X1 U5038 ( .A1(n5672), .A2(n5671), .A3(n5670), .ZN(n5674) );
  OR2_X1 U5039 ( .A1(n6958), .A2(n6961), .ZN(n6959) );
  INV_X1 U5040 ( .A(n5683), .ZN(n6185) );
  NAND4_X1 U5041 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n8539)
         );
  AND2_X2 U5042 ( .A1(n5638), .A2(n5639), .ZN(n9184) );
  AND3_X1 U5043 ( .A1(n6370), .A2(n6369), .A3(n6368), .ZN(n7310) );
  OR2_X1 U5044 ( .A1(n8297), .A2(n6788), .ZN(n6398) );
  AND3_X1 U5045 ( .A1(n6361), .A2(n6360), .A3(n5037), .ZN(n6371) );
  NAND2_X1 U5046 ( .A1(n6224), .A2(n5610), .ZN(n5680) );
  INV_X2 U5047 ( .A(n6383), .ZN(n8296) );
  INV_X1 U5048 ( .A(n6684), .ZN(n8339) );
  AND2_X2 U5049 ( .A1(n5639), .A2(n10022), .ZN(n5786) );
  XNOR2_X1 U5050 ( .A(n6672), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U5051 ( .A1(n6357), .A2(n8286), .ZN(n6383) );
  NAND2_X1 U5052 ( .A1(n5635), .A2(n5636), .ZN(n10022) );
  XNOR2_X1 U5053 ( .A(n5637), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U5054 ( .A(n6237), .B(n5653), .ZN(n9550) );
  NAND2_X1 U5055 ( .A1(n6845), .A2(n8619), .ZN(n6357) );
  NAND2_X1 U5056 ( .A1(n5636), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5637) );
  XNOR2_X1 U5057 ( .A(n5652), .B(n5614), .ZN(n9544) );
  XNOR2_X1 U5058 ( .A(n6311), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U5059 ( .A1(n6300), .A2(n6299), .ZN(n6302) );
  OR2_X1 U5060 ( .A1(n6500), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6513) );
  OR2_X1 U5061 ( .A1(n6489), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6500) );
  INV_X2 U5062 ( .A(n9141), .ZN(n9153) );
  XNOR2_X1 U5063 ( .A(n5000), .B(n6307), .ZN(n8204) );
  NAND2_X1 U5064 ( .A1(n6310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6311) );
  CLKBUF_X3 U5065 ( .A(n5506), .Z(n6656) );
  NAND2_X1 U5066 ( .A1(n9138), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5000) );
  CLKBUF_X3 U5067 ( .A(n5506), .Z(n8141) );
  NOR2_X1 U5068 ( .A1(n5377), .A2(n5376), .ZN(n5375) );
  AND3_X1 U5069 ( .A1(n5413), .A2(n6293), .A3(n6298), .ZN(n6309) );
  CLKBUF_X1 U5070 ( .A(n5600), .Z(n8286) );
  NOR2_X1 U5071 ( .A1(n6442), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6461) );
  AND3_X2 U5072 ( .A1(n6291), .A2(n6290), .A3(n5377), .ZN(n6293) );
  AND2_X1 U5073 ( .A1(n5463), .A2(n5145), .ZN(n5290) );
  NAND2_X1 U5074 ( .A1(n5494), .A2(n5495), .ZN(n5600) );
  OR2_X1 U5075 ( .A1(n5592), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4910) );
  OR2_X1 U5076 ( .A1(n6428), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6442) );
  AND2_X1 U5077 ( .A1(n5464), .A2(n5588), .ZN(n5463) );
  CLKBUF_X1 U5078 ( .A(n6364), .Z(n6860) );
  AND2_X1 U5079 ( .A1(n5586), .A2(n5587), .ZN(n5464) );
  OAI21_X1 U5080 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5491), .ZN(n5495) );
  AND4_X1 U5081 ( .A1(n6325), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n6291)
         );
  AND4_X1 U5082 ( .A1(n6288), .A2(n6287), .A3(n6286), .A4(n6333), .ZN(n6290)
         );
  INV_X1 U5083 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6689) );
  INV_X1 U5084 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6696) );
  INV_X1 U5085 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6719) );
  INV_X1 U5086 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6307) );
  NOR2_X1 U5087 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6285) );
  NOR2_X1 U5088 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6284) );
  NOR2_X1 U5089 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6283) );
  NOR2_X1 U5090 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6287) );
  NOR2_X1 U5091 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6286) );
  NOR2_X1 U5092 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6364) );
  INV_X1 U5093 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5492) );
  INV_X1 U5094 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6333) );
  NOR2_X1 U5095 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6325) );
  NOR2_X1 U5096 ( .A1(n6027), .A2(n6026), .ZN(n9256) );
  AOI21_X2 U5097 ( .B1(n8060), .B2(n5988), .A(n5472), .ZN(n8122) );
  AOI21_X2 U5098 ( .B1(n7719), .B2(n5136), .A(n7718), .ZN(n7840) );
  OR2_X1 U5099 ( .A1(n10649), .A2(n8222), .ZN(n8428) );
  OR2_X1 U5100 ( .A1(n9907), .A2(n9276), .ZN(n9458) );
  NAND2_X1 U5101 ( .A1(n4961), .A2(n5451), .ZN(n5445) );
  OAI21_X1 U5102 ( .B1(n6166), .B2(n6165), .A(n6168), .ZN(n6198) );
  INV_X1 U5103 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5589) );
  AND2_X1 U5104 ( .A1(n6684), .A2(n8518), .ZN(n8473) );
  NAND2_X1 U5105 ( .A1(n8268), .A2(n8191), .ZN(n8207) );
  AND2_X1 U5106 ( .A1(n8204), .A2(n6312), .ZN(n8300) );
  INV_X1 U5107 ( .A(n8771), .ZN(n8801) );
  NAND2_X1 U5108 ( .A1(n7059), .A2(n8473), .ZN(n8786) );
  AND2_X1 U5109 ( .A1(n8369), .A2(n8368), .ZN(n8378) );
  NAND2_X1 U5110 ( .A1(n6991), .A2(n6372), .ZN(n8335) );
  INV_X1 U5111 ( .A(n8168), .ZN(n5422) );
  AOI21_X1 U5112 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8590), .A(n10333), .ZN(
        n8591) );
  AOI21_X1 U5113 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8594), .A(n10365), .ZN(
        n8595) );
  NAND2_X1 U5114 ( .A1(n8866), .A2(n8527), .ZN(n5250) );
  NAND2_X1 U5115 ( .A1(n5229), .A2(n6740), .ZN(n5226) );
  OR2_X1 U5116 ( .A1(n8680), .A2(n8272), .ZN(n8474) );
  OR2_X1 U5117 ( .A1(n8858), .A2(n10643), .ZN(n8425) );
  OR2_X1 U5118 ( .A1(n8862), .A2(n8802), .ZN(n8331) );
  AND2_X1 U5119 ( .A1(n8401), .A2(n8400), .ZN(n8398) );
  AND2_X1 U5120 ( .A1(n5223), .A2(n5222), .ZN(n5415) );
  NOR2_X1 U5121 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5223) );
  NOR2_X1 U5122 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5222) );
  OR2_X1 U5123 ( .A1(n9916), .A2(n9750), .ZN(n9459) );
  NAND2_X1 U5124 ( .A1(n7803), .A2(n7776), .ZN(n9317) );
  OAI21_X1 U5125 ( .B1(n7431), .B2(n7665), .A(n7430), .ZN(n7669) );
  NOR2_X1 U5126 ( .A1(n4910), .A2(n5159), .ZN(n5155) );
  NAND2_X1 U5127 ( .A1(n6150), .A2(n6149), .ZN(n6166) );
  NOR2_X1 U5128 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5649) );
  NAND2_X1 U5129 ( .A1(n6122), .A2(n6121), .ZN(n6148) );
  INV_X1 U5130 ( .A(n5334), .ZN(n5333) );
  OAI21_X1 U5131 ( .B1(n5337), .B2(n4969), .A(n5573), .ZN(n5334) );
  INV_X1 U5132 ( .A(SI_18_), .ZN(n5566) );
  INV_X1 U5133 ( .A(n5743), .ZN(n5145) );
  OAI21_X1 U5134 ( .B1(n5901), .B2(n5544), .A(n5543), .ZN(n5930) );
  OR2_X1 U5135 ( .A1(n8082), .A2(n8802), .ZN(n5473) );
  NAND2_X1 U5136 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U5137 ( .A1(n5413), .A2(n6293), .ZN(n6296) );
  AND4_X1 U5138 ( .A1(n6575), .A2(n6574), .A3(n6573), .A4(n6572), .ZN(n8222)
         );
  XNOR2_X1 U5139 ( .A(n8591), .B(n10341), .ZN(n10350) );
  XNOR2_X1 U5140 ( .A(n8595), .B(n10372), .ZN(n10381) );
  OAI21_X1 U5141 ( .B1(n8720), .B2(n6613), .A(n5276), .ZN(n8710) );
  INV_X1 U5142 ( .A(n5278), .ZN(n5276) );
  AND2_X1 U5143 ( .A1(n8442), .A2(n8439), .ZN(n8737) );
  NAND2_X1 U5144 ( .A1(n5059), .A2(n5058), .ZN(n8743) );
  AOI21_X1 U5145 ( .B1(n5060), .B2(n8768), .A(n4950), .ZN(n5058) );
  OR2_X1 U5146 ( .A1(n8074), .A2(n8802), .ZN(n5474) );
  NAND2_X1 U5147 ( .A1(n7637), .A2(n8393), .ZN(n6733) );
  INV_X1 U5148 ( .A(n8297), .ZN(n6565) );
  BUF_X1 U5149 ( .A(n6384), .Z(n8297) );
  NAND2_X1 U5150 ( .A1(n6357), .A2(n6656), .ZN(n6384) );
  NAND2_X1 U5151 ( .A1(n5230), .A2(n8459), .ZN(n5229) );
  INV_X1 U5152 ( .A(n8686), .ZN(n5230) );
  NAND2_X1 U5153 ( .A1(n5228), .A2(n8459), .ZN(n8683) );
  NAND2_X1 U5154 ( .A1(n6301), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U5155 ( .A1(n8154), .A2(n8153), .ZN(n9907) );
  AND2_X1 U5156 ( .A1(n9458), .A2(n9531), .ZN(n9704) );
  OAI21_X1 U5157 ( .B1(n5461), .B2(n5462), .A(n5458), .ZN(n5455) );
  AOI21_X1 U5158 ( .B1(n5460), .B2(n9380), .A(n4946), .ZN(n5458) );
  INV_X1 U5159 ( .A(n9681), .ZN(n9798) );
  NAND2_X1 U5160 ( .A1(n5097), .A2(n5093), .ZN(n9790) );
  AND2_X1 U5161 ( .A1(n9791), .A2(n5096), .ZN(n5093) );
  AND2_X1 U5162 ( .A1(n9370), .A2(n9371), .ZN(n9814) );
  OR2_X1 U5163 ( .A1(n9950), .A2(n9851), .ZN(n5440) );
  OAI21_X1 U5164 ( .B1(n5073), .B2(n5071), .A(n5069), .ZN(n9827) );
  AOI21_X1 U5165 ( .B1(n5070), .B2(n5074), .A(n4952), .ZN(n5069) );
  NAND2_X1 U5166 ( .A1(n5074), .A2(n5072), .ZN(n5071) );
  AOI21_X1 U5167 ( .B1(n8098), .B2(n5443), .A(n4945), .ZN(n5442) );
  INV_X1 U5168 ( .A(n5445), .ZN(n5443) );
  INV_X2 U5169 ( .A(n5703), .ZN(n9273) );
  INV_X1 U5170 ( .A(n5778), .ZN(n6032) );
  INV_X1 U5171 ( .A(n6820), .ZN(n6031) );
  OR2_X1 U5172 ( .A1(n10444), .A2(n7244), .ZN(n10512) );
  NOR2_X1 U5173 ( .A1(n4910), .A2(n5630), .ZN(n5466) );
  INV_X1 U5174 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5306) );
  XNOR2_X1 U5175 ( .A(n6198), .B(n6197), .ZN(n8015) );
  INV_X1 U5176 ( .A(n8715), .ZN(n8828) );
  XNOR2_X1 U5177 ( .A(n6668), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8633) );
  AOI21_X1 U5178 ( .B1(n6683), .B2(n8793), .A(n6682), .ZN(n8674) );
  INV_X1 U5179 ( .A(n9181), .ZN(n9182) );
  OAI21_X1 U5180 ( .B1(n9757), .B2(n9243), .A(n6278), .ZN(n6279) );
  NAND2_X1 U5181 ( .A1(n8385), .A2(n8473), .ZN(n5126) );
  NAND2_X1 U5182 ( .A1(n5128), .A2(n8477), .ZN(n5127) );
  OAI21_X1 U5183 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(n5128) );
  INV_X1 U5184 ( .A(n5141), .ZN(n5140) );
  OAI211_X1 U5185 ( .C1(n8423), .C2(n8424), .A(n8792), .B(n4942), .ZN(n5141)
         );
  OAI21_X1 U5186 ( .B1(n5144), .B2(n5143), .A(n8737), .ZN(n5330) );
  NAND2_X1 U5187 ( .A1(n8750), .A2(n4934), .ZN(n5143) );
  AOI21_X1 U5188 ( .B1(n8436), .B2(n8435), .A(n8434), .ZN(n5144) );
  NAND2_X1 U5189 ( .A1(n5114), .A2(n9365), .ZN(n9368) );
  NAND2_X1 U5190 ( .A1(n9368), .A2(n5112), .ZN(n5111) );
  NOR2_X1 U5191 ( .A1(n5113), .A2(n9394), .ZN(n5112) );
  INV_X1 U5192 ( .A(n9426), .ZN(n5113) );
  AOI21_X1 U5193 ( .B1(n5254), .B2(n5253), .A(n4947), .ZN(n5252) );
  INV_X1 U5194 ( .A(n5487), .ZN(n5253) );
  INV_X1 U5195 ( .A(n9382), .ZN(n5120) );
  NAND2_X1 U5196 ( .A1(n5122), .A2(n9394), .ZN(n5119) );
  AOI211_X1 U5197 ( .C1(n5123), .C2(n9379), .A(n9378), .B(n5122), .ZN(n5121)
         );
  OAI21_X1 U5198 ( .B1(n9375), .B2(n9374), .A(n5124), .ZN(n5123) );
  NAND2_X1 U5199 ( .A1(n8096), .A2(n8126), .ZN(n5451) );
  INV_X1 U5200 ( .A(n9500), .ZN(n5286) );
  AND2_X1 U5201 ( .A1(n7044), .A2(n8339), .ZN(n7046) );
  AND2_X1 U5202 ( .A1(n7043), .A2(n8507), .ZN(n7044) );
  OAI21_X1 U5203 ( .B1(n8470), .B2(n8469), .A(n5349), .ZN(n5348) );
  NOR2_X1 U5204 ( .A1(n5351), .A2(n5350), .ZN(n5349) );
  OR2_X1 U5205 ( .A1(n8475), .A2(n8476), .ZN(n5347) );
  INV_X1 U5206 ( .A(n5034), .ZN(n5033) );
  OAI21_X1 U5207 ( .B1(n8204), .B2(P2_REG3_REG_1__SCAN_IN), .A(n6312), .ZN(
        n5034) );
  NAND2_X1 U5208 ( .A1(n8204), .A2(n5036), .ZN(n5035) );
  NAND2_X1 U5209 ( .A1(n7146), .A2(n7145), .ZN(n7147) );
  AOI21_X1 U5210 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8586), .A(n10301), .ZN(
        n8587) );
  NOR2_X1 U5211 ( .A1(n10288), .A2(n8609), .ZN(n5384) );
  INV_X1 U5212 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8604) );
  OAI21_X1 U5213 ( .B1(n7626), .B2(n5055), .A(n5053), .ZN(n6534) );
  INV_X1 U5214 ( .A(n5256), .ZN(n5055) );
  AOI21_X1 U5215 ( .B1(n5054), .B2(n5256), .A(n7877), .ZN(n5053) );
  NOR2_X1 U5216 ( .A1(n5259), .A2(n5057), .ZN(n5056) );
  INV_X1 U5217 ( .A(n7622), .ZN(n5057) );
  INV_X1 U5218 ( .A(n5264), .ZN(n5259) );
  AND2_X1 U5219 ( .A1(n5261), .A2(n5257), .ZN(n5256) );
  INV_X1 U5220 ( .A(n5262), .ZN(n5261) );
  NAND2_X1 U5221 ( .A1(n5264), .A2(n5258), .ZN(n5257) );
  OAI21_X1 U5222 ( .B1(n6520), .B2(n5263), .A(n5266), .ZN(n5262) );
  NAND2_X1 U5223 ( .A1(n5241), .A2(n8380), .ZN(n5240) );
  NAND2_X1 U5224 ( .A1(n8376), .A2(n5243), .ZN(n5241) );
  AND2_X1 U5225 ( .A1(n8376), .A2(n5247), .ZN(n5244) );
  NAND2_X1 U5226 ( .A1(n5014), .A2(n8491), .ZN(n5012) );
  NAND2_X1 U5227 ( .A1(n5137), .A2(n5136), .ZN(n8369) );
  INV_X1 U5228 ( .A(n7703), .ZN(n5137) );
  NAND2_X1 U5229 ( .A1(n7703), .A2(n7627), .ZN(n8382) );
  NAND2_X1 U5230 ( .A1(n6427), .A2(n5275), .ZN(n5269) );
  INV_X1 U5231 ( .A(n8486), .ZN(n5247) );
  NAND2_X1 U5232 ( .A1(n6702), .A2(n6701), .ZN(n7045) );
  OR2_X1 U5233 ( .A1(n8835), .A2(n8724), .ZN(n8442) );
  OR2_X1 U5234 ( .A1(n5232), .A2(n5007), .ZN(n5006) );
  INV_X1 U5235 ( .A(n8413), .ZN(n5007) );
  AND2_X1 U5236 ( .A1(n6735), .A2(n8478), .ZN(n5232) );
  NAND2_X1 U5237 ( .A1(n6688), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U5238 ( .A1(n6669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6673) );
  INV_X1 U5239 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U5240 ( .A1(n5213), .A2(n5210), .ZN(n5209) );
  INV_X1 U5241 ( .A(n9202), .ZN(n5210) );
  NAND2_X1 U5242 ( .A1(n6063), .A2(n6062), .ZN(n5217) );
  AND2_X1 U5243 ( .A1(n5679), .A2(n5678), .ZN(n5687) );
  INV_X1 U5244 ( .A(n4976), .ZN(n5196) );
  NAND2_X1 U5245 ( .A1(n5198), .A2(n4976), .ZN(n5197) );
  OAI211_X1 U5246 ( .C1(n7237), .C2(n9550), .A(n5680), .B(n7472), .ZN(n5683)
         );
  NAND2_X1 U5247 ( .A1(n6777), .A2(n5171), .ZN(n5797) );
  NOR2_X1 U5248 ( .A1(n7528), .A2(n5172), .ZN(n5171) );
  AND2_X1 U5249 ( .A1(n6777), .A2(n5794), .ZN(n7522) );
  NOR2_X1 U5250 ( .A1(n9764), .A2(n5315), .ZN(n5314) );
  NAND2_X1 U5251 ( .A1(n5325), .A2(n9370), .ZN(n5324) );
  INV_X1 U5252 ( .A(n5323), .ZN(n5321) );
  NOR2_X1 U5253 ( .A1(n9519), .A2(n5300), .ZN(n5299) );
  INV_X1 U5254 ( .A(n9517), .ZN(n5297) );
  NOR3_X2 U5255 ( .A1(n7777), .A2(n5152), .A3(n5153), .ZN(n8006) );
  OR2_X1 U5256 ( .A1(n7981), .A2(n8002), .ZN(n5152) );
  INV_X1 U5257 ( .A(n7949), .ZN(n5083) );
  NAND2_X1 U5258 ( .A1(n10511), .A2(n9569), .ZN(n9303) );
  NAND2_X1 U5259 ( .A1(n7562), .A2(n7547), .ZN(n9494) );
  NOR2_X1 U5260 ( .A1(n7480), .A2(n9404), .ZN(n5161) );
  NAND2_X1 U5261 ( .A1(n9544), .A2(n6030), .ZN(n7237) );
  OR2_X1 U5262 ( .A1(n6086), .A2(n6085), .ZN(n6090) );
  AND2_X1 U5263 ( .A1(n5577), .A2(n5576), .ZN(n6049) );
  NOR2_X1 U5264 ( .A1(n5569), .A2(n5338), .ZN(n5337) );
  INV_X1 U5265 ( .A(n5564), .ZN(n5338) );
  INV_X1 U5266 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5645) );
  AND2_X1 U5267 ( .A1(n5564), .A2(n5563), .ZN(n6007) );
  INV_X1 U5268 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5992) );
  NOR2_X1 U5269 ( .A1(n5293), .A2(n5292), .ZN(n5291) );
  NAND2_X1 U5270 ( .A1(n5583), .A2(n5584), .ZN(n5293) );
  OR2_X1 U5271 ( .A1(n5847), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5906) );
  NOR2_X1 U5272 ( .A1(n5536), .A2(n5345), .ZN(n5344) );
  INV_X1 U5273 ( .A(n5532), .ZN(n5345) );
  NAND2_X1 U5274 ( .A1(n5102), .A2(n5104), .ZN(n5533) );
  INV_X1 U5275 ( .A(n5105), .ZN(n5104) );
  OAI21_X1 U5276 ( .B1(n5107), .B2(n5106), .A(n5488), .ZN(n5105) );
  OR2_X1 U5277 ( .A1(n5824), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U5278 ( .A1(n5600), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U5279 ( .A1(n7923), .A2(n5412), .ZN(n5411) );
  NAND2_X1 U5280 ( .A1(n7922), .A2(n7871), .ZN(n5412) );
  AOI21_X1 U5281 ( .B1(n8206), .B2(n5399), .A(n8193), .ZN(n5398) );
  INV_X1 U5282 ( .A(n8191), .ZN(n5399) );
  INV_X1 U5283 ( .A(n8195), .ZN(n5396) );
  INV_X1 U5284 ( .A(n5429), .ZN(n5428) );
  OAI21_X1 U5285 ( .B1(n7698), .B2(n5432), .A(n5431), .ZN(n5429) );
  OR2_X1 U5286 ( .A1(n7698), .A2(n7380), .ZN(n5430) );
  OAI21_X1 U5287 ( .B1(n8169), .B2(n5418), .A(n5416), .ZN(n10659) );
  AOI21_X1 U5288 ( .B1(n5417), .B2(n5421), .A(n4912), .ZN(n5416) );
  INV_X1 U5289 ( .A(n8267), .ZN(n8188) );
  INV_X1 U5290 ( .A(n5410), .ZN(n5409) );
  OAI21_X1 U5291 ( .B1(n5411), .B2(n7922), .A(n7987), .ZN(n5410) );
  OR2_X1 U5292 ( .A1(n7986), .A2(n8528), .ZN(n7987) );
  OR2_X1 U5293 ( .A1(n6374), .A2(n6390), .ZN(n6393) );
  INV_X1 U5294 ( .A(n10273), .ZN(n5357) );
  AND2_X1 U5295 ( .A1(n5355), .A2(n10272), .ZN(n5356) );
  OR2_X1 U5296 ( .A1(n6865), .A2(n6949), .ZN(n6866) );
  NAND2_X1 U5297 ( .A1(n6865), .A2(n6949), .ZN(n10273) );
  OR2_X1 U5298 ( .A1(n7147), .A2(n7209), .ZN(n7148) );
  NOR2_X1 U5299 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  OAI21_X1 U5300 ( .B1(n10350), .B2(n5359), .A(n5358), .ZN(n10365) );
  NAND2_X1 U5301 ( .A1(n8593), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5359) );
  OR2_X1 U5302 ( .A1(n10350), .A2(n6529), .ZN(n5361) );
  NAND2_X1 U5303 ( .A1(n8597), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5368) );
  OR2_X1 U5304 ( .A1(n10381), .A2(n7968), .ZN(n5370) );
  NOR2_X1 U5305 ( .A1(n10416), .A2(n10417), .ZN(n10415) );
  NAND2_X1 U5306 ( .A1(n4998), .A2(n8295), .ZN(n8652) );
  NAND2_X1 U5307 ( .A1(n8294), .A2(n8503), .ZN(n4998) );
  OR2_X1 U5308 ( .A1(n6651), .A2(n5051), .ZN(n5050) );
  NAND2_X1 U5309 ( .A1(n8656), .A2(n5254), .ZN(n5051) );
  AOI21_X1 U5310 ( .B1(n6651), .B2(n5048), .A(n5044), .ZN(n5043) );
  NOR2_X1 U5311 ( .A1(n8656), .A2(n5049), .ZN(n5048) );
  NAND2_X1 U5312 ( .A1(n5045), .A2(n8660), .ZN(n5044) );
  OAI21_X1 U5313 ( .B1(n8656), .B2(n5047), .A(n5046), .ZN(n5045) );
  NAND2_X1 U5314 ( .A1(n8657), .A2(n8797), .ZN(n6763) );
  OAI21_X1 U5315 ( .B1(n8720), .B2(n5279), .A(n5277), .ZN(n8687) );
  NAND2_X1 U5316 ( .A1(n5281), .A2(n5280), .ZN(n5279) );
  OAI21_X1 U5317 ( .B1(n5282), .B2(n5278), .A(n5281), .ZN(n5277) );
  INV_X1 U5318 ( .A(n6613), .ZN(n5280) );
  AOI21_X1 U5319 ( .B1(n8743), .B2(n8742), .A(n6595), .ZN(n8731) );
  NOR2_X1 U5320 ( .A1(n8749), .A2(n6594), .ZN(n6595) );
  AOI21_X1 U5321 ( .B1(n5028), .B2(n8328), .A(n8329), .ZN(n5027) );
  INV_X1 U5322 ( .A(n5063), .ZN(n5062) );
  OAI21_X1 U5323 ( .B1(n8768), .B2(n8767), .A(n4957), .ZN(n5063) );
  AND2_X1 U5324 ( .A1(n5062), .A2(n8758), .ZN(n5060) );
  OR2_X1 U5325 ( .A1(n8766), .A2(n8768), .ZN(n5061) );
  OR2_X1 U5326 ( .A1(n6562), .A2(n10643), .ZN(n5482) );
  NAND2_X1 U5327 ( .A1(n6495), .A2(n7623), .ZN(n7635) );
  NAND2_X1 U5328 ( .A1(n7626), .A2(n7622), .ZN(n6495) );
  AND2_X1 U5329 ( .A1(n6461), .A2(n9078), .ZN(n6475) );
  NAND2_X1 U5330 ( .A1(n5248), .A2(n5247), .ZN(n5246) );
  NAND2_X1 U5331 ( .A1(n5246), .A2(n5245), .ZN(n7592) );
  INV_X1 U5332 ( .A(n5243), .ZN(n5245) );
  AND4_X1 U5333 ( .A1(n6447), .A2(n6446), .A3(n6445), .A4(n6444), .ZN(n7554)
         );
  NOR2_X1 U5334 ( .A1(n6426), .A2(n5272), .ZN(n5271) );
  INV_X1 U5335 ( .A(n6411), .ZN(n5272) );
  INV_X1 U5336 ( .A(n8538), .ZN(n7140) );
  INV_X1 U5337 ( .A(n8536), .ZN(n7289) );
  NAND2_X1 U5338 ( .A1(n6744), .A2(n6753), .ZN(n8661) );
  INV_X1 U5339 ( .A(n8786), .ZN(n8797) );
  AND2_X1 U5340 ( .A1(n6990), .A2(n8473), .ZN(n8771) );
  NAND2_X1 U5341 ( .A1(n5017), .A2(n4920), .ZN(n5016) );
  AND2_X1 U5342 ( .A1(n8474), .A2(n8467), .ZN(n8505) );
  AND2_X1 U5343 ( .A1(n6639), .A2(n6638), .ZN(n8686) );
  INV_X1 U5344 ( .A(n8704), .ZN(n5231) );
  NAND2_X1 U5345 ( .A1(n5237), .A2(n8449), .ZN(n5236) );
  AOI21_X1 U5346 ( .B1(n4958), .B2(n5237), .A(n8444), .ZN(n5235) );
  INV_X1 U5347 ( .A(n8737), .ZN(n5239) );
  AOI21_X1 U5348 ( .B1(n8737), .B2(n8440), .A(n5238), .ZN(n5237) );
  INV_X1 U5349 ( .A(n8442), .ZN(n5238) );
  NAND2_X1 U5350 ( .A1(n5031), .A2(n8327), .ZN(n5030) );
  NAND2_X1 U5351 ( .A1(n6738), .A2(n8428), .ZN(n8765) );
  NAND2_X1 U5352 ( .A1(n6338), .A2(n6337), .ZN(n8866) );
  NAND2_X1 U5353 ( .A1(n6734), .A2(n4939), .ZN(n5233) );
  NAND2_X1 U5354 ( .A1(n5233), .A2(n5232), .ZN(n7897) );
  OR3_X1 U5355 ( .A1(n6684), .A2(n8322), .A3(n6749), .ZN(n6983) );
  NOR2_X2 U5356 ( .A1(n5476), .A2(n5414), .ZN(n5413) );
  AND2_X1 U5357 ( .A1(n6293), .A2(n5415), .ZN(n6692) );
  INV_X1 U5358 ( .A(n6324), .ZN(n5377) );
  AND2_X1 U5359 ( .A1(n9139), .A2(n6289), .ZN(n5376) );
  AND2_X1 U5360 ( .A1(n5187), .A2(n4911), .ZN(n5183) );
  NAND2_X1 U5361 ( .A1(n5186), .A2(n5185), .ZN(n5184) );
  AND2_X1 U5362 ( .A1(n5218), .A2(n5217), .ZN(n5212) );
  NAND2_X1 U5363 ( .A1(n9163), .A2(n5211), .ZN(n5207) );
  AND2_X1 U5364 ( .A1(n9202), .A2(n5212), .ZN(n5211) );
  INV_X1 U5365 ( .A(n5209), .ZN(n5205) );
  OR2_X1 U5366 ( .A1(n5215), .A2(n5214), .ZN(n5213) );
  INV_X1 U5367 ( .A(n5217), .ZN(n5214) );
  AOI21_X1 U5368 ( .B1(n9164), .B2(n5218), .A(n5216), .ZN(n5215) );
  INV_X1 U5369 ( .A(n9234), .ZN(n5216) );
  NAND2_X1 U5370 ( .A1(n7522), .A2(n5795), .ZN(n7542) );
  NAND2_X1 U5371 ( .A1(n7533), .A2(n7534), .ZN(n6775) );
  OR2_X1 U5372 ( .A1(n6048), .A2(n6047), .ZN(n5218) );
  NAND2_X1 U5373 ( .A1(n5189), .A2(n4938), .ZN(n7975) );
  AND2_X1 U5374 ( .A1(n5194), .A2(n5864), .ZN(n5193) );
  OAI21_X1 U5375 ( .B1(n10511), .B2(n6183), .A(n5791), .ZN(n5792) );
  AOI21_X1 U5376 ( .B1(n5187), .B2(n5949), .A(n4911), .ZN(n5180) );
  NAND2_X1 U5377 ( .A1(n5652), .A2(n5651), .ZN(n6237) );
  NAND2_X1 U5378 ( .A1(n4916), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5092) );
  AND2_X1 U5379 ( .A1(n6820), .A2(n6819), .ZN(n7340) );
  NAND2_X1 U5380 ( .A1(n9732), .A2(n9740), .ZN(n5068) );
  AOI21_X1 U5381 ( .B1(n5316), .B2(n9700), .A(n5312), .ZN(n5311) );
  AND2_X1 U5382 ( .A1(n6182), .A2(n6181), .ZN(n9763) );
  NAND2_X1 U5383 ( .A1(n9780), .A2(n5314), .ZN(n5313) );
  AND2_X1 U5384 ( .A1(n9698), .A2(n9446), .ZN(n9781) );
  NAND2_X1 U5385 ( .A1(n9943), .A2(n9680), .ZN(n5096) );
  NOR2_X1 U5386 ( .A1(n9814), .A2(n5095), .ZN(n5094) );
  INV_X1 U5387 ( .A(n5440), .ZN(n5095) );
  NAND2_X1 U5388 ( .A1(n9693), .A2(n9451), .ZN(n5323) );
  NAND2_X1 U5389 ( .A1(n9695), .A2(n4922), .ZN(n5322) );
  AND2_X1 U5390 ( .A1(n5322), .A2(n5320), .ZN(n9805) );
  NAND2_X1 U5391 ( .A1(n9827), .A2(n9832), .ZN(n9826) );
  NOR2_X1 U5392 ( .A1(n5075), .A2(n4949), .ZN(n5074) );
  NOR2_X1 U5393 ( .A1(n5076), .A2(n4917), .ZN(n5075) );
  AND2_X1 U5394 ( .A1(n9694), .A2(n9829), .ZN(n9850) );
  OR2_X1 U5395 ( .A1(n9675), .A2(n9674), .ZN(n5483) );
  NOR2_X1 U5396 ( .A1(n5444), .A2(n5448), .ZN(n5441) );
  NAND2_X1 U5397 ( .A1(n8010), .A2(n5302), .ZN(n5301) );
  OR2_X1 U5398 ( .A1(n5871), .A2(n5870), .ZN(n5890) );
  NAND2_X1 U5399 ( .A1(n5435), .A2(n5434), .ZN(n7805) );
  AOI21_X1 U5400 ( .B1(n5437), .B2(n5439), .A(n4944), .ZN(n5434) );
  INV_X1 U5401 ( .A(n9569), .ZN(n10534) );
  OR2_X1 U5402 ( .A1(n7672), .A2(n7665), .ZN(n7666) );
  NAND2_X1 U5403 ( .A1(n4908), .A2(n9471), .ZN(n10531) );
  XNOR2_X1 U5404 ( .A(n7234), .B(n5284), .ZN(n9406) );
  INV_X1 U5405 ( .A(n10531), .ZN(n9887) );
  OR2_X1 U5406 ( .A1(n10512), .A2(n6030), .ZN(n7253) );
  NAND2_X1 U5407 ( .A1(n6203), .A2(n6202), .ZN(n9916) );
  INV_X1 U5408 ( .A(n9849), .ZN(n9953) );
  INV_X1 U5409 ( .A(n7576), .ZN(n10511) );
  INV_X1 U5410 ( .A(n7547), .ZN(n10503) );
  NAND2_X1 U5411 ( .A1(n6224), .A2(n6223), .ZN(n6823) );
  INV_X1 U5412 ( .A(n5160), .ZN(n5465) );
  NOR2_X1 U5413 ( .A1(n4910), .A2(n5157), .ZN(n5156) );
  NAND2_X1 U5414 ( .A1(n5594), .A2(n5477), .ZN(n5157) );
  AND2_X1 U5415 ( .A1(n5594), .A2(n5307), .ZN(n5158) );
  NAND2_X1 U5416 ( .A1(n5160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5605) );
  INV_X1 U5417 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U5418 ( .A1(n5590), .A2(n5477), .ZN(n5611) );
  NAND2_X1 U5419 ( .A1(n6101), .A2(n6099), .ZN(n6122) );
  NAND2_X1 U5420 ( .A1(n6089), .A2(n6087), .ZN(n6068) );
  XNOR2_X1 U5421 ( .A(n5332), .B(n6087), .ZN(n7732) );
  INV_X1 U5422 ( .A(n6089), .ZN(n5332) );
  OAI21_X2 U5423 ( .B1(n5611), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  INV_X1 U5424 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U5425 ( .A1(n5103), .A2(n5527), .ZN(n5846) );
  NAND2_X1 U5426 ( .A1(n5109), .A2(n5107), .ZN(n5103) );
  NAND2_X1 U5427 ( .A1(n5202), .A2(n5513), .ZN(n5758) );
  NAND2_X1 U5428 ( .A1(n5742), .A2(n5741), .ZN(n5202) );
  AND2_X1 U5429 ( .A1(n5762), .A2(n5761), .ZN(n7353) );
  NAND2_X1 U5430 ( .A1(n4987), .A2(n5400), .ZN(n4991) );
  INV_X1 U5431 ( .A(n8207), .ZN(n4987) );
  NAND2_X1 U5432 ( .A1(n6545), .A2(n6544), .ZN(n8862) );
  NAND2_X1 U5433 ( .A1(n8212), .A2(n8180), .ZN(n8246) );
  AND2_X1 U5434 ( .A1(n7116), .A2(n5402), .ZN(n5401) );
  INV_X1 U5435 ( .A(n5479), .ZN(n5402) );
  INV_X1 U5436 ( .A(n8326), .ZN(n8657) );
  INV_X1 U5437 ( .A(n10642), .ZN(n10656) );
  INV_X1 U5438 ( .A(n8222), .ZN(n8798) );
  OAI21_X1 U5439 ( .B1(n8611), .B2(n8639), .A(n5381), .ZN(n5380) );
  AOI21_X1 U5440 ( .B1(n8610), .B2(n8617), .A(n5382), .ZN(n5381) );
  NAND2_X1 U5441 ( .A1(n6892), .A2(n6859), .ZN(n10418) );
  OAI21_X1 U5442 ( .B1(n8640), .B2(n8639), .A(n4985), .ZN(n4984) );
  NAND2_X1 U5443 ( .A1(n8638), .A2(n10412), .ZN(n4985) );
  XNOR2_X1 U5444 ( .A(n8652), .B(n8655), .ZN(n8815) );
  NAND2_X1 U5445 ( .A1(n6642), .A2(n6641), .ZN(n8680) );
  OAI21_X1 U5446 ( .B1(n8710), .B2(n8446), .A(n8445), .ZN(n8697) );
  OAI21_X1 U5447 ( .B1(n8765), .B2(n5024), .A(n5026), .ZN(n8840) );
  AOI21_X1 U5448 ( .B1(n5027), .B2(n5029), .A(n8742), .ZN(n5026) );
  INV_X1 U5449 ( .A(n5027), .ZN(n5024) );
  AND3_X1 U5450 ( .A1(n6388), .A2(n6387), .A3(n6386), .ZN(n10470) );
  OR2_X1 U5451 ( .A1(n6384), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U5452 ( .A1(n6706), .A2(n6705), .ZN(n7000) );
  INV_X1 U5453 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U5454 ( .A1(n5959), .A2(n5958), .ZN(n9986) );
  NAND2_X1 U5455 ( .A1(n6833), .A2(n9273), .ZN(n5125) );
  NAND2_X1 U5456 ( .A1(n6034), .A2(n6033), .ZN(n9960) );
  NAND2_X1 U5457 ( .A1(n6274), .A2(n5470), .ZN(n9181) );
  AND2_X1 U5458 ( .A1(n6115), .A2(n6114), .ZN(n9809) );
  INV_X1 U5459 ( .A(n8002), .ZN(n10626) );
  AND4_X1 U5460 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n8004)
         );
  AND3_X1 U5461 ( .A1(n5642), .A2(n5641), .A3(n5640), .ZN(n9808) );
  NAND2_X1 U5462 ( .A1(n5664), .A2(n5663), .ZN(n9964) );
  NAND2_X1 U5463 ( .A1(n6270), .A2(n6192), .ZN(n6274) );
  AND2_X1 U5464 ( .A1(n6272), .A2(n6271), .ZN(n6192) );
  AND4_X1 U5465 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(n8108)
         );
  NAND2_X1 U5466 ( .A1(n6263), .A2(n4908), .ZN(n9264) );
  NAND2_X1 U5467 ( .A1(n5974), .A2(n5973), .ZN(n9980) );
  INV_X1 U5468 ( .A(n9763), .ZN(n9684) );
  NAND2_X1 U5469 ( .A1(n6136), .A2(n6135), .ZN(n9681) );
  OR2_X1 U5470 ( .A1(n9777), .A2(n6207), .ZN(n6136) );
  INV_X1 U5471 ( .A(n9834), .ZN(n9680) );
  INV_X1 U5472 ( .A(n9808), .ZN(n9851) );
  INV_X1 U5473 ( .A(n8004), .ZN(n9561) );
  OR2_X1 U5474 ( .A1(n8157), .A2(n10512), .ZN(n5150) );
  NAND2_X1 U5475 ( .A1(n9712), .A2(n9711), .ZN(n5295) );
  AOI21_X1 U5476 ( .B1(n9710), .B2(n9889), .A(n9709), .ZN(n9711) );
  INV_X1 U5477 ( .A(n5455), .ZN(n5454) );
  AND2_X1 U5478 ( .A1(n6174), .A2(n6173), .ZN(n9757) );
  INV_X1 U5479 ( .A(n6030), .ZN(n9778) );
  NAND2_X1 U5480 ( .A1(n9868), .A2(n7399), .ZN(n9896) );
  AND2_X1 U5481 ( .A1(n5150), .A2(n5149), .ZN(n9992) );
  AOI21_X1 U5482 ( .B1(n9902), .B2(n10490), .A(n9901), .ZN(n5149) );
  INV_X1 U5483 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U5484 ( .A1(n5135), .A2(n5134), .ZN(n8374) );
  NAND2_X1 U5485 ( .A1(n8378), .A2(n8473), .ZN(n5135) );
  NAND2_X1 U5486 ( .A1(n5127), .A2(n4931), .ZN(n8399) );
  NAND2_X1 U5487 ( .A1(n5101), .A2(n5100), .ZN(n9337) );
  OR2_X1 U5488 ( .A1(n9330), .A2(n9394), .ZN(n5101) );
  AND2_X1 U5489 ( .A1(n9332), .A2(n4959), .ZN(n5100) );
  OAI21_X1 U5490 ( .B1(n8422), .B2(n5142), .A(n5140), .ZN(n5139) );
  INV_X1 U5491 ( .A(n8421), .ZN(n5142) );
  NAND2_X1 U5492 ( .A1(n5098), .A2(n9336), .ZN(n9334) );
  NAND2_X1 U5493 ( .A1(n9337), .A2(n5099), .ZN(n5098) );
  AND2_X1 U5494 ( .A1(n9510), .A2(n9333), .ZN(n5099) );
  OAI21_X1 U5495 ( .B1(n5330), .B2(n8443), .A(n8442), .ZN(n5327) );
  NAND2_X1 U5496 ( .A1(n5328), .A2(n5326), .ZN(n8454) );
  NAND2_X1 U5497 ( .A1(n5329), .A2(n8477), .ZN(n5328) );
  NAND2_X1 U5498 ( .A1(n5327), .A2(n8473), .ZN(n5326) );
  OAI21_X1 U5499 ( .B1(n5330), .B2(n8440), .A(n8439), .ZN(n5329) );
  NAND2_X1 U5500 ( .A1(n9360), .A2(n9394), .ZN(n5116) );
  NAND2_X1 U5501 ( .A1(n9359), .A2(n9383), .ZN(n5117) );
  INV_X1 U5502 ( .A(n9366), .ZN(n5115) );
  INV_X1 U5503 ( .A(n9317), .ZN(n9318) );
  NAND2_X1 U5504 ( .A1(n5111), .A2(n5110), .ZN(n9367) );
  NAND2_X1 U5505 ( .A1(n9451), .A2(n9394), .ZN(n5110) );
  AND2_X1 U5506 ( .A1(n9781), .A2(n9373), .ZN(n5124) );
  INV_X1 U5507 ( .A(SI_20_), .ZN(n9020) );
  INV_X1 U5508 ( .A(SI_16_), .ZN(n9030) );
  INV_X1 U5509 ( .A(SI_14_), .ZN(n9034) );
  INV_X1 U5510 ( .A(SI_11_), .ZN(n9035) );
  NOR2_X1 U5511 ( .A1(n8471), .A2(n8472), .ZN(n5351) );
  NOR2_X1 U5512 ( .A1(n8474), .A2(n8473), .ZN(n5350) );
  INV_X1 U5513 ( .A(n5056), .ZN(n5054) );
  NAND2_X1 U5514 ( .A1(n6508), .A2(n6507), .ZN(n5263) );
  NAND2_X1 U5515 ( .A1(n5267), .A2(n7868), .ZN(n5266) );
  INV_X1 U5516 ( .A(n8870), .ZN(n5267) );
  NOR2_X1 U5517 ( .A1(n6520), .A2(n5265), .ZN(n5264) );
  INV_X1 U5518 ( .A(n6507), .ZN(n5265) );
  INV_X1 U5519 ( .A(n7623), .ZN(n5258) );
  OR2_X1 U5520 ( .A1(n8123), .A2(n6006), .ZN(n5199) );
  INV_X1 U5521 ( .A(n5794), .ZN(n5172) );
  NAND2_X1 U5522 ( .A1(n10617), .A2(n5154), .ZN(n5153) );
  INV_X1 U5523 ( .A(n5568), .ZN(n5335) );
  INV_X1 U5524 ( .A(SI_12_), .ZN(n9037) );
  INV_X1 U5525 ( .A(n5882), .ZN(n5343) );
  INV_X1 U5526 ( .A(n5513), .ZN(n5203) );
  INV_X1 U5527 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5581) );
  OR2_X1 U5528 ( .A1(n7867), .A2(n8530), .ZN(n7865) );
  AND2_X1 U5529 ( .A1(n5388), .A2(n8240), .ZN(n5387) );
  NAND2_X1 U5530 ( .A1(n8249), .A2(n8183), .ZN(n5388) );
  AND2_X1 U5531 ( .A1(n5353), .A2(n6957), .ZN(n5352) );
  AOI21_X1 U5532 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8598), .A(n10396), .ZN(
        n8599) );
  OR2_X1 U5533 ( .A1(n10405), .A2(n8599), .ZN(n8624) );
  NAND2_X1 U5534 ( .A1(n5487), .A2(n4925), .ZN(n5255) );
  INV_X1 U5535 ( .A(n5252), .ZN(n5049) );
  NOR2_X1 U5536 ( .A1(n5049), .A2(n5254), .ZN(n5047) );
  NAND2_X1 U5537 ( .A1(n8656), .A2(n5252), .ZN(n5046) );
  NAND2_X1 U5538 ( .A1(n8703), .A2(n5283), .ZN(n5282) );
  INV_X1 U5539 ( .A(n8446), .ZN(n5283) );
  AOI21_X1 U5540 ( .B1(n8703), .B2(n8447), .A(n5484), .ZN(n5281) );
  NOR2_X1 U5541 ( .A1(n8218), .A2(n8713), .ZN(n5278) );
  NAND2_X1 U5542 ( .A1(n5242), .A2(n8362), .ZN(n5243) );
  NAND2_X1 U5543 ( .A1(n8322), .A2(n7611), .ZN(n7047) );
  INV_X1 U5544 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6308) );
  OR2_X1 U5545 ( .A1(n6408), .A2(n6326), .ZN(n6468) );
  NOR2_X1 U5546 ( .A1(n4914), .A2(n4936), .ZN(n5219) );
  NAND2_X1 U5547 ( .A1(n5817), .A2(n7521), .ZN(n5220) );
  NAND2_X1 U5548 ( .A1(n5207), .A2(n5206), .ZN(n6082) );
  NOR2_X1 U5549 ( .A1(n5209), .A2(n4951), .ZN(n5206) );
  NOR2_X1 U5550 ( .A1(n7764), .A2(n7765), .ZN(n5192) );
  NAND2_X1 U5551 ( .A1(n7764), .A2(n7765), .ZN(n5194) );
  NOR2_X1 U5552 ( .A1(n5192), .A2(n5191), .ZN(n5190) );
  INV_X1 U5553 ( .A(n5861), .ZN(n5191) );
  AND2_X1 U5554 ( .A1(n5680), .A2(n5615), .ZN(n6046) );
  OAI21_X1 U5556 ( .B1(n5121), .B2(n5118), .A(n4948), .ZN(n9385) );
  NAND2_X1 U5557 ( .A1(n5120), .A2(n5119), .ZN(n5118) );
  NOR2_X1 U5558 ( .A1(n9748), .A2(n5310), .ZN(n5309) );
  INV_X1 U5559 ( .A(n5314), .ZN(n5310) );
  INV_X1 U5560 ( .A(n9701), .ZN(n5312) );
  NOR2_X1 U5561 ( .A1(n5167), .A2(n9934), .ZN(n5165) );
  INV_X1 U5562 ( .A(n9850), .ZN(n5072) );
  NOR2_X1 U5563 ( .A1(n9850), .A2(n9677), .ZN(n5070) );
  OR2_X1 U5564 ( .A1(n5442), .A2(n9353), .ZN(n5078) );
  INV_X1 U5565 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5996) );
  NOR2_X1 U5566 ( .A1(n5087), .A2(n7949), .ZN(n5081) );
  OR2_X1 U5567 ( .A1(n5914), .A2(n5913), .ZN(n5936) );
  INV_X1 U5568 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5870) );
  INV_X1 U5569 ( .A(n5438), .ZN(n5437) );
  OAI21_X1 U5570 ( .B1(n7744), .B2(n5439), .A(n7773), .ZN(n5438) );
  INV_X1 U5571 ( .A(n7747), .ZN(n5439) );
  NAND2_X1 U5572 ( .A1(n10536), .A2(n7674), .ZN(n7677) );
  NAND2_X1 U5573 ( .A1(n5289), .A2(n9405), .ZN(n10535) );
  INV_X1 U5574 ( .A(n7680), .ZN(n5289) );
  NAND2_X1 U5575 ( .A1(n7395), .A2(n7496), .ZN(n9489) );
  INV_X1 U5576 ( .A(n6251), .ZN(n9471) );
  AND2_X1 U5577 ( .A1(n9499), .A2(n9496), .ZN(n5285) );
  INV_X1 U5578 ( .A(n9544), .ZN(n7244) );
  NAND2_X1 U5579 ( .A1(n7394), .A2(n7393), .ZN(n7485) );
  NAND2_X1 U5580 ( .A1(n7485), .A2(n7484), .ZN(n7663) );
  NAND2_X1 U5581 ( .A1(n7300), .A2(n7235), .ZN(n7236) );
  NAND2_X1 U5582 ( .A1(n7236), .A2(n9399), .ZN(n7394) );
  NOR2_X1 U5583 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5629) );
  XNOR2_X1 U5584 ( .A(n8144), .B(n8142), .ZN(n8152) );
  OAI21_X1 U5585 ( .B1(n6198), .B2(n6197), .A(n6196), .ZN(n6653) );
  AND2_X1 U5586 ( .A1(n6654), .A2(n6201), .ZN(n6652) );
  AND2_X1 U5587 ( .A1(n6149), .A2(n6125), .ZN(n6147) );
  INV_X1 U5588 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U5589 ( .A1(n5331), .A2(n5547), .ZN(n5953) );
  NAND2_X1 U5590 ( .A1(n5930), .A2(n5545), .ZN(n5331) );
  OAI21_X1 U5591 ( .B1(n5533), .B2(n5342), .A(n5340), .ZN(n5901) );
  INV_X1 U5592 ( .A(n5341), .ZN(n5340) );
  OAI21_X1 U5593 ( .B1(n5344), .B2(n5342), .A(n5541), .ZN(n5341) );
  NAND2_X1 U5594 ( .A1(n5343), .A2(n5535), .ZN(n5342) );
  NOR2_X1 U5595 ( .A1(n5826), .A2(n5108), .ZN(n5107) );
  INV_X1 U5596 ( .A(n5523), .ZN(n5108) );
  OAI21_X1 U5597 ( .B1(n6656), .B2(n4993), .A(n4992), .ZN(n5512) );
  NAND2_X1 U5598 ( .A1(n6656), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4992) );
  NOR2_X1 U5599 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5704) );
  NAND2_X1 U5600 ( .A1(n5499), .A2(n6355), .ZN(n5691) );
  NAND2_X1 U5601 ( .A1(n5493), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5494) );
  OR2_X1 U5602 ( .A1(n8170), .A2(n8798), .ZN(n5424) );
  NAND2_X1 U5603 ( .A1(n8169), .A2(n5420), .ZN(n5419) );
  NAND2_X1 U5604 ( .A1(n7553), .A2(n7554), .ZN(n5432) );
  OR2_X1 U5605 ( .A1(n7379), .A2(n7380), .ZN(n5433) );
  INV_X1 U5606 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U5607 ( .A1(n5389), .A2(n8181), .ZN(n8247) );
  NAND2_X1 U5608 ( .A1(n5346), .A2(n8477), .ZN(n5132) );
  OR2_X1 U5609 ( .A1(n5346), .A2(n4962), .ZN(n5133) );
  AOI21_X1 U5610 ( .B1(n5348), .B2(n5347), .A(n8318), .ZN(n5346) );
  OR2_X1 U5611 ( .A1(n8508), .A2(n8322), .ZN(n5129) );
  AND2_X1 U5612 ( .A1(n8510), .A2(n8651), .ZN(n5130) );
  INV_X1 U5613 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U5614 ( .A1(n5035), .A2(n5033), .ZN(n5037) );
  OR2_X1 U5615 ( .A1(n6374), .A2(n6358), .ZN(n6361) );
  OR2_X1 U5616 ( .A1(n6677), .A2(n6839), .ZN(n6351) );
  OR2_X1 U5617 ( .A1(n6376), .A2(n6997), .ZN(n5022) );
  OR2_X1 U5618 ( .A1(n6378), .A2(n6349), .ZN(n6352) );
  NAND2_X1 U5619 ( .A1(n6867), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U5620 ( .A1(n5366), .A2(n6959), .ZN(n7033) );
  AND2_X1 U5621 ( .A1(n7032), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5366) );
  NOR2_X1 U5622 ( .A1(n8582), .A2(n4997), .ZN(n10303) );
  AND2_X1 U5623 ( .A1(n8583), .A2(n8584), .ZN(n4997) );
  NOR2_X1 U5624 ( .A1(n8588), .A2(n10317), .ZN(n10335) );
  NAND2_X1 U5625 ( .A1(n8608), .A2(n5383), .ZN(n5382) );
  NOR2_X1 U5626 ( .A1(n8605), .A2(n5384), .ZN(n5383) );
  OR2_X1 U5627 ( .A1(n8211), .A2(n8272), .ZN(n5487) );
  INV_X1 U5628 ( .A(n6644), .ZN(n6645) );
  AND2_X1 U5629 ( .A1(n8828), .A2(n8524), .ZN(n8446) );
  INV_X1 U5630 ( .A(n8732), .ZN(n8713) );
  INV_X1 U5631 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9075) );
  AND4_X1 U5632 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n8724)
         );
  AND4_X1 U5633 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n8725)
         );
  INV_X1 U5634 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8258) );
  AND2_X1 U5635 ( .A1(n6599), .A2(n8258), .ZN(n6607) );
  INV_X1 U5636 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8974) );
  AND2_X1 U5637 ( .A1(n6588), .A2(n8974), .ZN(n6599) );
  INV_X1 U5638 ( .A(n6578), .ZN(n6579) );
  AND2_X1 U5639 ( .A1(n6577), .A2(n6576), .ZN(n8171) );
  AND4_X1 U5640 ( .A1(n6552), .A2(n6551), .A3(n6550), .A4(n6549), .ZN(n8802)
         );
  NAND2_X1 U5641 ( .A1(n5251), .A2(n5250), .ZN(n5039) );
  NAND2_X1 U5642 ( .A1(n6537), .A2(n6536), .ZN(n7898) );
  NAND2_X1 U5643 ( .A1(n7626), .A2(n5056), .ZN(n5052) );
  AOI21_X1 U5644 ( .B1(n5010), .B2(n8491), .A(n5009), .ZN(n5008) );
  INV_X1 U5645 ( .A(n8375), .ZN(n5009) );
  NOR2_X1 U5646 ( .A1(n5240), .A2(n5244), .ZN(n5010) );
  INV_X1 U5647 ( .A(n8531), .ZN(n7843) );
  INV_X1 U5648 ( .A(n5240), .ZN(n5014) );
  NAND2_X1 U5649 ( .A1(n5248), .A2(n5244), .ZN(n5013) );
  NAND2_X1 U5650 ( .A1(n5013), .A2(n5011), .ZN(n7624) );
  INV_X1 U5651 ( .A(n5012), .ZN(n5011) );
  INV_X1 U5652 ( .A(n8532), .ZN(n7841) );
  AND4_X1 U5653 ( .A1(n6466), .A2(n6465), .A3(n6464), .A4(n6463), .ZN(n7598)
         );
  OAI22_X1 U5654 ( .A1(n7138), .A2(n5269), .B1(n5271), .B2(n5268), .ZN(n6440)
         );
  NAND2_X1 U5655 ( .A1(n6732), .A2(n8361), .ZN(n7286) );
  OR2_X1 U5656 ( .A1(n7178), .A2(n8354), .ZN(n6732) );
  NAND2_X1 U5657 ( .A1(n5273), .A2(n6411), .ZN(n7181) );
  NAND2_X1 U5658 ( .A1(n5274), .A2(n5275), .ZN(n5273) );
  INV_X1 U5659 ( .A(n7138), .ZN(n5274) );
  CLKBUF_X1 U5660 ( .A(n6357), .Z(n8643) );
  AND2_X1 U5661 ( .A1(n8351), .A2(n8356), .ZN(n8479) );
  NAND2_X1 U5662 ( .A1(n7129), .A2(n8343), .ZN(n7099) );
  NAND2_X1 U5663 ( .A1(n5023), .A2(n5021), .ZN(n7129) );
  NAND2_X1 U5664 ( .A1(n6739), .A2(n8455), .ZN(n8704) );
  NOR2_X1 U5665 ( .A1(n8447), .A2(n8446), .ZN(n8709) );
  INV_X1 U5666 ( .A(n8782), .ZN(n8781) );
  INV_X1 U5667 ( .A(n8795), .ZN(n8792) );
  AOI21_X1 U5668 ( .B1(n5004), .B2(n5007), .A(n5003), .ZN(n5002) );
  INV_X1 U5669 ( .A(n8414), .ZN(n5003) );
  NAND2_X1 U5670 ( .A1(n5260), .A2(n6507), .ZN(n7823) );
  OR2_X1 U5671 ( .A1(n7635), .A2(n6508), .ZN(n5260) );
  NAND2_X1 U5672 ( .A1(n8339), .A2(n7820), .ZN(n8844) );
  NAND2_X1 U5673 ( .A1(n6687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6718) );
  NAND2_X1 U5674 ( .A1(n6692), .A2(n6686), .ZN(n6687) );
  OR2_X1 U5675 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  INV_X1 U5676 ( .A(n6973), .ZN(n7750) );
  NAND2_X1 U5677 ( .A1(n6671), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6672) );
  INV_X1 U5678 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6670) );
  AND2_X1 U5679 ( .A1(n6456), .A2(n6453), .ZN(n7150) );
  INV_X1 U5680 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6435) );
  INV_X1 U5681 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6420) );
  OR2_X1 U5682 ( .A1(n6324), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U5683 ( .A1(n5842), .A2(n5843), .ZN(n7706) );
  NAND2_X1 U5684 ( .A1(n8122), .A2(n8123), .ZN(n8121) );
  NOR2_X1 U5685 ( .A1(n6780), .A2(n5174), .ZN(n5173) );
  INV_X1 U5686 ( .A(n6776), .ZN(n5174) );
  INV_X1 U5687 ( .A(n5183), .ZN(n5178) );
  AOI21_X1 U5688 ( .B1(n5187), .B2(n5182), .A(n8049), .ZN(n5181) );
  AND2_X1 U5689 ( .A1(n5949), .A2(n4911), .ZN(n5182) );
  AND2_X1 U5690 ( .A1(n9191), .A2(n9190), .ZN(n9276) );
  AND4_X1 U5691 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n7734)
         );
  NOR2_X1 U5692 ( .A1(n5461), .A2(n5457), .ZN(n5456) );
  INV_X1 U5693 ( .A(n9685), .ZN(n5457) );
  AOI21_X1 U5694 ( .B1(n9747), .B2(n9685), .A(n5459), .ZN(n9732) );
  OR2_X1 U5695 ( .A1(n9734), .A2(n6207), .ZN(n6213) );
  NAND2_X1 U5696 ( .A1(n9835), .A2(n5165), .ZN(n9775) );
  AND2_X1 U5697 ( .A1(n6160), .A2(n6159), .ZN(n9786) );
  OR2_X1 U5698 ( .A1(n6108), .A2(n6107), .ZN(n6129) );
  INV_X1 U5699 ( .A(n5319), .ZN(n5317) );
  INV_X1 U5700 ( .A(n9695), .ZN(n5318) );
  AOI21_X1 U5701 ( .B1(n5320), .B2(n9452), .A(n5324), .ZN(n5319) );
  NAND2_X1 U5702 ( .A1(n9835), .A2(n9819), .ZN(n9816) );
  OR2_X1 U5703 ( .A1(n6055), .A2(n5626), .ZN(n6073) );
  AND2_X1 U5704 ( .A1(n6079), .A2(n6078), .ZN(n9834) );
  OR2_X1 U5705 ( .A1(n5997), .A2(n5996), .ZN(n6014) );
  NAND2_X1 U5706 ( .A1(n5623), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6037) );
  INV_X1 U5707 ( .A(n6014), .ZN(n5623) );
  NAND2_X1 U5708 ( .A1(n5301), .A2(n5299), .ZN(n8112) );
  AOI21_X1 U5709 ( .B1(n5299), .B2(n9339), .A(n5297), .ZN(n5296) );
  INV_X1 U5710 ( .A(n5299), .ZN(n5298) );
  NAND2_X1 U5711 ( .A1(n5446), .A2(n5445), .ZN(n8099) );
  NAND2_X1 U5712 ( .A1(n8024), .A2(n5447), .ZN(n5446) );
  AOI21_X1 U5713 ( .B1(n7806), .B2(n5087), .A(n4953), .ZN(n5084) );
  NOR2_X1 U5714 ( .A1(n7777), .A2(n7803), .ZN(n7813) );
  NOR3_X1 U5715 ( .A1(n7777), .A2(n7981), .A3(n7803), .ZN(n7889) );
  OR2_X1 U5716 ( .A1(n7672), .A2(n7671), .ZN(n10522) );
  NAND2_X1 U5717 ( .A1(n9405), .A2(n9303), .ZN(n9300) );
  AND2_X1 U5718 ( .A1(n5161), .A2(n7415), .ZN(n5162) );
  AND2_X1 U5719 ( .A1(n9491), .A2(n9493), .ZN(n9400) );
  NAND2_X1 U5720 ( .A1(n5163), .A2(n9279), .ZN(n7492) );
  NAND2_X1 U5721 ( .A1(n7242), .A2(n7243), .ZN(n7400) );
  NAND2_X1 U5722 ( .A1(n7240), .A2(n10450), .ZN(n8025) );
  NAND2_X1 U5723 ( .A1(n9395), .A2(n7831), .ZN(n10444) );
  AND2_X1 U5724 ( .A1(n9907), .A2(n10490), .ZN(n5294) );
  NAND2_X1 U5725 ( .A1(n8156), .A2(n8155), .ZN(n9910) );
  INV_X1 U5726 ( .A(n9757), .ZN(n9922) );
  OR2_X1 U5727 ( .A1(n9383), .A2(n7244), .ZN(n9990) );
  AND3_X1 U5728 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n10530) );
  AND2_X1 U5729 ( .A1(n10451), .A2(n7237), .ZN(n10490) );
  NAND2_X1 U5730 ( .A1(n8025), .A2(n9990), .ZN(n10628) );
  AND2_X1 U5731 ( .A1(n5680), .A2(n6825), .ZN(n6824) );
  XNOR2_X1 U5732 ( .A(n5603), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U5733 ( .A1(n5607), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5603) );
  OR2_X1 U5734 ( .A1(n6094), .A2(n6093), .ZN(n6100) );
  NAND2_X1 U5735 ( .A1(n6089), .A2(n6088), .ZN(n6101) );
  AND2_X1 U5736 ( .A1(n6087), .A2(n6090), .ZN(n6088) );
  XNOR2_X1 U5737 ( .A(n6239), .B(n6238), .ZN(n6821) );
  OAI21_X1 U5738 ( .B1(n6237), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U5739 ( .A1(n5612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5613) );
  INV_X1 U5740 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U5741 ( .A1(n5336), .A2(n5568), .ZN(n6029) );
  NAND2_X1 U5742 ( .A1(n5565), .A2(n5337), .ZN(n5336) );
  AND2_X1 U5743 ( .A1(n6009), .A2(n5993), .ZN(n9656) );
  AND2_X1 U5744 ( .A1(n5910), .A2(n5909), .ZN(n9634) );
  NAND2_X1 U5745 ( .A1(n5339), .A2(n5535), .ZN(n5883) );
  NAND2_X1 U5746 ( .A1(n5533), .A2(n5344), .ZN(n5339) );
  NAND2_X1 U5747 ( .A1(n5109), .A2(n5523), .ZN(n5827) );
  INV_X1 U5748 ( .A(n5405), .ZN(n7114) );
  NAND2_X1 U5749 ( .A1(n5419), .A2(n5417), .ZN(n8220) );
  NOR2_X1 U5750 ( .A1(n5392), .A2(n8195), .ZN(n5391) );
  INV_X1 U5751 ( .A(n5398), .ZN(n5392) );
  NAND2_X1 U5752 ( .A1(n5394), .A2(n4927), .ZN(n5393) );
  NAND2_X1 U5753 ( .A1(n5398), .A2(n5395), .ZN(n5394) );
  NAND2_X1 U5754 ( .A1(n5396), .A2(n5400), .ZN(n5395) );
  NAND2_X1 U5755 ( .A1(n8206), .A2(n8195), .ZN(n5397) );
  CLKBUF_X1 U5756 ( .A(n7054), .Z(n7091) );
  NAND2_X1 U5757 ( .A1(n6623), .A2(n6622), .ZN(n8824) );
  NAND2_X1 U5758 ( .A1(n7169), .A2(n7168), .ZN(n7198) );
  NOR2_X1 U5759 ( .A1(n7114), .A2(n5479), .ZN(n7117) );
  AND2_X1 U5760 ( .A1(n5428), .A2(n5426), .ZN(n5425) );
  INV_X1 U5761 ( .A(n7700), .ZN(n5426) );
  NAND2_X1 U5762 ( .A1(n5427), .A2(n5428), .ZN(n7699) );
  CLKBUF_X1 U5763 ( .A(n10659), .Z(n10664) );
  NOR2_X1 U5764 ( .A1(n4995), .A2(n7871), .ZN(n7925) );
  CLKBUF_X1 U5765 ( .A(n7870), .Z(n4995) );
  NAND2_X1 U5766 ( .A1(n8257), .A2(n8256), .ZN(n8255) );
  INV_X1 U5767 ( .A(n10641), .ZN(n10657) );
  AND4_X1 U5768 ( .A1(n6561), .A2(n6560), .A3(n6559), .A4(n6558), .ZN(n10643)
         );
  OR2_X1 U5769 ( .A1(n7060), .A2(n6990), .ZN(n10641) );
  NAND2_X1 U5770 ( .A1(n8169), .A2(n8168), .ZN(n10648) );
  AND2_X1 U5771 ( .A1(n7852), .A2(n8871), .ZN(n10667) );
  AND2_X1 U5772 ( .A1(n6981), .A2(n6980), .ZN(n10653) );
  INV_X1 U5773 ( .A(n7988), .ZN(n5406) );
  NAND2_X1 U5774 ( .A1(n5407), .A2(n5409), .ZN(n7989) );
  NAND2_X1 U5775 ( .A1(n6298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6299) );
  XNOR2_X1 U5776 ( .A(n6674), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8518) );
  INV_X1 U5777 ( .A(n8724), .ZN(n8744) );
  INV_X1 U5778 ( .A(n10643), .ZN(n8525) );
  INV_X1 U5779 ( .A(n7598), .ZN(n8533) );
  NAND4_X1 U5780 ( .A1(n6395), .A2(n6394), .A3(n6393), .A4(n6392), .ZN(n8538)
         );
  INV_X2 U5781 ( .A(P2_U3893), .ZN(n8580) );
  OAI21_X1 U5782 ( .B1(n6867), .B2(n5357), .A(n5356), .ZN(n10277) );
  NAND2_X1 U5783 ( .A1(n4980), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7215) );
  AOI21_X1 U5784 ( .B1(n7214), .B2(n5374), .A(n5373), .ZN(n5371) );
  INV_X1 U5785 ( .A(n5361), .ZN(n10349) );
  INV_X1 U5786 ( .A(n8592), .ZN(n5360) );
  INV_X1 U5787 ( .A(n5370), .ZN(n10380) );
  INV_X1 U5788 ( .A(n8596), .ZN(n5369) );
  AND2_X1 U5789 ( .A1(n6553), .A2(n6543), .ZN(n10387) );
  NAND2_X1 U5790 ( .A1(n6849), .A2(n6848), .ZN(n10404) );
  INV_X1 U5791 ( .A(n8642), .ZN(n8662) );
  INV_X1 U5792 ( .A(n5225), .ZN(n5224) );
  AOI21_X1 U5793 ( .B1(n5050), .B2(n5043), .A(n4913), .ZN(n5225) );
  NAND2_X1 U5794 ( .A1(n6763), .A2(n6762), .ZN(n6764) );
  XNOR2_X1 U5795 ( .A(n6761), .B(n8505), .ZN(n6765) );
  NAND2_X1 U5796 ( .A1(n6632), .A2(n6631), .ZN(n8820) );
  AND2_X1 U5797 ( .A1(n6615), .A2(n6614), .ZN(n8715) );
  NAND2_X1 U5798 ( .A1(n6606), .A2(n6605), .ZN(n8832) );
  NAND2_X1 U5799 ( .A1(n8738), .A2(n8737), .ZN(n8736) );
  NAND2_X1 U5800 ( .A1(n8840), .A2(n8438), .ZN(n8738) );
  NAND2_X1 U5801 ( .A1(n6597), .A2(n6596), .ZN(n8835) );
  NAND2_X1 U5802 ( .A1(n5025), .A2(n5027), .ZN(n8751) );
  OR2_X1 U5803 ( .A1(n5031), .A2(n5029), .ZN(n5025) );
  NAND2_X1 U5804 ( .A1(n6586), .A2(n6585), .ZN(n8749) );
  NAND2_X1 U5805 ( .A1(n7732), .A2(n8296), .ZN(n6586) );
  NAND2_X1 U5806 ( .A1(n5061), .A2(n5060), .ZN(n8755) );
  INV_X1 U5807 ( .A(n8171), .ZN(n10668) );
  AOI21_X1 U5808 ( .B1(n8766), .B2(n8767), .A(n8768), .ZN(n8774) );
  NAND2_X1 U5809 ( .A1(n6567), .A2(n6566), .ZN(n10649) );
  NAND2_X1 U5810 ( .A1(n6556), .A2(n6555), .ZN(n8858) );
  NAND2_X1 U5811 ( .A1(n7897), .A2(n8413), .ZN(n7967) );
  NAND2_X1 U5812 ( .A1(n6473), .A2(n6472), .ZN(n7703) );
  NAND2_X1 U5813 ( .A1(n5246), .A2(n8362), .ZN(n7590) );
  NAND2_X1 U5814 ( .A1(n5270), .A2(n6427), .ZN(n7287) );
  OAI21_X1 U5815 ( .B1(n7138), .B2(n6412), .A(n5271), .ZN(n5270) );
  OR2_X1 U5816 ( .A1(n7010), .A2(n10469), .ZN(n8649) );
  INV_X2 U5817 ( .A(n7621), .ZN(n8876) );
  OAI21_X1 U5818 ( .B1(n6739), .B2(n4920), .A(n5017), .ZN(n6768) );
  INV_X1 U5819 ( .A(n5229), .ZN(n5227) );
  OAI21_X1 U5820 ( .B1(n8840), .B2(n5239), .A(n5237), .ZN(n8719) );
  NAND2_X1 U5821 ( .A1(n5030), .A2(n5028), .ZN(n8761) );
  NAND2_X1 U5822 ( .A1(n5030), .A2(n8433), .ZN(n8759) );
  XNOR2_X1 U5823 ( .A(n6718), .B(n6719), .ZN(n6973) );
  AND2_X1 U5824 ( .A1(n6298), .A2(n6306), .ZN(n4999) );
  NAND2_X1 U5825 ( .A1(n6693), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6694) );
  BUF_X1 U5826 ( .A(n6698), .Z(n7920) );
  INV_X1 U5827 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7752) );
  INV_X1 U5828 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7692) );
  INV_X1 U5829 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7612) );
  INV_X1 U5830 ( .A(n8633), .ZN(n7611) );
  INV_X1 U5831 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7392) );
  INV_X1 U5832 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7319) );
  INV_X1 U5833 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7194) );
  INV_X1 U5834 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7125) );
  INV_X1 U5835 ( .A(n10290), .ZN(n8586) );
  INV_X1 U5836 ( .A(n7150), .ZN(n7209) );
  NOR2_X1 U5837 ( .A1(n8286), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9141) );
  XNOR2_X1 U5838 ( .A(n6421), .B(n6420), .ZN(n10270) );
  NAND2_X1 U5839 ( .A1(n6385), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5378) );
  CLKBUF_X1 U5840 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n4996) );
  AND4_X1 U5841 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n10532)
         );
  NAND2_X1 U5842 ( .A1(n5175), .A2(n5180), .ZN(n8048) );
  NAND2_X1 U5843 ( .A1(n7909), .A2(n5187), .ZN(n5175) );
  NAND2_X1 U5844 ( .A1(n7651), .A2(n5861), .ZN(n5195) );
  AND4_X1 U5845 ( .A1(n5752), .A2(n5751), .A3(n5750), .A4(n5749), .ZN(n7665)
         );
  NAND2_X1 U5846 ( .A1(n5700), .A2(n5699), .ZN(n7260) );
  INV_X1 U5847 ( .A(n5697), .ZN(n5700) );
  NAND2_X1 U5848 ( .A1(n5208), .A2(n5213), .ZN(n9203) );
  AND2_X1 U5849 ( .A1(n5207), .A2(n5205), .ZN(n9201) );
  NAND2_X1 U5850 ( .A1(n9163), .A2(n5212), .ZN(n5208) );
  INV_X1 U5851 ( .A(n9564), .ZN(n7914) );
  INV_X1 U5852 ( .A(n9975), .ZN(n8130) );
  NAND3_X1 U5853 ( .A1(n5765), .A2(n5764), .A3(n5763), .ZN(n7547) );
  INV_X1 U5854 ( .A(n9251), .ZN(n9262) );
  NAND2_X1 U5855 ( .A1(n8121), .A2(n5198), .ZN(n9218) );
  NAND2_X1 U5856 ( .A1(n6012), .A2(n6011), .ZN(n9970) );
  AND4_X1 U5857 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n7776)
         );
  OAI21_X1 U5858 ( .B1(n9163), .B2(n9164), .A(n5218), .ZN(n9233) );
  NAND2_X1 U5859 ( .A1(n7081), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9251) );
  INV_X1 U5860 ( .A(n9261), .ZN(n9250) );
  XNOR2_X1 U5861 ( .A(n5819), .B(n5818), .ZN(n7528) );
  NAND2_X1 U5862 ( .A1(n5221), .A2(n5782), .ZN(n7576) );
  AND2_X1 U5863 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  NAND2_X1 U5864 ( .A1(n6434), .A2(n9273), .ZN(n5221) );
  OAI211_X1 U5865 ( .C1(n5179), .C2(n7909), .A(n5177), .B(n5176), .ZN(n8060)
         );
  NAND2_X1 U5866 ( .A1(n5178), .A2(n5181), .ZN(n5177) );
  NAND2_X1 U5867 ( .A1(n5188), .A2(n5180), .ZN(n5176) );
  NOR2_X1 U5868 ( .A1(n5180), .A2(n5181), .ZN(n5179) );
  INV_X1 U5869 ( .A(n9243), .ZN(n9266) );
  OR2_X1 U5870 ( .A1(n5654), .A2(n7238), .ZN(n10450) );
  INV_X1 U5871 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5653) );
  AND2_X1 U5872 ( .A1(n6261), .A2(n6260), .ZN(n9741) );
  INV_X1 U5873 ( .A(n9809), .ZN(n9783) );
  INV_X1 U5874 ( .A(n7734), .ZN(n9566) );
  NAND4_X1 U5875 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .ZN(n9568)
         );
  NAND4_X1 U5876 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n9569)
         );
  NAND4_X1 U5877 ( .A1(n5734), .A2(n5733), .A3(n5732), .A4(n5731), .ZN(n9572)
         );
  NAND2_X1 U5878 ( .A1(n5786), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U5879 ( .A1(n9184), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5091) );
  INV_X1 U5880 ( .A(n10218), .ZN(n10431) );
  INV_X1 U5881 ( .A(n10222), .ZN(n10427) );
  INV_X1 U5882 ( .A(n9910), .ZN(n9722) );
  NAND2_X1 U5883 ( .A1(n5066), .A2(n5065), .ZN(n9914) );
  NAND2_X1 U5884 ( .A1(n5068), .A2(n5460), .ZN(n5065) );
  INV_X1 U5885 ( .A(n5067), .ZN(n5066) );
  AOI21_X1 U5886 ( .B1(n5068), .B2(n4921), .A(n9716), .ZN(n5067) );
  AND2_X1 U5887 ( .A1(n6205), .A2(n6176), .ZN(n9754) );
  INV_X1 U5888 ( .A(n5313), .ZN(n9760) );
  NAND2_X1 U5889 ( .A1(n9780), .A2(n9698), .ZN(n9761) );
  AND2_X1 U5890 ( .A1(n5097), .A2(n5096), .ZN(n9792) );
  NAND2_X1 U5891 ( .A1(n9826), .A2(n5440), .ZN(n9813) );
  NAND2_X1 U5892 ( .A1(n5322), .A2(n5323), .ZN(n9807) );
  AND2_X1 U5893 ( .A1(n6052), .A2(n6051), .ZN(n9849) );
  OAI21_X1 U5894 ( .B1(n9871), .B2(n5076), .A(n5074), .ZN(n9842) );
  NAND2_X1 U5895 ( .A1(n9871), .A2(n4917), .ZN(n9857) );
  INV_X1 U5896 ( .A(n9964), .ZN(n9880) );
  NAND2_X1 U5897 ( .A1(n8109), .A2(n9423), .ZN(n9676) );
  NAND2_X1 U5898 ( .A1(n5079), .A2(n5442), .ZN(n8109) );
  NAND2_X1 U5899 ( .A1(n8024), .A2(n5441), .ZN(n5079) );
  NAND2_X1 U5900 ( .A1(n8099), .A2(n8098), .ZN(n9973) );
  NAND2_X1 U5901 ( .A1(n5301), .A2(n9346), .ZN(n8110) );
  NAND2_X1 U5902 ( .A1(n8010), .A2(n9511), .ZN(n8094) );
  AND2_X1 U5903 ( .A1(n5449), .A2(n5452), .ZN(n8097) );
  NAND2_X1 U5904 ( .A1(n8024), .A2(n8023), .ZN(n5449) );
  NAND2_X1 U5905 ( .A1(n5935), .A2(n5934), .ZN(n8002) );
  INV_X1 U5906 ( .A(n7804), .ZN(n5086) );
  NAND2_X1 U5907 ( .A1(n7805), .A2(n9412), .ZN(n5088) );
  NAND2_X1 U5908 ( .A1(n5436), .A2(n7747), .ZN(n7774) );
  NAND2_X1 U5909 ( .A1(n7745), .A2(n7744), .ZN(n5436) );
  AND3_X1 U5910 ( .A1(n5747), .A2(n5746), .A3(n5745), .ZN(n7430) );
  OR2_X1 U5911 ( .A1(n5778), .A2(n6796), .ZN(n5746) );
  INV_X1 U5912 ( .A(n7234), .ZN(n7415) );
  AND3_X2 U5913 ( .A1(n7396), .A2(n7321), .A3(n7320), .ZN(n10632) );
  NAND2_X1 U5914 ( .A1(n6824), .A2(n6823), .ZN(n10027) );
  XNOR2_X1 U5915 ( .A(n8290), .B(n8289), .ZN(n10016) );
  MUX2_X1 U5916 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5632), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5635) );
  NAND2_X1 U5917 ( .A1(n5631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5632) );
  INV_X1 U5918 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U5919 ( .A1(n5305), .A2(n5304), .ZN(n5596) );
  AOI21_X1 U5920 ( .B1(n4926), .B2(n5307), .A(n5307), .ZN(n5304) );
  NAND2_X1 U5921 ( .A1(n5599), .A2(n5598), .ZN(n8162) );
  OR2_X1 U5922 ( .A1(n5597), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U5923 ( .A1(n5607), .A2(n5606), .ZN(n7896) );
  XNOR2_X1 U5924 ( .A(n5609), .B(n5608), .ZN(n7863) );
  NAND2_X1 U5925 ( .A1(n4923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5609) );
  INV_X1 U5926 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7757) );
  INV_X1 U5927 ( .A(n9550), .ZN(n7831) );
  INV_X1 U5928 ( .A(n6236), .ZN(n9395) );
  INV_X1 U5929 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U5930 ( .A1(n5662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5648) );
  AND2_X1 U5931 ( .A1(n5662), .A2(n5661), .ZN(n10214) );
  INV_X1 U5932 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7317) );
  INV_X1 U5933 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7192) );
  INV_X1 U5934 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7127) );
  INV_X1 U5935 ( .A(n6434), .ZN(n8133) );
  AND2_X1 U5936 ( .A1(n8210), .A2(n4975), .ZN(n4989) );
  NAND2_X1 U5937 ( .A1(n5385), .A2(n5379), .ZN(P2_U3200) );
  NAND2_X1 U5938 ( .A1(n8606), .A2(n8607), .ZN(n5385) );
  INV_X1 U5939 ( .A(n5380), .ZN(n5379) );
  NAND2_X1 U5940 ( .A1(n4986), .A2(n4983), .ZN(P2_U3201) );
  INV_X1 U5941 ( .A(n8637), .ZN(n4986) );
  INV_X1 U5942 ( .A(n4984), .ZN(n4983) );
  OR2_X1 U5943 ( .A1(n8669), .A2(n8865), .ZN(n6745) );
  OAI21_X1 U5944 ( .B1(n6241), .B2(n9182), .A(n9235), .ZN(n6269) );
  NOR2_X1 U5945 ( .A1(n6273), .A2(n6272), .ZN(n6282) );
  INV_X1 U5946 ( .A(n5150), .ZN(n9900) );
  NAND2_X1 U5947 ( .A1(n5295), .A2(n9868), .ZN(n9713) );
  OAI21_X1 U5948 ( .B1(n9992), .B2(n10633), .A(n5148), .ZN(P1_U3520) );
  OR2_X1 U5949 ( .A1(n10636), .A2(n9993), .ZN(n5148) );
  INV_X1 U5950 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7518) );
  OAI21_X1 U5951 ( .B1(n5949), .B2(n5928), .A(n4940), .ZN(n5188) );
  AND2_X4 U5952 ( .A1(n10021), .A2(n10022), .ZN(n4918) );
  INV_X1 U5953 ( .A(n4916), .ZN(n9187) );
  INV_X1 U5954 ( .A(n5461), .ZN(n5460) );
  NAND2_X1 U5955 ( .A1(n9716), .A2(n4921), .ZN(n5461) );
  XOR2_X1 U5956 ( .A(n5969), .B(n6216), .Z(n4911) );
  INV_X1 U5957 ( .A(n8098), .ZN(n5444) );
  INV_X1 U5958 ( .A(n5029), .ZN(n5028) );
  NAND2_X1 U5959 ( .A1(n5032), .A2(n8433), .ZN(n5029) );
  NAND2_X1 U5960 ( .A1(n6820), .A2(n8141), .ZN(n5703) );
  INV_X1 U5961 ( .A(n9346), .ZN(n5300) );
  AND2_X1 U5962 ( .A1(n8219), .A2(n10656), .ZN(n4912) );
  INV_X1 U5963 ( .A(n8488), .ZN(n5242) );
  NAND2_X1 U5964 ( .A1(n9459), .A2(n9462), .ZN(n9740) );
  AND2_X1 U5965 ( .A1(n8660), .A2(n8723), .ZN(n4913) );
  INV_X1 U5966 ( .A(n9791), .ZN(n5325) );
  AND2_X1 U5967 ( .A1(n5823), .A2(n5822), .ZN(n4914) );
  NOR2_X1 U5968 ( .A1(n9514), .A2(n5303), .ZN(n5302) );
  NAND2_X1 U5969 ( .A1(n6127), .A2(n6126), .ZN(n9934) );
  XNOR2_X1 U5970 ( .A(n6694), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6700) );
  OR2_X1 U5971 ( .A1(n9950), .A2(n9808), .ZN(n9451) );
  AND2_X1 U5972 ( .A1(n5165), .A2(n5164), .ZN(n4915) );
  INV_X1 U5973 ( .A(n5018), .ZN(n5017) );
  OAI21_X1 U5974 ( .B1(n4920), .B2(n8455), .A(n5226), .ZN(n5018) );
  OR2_X1 U5975 ( .A1(n8851), .A2(n10642), .ZN(n8327) );
  INV_X1 U5976 ( .A(n8219), .ZN(n5423) );
  INV_X1 U5977 ( .A(n6006), .ZN(n5198) );
  INV_X1 U5978 ( .A(n5188), .ZN(n5187) );
  NAND2_X1 U5979 ( .A1(n10534), .A2(n7576), .ZN(n9405) );
  AND3_X1 U5980 ( .A1(n5707), .A2(n5706), .A3(n5705), .ZN(n9279) );
  INV_X2 U5981 ( .A(n6357), .ZN(n6367) );
  OR2_X1 U5982 ( .A1(n9880), .A2(n9866), .ZN(n4917) );
  NAND2_X1 U5983 ( .A1(n5634), .A2(n5633), .ZN(n5636) );
  INV_X1 U5984 ( .A(n8765), .ZN(n5031) );
  OR2_X1 U5985 ( .A1(n8086), .A2(n8525), .ZN(n4919) );
  OR2_X1 U5986 ( .A1(n8703), .A2(n6741), .ZN(n4920) );
  INV_X1 U5987 ( .A(n8530), .ZN(n7868) );
  NAND2_X1 U5988 ( .A1(n5145), .A2(n5581), .ZN(n5759) );
  OR2_X1 U5989 ( .A1(n9916), .A2(n9726), .ZN(n4921) );
  AND2_X1 U5990 ( .A1(n9451), .A2(n9694), .ZN(n4922) );
  OR2_X1 U5991 ( .A1(n5611), .A2(n5592), .ZN(n4923) );
  NAND2_X1 U5992 ( .A1(n8247), .A2(n8183), .ZN(n8239) );
  AND2_X1 U5993 ( .A1(n5313), .A2(n9699), .ZN(n4924) );
  NOR2_X1 U5994 ( .A1(n8680), .A2(n8688), .ZN(n4925) );
  AND2_X1 U5995 ( .A1(n5594), .A2(n5306), .ZN(n4926) );
  INV_X1 U5996 ( .A(n6371), .ZN(n6991) );
  OR2_X1 U5997 ( .A1(n5398), .A2(n8195), .ZN(n4927) );
  INV_X1 U5998 ( .A(n8206), .ZN(n5400) );
  AND2_X1 U5999 ( .A1(n5082), .A2(n5080), .ZN(n4928) );
  AND4_X1 U6000 ( .A1(n6686), .A2(n6696), .A3(n6689), .A4(n6719), .ZN(n4929)
         );
  OR2_X1 U6001 ( .A1(n9906), .A2(n5294), .ZN(n4930) );
  INV_X1 U6002 ( .A(n8535), .ZN(n7599) );
  OR2_X1 U6003 ( .A1(n8749), .A2(n8259), .ZN(n8438) );
  AND3_X1 U6004 ( .A1(n8386), .A2(n8492), .A3(n5126), .ZN(n4931) );
  INV_X1 U6005 ( .A(n5949), .ZN(n5185) );
  AND2_X1 U6006 ( .A1(n5084), .A2(n5083), .ZN(n4932) );
  AND2_X1 U6007 ( .A1(n8327), .A2(n8433), .ZN(n8768) );
  INV_X1 U6008 ( .A(n8768), .ZN(n5064) );
  AND2_X1 U6009 ( .A1(n9980), .A2(n9560), .ZN(n4933) );
  INV_X1 U6010 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6298) );
  AND2_X1 U6011 ( .A1(n8413), .A2(n8412), .ZN(n8478) );
  INV_X1 U6012 ( .A(n8478), .ZN(n5040) );
  OR2_X1 U6013 ( .A1(n9934), .A2(n9798), .ZN(n9698) );
  INV_X1 U6014 ( .A(n9698), .ZN(n5315) );
  OR2_X1 U6015 ( .A1(n8437), .A2(n8477), .ZN(n4934) );
  INV_X1 U6016 ( .A(n9748), .ZN(n5316) );
  AND4_X1 U6017 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n7627)
         );
  INV_X1 U6018 ( .A(n7627), .ZN(n5136) );
  INV_X1 U6019 ( .A(n5527), .ZN(n5106) );
  NOR2_X1 U6020 ( .A1(n7981), .A2(n9564), .ZN(n4935) );
  NOR2_X1 U6021 ( .A1(n5820), .A2(n7602), .ZN(n4936) );
  OR2_X1 U6022 ( .A1(n7869), .A2(n7868), .ZN(n4937) );
  NAND2_X1 U6023 ( .A1(n9835), .A2(n5166), .ZN(n5169) );
  OR2_X1 U6024 ( .A1(n5193), .A2(n5192), .ZN(n4938) );
  INV_X1 U6025 ( .A(n5087), .ZN(n5085) );
  NOR2_X1 U6026 ( .A1(n4935), .A2(n7804), .ZN(n5087) );
  AND2_X1 U6027 ( .A1(n5471), .A2(n8401), .ZN(n4939) );
  OR2_X1 U6028 ( .A1(n5951), .A2(n5950), .ZN(n4940) );
  AND2_X1 U6029 ( .A1(n5061), .A2(n5062), .ZN(n4941) );
  OR2_X1 U6030 ( .A1(n8421), .A2(n8473), .ZN(n4942) );
  INV_X1 U6031 ( .A(n5421), .ZN(n5420) );
  OR2_X1 U6032 ( .A1(n10647), .A2(n5422), .ZN(n5421) );
  AND2_X1 U6033 ( .A1(n5370), .A2(n5369), .ZN(n4943) );
  OR2_X1 U6034 ( .A1(n9943), .A2(n9834), .ZN(n9370) );
  NOR2_X1 U6035 ( .A1(n7775), .A2(n9566), .ZN(n4944) );
  NOR2_X1 U6036 ( .A1(n8130), .A2(n8108), .ZN(n4945) );
  NOR2_X1 U6037 ( .A1(n9722), .A2(n9741), .ZN(n4946) );
  AND2_X1 U6038 ( .A1(n8672), .A2(n8657), .ZN(n4947) );
  INV_X1 U6039 ( .A(n8742), .ZN(n8750) );
  INV_X1 U6040 ( .A(n5167), .ZN(n5166) );
  NAND2_X1 U6041 ( .A1(n9819), .A2(n5168), .ZN(n5167) );
  AND2_X1 U6042 ( .A1(n9725), .A2(n9381), .ZN(n4948) );
  AND2_X1 U6043 ( .A1(n6523), .A2(n6522), .ZN(n8406) );
  NOR2_X1 U6044 ( .A1(n9859), .A2(n9678), .ZN(n4949) );
  NOR2_X1 U6045 ( .A1(n10668), .A2(n8770), .ZN(n4950) );
  NOR2_X1 U6046 ( .A1(n6065), .A2(n6066), .ZN(n4951) );
  INV_X1 U6047 ( .A(n9677), .ZN(n5076) );
  OR2_X1 U6048 ( .A1(n9960), .A2(n9888), .ZN(n9677) );
  NOR2_X1 U6049 ( .A1(n9953), .A2(n9679), .ZN(n4952) );
  NOR2_X1 U6050 ( .A1(n10607), .A2(n7914), .ZN(n4953) );
  INV_X1 U6051 ( .A(n5448), .ZN(n5447) );
  NAND2_X1 U6052 ( .A1(n5451), .A2(n8023), .ZN(n5448) );
  NAND2_X1 U6053 ( .A1(n5228), .A2(n5227), .ZN(n4954) );
  AND2_X1 U6054 ( .A1(n5199), .A2(n9216), .ZN(n4955) );
  INV_X1 U6055 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5608) );
  OR2_X1 U6056 ( .A1(n8866), .A2(n8527), .ZN(n4956) );
  NAND2_X1 U6057 ( .A1(n8851), .A2(n10656), .ZN(n4957) );
  INV_X1 U6058 ( .A(n5418), .ZN(n5417) );
  NAND2_X1 U6059 ( .A1(n5423), .A2(n5424), .ZN(n5418) );
  AND2_X1 U6060 ( .A1(n5239), .A2(n8449), .ZN(n4958) );
  OR2_X1 U6061 ( .A1(n9331), .A2(n9383), .ZN(n4959) );
  AND3_X1 U6062 ( .A1(n5730), .A2(n5729), .A3(n5728), .ZN(n10478) );
  INV_X1 U6063 ( .A(n5251), .ZN(n5041) );
  NOR2_X1 U6064 ( .A1(n8528), .A2(n7934), .ZN(n5251) );
  AND2_X1 U6065 ( .A1(n6351), .A2(n7051), .ZN(n4960) );
  OR2_X1 U6066 ( .A1(n4933), .A2(n5450), .ZN(n4961) );
  OR2_X1 U6067 ( .A1(n5231), .A2(n8703), .ZN(n5228) );
  OR2_X1 U6068 ( .A1(n9986), .A2(n8004), .ZN(n9511) );
  INV_X1 U6069 ( .A(n9511), .ZN(n5303) );
  OR2_X1 U6070 ( .A1(n9922), .A2(n9763), .ZN(n9460) );
  INV_X1 U6071 ( .A(n9460), .ZN(n5122) );
  AND2_X1 U6072 ( .A1(n8650), .A2(n8477), .ZN(n4962) );
  AND2_X1 U6073 ( .A1(n10617), .A2(n7974), .ZN(n4963) );
  INV_X1 U6074 ( .A(n8758), .ZN(n5032) );
  AND2_X1 U6075 ( .A1(n9423), .A2(n5441), .ZN(n4964) );
  AND3_X1 U6076 ( .A1(n5589), .A2(n5992), .A3(n5647), .ZN(n5477) );
  INV_X1 U6077 ( .A(n5477), .ZN(n5159) );
  AND2_X1 U6078 ( .A1(n5521), .A2(n5527), .ZN(n4965) );
  AND2_X1 U6079 ( .A1(n5016), .A2(n8505), .ZN(n4966) );
  AND2_X1 U6080 ( .A1(n5409), .A2(n5406), .ZN(n4967) );
  AND2_X1 U6081 ( .A1(n5078), .A2(n5483), .ZN(n4968) );
  INV_X1 U6082 ( .A(n5005), .ZN(n5004) );
  NAND2_X1 U6083 ( .A1(n5006), .A2(n8417), .ZN(n5005) );
  NAND2_X1 U6084 ( .A1(n6106), .A2(n6105), .ZN(n9939) );
  INV_X1 U6085 ( .A(n9939), .ZN(n5168) );
  NAND2_X1 U6086 ( .A1(n9826), .A2(n5094), .ZN(n5097) );
  NAND2_X1 U6087 ( .A1(n6152), .A2(n6151), .ZN(n9929) );
  INV_X1 U6088 ( .A(n9929), .ZN(n5164) );
  NAND2_X1 U6089 ( .A1(n5908), .A2(n5464), .ZN(n5955) );
  AND2_X1 U6090 ( .A1(n7909), .A2(n5928), .ZN(n7911) );
  AOI21_X2 U6091 ( .B1(n7437), .B2(n6483), .A(n5468), .ZN(n7626) );
  OR2_X1 U6092 ( .A1(n6028), .A2(n5335), .ZN(n4969) );
  AND2_X1 U6093 ( .A1(n5908), .A2(n5586), .ZN(n5932) );
  INV_X1 U6094 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5364) );
  INV_X1 U6095 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6096 ( .A1(n6734), .A2(n8401), .ZN(n7833) );
  AND4_X1 U6097 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(n7994)
         );
  INV_X1 U6098 ( .A(n7909), .ZN(n5186) );
  AOI21_X1 U6099 ( .B1(n4995), .B2(n7922), .A(n5411), .ZN(n5408) );
  AND2_X1 U6100 ( .A1(n5361), .A2(n5360), .ZN(n4970) );
  OR2_X1 U6101 ( .A1(n7911), .A2(n5949), .ZN(n4971) );
  INV_X1 U6102 ( .A(n8249), .ZN(n8181) );
  AND2_X1 U6103 ( .A1(n5419), .A2(n5424), .ZN(n4972) );
  NAND2_X1 U6104 ( .A1(n5184), .A2(n5183), .ZN(n4973) );
  INV_X1 U6105 ( .A(n5462), .ZN(n5459) );
  NAND2_X1 U6106 ( .A1(n9922), .A2(n9684), .ZN(n5462) );
  AND2_X1 U6107 ( .A1(n5042), .A2(n5041), .ZN(n4974) );
  OR2_X1 U6108 ( .A1(n8211), .A2(n8277), .ZN(n4975) );
  NAND2_X1 U6109 ( .A1(n5125), .A2(n5869), .ZN(n7803) );
  INV_X1 U6110 ( .A(n7803), .ZN(n5154) );
  INV_X1 U6111 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6112 ( .A1(n5195), .A2(n5864), .ZN(n7763) );
  INV_X1 U6113 ( .A(n6702), .ZN(n6703) );
  NAND2_X1 U6114 ( .A1(n7663), .A2(n7661), .ZN(n7431) );
  INV_X1 U6115 ( .A(n5151), .ZN(n7953) );
  NOR3_X1 U6116 ( .A1(n7777), .A2(n5153), .A3(n7981), .ZN(n5151) );
  INV_X1 U6117 ( .A(n6412), .ZN(n5275) );
  NAND2_X1 U6118 ( .A1(n6024), .A2(n6023), .ZN(n4976) );
  AND2_X1 U6119 ( .A1(n5088), .A2(n5086), .ZN(n4977) );
  AND2_X1 U6120 ( .A1(n5433), .A2(n5432), .ZN(n4978) );
  AND2_X1 U6121 ( .A1(n5233), .A2(n6735), .ZN(n4979) );
  INV_X1 U6122 ( .A(n5452), .ZN(n5450) );
  NAND2_X1 U6123 ( .A1(n9986), .A2(n9561), .ZN(n5452) );
  INV_X1 U6124 ( .A(n10636), .ZN(n10633) );
  AND2_X1 U6125 ( .A1(n7148), .A2(n7214), .ZN(n4980) );
  NAND2_X1 U6126 ( .A1(n8320), .A2(n6749), .ZN(n8793) );
  NAND2_X1 U6127 ( .A1(n5162), .A2(n10478), .ZN(n4981) );
  NAND4_X1 U6128 ( .A1(n5092), .A2(n5091), .A3(n5090), .A4(n5089), .ZN(n5284)
         );
  INV_X1 U6129 ( .A(n7031), .ZN(n5365) );
  INV_X1 U6130 ( .A(n7213), .ZN(n5373) );
  NAND2_X1 U6131 ( .A1(n7415), .A2(n10445), .ZN(n7412) );
  INV_X1 U6132 ( .A(n7412), .ZN(n5163) );
  NAND2_X1 U6133 ( .A1(n4960), .A2(n5019), .ZN(n8340) );
  INV_X1 U6134 ( .A(n8340), .ZN(n5021) );
  AND2_X1 U6135 ( .A1(n6959), .A2(n7032), .ZN(n4982) );
  XNOR2_X1 U6136 ( .A(n6673), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8507) );
  INV_X1 U6137 ( .A(n8507), .ZN(n8322) );
  INV_X1 U6138 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5036) );
  XNOR2_X1 U6139 ( .A(n8587), .B(n10309), .ZN(n10318) );
  OAI21_X1 U6140 ( .B1(n5372), .B2(n7148), .A(n5371), .ZN(n7449) );
  NAND2_X1 U6141 ( .A1(n6904), .A2(n6903), .ZN(n6902) );
  OAI21_X1 U6142 ( .B1(n5363), .B2(n6959), .A(n5362), .ZN(n7146) );
  NAND2_X1 U6143 ( .A1(n8592), .A2(n8593), .ZN(n5358) );
  NAND2_X1 U6144 ( .A1(n8596), .A2(n8597), .ZN(n5367) );
  AOI22_X1 U6145 ( .A1(n7198), .A2(n7197), .B1(n7196), .B2(n7289), .ZN(n7201)
         );
  NAND2_X1 U6146 ( .A1(n7378), .A2(n7377), .ZN(n7379) );
  OR2_X1 U6147 ( .A1(n8232), .A2(n8228), .ZN(n8174) );
  NAND2_X1 U6148 ( .A1(n4988), .A2(n4937), .ZN(n7870) );
  NAND2_X1 U6149 ( .A1(n4990), .A2(n4989), .ZN(P2_U3154) );
  NAND2_X1 U6150 ( .A1(n7866), .A2(n7865), .ZN(n4988) );
  INV_X1 U6151 ( .A(n6692), .ZN(n6685) );
  NAND3_X1 U6152 ( .A1(n4991), .A2(n8205), .A3(n10665), .ZN(n4990) );
  AOI21_X2 U6153 ( .B1(n6699), .B2(n6704), .A(n8018), .ZN(n6702) );
  NAND2_X1 U6154 ( .A1(n8174), .A2(n8229), .ZN(n8257) );
  NAND2_X1 U6155 ( .A1(n5204), .A2(n5516), .ZN(n5777) );
  NOR2_X2 U6156 ( .A1(n9538), .A2(n9392), .ZN(n9469) );
  NAND2_X4 U6157 ( .A1(n4994), .A2(n7049), .ZN(n7050) );
  NAND2_X2 U6158 ( .A1(n7045), .A2(n7046), .ZN(n4994) );
  INV_X1 U6159 ( .A(n6293), .ZN(n6563) );
  NAND2_X1 U6160 ( .A1(n5407), .A2(n4967), .ZN(n8039) );
  OAI21_X1 U6161 ( .B1(n7069), .B2(n8539), .A(n7068), .ZN(n7070) );
  NAND2_X1 U6162 ( .A1(n5405), .A2(n5401), .ZN(n7169) );
  OAI21_X1 U6163 ( .B1(n8084), .B2(n8083), .A(n5473), .ZN(n8167) );
  XNOR2_X2 U6164 ( .A(n7050), .B(n7310), .ZN(n7052) );
  XNOR2_X1 U6165 ( .A(n8583), .B(n8584), .ZN(n7450) );
  NAND2_X1 U6166 ( .A1(n8207), .A2(n8206), .ZN(n8205) );
  NAND3_X1 U6167 ( .A1(n5413), .A2(n6293), .A3(n4999), .ZN(n9138) );
  INV_X1 U6168 ( .A(n5233), .ZN(n5001) );
  OAI21_X1 U6169 ( .B1(n5001), .B2(n5005), .A(n5002), .ZN(n8072) );
  OAI21_X1 U6170 ( .B1(n5012), .B2(n5248), .A(n5008), .ZN(n7637) );
  AND2_X1 U6171 ( .A1(n5013), .A2(n5014), .ZN(n5490) );
  INV_X1 U6172 ( .A(n6739), .ZN(n5015) );
  OAI21_X1 U6173 ( .B1(n5015), .B2(n5018), .A(n4966), .ZN(n6767) );
  INV_X1 U6174 ( .A(n7128), .ZN(n5023) );
  AND2_X1 U6175 ( .A1(n5022), .A2(n5020), .ZN(n5019) );
  NAND2_X1 U6176 ( .A1(n5019), .A2(n6351), .ZN(n7132) );
  AND2_X1 U6177 ( .A1(n6352), .A2(n6350), .ZN(n5020) );
  OR2_X2 U6178 ( .A1(n8204), .A2(n9146), .ZN(n6376) );
  INV_X1 U6179 ( .A(n8204), .ZN(n6313) );
  AND2_X1 U6180 ( .A1(n5038), .A2(n5039), .ZN(n5249) );
  NAND4_X1 U6181 ( .A1(n6537), .A2(n6536), .A3(n5250), .A4(n5040), .ZN(n5038)
         );
  NAND3_X1 U6182 ( .A1(n6537), .A2(n5040), .A3(n6536), .ZN(n5042) );
  INV_X1 U6183 ( .A(n5042), .ZN(n7900) );
  NAND2_X1 U6184 ( .A1(n8766), .A2(n5060), .ZN(n5059) );
  NAND2_X1 U6185 ( .A1(n7302), .A2(n7301), .ZN(n7300) );
  INV_X1 U6186 ( .A(n9871), .ZN(n5073) );
  NAND2_X1 U6187 ( .A1(n8024), .A2(n4964), .ZN(n5077) );
  NAND2_X1 U6188 ( .A1(n5077), .A2(n4968), .ZN(n9872) );
  OAI21_X1 U6189 ( .B1(n7805), .B2(n5085), .A(n5084), .ZN(n7950) );
  AOI21_X1 U6190 ( .B1(n5084), .B2(n5081), .A(n4963), .ZN(n5080) );
  NAND2_X1 U6191 ( .A1(n7805), .A2(n4932), .ZN(n5082) );
  NAND2_X1 U6192 ( .A1(n4918), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5089) );
  INV_X1 U6193 ( .A(n5097), .ZN(n9812) );
  NAND2_X1 U6194 ( .A1(n5799), .A2(n5521), .ZN(n5109) );
  NAND2_X1 U6195 ( .A1(n5799), .A2(n4965), .ZN(n5102) );
  NAND3_X1 U6196 ( .A1(n5117), .A2(n5116), .A3(n5115), .ZN(n5114) );
  NAND3_X1 U6197 ( .A1(n5131), .A2(n5130), .A3(n5129), .ZN(n8512) );
  NAND3_X1 U6198 ( .A1(n5133), .A2(n5132), .A3(n8322), .ZN(n5131) );
  NAND3_X1 U6199 ( .A1(n8382), .A2(n8380), .A3(n8477), .ZN(n5134) );
  NAND3_X1 U6200 ( .A1(n5138), .A2(n8768), .A3(n8430), .ZN(n8431) );
  NAND3_X1 U6201 ( .A1(n5139), .A2(n8781), .A3(n8427), .ZN(n5138) );
  AND2_X1 U6202 ( .A1(n5291), .A2(n5145), .ZN(n5908) );
  OR2_X1 U6203 ( .A1(n6820), .A2(n7344), .ZN(n5146) );
  OR2_X1 U6204 ( .A1(n5778), .A2(n5497), .ZN(n5147) );
  NAND2_X2 U6205 ( .A1(n6820), .A2(n8286), .ZN(n5778) );
  NAND2_X2 U6206 ( .A1(n8162), .A2(n6245), .ZN(n6820) );
  NAND2_X1 U6207 ( .A1(n5590), .A2(n5155), .ZN(n5160) );
  AOI21_X1 U6208 ( .B1(n5590), .B2(n5156), .A(n5158), .ZN(n5597) );
  NAND4_X1 U6209 ( .A1(n10478), .A2(n5161), .A3(n7415), .A4(n7430), .ZN(n7425)
         );
  INV_X1 U6210 ( .A(n5169), .ZN(n9799) );
  NAND2_X1 U6211 ( .A1(n5702), .A2(n5701), .ZN(n5505) );
  NAND2_X1 U6212 ( .A1(n5170), .A2(n5502), .ZN(n5702) );
  NAND2_X1 U6213 ( .A1(n5691), .A2(n5500), .ZN(n5170) );
  NAND2_X1 U6214 ( .A1(n5720), .A2(n5719), .ZN(n7533) );
  NAND2_X1 U6215 ( .A1(n7651), .A2(n5190), .ZN(n5189) );
  OAI21_X1 U6216 ( .B1(n5742), .B2(n5203), .A(n5200), .ZN(n5204) );
  INV_X1 U6217 ( .A(n5201), .ZN(n5200) );
  OAI21_X1 U6218 ( .B1(n5203), .B2(n5741), .A(n5514), .ZN(n5201) );
  INV_X1 U6219 ( .A(n7132), .ZN(n7092) );
  OAI21_X1 U6220 ( .B1(n8815), .B2(n8661), .A(n5224), .ZN(n8811) );
  INV_X1 U6221 ( .A(n8840), .ZN(n5234) );
  OAI21_X1 U6222 ( .B1(n5234), .B2(n5236), .A(n5235), .ZN(n8708) );
  INV_X1 U6223 ( .A(n7286), .ZN(n5248) );
  NAND2_X1 U6224 ( .A1(n6733), .A2(n8391), .ZN(n7822) );
  NAND2_X1 U6225 ( .A1(n6731), .A2(n8357), .ZN(n7178) );
  NAND2_X1 U6226 ( .A1(n6767), .A2(n8467), .ZN(n8294) );
  NAND2_X1 U6227 ( .A1(n6729), .A2(n8346), .ZN(n7106) );
  NAND2_X1 U6228 ( .A1(n9156), .A2(n9157), .ZN(n9155) );
  NAND2_X1 U6229 ( .A1(n7258), .A2(n7257), .ZN(n7256) );
  INV_X1 U6230 ( .A(n5415), .ZN(n5414) );
  OAI21_X1 U6231 ( .B1(n6651), .B2(n4925), .A(n5487), .ZN(n8654) );
  INV_X1 U6232 ( .A(n6427), .ZN(n5268) );
  INV_X1 U6233 ( .A(n9406), .ZN(n7302) );
  NAND2_X1 U6234 ( .A1(n7305), .A2(n9406), .ZN(n7304) );
  NOR2_X1 U6235 ( .A1(n5286), .A2(n5285), .ZN(n5287) );
  NAND2_X1 U6236 ( .A1(n7680), .A2(n9499), .ZN(n5288) );
  INV_X2 U6237 ( .A(n5643), .ZN(n5590) );
  NAND3_X1 U6238 ( .A1(n5585), .A2(n5582), .A3(n5581), .ZN(n5292) );
  OAI21_X1 U6239 ( .B1(n8010), .B2(n5298), .A(n5296), .ZN(n8111) );
  NAND2_X1 U6240 ( .A1(n5465), .A2(n4926), .ZN(n5305) );
  INV_X1 U6241 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6242 ( .A1(n9780), .A2(n5309), .ZN(n5308) );
  NAND2_X1 U6243 ( .A1(n5308), .A2(n5311), .ZN(n9739) );
  NOR2_X2 U6244 ( .A1(n9806), .A2(n5321), .ZN(n5320) );
  OAI21_X2 U6245 ( .B1(n5953), .B2(n5952), .A(n5551), .ZN(n5971) );
  NAND2_X1 U6246 ( .A1(n5565), .A2(n5564), .ZN(n5659) );
  OAI21_X2 U6247 ( .B1(n5565), .B2(n4969), .A(n5333), .ZN(n6050) );
  NAND2_X1 U6248 ( .A1(n5533), .A2(n5532), .ZN(n5866) );
  NAND2_X1 U6249 ( .A1(n6867), .A2(n5356), .ZN(n5354) );
  NAND2_X1 U6250 ( .A1(n10273), .A2(n6390), .ZN(n5355) );
  NAND2_X1 U6251 ( .A1(n5354), .A2(n5352), .ZN(n6958) );
  NAND3_X1 U6252 ( .A1(n5355), .A2(n10272), .A3(n5357), .ZN(n5353) );
  AOI21_X1 U6253 ( .B1(n7032), .B2(n5364), .A(n5365), .ZN(n5362) );
  INV_X1 U6254 ( .A(n7032), .ZN(n5363) );
  OAI21_X1 U6255 ( .B1(n10381), .B2(n5368), .A(n5367), .ZN(n10396) );
  INV_X1 U6256 ( .A(n7214), .ZN(n5372) );
  MUX2_X1 U6257 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10476), .S(n6863), .Z(n6904)
         );
  INV_X1 U6258 ( .A(n8246), .ZN(n5389) );
  NAND2_X1 U6259 ( .A1(n5386), .A2(n5387), .ZN(n8187) );
  NAND2_X1 U6260 ( .A1(n8246), .A2(n8183), .ZN(n5386) );
  NAND2_X1 U6261 ( .A1(n8268), .A2(n5391), .ZN(n5390) );
  OAI211_X1 U6262 ( .C1(n8269), .C2(n5397), .A(n5393), .B(n5390), .ZN(n8200)
         );
  INV_X1 U6263 ( .A(n7071), .ZN(n5403) );
  INV_X1 U6264 ( .A(n7070), .ZN(n5404) );
  OR2_X2 U6265 ( .A1(n7870), .A2(n5411), .ZN(n5407) );
  NAND2_X1 U6266 ( .A1(n6293), .A2(n6292), .ZN(n6303) );
  AND2_X2 U6267 ( .A1(n5427), .A2(n5425), .ZN(n7718) );
  OR2_X2 U6268 ( .A1(n7379), .A2(n5430), .ZN(n5427) );
  INV_X1 U6269 ( .A(n5433), .ZN(n7552) );
  OR2_X1 U6270 ( .A1(n7697), .A2(n8533), .ZN(n5431) );
  NAND2_X1 U6271 ( .A1(n7745), .A2(n5437), .ZN(n5435) );
  NAND2_X1 U6272 ( .A1(n9747), .A2(n5456), .ZN(n5453) );
  NAND2_X1 U6273 ( .A1(n5453), .A2(n5454), .ZN(n9686) );
  NAND2_X1 U6274 ( .A1(n6695), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U6275 ( .A1(n6269), .A2(n6268), .ZN(P1_U3214) );
  NAND2_X1 U6276 ( .A1(n7542), .A2(n7544), .ZN(n7521) );
  INV_X1 U6277 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U6278 ( .A1(n5605), .A2(n5604), .ZN(n5607) );
  INV_X1 U6279 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6451) );
  CLKBUF_X1 U6280 ( .A(n8079), .Z(n8040) );
  NAND2_X1 U6281 ( .A1(n6691), .A2(n6695), .ZN(n6698) );
  INV_X1 U6282 ( .A(n5786), .ZN(n6257) );
  INV_X1 U6283 ( .A(n9184), .ZN(n6207) );
  NAND2_X1 U6284 ( .A1(n9184), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U6285 ( .A(n7050), .B(n10470), .ZN(n7069) );
  NOR2_X1 U6286 ( .A1(n9796), .A2(n9697), .ZN(n9782) );
  AOI22_X1 U6287 ( .A1(n9774), .A2(n9683), .B1(n9682), .B2(n9798), .ZN(n9765)
         );
  NOR2_X1 U6288 ( .A1(n6475), .A2(n6462), .ZN(n5467) );
  NOR2_X1 U6289 ( .A1(n6482), .A2(n7581), .ZN(n5468) );
  AND2_X1 U6290 ( .A1(n6759), .A2(n6758), .ZN(n5469) );
  AND2_X1 U6291 ( .A1(n6220), .A2(n6219), .ZN(n5470) );
  AND2_X1 U6292 ( .A1(n9396), .A2(n9435), .ZN(n10539) );
  INV_X1 U6293 ( .A(n10539), .ZN(n9892) );
  OR2_X1 U6294 ( .A1(n7877), .A2(n8405), .ZN(n5471) );
  AND2_X1 U6295 ( .A1(n5987), .A2(n8057), .ZN(n5472) );
  OR2_X1 U6296 ( .A1(n8677), .A2(n9134), .ZN(n5475) );
  NAND2_X1 U6297 ( .A1(n4929), .A2(n6294), .ZN(n5476) );
  AND2_X1 U6298 ( .A1(n8629), .A2(n8628), .ZN(n5478) );
  AND4_X1 U6299 ( .A1(n6593), .A2(n6592), .A3(n6591), .A4(n6590), .ZN(n8259)
         );
  AND2_X1 U6300 ( .A1(n7113), .A2(n8538), .ZN(n5479) );
  AND2_X1 U6301 ( .A1(n8535), .A2(n7199), .ZN(n5480) );
  OR2_X1 U6302 ( .A1(n8535), .A2(n7199), .ZN(n5481) );
  INV_X1 U6303 ( .A(n9986), .ZN(n8005) );
  AND2_X1 U6304 ( .A1(n8701), .A2(n8712), .ZN(n5484) );
  OR2_X1 U6305 ( .A1(n8325), .A2(n8844), .ZN(n5485) );
  OR2_X1 U6306 ( .A1(n8677), .A2(n8865), .ZN(n5486) );
  INV_X1 U6307 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5497) );
  INV_X1 U6308 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U6309 ( .A1(n9588), .A2(n9471), .ZN(n10533) );
  INV_X1 U6310 ( .A(n10533), .ZN(n9889) );
  INV_X1 U6311 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6525) );
  INV_X1 U6312 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6474) );
  INV_X1 U6313 ( .A(SI_28_), .ZN(n8137) );
  AND2_X1 U6314 ( .A1(n5532), .A2(n5531), .ZN(n5488) );
  XOR2_X1 U6315 ( .A(n8633), .B(P2_REG2_REG_19__SCAN_IN), .Z(n5489) );
  INV_X1 U6316 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6294) );
  OAI21_X1 U6317 ( .B1(n8339), .B2(n8507), .A(n7047), .ZN(n7048) );
  INV_X1 U6318 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U6319 ( .A1(n9300), .A2(n7660), .ZN(n7664) );
  NOR2_X1 U6320 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5591) );
  INV_X1 U6321 ( .A(n7048), .ZN(n7049) );
  INV_X1 U6322 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6686) );
  INV_X1 U6323 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6107) );
  INV_X1 U6324 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5830) );
  INV_X1 U6325 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9078) );
  INV_X1 U6326 ( .A(n8259), .ZN(n6594) );
  INV_X1 U6327 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U6328 ( .A1(n5656), .A2(n5683), .ZN(n5708) );
  INV_X1 U6329 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6275) );
  INV_X1 U6330 ( .A(n6053), .ZN(n5625) );
  INV_X1 U6331 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5913) );
  OR2_X1 U6332 ( .A1(n6175), .A2(n6275), .ZN(n6205) );
  OR2_X1 U6333 ( .A1(n5831), .A2(n5830), .ZN(n5851) );
  INV_X1 U6334 ( .A(SI_30_), .ZN(n9010) );
  INV_X1 U6335 ( .A(SI_24_), .ZN(n9017) );
  INV_X1 U6336 ( .A(SI_17_), .ZN(n8930) );
  INV_X1 U6337 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5586) );
  INV_X1 U6338 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5491) );
  AND2_X1 U6339 ( .A1(n6661), .A2(n6660), .ZN(n8642) );
  NAND2_X1 U6340 ( .A1(n6607), .A2(n9075), .ZN(n6616) );
  INV_X1 U6341 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U6342 ( .A1(n7043), .A2(n7045), .ZN(n7002) );
  OR2_X1 U6343 ( .A1(n8477), .A2(n7047), .ZN(n6753) );
  INV_X1 U6344 ( .A(n10177), .ZN(n9637) );
  NAND2_X1 U6345 ( .A1(n7078), .A2(n5688), .ZN(n5697) );
  NAND2_X1 U6346 ( .A1(n6117), .A2(n6119), .ZN(n6120) );
  OR2_X1 U6347 ( .A1(n7958), .A2(n7959), .ZN(n5949) );
  NAND2_X1 U6348 ( .A1(n5625), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6055) );
  OR2_X1 U6349 ( .A1(n5936), .A2(n7961), .ZN(n5961) );
  INV_X1 U6350 ( .A(n9741), .ZN(n9710) );
  OR2_X1 U6351 ( .A1(n6154), .A2(n6153), .ZN(n6175) );
  AND2_X1 U6352 ( .A1(n6100), .A2(n6098), .ZN(n6099) );
  INV_X1 U6353 ( .A(SI_10_), .ZN(n8940) );
  NAND2_X1 U6354 ( .A1(n7376), .A2(n8535), .ZN(n7377) );
  INV_X1 U6355 ( .A(n8167), .ZN(n8085) );
  NOR2_X1 U6356 ( .A1(n6557), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6568) );
  INV_X1 U6357 ( .A(n10655), .ZN(n10644) );
  NAND2_X1 U6358 ( .A1(n8522), .A2(n8771), .ZN(n6762) );
  NAND2_X1 U6359 ( .A1(n8999), .A2(n6546), .ZN(n6557) );
  OR2_X1 U6360 ( .A1(n8844), .A2(n6992), .ZN(n7006) );
  AND2_X1 U6361 ( .A1(n8391), .A2(n8389), .ZN(n8492) );
  INV_X1 U6362 ( .A(n8793), .ZN(n8723) );
  NOR2_X1 U6363 ( .A1(n6468), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6484) );
  OR2_X1 U6364 ( .A1(n5740), .A2(n5739), .ZN(n6776) );
  INV_X1 U6365 ( .A(n7253), .ZN(n6243) );
  INV_X1 U6366 ( .A(n9468), .ZN(n9542) );
  OR2_X1 U6367 ( .A1(n9768), .A2(n6207), .ZN(n6160) );
  OR2_X1 U6368 ( .A1(n6037), .A2(n5624), .ZN(n6053) );
  INV_X1 U6369 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7961) );
  OR2_X1 U6370 ( .A1(n10090), .A2(n9587), .ZN(n10218) );
  INV_X1 U6371 ( .A(n9562), .ZN(n8053) );
  AND2_X1 U6372 ( .A1(n9325), .A2(n9327), .ZN(n9415) );
  OR2_X1 U6373 ( .A1(n7404), .A2(n9778), .ZN(n8103) );
  INV_X1 U6374 ( .A(n10512), .ZN(n10527) );
  INV_X1 U6375 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6238) );
  OR3_X1 U6376 ( .A1(n6704), .A2(n7920), .A3(n8018), .ZN(n6976) );
  INV_X1 U6377 ( .A(n8406), .ZN(n7877) );
  AND2_X1 U6378 ( .A1(n6994), .A2(n7008), .ZN(n7852) );
  INV_X1 U6379 ( .A(n8266), .ZN(n10665) );
  OR2_X1 U6380 ( .A1(n6376), .A2(n8662), .ZN(n8312) );
  AND4_X1 U6381 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n8712)
         );
  AND4_X1 U6382 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n10642)
         );
  NAND2_X1 U6383 ( .A1(n8300), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6380) );
  INV_X1 U6384 ( .A(n8619), .ZN(n6859) );
  INV_X1 U6385 ( .A(n8639), .ZN(n10413) );
  AND2_X1 U6386 ( .A1(P2_U3893), .A2(n6845), .ZN(n10412) );
  INV_X1 U6387 ( .A(n8496), .ZN(n8403) );
  INV_X1 U6388 ( .A(n8649), .ZN(n10568) );
  INV_X2 U6389 ( .A(n10572), .ZN(n10468) );
  AND2_X1 U6390 ( .A1(n7008), .A2(n7007), .ZN(n10572) );
  NAND2_X1 U6391 ( .A1(n6747), .A2(n6721), .ZN(n6998) );
  INV_X1 U6392 ( .A(n8067), .ZN(n8499) );
  INV_X1 U6393 ( .A(n8844), .ZN(n8871) );
  AND2_X1 U6394 ( .A1(n7592), .A2(n7591), .ZN(n10571) );
  NAND2_X1 U6395 ( .A1(n8661), .A2(n8814), .ZN(n8872) );
  AND2_X1 U6396 ( .A1(n6976), .A2(n6720), .ZN(n7008) );
  AND2_X1 U6397 ( .A1(n8286), .A2(P2_U3151), .ZN(n9148) );
  NAND2_X1 U6398 ( .A1(n6824), .A2(n6243), .ZN(n10448) );
  INV_X1 U6399 ( .A(n9264), .ZN(n9213) );
  INV_X1 U6400 ( .A(n9268), .ZN(n9235) );
  INV_X1 U6401 ( .A(n9551), .ZN(n9546) );
  AND2_X1 U6402 ( .A1(n6213), .A2(n6212), .ZN(n9750) );
  AND4_X1 U6403 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n9674)
         );
  NAND2_X1 U6404 ( .A1(n4916), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5712) );
  INV_X1 U6405 ( .A(n7085), .ZN(n10228) );
  INV_X1 U6406 ( .A(n10437), .ZN(n10229) );
  INV_X1 U6407 ( .A(n10448), .ZN(n10551) );
  INV_X1 U6408 ( .A(n8103), .ZN(n10556) );
  INV_X1 U6409 ( .A(n9896), .ZN(n9815) );
  AOI21_X1 U6410 ( .B1(n6233), .B2(n6827), .A(n6826), .ZN(n7320) );
  INV_X1 U6411 ( .A(n10628), .ZN(n10494) );
  INV_X1 U6412 ( .A(n9990), .ZN(n10609) );
  AND2_X1 U6413 ( .A1(n7252), .A2(n7251), .ZN(n7396) );
  INV_X1 U6414 ( .A(n4908), .ZN(n9588) );
  NOR2_X1 U6415 ( .A1(n8286), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10015) );
  NOR2_X1 U6416 ( .A1(n6976), .A2(n7750), .ZN(n6847) );
  INV_X1 U6417 ( .A(n8680), .ZN(n8211) );
  NAND2_X1 U6418 ( .A1(n6987), .A2(n6986), .ZN(n8266) );
  INV_X1 U6419 ( .A(n10667), .ZN(n8277) );
  AND4_X1 U6420 ( .A1(n8312), .A2(n6681), .A3(n6680), .A4(n6679), .ZN(n8317)
         );
  INV_X1 U6421 ( .A(n7554), .ZN(n8534) );
  INV_X1 U6422 ( .A(n10412), .ZN(n10282) );
  INV_X1 U6423 ( .A(n8314), .ZN(n8810) );
  NAND2_X1 U6424 ( .A1(n10575), .A2(n10474), .ZN(n8807) );
  NAND2_X2 U6425 ( .A1(n7010), .A2(n10468), .ZN(n10575) );
  INV_X1 U6426 ( .A(n10575), .ZN(n10577) );
  NAND2_X1 U6427 ( .A1(n8876), .A2(n8872), .ZN(n8865) );
  OR2_X1 U6428 ( .A1(n6998), .A2(n6726), .ZN(n7621) );
  OR2_X1 U6429 ( .A1(n8669), .A2(n9134), .ZN(n6760) );
  OR2_X1 U6430 ( .A1(n10637), .A2(n8839), .ZN(n9134) );
  AND2_X1 U6431 ( .A1(n6756), .A2(n6755), .ZN(n10637) );
  INV_X2 U6432 ( .A(n10637), .ZN(n10640) );
  NOR2_X1 U6433 ( .A1(n6807), .A2(n6702), .ZN(n6917) );
  INV_X1 U6434 ( .A(n6700), .ZN(n8018) );
  INV_X1 U6435 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6970) );
  AND2_X1 U6436 ( .A1(n6822), .A2(n7341), .ZN(n10439) );
  INV_X1 U6437 ( .A(n7948), .ZN(n10617) );
  AND2_X1 U6438 ( .A1(n6244), .A2(n10448), .ZN(n9243) );
  OR2_X1 U6439 ( .A1(n6250), .A2(n6240), .ZN(n9268) );
  INV_X1 U6440 ( .A(n9750), .ZN(n9726) );
  AND4_X1 U6441 ( .A1(n5668), .A2(n5667), .A3(n5666), .A4(n5665), .ZN(n9866)
         );
  INV_X1 U6442 ( .A(n7776), .ZN(n9565) );
  INV_X1 U6443 ( .A(n10439), .ZN(n10264) );
  NAND2_X1 U6444 ( .A1(n9868), .A2(n7406), .ZN(n9879) );
  AND2_X1 U6445 ( .A1(n7572), .A2(n7571), .ZN(n10517) );
  INV_X1 U6446 ( .A(n10632), .ZN(n10630) );
  AND2_X1 U6447 ( .A1(n10517), .A2(n10516), .ZN(n10520) );
  AND3_X2 U6448 ( .A1(n7398), .A2(n7321), .A3(n7396), .ZN(n10636) );
  AND2_X1 U6449 ( .A1(n6821), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6825) );
  INV_X1 U6450 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7614) );
  NAND2_X1 U6451 ( .A1(n8286), .A2(P1_U3086), .ZN(n10025) );
  AND2_X1 U6452 ( .A1(n6847), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3893) );
  AND2_X1 U6453 ( .A1(n6774), .A2(n6825), .ZN(P1_U3973) );
  NAND2_X1 U6454 ( .A1(n5492), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5493) );
  OAI21_X1 U6455 ( .B1(n5600), .B2(n5497), .A(n5496), .ZN(n5501) );
  XNOR2_X1 U6456 ( .A(n5501), .B(SI_1_), .ZN(n5692) );
  INV_X1 U6457 ( .A(n5692), .ZN(n5500) );
  INV_X2 U6458 ( .A(n5600), .ZN(n5506) );
  NAND3_X1 U6459 ( .A1(n6656), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n5499) );
  AND2_X1 U6460 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6461 ( .A1(n5600), .A2(n5498), .ZN(n6355) );
  NAND2_X1 U6462 ( .A1(n5501), .A2(SI_1_), .ZN(n5502) );
  MUX2_X1 U6463 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5506), .Z(n5503) );
  INV_X1 U6464 ( .A(SI_2_), .ZN(n9055) );
  XNOR2_X1 U6465 ( .A(n5503), .B(n9055), .ZN(n5701) );
  NAND2_X1 U6466 ( .A1(n5503), .A2(SI_2_), .ZN(n5504) );
  NAND2_X1 U6467 ( .A1(n5505), .A2(n5504), .ZN(n5722) );
  MUX2_X1 U6468 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n8141), .Z(n5508) );
  INV_X1 U6469 ( .A(SI_3_), .ZN(n5507) );
  XNOR2_X1 U6470 ( .A(n5508), .B(n5507), .ZN(n5721) );
  NAND2_X1 U6471 ( .A1(n5722), .A2(n5721), .ZN(n5510) );
  NAND2_X1 U6472 ( .A1(n5508), .A2(SI_3_), .ZN(n5509) );
  NAND2_X1 U6473 ( .A1(n5510), .A2(n5509), .ZN(n5742) );
  INV_X1 U6474 ( .A(SI_4_), .ZN(n5511) );
  XNOR2_X1 U6475 ( .A(n5512), .B(n5511), .ZN(n5741) );
  NAND2_X1 U6476 ( .A1(n5512), .A2(SI_4_), .ZN(n5513) );
  MUX2_X1 U6477 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8141), .Z(n5515) );
  INV_X1 U6478 ( .A(n5757), .ZN(n5514) );
  NAND2_X1 U6479 ( .A1(n5515), .A2(SI_5_), .ZN(n5516) );
  MUX2_X1 U6480 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8141), .Z(n5518) );
  XNOR2_X1 U6481 ( .A(n5518), .B(SI_6_), .ZN(n5776) );
  INV_X1 U6482 ( .A(n5776), .ZN(n5517) );
  NAND2_X1 U6483 ( .A1(n5777), .A2(n5517), .ZN(n5520) );
  NAND2_X1 U6484 ( .A1(n5518), .A2(SI_6_), .ZN(n5519) );
  NAND2_X1 U6485 ( .A1(n5520), .A2(n5519), .ZN(n5799) );
  MUX2_X1 U6486 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6656), .Z(n5522) );
  XNOR2_X1 U6487 ( .A(n5522), .B(SI_7_), .ZN(n5798) );
  INV_X1 U6488 ( .A(n5798), .ZN(n5521) );
  NAND2_X1 U6489 ( .A1(n5522), .A2(SI_7_), .ZN(n5523) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6816) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6814) );
  MUX2_X1 U6492 ( .A(n6816), .B(n6814), .S(n6656), .Z(n5524) );
  INV_X1 U6493 ( .A(SI_8_), .ZN(n8907) );
  NAND2_X1 U6494 ( .A1(n5524), .A2(n8907), .ZN(n5527) );
  INV_X1 U6495 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U6496 ( .A1(n5525), .A2(SI_8_), .ZN(n5526) );
  NAND2_X1 U6497 ( .A1(n5527), .A2(n5526), .ZN(n5826) );
  INV_X1 U6498 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6831) );
  INV_X1 U6499 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6829) );
  MUX2_X1 U6500 ( .A(n6831), .B(n6829), .S(n6656), .Z(n5529) );
  INV_X1 U6501 ( .A(SI_9_), .ZN(n5528) );
  NAND2_X1 U6502 ( .A1(n5529), .A2(n5528), .ZN(n5532) );
  INV_X1 U6503 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U6504 ( .A1(n5530), .A2(SI_9_), .ZN(n5531) );
  MUX2_X1 U6505 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6656), .Z(n5534) );
  XNOR2_X1 U6506 ( .A(n5534), .B(n8940), .ZN(n5865) );
  INV_X1 U6507 ( .A(n5865), .ZN(n5536) );
  NAND2_X1 U6508 ( .A1(n5534), .A2(SI_10_), .ZN(n5535) );
  INV_X1 U6509 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5537) );
  MUX2_X1 U6510 ( .A(n6970), .B(n5537), .S(n8141), .Z(n5538) );
  NAND2_X1 U6511 ( .A1(n5538), .A2(n9035), .ZN(n5541) );
  INV_X1 U6512 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U6513 ( .A1(n5539), .A2(SI_11_), .ZN(n5540) );
  NAND2_X1 U6514 ( .A1(n5541), .A2(n5540), .ZN(n5882) );
  MUX2_X1 U6515 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8141), .Z(n5542) );
  XNOR2_X1 U6516 ( .A(n5542), .B(n9037), .ZN(n5900) );
  INV_X1 U6517 ( .A(n5900), .ZN(n5544) );
  NAND2_X1 U6518 ( .A1(n5542), .A2(SI_12_), .ZN(n5543) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8141), .Z(n5546) );
  XNOR2_X1 U6520 ( .A(n5546), .B(SI_13_), .ZN(n5929) );
  INV_X1 U6521 ( .A(n5929), .ZN(n5545) );
  NAND2_X1 U6522 ( .A1(n5546), .A2(SI_13_), .ZN(n5547) );
  MUX2_X1 U6523 ( .A(n7125), .B(n7127), .S(n6656), .Z(n5548) );
  NAND2_X1 U6524 ( .A1(n5548), .A2(n9034), .ZN(n5551) );
  INV_X1 U6525 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U6526 ( .A1(n5549), .A2(SI_14_), .ZN(n5550) );
  NAND2_X1 U6527 ( .A1(n5551), .A2(n5550), .ZN(n5952) );
  MUX2_X1 U6528 ( .A(n7194), .B(n7192), .S(n8141), .Z(n5552) );
  XNOR2_X1 U6529 ( .A(n5552), .B(SI_15_), .ZN(n5970) );
  INV_X1 U6530 ( .A(n5970), .ZN(n5555) );
  INV_X1 U6531 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U6532 ( .A1(n5553), .A2(SI_15_), .ZN(n5554) );
  MUX2_X1 U6533 ( .A(n7319), .B(n7317), .S(n6656), .Z(n5556) );
  NAND2_X1 U6534 ( .A1(n5556), .A2(n9030), .ZN(n5559) );
  INV_X1 U6535 ( .A(n5556), .ZN(n5557) );
  NAND2_X1 U6536 ( .A1(n5557), .A2(SI_16_), .ZN(n5558) );
  NAND2_X1 U6537 ( .A1(n5559), .A2(n5558), .ZN(n5989) );
  OAI21_X2 U6538 ( .B1(n5990), .B2(n5989), .A(n5559), .ZN(n6008) );
  INV_X1 U6539 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5560) );
  MUX2_X1 U6540 ( .A(n7392), .B(n5560), .S(n8141), .Z(n5561) );
  NAND2_X1 U6541 ( .A1(n5561), .A2(n8930), .ZN(n5564) );
  INV_X1 U6542 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U6543 ( .A1(n5562), .A2(SI_17_), .ZN(n5563) );
  NAND2_X1 U6544 ( .A1(n6008), .A2(n6007), .ZN(n5565) );
  MUX2_X1 U6545 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6656), .Z(n5567) );
  XNOR2_X1 U6546 ( .A(n5567), .B(n5566), .ZN(n5658) );
  INV_X1 U6547 ( .A(n5658), .ZN(n5569) );
  NAND2_X1 U6548 ( .A1(n5567), .A2(SI_18_), .ZN(n5568) );
  MUX2_X1 U6549 ( .A(n7612), .B(n7614), .S(n8141), .Z(n5570) );
  INV_X1 U6550 ( .A(SI_19_), .ZN(n9025) );
  NAND2_X1 U6551 ( .A1(n5570), .A2(n9025), .ZN(n5573) );
  INV_X1 U6552 ( .A(n5570), .ZN(n5571) );
  NAND2_X1 U6553 ( .A1(n5571), .A2(SI_19_), .ZN(n5572) );
  NAND2_X1 U6554 ( .A1(n5573), .A2(n5572), .ZN(n6028) );
  MUX2_X1 U6555 ( .A(n7692), .B(n7650), .S(n8141), .Z(n5574) );
  NAND2_X1 U6556 ( .A1(n5574), .A2(n9020), .ZN(n5577) );
  INV_X1 U6557 ( .A(n5574), .ZN(n5575) );
  NAND2_X1 U6558 ( .A1(n5575), .A2(SI_20_), .ZN(n5576) );
  NAND2_X1 U6559 ( .A1(n6050), .A2(n6049), .ZN(n5578) );
  MUX2_X1 U6560 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6656), .Z(n6067) );
  INV_X1 U6561 ( .A(SI_21_), .ZN(n5579) );
  XNOR2_X1 U6562 ( .A(n6067), .B(n5579), .ZN(n6087) );
  NOR2_X1 U6563 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5580) );
  NAND2_X1 U6564 ( .A1(n5704), .A2(n5580), .ZN(n5743) );
  NOR2_X1 U6565 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5585) );
  NOR2_X1 U6566 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5584) );
  NOR2_X1 U6567 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5583) );
  NOR2_X1 U6568 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5582) );
  INV_X1 U6569 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5588) );
  NAND3_X1 U6570 ( .A1(n5649), .A2(n5591), .A3(n5645), .ZN(n5592) );
  INV_X1 U6571 ( .A(n5629), .ZN(n5593) );
  NAND2_X1 U6572 ( .A1(n5593), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U6573 ( .A1(n5597), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6574 ( .A1(n7732), .A2(n9273), .ZN(n5602) );
  INV_X1 U6575 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7733) );
  OR2_X1 U6576 ( .A1(n5778), .A2(n7733), .ZN(n5601) );
  INV_X1 U6577 ( .A(n9950), .ZN(n9839) );
  OR2_X1 U6578 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  NOR2_X1 U6579 ( .A1(n7896), .A2(n7863), .ZN(n5610) );
  NAND2_X1 U6580 ( .A1(n5652), .A2(n5614), .ZN(n5612) );
  XNOR2_X2 U6581 ( .A(n5613), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6236) );
  INV_X1 U6582 ( .A(n5654), .ZN(n5615) );
  NAND2_X1 U6583 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5767) );
  INV_X1 U6584 ( .A(n5767), .ZN(n5616) );
  NAND2_X1 U6585 ( .A1(n5616), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5784) );
  INV_X1 U6586 ( .A(n5784), .ZN(n5617) );
  NAND2_X1 U6587 ( .A1(n5617), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5807) );
  INV_X1 U6588 ( .A(n5807), .ZN(n5618) );
  NAND2_X1 U6589 ( .A1(n5618), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5831) );
  INV_X1 U6590 ( .A(n5851), .ZN(n5619) );
  NAND2_X1 U6591 ( .A1(n5619), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5871) );
  INV_X1 U6592 ( .A(n5890), .ZN(n5620) );
  NAND2_X1 U6593 ( .A1(n5620), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5914) );
  INV_X1 U6594 ( .A(n5961), .ZN(n5621) );
  NAND2_X1 U6595 ( .A1(n5621), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5976) );
  INV_X1 U6596 ( .A(n5976), .ZN(n5622) );
  NAND2_X1 U6597 ( .A1(n5622), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U6598 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5624) );
  INV_X1 U6599 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U6600 ( .A1(n6055), .A2(n5626), .ZN(n5627) );
  AND2_X1 U6601 ( .A1(n6073), .A2(n5627), .ZN(n9836) );
  NOR2_X1 U6602 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5628) );
  NAND2_X1 U6603 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  INV_X1 U6604 ( .A(n5634), .ZN(n5631) );
  NAND2_X1 U6605 ( .A1(n9836), .A2(n9184), .ZN(n5642) );
  AOI22_X1 U6606 ( .A1(n4916), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5786), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U6607 ( .A1(n4918), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U6608 ( .A1(n5643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5991) );
  OAI21_X1 U6609 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U6610 ( .A1(n5991), .A2(n5644), .ZN(n5660) );
  INV_X1 U6611 ( .A(n5660), .ZN(n5646) );
  NAND2_X1 U6612 ( .A1(n5646), .A2(n5645), .ZN(n5662) );
  XNOR2_X2 U6613 ( .A(n5648), .B(n5647), .ZN(n6030) );
  INV_X1 U6614 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U6615 ( .A1(n5650), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5651) );
  OR2_X1 U6616 ( .A1(n5654), .A2(n6030), .ZN(n7472) );
  OAI22_X1 U6617 ( .A1(n9839), .A2(n9170), .B1(n9808), .B2(n9176), .ZN(n6064)
         );
  INV_X1 U6618 ( .A(n6064), .ZN(n6066) );
  NAND2_X1 U6619 ( .A1(n9550), .A2(n6030), .ZN(n7238) );
  AND2_X1 U6620 ( .A1(n7238), .A2(n5654), .ZN(n5655) );
  NAND2_X1 U6621 ( .A1(n5680), .A2(n5655), .ZN(n5656) );
  AOI22_X1 U6622 ( .A1(n9950), .A2(n9169), .B1(n6214), .B2(n9851), .ZN(n5657)
         );
  CLKBUF_X3 U6623 ( .A(n5656), .Z(n6216) );
  XNOR2_X1 U6624 ( .A(n5657), .B(n6216), .ZN(n6065) );
  XNOR2_X1 U6625 ( .A(n5659), .B(n5658), .ZN(n7388) );
  NAND2_X1 U6626 ( .A1(n7388), .A2(n9273), .ZN(n5664) );
  NAND2_X1 U6627 ( .A1(n5660), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5661) );
  AOI22_X1 U6628 ( .A1(n6032), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6031), .B2(
        n10214), .ZN(n5663) );
  XNOR2_X1 U6629 ( .A(n6037), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U6630 ( .A1(n9877), .A2(n9184), .ZN(n5668) );
  NAND2_X1 U6631 ( .A1(n4916), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U6632 ( .A1(n5786), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U6633 ( .A1(n4918), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5665) );
  NOR2_X1 U6634 ( .A1(n9866), .A2(n9176), .ZN(n5669) );
  AOI21_X1 U6635 ( .B1(n9964), .B2(n6214), .A(n5669), .ZN(n9259) );
  NAND2_X1 U6636 ( .A1(n4916), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6637 ( .A1(n4918), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6638 ( .A1(n5786), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U6639 ( .A1(n9574), .A2(n4909), .ZN(n5679) );
  INV_X1 U6640 ( .A(SI_0_), .ZN(n5675) );
  NOR2_X1 U6641 ( .A1(n8286), .A2(n5675), .ZN(n5677) );
  INV_X1 U6642 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U6643 ( .A(n5677), .B(n5676), .ZN(n10026) );
  MUX2_X1 U6644 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10026), .S(n6820), .Z(n9404)
         );
  NAND2_X1 U6645 ( .A1(n9404), .A2(n5708), .ZN(n5678) );
  INV_X1 U6646 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5681) );
  OR2_X1 U6647 ( .A1(n5680), .A2(n5681), .ZN(n5682) );
  NAND2_X1 U6648 ( .A1(n5687), .A2(n5682), .ZN(n7080) );
  INV_X1 U6649 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U6650 ( .A1(n9404), .A2(n4909), .ZN(n5685) );
  NAND2_X1 U6651 ( .A1(n9574), .A2(n6185), .ZN(n5684) );
  OAI211_X1 U6652 ( .C1(n5680), .C2(n5686), .A(n5685), .B(n5684), .ZN(n7079)
         );
  NAND2_X1 U6653 ( .A1(n7080), .A2(n7079), .ZN(n7078) );
  INV_X2 U6654 ( .A(n6216), .ZN(n9173) );
  NAND2_X1 U6655 ( .A1(n5687), .A2(n9173), .ZN(n5688) );
  INV_X1 U6656 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U6657 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5689) );
  XNOR2_X1 U6658 ( .A(n5690), .B(n5689), .ZN(n7344) );
  XNOR2_X1 U6659 ( .A(n5692), .B(n5691), .ZN(n6362) );
  INV_X1 U6660 ( .A(n6362), .ZN(n6792) );
  NAND2_X1 U6661 ( .A1(n7234), .A2(n5708), .ZN(n5693) );
  OAI21_X1 U6662 ( .B1(n10446), .B2(n9170), .A(n5693), .ZN(n5694) );
  XNOR2_X1 U6663 ( .A(n5694), .B(n6216), .ZN(n5698) );
  NAND2_X1 U6664 ( .A1(n5697), .A2(n5698), .ZN(n7258) );
  OR2_X1 U6665 ( .A1(n10446), .A2(n9176), .ZN(n5696) );
  NAND2_X1 U6666 ( .A1(n7234), .A2(n4909), .ZN(n5695) );
  AND2_X1 U6667 ( .A1(n5696), .A2(n5695), .ZN(n7257) );
  NAND2_X1 U6668 ( .A1(n7256), .A2(n7260), .ZN(n7266) );
  INV_X1 U6669 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6794) );
  OR2_X1 U6670 ( .A1(n5778), .A2(n6794), .ZN(n5707) );
  XNOR2_X1 U6671 ( .A(n5702), .B(n5701), .ZN(n6793) );
  OR2_X1 U6672 ( .A1(n5703), .A2(n6793), .ZN(n5706) );
  OR2_X1 U6673 ( .A1(n5704), .A2(n5307), .ZN(n5724) );
  INV_X1 U6674 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5723) );
  XNOR2_X1 U6675 ( .A(n5724), .B(n5723), .ZN(n9596) );
  OR2_X1 U6676 ( .A1(n6820), .A2(n9596), .ZN(n5705) );
  NAND2_X1 U6678 ( .A1(n9184), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6679 ( .A1(n4918), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U6680 ( .A1(n5786), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6681 ( .A1(n9573), .A2(n4909), .ZN(n5713) );
  OAI21_X1 U6682 ( .B1(n9279), .B2(n6183), .A(n5713), .ZN(n5714) );
  XNOR2_X1 U6683 ( .A(n5714), .B(n9173), .ZN(n5716) );
  NAND2_X1 U6684 ( .A1(n9573), .A2(n6185), .ZN(n5715) );
  OAI21_X1 U6685 ( .B1(n9279), .B2(n9170), .A(n5715), .ZN(n5717) );
  XNOR2_X1 U6686 ( .A(n5716), .B(n5717), .ZN(n7265) );
  NAND2_X1 U6687 ( .A1(n7266), .A2(n7265), .ZN(n5720) );
  INV_X1 U6688 ( .A(n5716), .ZN(n5718) );
  OR2_X1 U6689 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  INV_X1 U6690 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6800) );
  OR2_X1 U6691 ( .A1(n5778), .A2(n6800), .ZN(n5730) );
  XNOR2_X1 U6692 ( .A(n5721), .B(n5722), .ZN(n6799) );
  OR2_X1 U6693 ( .A1(n5703), .A2(n6799), .ZN(n5729) );
  NAND2_X1 U6694 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  NAND2_X1 U6695 ( .A1(n5725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5727) );
  INV_X1 U6696 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5726) );
  XNOR2_X1 U6697 ( .A(n5727), .B(n5726), .ZN(n7348) );
  OR2_X1 U6698 ( .A1(n6820), .A2(n7348), .ZN(n5728) );
  NAND2_X1 U6699 ( .A1(n4916), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5734) );
  INV_X1 U6700 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7538) );
  NAND2_X1 U6701 ( .A1(n9184), .A2(n7538), .ZN(n5733) );
  NAND2_X1 U6702 ( .A1(n5786), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U6703 ( .A1(n4918), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6704 ( .A1(n9572), .A2(n4909), .ZN(n5735) );
  OAI21_X1 U6705 ( .B1(n10478), .B2(n6183), .A(n5735), .ZN(n5736) );
  XNOR2_X1 U6706 ( .A(n5736), .B(n9173), .ZN(n5738) );
  NAND2_X1 U6707 ( .A1(n9572), .A2(n6185), .ZN(n5737) );
  OAI21_X1 U6708 ( .B1(n10478), .B2(n9170), .A(n5737), .ZN(n5739) );
  XNOR2_X1 U6709 ( .A(n5738), .B(n5739), .ZN(n7534) );
  INV_X1 U6710 ( .A(n5738), .ZN(n5740) );
  XNOR2_X1 U6711 ( .A(n5742), .B(n5741), .ZN(n6795) );
  OR2_X1 U6712 ( .A1(n5703), .A2(n6795), .ZN(n5747) );
  INV_X1 U6713 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U6714 ( .A1(n5743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5744) );
  XNOR2_X1 U6715 ( .A(n5744), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7350) );
  INV_X1 U6716 ( .A(n7350), .ZN(n10436) );
  OR2_X1 U6717 ( .A1(n6820), .A2(n10436), .ZN(n5745) );
  NAND2_X1 U6718 ( .A1(n5786), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U6719 ( .A1(n4916), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5751) );
  OAI21_X1 U6720 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n5767), .ZN(n7407) );
  INV_X1 U6721 ( .A(n7407), .ZN(n5748) );
  NAND2_X1 U6722 ( .A1(n9184), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U6723 ( .A1(n4918), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5749) );
  OAI22_X1 U6724 ( .A1(n7430), .A2(n6183), .B1(n7665), .B2(n9170), .ZN(n5753)
         );
  XNOR2_X1 U6725 ( .A(n5753), .B(n6216), .ZN(n5756) );
  OR2_X1 U6726 ( .A1(n7665), .A2(n9176), .ZN(n5754) );
  OAI21_X1 U6727 ( .B1(n7430), .B2(n9170), .A(n5754), .ZN(n5755) );
  XNOR2_X1 U6728 ( .A(n5756), .B(n5755), .ZN(n6780) );
  NAND2_X1 U6729 ( .A1(n5756), .A2(n5755), .ZN(n5794) );
  INV_X1 U6730 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6798) );
  OR2_X1 U6731 ( .A1(n5778), .A2(n6798), .ZN(n5765) );
  XNOR2_X1 U6732 ( .A(n5758), .B(n5757), .ZN(n6423) );
  INV_X1 U6733 ( .A(n6423), .ZN(n6797) );
  OR2_X1 U6734 ( .A1(n5703), .A2(n6797), .ZN(n5764) );
  NAND2_X1 U6735 ( .A1(n5759), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5760) );
  MUX2_X1 U6736 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5760), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5762) );
  NOR2_X1 U6737 ( .A1(n5759), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5801) );
  INV_X1 U6738 ( .A(n5801), .ZN(n5761) );
  INV_X1 U6739 ( .A(n7353), .ZN(n10101) );
  OR2_X1 U6740 ( .A1(n6820), .A2(n10101), .ZN(n5763) );
  NAND2_X1 U6741 ( .A1(n4916), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5772) );
  INV_X1 U6742 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U6743 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  AND2_X1 U6744 ( .A1(n5784), .A2(n5768), .ZN(n7545) );
  NAND2_X1 U6745 ( .A1(n9184), .A2(n7545), .ZN(n5771) );
  NAND2_X1 U6746 ( .A1(n5786), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U6747 ( .A1(n4918), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5769) );
  NAND4_X1 U6748 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n9570)
         );
  NAND2_X1 U6749 ( .A1(n9570), .A2(n4909), .ZN(n5773) );
  OAI21_X1 U6750 ( .B1(n10503), .B2(n6183), .A(n5773), .ZN(n5774) );
  XNOR2_X1 U6751 ( .A(n5774), .B(n9173), .ZN(n5795) );
  NAND2_X1 U6752 ( .A1(n9570), .A2(n6185), .ZN(n5775) );
  OAI21_X1 U6753 ( .B1(n10503), .B2(n9170), .A(n5775), .ZN(n7544) );
  XNOR2_X1 U6754 ( .A(n5777), .B(n5776), .ZN(n6434) );
  INV_X1 U6755 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6802) );
  OR2_X1 U6756 ( .A1(n5778), .A2(n6802), .ZN(n5781) );
  OR2_X1 U6757 ( .A1(n5801), .A2(n5307), .ZN(n5779) );
  XNOR2_X1 U6758 ( .A(n5779), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7356) );
  INV_X1 U6759 ( .A(n7356), .ZN(n10116) );
  OR2_X1 U6760 ( .A1(n6820), .A2(n10116), .ZN(n5780) );
  NAND2_X1 U6761 ( .A1(n4916), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5790) );
  INV_X1 U6762 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6763 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  AND2_X1 U6764 ( .A1(n5807), .A2(n5785), .ZN(n7575) );
  NAND2_X1 U6765 ( .A1(n9184), .A2(n7575), .ZN(n5789) );
  NAND2_X1 U6766 ( .A1(n4918), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U6767 ( .A1(n5786), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U6768 ( .A1(n9569), .A2(n4909), .ZN(n5791) );
  XNOR2_X1 U6769 ( .A(n5792), .B(n6216), .ZN(n5819) );
  NAND2_X1 U6770 ( .A1(n9569), .A2(n6185), .ZN(n5793) );
  OAI21_X1 U6771 ( .B1(n10511), .B2(n9170), .A(n5793), .ZN(n5818) );
  INV_X1 U6772 ( .A(n5795), .ZN(n7523) );
  OR2_X1 U6773 ( .A1(n7528), .A2(n7523), .ZN(n5796) );
  NAND2_X1 U6774 ( .A1(n5797), .A2(n5796), .ZN(n7525) );
  XNOR2_X1 U6775 ( .A(n5799), .B(n5798), .ZN(n6803) );
  NAND2_X1 U6776 ( .A1(n9273), .A2(n6803), .ZN(n5805) );
  INV_X1 U6777 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U6778 ( .A1(n5801), .A2(n5800), .ZN(n5824) );
  NAND2_X1 U6779 ( .A1(n5824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U6780 ( .A(n5802), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7359) );
  INV_X1 U6781 ( .A(n7359), .ZN(n10131) );
  OR2_X1 U6782 ( .A1(n6820), .A2(n10131), .ZN(n5804) );
  INV_X1 U6783 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6804) );
  OR2_X1 U6784 ( .A1(n5778), .A2(n6804), .ZN(n5803) );
  NAND2_X1 U6785 ( .A1(n4916), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5812) );
  INV_X1 U6786 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U6787 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  AND2_X1 U6788 ( .A1(n5831), .A2(n5808), .ZN(n10550) );
  NAND2_X1 U6789 ( .A1(n9184), .A2(n10550), .ZN(n5811) );
  NAND2_X1 U6790 ( .A1(n4918), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6791 ( .A1(n5786), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U6792 ( .A1(n9568), .A2(n4909), .ZN(n5813) );
  OAI21_X1 U6793 ( .B1(n10530), .B2(n6183), .A(n5813), .ZN(n5814) );
  XNOR2_X1 U6794 ( .A(n5814), .B(n9173), .ZN(n5823) );
  OR2_X1 U6795 ( .A1(n10530), .A2(n9170), .ZN(n5816) );
  NAND2_X1 U6796 ( .A1(n9568), .A2(n6185), .ZN(n5815) );
  NAND2_X1 U6797 ( .A1(n5816), .A2(n5815), .ZN(n5821) );
  XNOR2_X1 U6798 ( .A(n5823), .B(n5821), .ZN(n7605) );
  AND2_X1 U6799 ( .A1(n7525), .A2(n7605), .ZN(n5817) );
  INV_X1 U6800 ( .A(n7605), .ZN(n5820) );
  OR2_X1 U6801 ( .A1(n5819), .A2(n5818), .ZN(n7602) );
  INV_X1 U6802 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U6803 ( .A1(n5847), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U6804 ( .A(n5825), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7361) );
  AOI22_X1 U6805 ( .A1(n6032), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6031), .B2(
        n7361), .ZN(n5829) );
  XNOR2_X1 U6806 ( .A(n5827), .B(n5826), .ZN(n6813) );
  NAND2_X1 U6807 ( .A1(n6813), .A2(n9273), .ZN(n5828) );
  NAND2_X1 U6808 ( .A1(n5829), .A2(n5828), .ZN(n7746) );
  NAND2_X1 U6809 ( .A1(n7746), .A2(n9169), .ZN(n5838) );
  NAND2_X1 U6810 ( .A1(n4916), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U6811 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  AND2_X1 U6812 ( .A1(n5851), .A2(n5832), .ZN(n7712) );
  NAND2_X1 U6813 ( .A1(n9184), .A2(n7712), .ZN(n5835) );
  NAND2_X1 U6814 ( .A1(n5786), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U6815 ( .A1(n4918), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5833) );
  OR2_X1 U6816 ( .A1(n10532), .A2(n9170), .ZN(n5837) );
  NAND2_X1 U6817 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  XNOR2_X1 U6818 ( .A(n5839), .B(n9173), .ZN(n5843) );
  NAND2_X1 U6819 ( .A1(n7746), .A2(n6214), .ZN(n5841) );
  OR2_X1 U6820 ( .A1(n10532), .A2(n9176), .ZN(n5840) );
  NAND2_X1 U6821 ( .A1(n5841), .A2(n5840), .ZN(n7705) );
  NAND2_X1 U6822 ( .A1(n7706), .A2(n7705), .ZN(n7710) );
  INV_X1 U6823 ( .A(n5842), .ZN(n5845) );
  INV_X1 U6824 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U6825 ( .A1(n5845), .A2(n5844), .ZN(n7707) );
  NAND2_X1 U6826 ( .A1(n7710), .A2(n7707), .ZN(n7651) );
  XNOR2_X1 U6827 ( .A(n5846), .B(n5488), .ZN(n6828) );
  NAND2_X1 U6828 ( .A1(n6828), .A2(n9273), .ZN(n5849) );
  NAND2_X1 U6829 ( .A1(n5906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5867) );
  XNOR2_X1 U6830 ( .A(n5867), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7362) );
  AOI22_X1 U6831 ( .A1(n6032), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6031), .B2(
        n7362), .ZN(n5848) );
  NAND2_X1 U6832 ( .A1(n5849), .A2(n5848), .ZN(n7775) );
  NAND2_X1 U6833 ( .A1(n7775), .A2(n9169), .ZN(n5858) );
  NAND2_X1 U6834 ( .A1(n4916), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5856) );
  INV_X1 U6835 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U6836 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  AND2_X1 U6837 ( .A1(n5871), .A2(n5852), .ZN(n7740) );
  NAND2_X1 U6838 ( .A1(n9184), .A2(n7740), .ZN(n5855) );
  NAND2_X1 U6839 ( .A1(n5786), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6840 ( .A1(n4918), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5853) );
  OR2_X1 U6841 ( .A1(n7734), .A2(n9170), .ZN(n5857) );
  NAND2_X1 U6842 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  XNOR2_X1 U6843 ( .A(n5859), .B(n9173), .ZN(n7653) );
  NOR2_X1 U6844 ( .A1(n7734), .A2(n9176), .ZN(n5860) );
  AOI21_X1 U6845 ( .B1(n7775), .B2(n6214), .A(n5860), .ZN(n5862) );
  NAND2_X1 U6846 ( .A1(n7653), .A2(n5862), .ZN(n5861) );
  INV_X1 U6847 ( .A(n7653), .ZN(n5863) );
  INV_X1 U6848 ( .A(n5862), .ZN(n7652) );
  NAND2_X1 U6849 ( .A1(n5863), .A2(n7652), .ZN(n5864) );
  XNOR2_X1 U6850 ( .A(n5866), .B(n5865), .ZN(n6833) );
  INV_X1 U6851 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U6852 ( .A1(n5867), .A2(n5904), .ZN(n5868) );
  NAND2_X1 U6853 ( .A1(n5868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5884) );
  XNOR2_X1 U6854 ( .A(n5884), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7363) );
  AOI22_X1 U6855 ( .A1(n6032), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6031), .B2(
        n7363), .ZN(n5869) );
  NAND2_X1 U6856 ( .A1(n7803), .A2(n6214), .ZN(n5878) );
  NAND2_X1 U6857 ( .A1(n4916), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U6858 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  AND2_X1 U6859 ( .A1(n5890), .A2(n5872), .ZN(n7784) );
  NAND2_X1 U6860 ( .A1(n9184), .A2(n7784), .ZN(n5875) );
  NAND2_X1 U6861 ( .A1(n5786), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U6862 ( .A1(n4918), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5873) );
  OR2_X1 U6863 ( .A1(n7776), .A2(n9176), .ZN(n5877) );
  NAND2_X1 U6864 ( .A1(n5878), .A2(n5877), .ZN(n7765) );
  NAND2_X1 U6865 ( .A1(n7803), .A2(n9169), .ZN(n5880) );
  OR2_X1 U6866 ( .A1(n7776), .A2(n9170), .ZN(n5879) );
  NAND2_X1 U6867 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XNOR2_X1 U6868 ( .A(n5881), .B(n6216), .ZN(n7764) );
  XNOR2_X1 U6869 ( .A(n5883), .B(n5882), .ZN(n6915) );
  NAND2_X1 U6870 ( .A1(n6915), .A2(n9273), .ZN(n5888) );
  INV_X1 U6871 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U6872 ( .A1(n5884), .A2(n5903), .ZN(n5885) );
  NAND2_X1 U6873 ( .A1(n5885), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5886) );
  XNOR2_X1 U6874 ( .A(n5886), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U6875 ( .A1(n6032), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6031), .B2(
        n10151), .ZN(n5887) );
  NAND2_X1 U6876 ( .A1(n5888), .A2(n5887), .ZN(n7981) );
  NAND2_X1 U6877 ( .A1(n7981), .A2(n9169), .ZN(n5897) );
  NAND2_X1 U6878 ( .A1(n4916), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5895) );
  INV_X1 U6879 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U6880 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  AND2_X1 U6881 ( .A1(n5914), .A2(n5891), .ZN(n7972) );
  NAND2_X1 U6882 ( .A1(n9184), .A2(n7972), .ZN(n5894) );
  NAND2_X1 U6883 ( .A1(n4918), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U6884 ( .A1(n5786), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5892) );
  NAND4_X1 U6885 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(n9564)
         );
  NAND2_X1 U6886 ( .A1(n9564), .A2(n6214), .ZN(n5896) );
  NAND2_X1 U6887 ( .A1(n5897), .A2(n5896), .ZN(n5898) );
  XNOR2_X1 U6888 ( .A(n5898), .B(n9173), .ZN(n5924) );
  AND2_X1 U6889 ( .A1(n9564), .A2(n6185), .ZN(n5899) );
  AOI21_X1 U6890 ( .B1(n7981), .B2(n6214), .A(n5899), .ZN(n5925) );
  NAND2_X1 U6891 ( .A1(n5924), .A2(n5925), .ZN(n7976) );
  NAND2_X1 U6892 ( .A1(n7975), .A2(n7976), .ZN(n7909) );
  XNOR2_X1 U6893 ( .A(n5901), .B(n5900), .ZN(n7064) );
  NAND2_X1 U6894 ( .A1(n7064), .A2(n9273), .ZN(n5912) );
  INV_X1 U6895 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5902) );
  NAND3_X1 U6896 ( .A1(n5904), .A2(n5903), .A3(n5902), .ZN(n5905) );
  OAI21_X1 U6897 ( .B1(n5906), .B2(n5905), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5907) );
  MUX2_X1 U6898 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5907), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5910) );
  INV_X1 U6899 ( .A(n5908), .ZN(n5909) );
  AOI22_X1 U6900 ( .A1(n6032), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6031), .B2(
        n9634), .ZN(n5911) );
  NAND2_X1 U6901 ( .A1(n5912), .A2(n5911), .ZN(n7948) );
  NAND2_X1 U6902 ( .A1(n7948), .A2(n9169), .ZN(n5921) );
  NAND2_X1 U6903 ( .A1(n4916), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U6904 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  AND2_X1 U6905 ( .A1(n5936), .A2(n5915), .ZN(n7887) );
  NAND2_X1 U6906 ( .A1(n9184), .A2(n7887), .ZN(n5918) );
  NAND2_X1 U6907 ( .A1(n4918), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U6908 ( .A1(n5786), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5916) );
  NAND4_X1 U6909 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n9563)
         );
  NAND2_X1 U6910 ( .A1(n9563), .A2(n6214), .ZN(n5920) );
  NAND2_X1 U6911 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  XNOR2_X1 U6912 ( .A(n5922), .B(n6216), .ZN(n5948) );
  AND2_X1 U6913 ( .A1(n9563), .A2(n6185), .ZN(n5923) );
  AOI21_X1 U6914 ( .B1(n7948), .B2(n6214), .A(n5923), .ZN(n5946) );
  XNOR2_X1 U6915 ( .A(n5948), .B(n5946), .ZN(n7910) );
  INV_X1 U6916 ( .A(n5924), .ZN(n5927) );
  INV_X1 U6917 ( .A(n5925), .ZN(n5926) );
  NAND2_X1 U6918 ( .A1(n5927), .A2(n5926), .ZN(n7978) );
  AND2_X1 U6919 ( .A1(n7910), .A2(n7978), .ZN(n5928) );
  XNOR2_X1 U6920 ( .A(n5930), .B(n5929), .ZN(n7084) );
  NAND2_X1 U6921 ( .A1(n7084), .A2(n9273), .ZN(n5935) );
  NOR2_X1 U6922 ( .A1(n5908), .A2(n5307), .ZN(n5931) );
  MUX2_X1 U6923 ( .A(n5307), .B(n5931), .S(P1_IR_REG_13__SCAN_IN), .Z(n5933)
         );
  OR2_X1 U6924 ( .A1(n5933), .A2(n5932), .ZN(n7085) );
  AOI22_X1 U6925 ( .A1(n6032), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6031), .B2(
        n10228), .ZN(n5934) );
  NAND2_X1 U6926 ( .A1(n8002), .A2(n9169), .ZN(n5943) );
  NAND2_X1 U6927 ( .A1(n4916), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U6928 ( .A1(n5936), .A2(n7961), .ZN(n5937) );
  AND2_X1 U6929 ( .A1(n5961), .A2(n5937), .ZN(n7951) );
  NAND2_X1 U6930 ( .A1(n9184), .A2(n7951), .ZN(n5940) );
  NAND2_X1 U6931 ( .A1(n5786), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U6932 ( .A1(n4918), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5938) );
  NAND4_X1 U6933 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(n9562)
         );
  NAND2_X1 U6934 ( .A1(n9562), .A2(n6214), .ZN(n5942) );
  NAND2_X1 U6935 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  XNOR2_X1 U6936 ( .A(n5944), .B(n9173), .ZN(n5951) );
  AND2_X1 U6937 ( .A1(n9562), .A2(n6185), .ZN(n5945) );
  AOI21_X1 U6938 ( .B1(n8002), .B2(n6214), .A(n5945), .ZN(n5950) );
  XNOR2_X1 U6939 ( .A(n5951), .B(n5950), .ZN(n7958) );
  INV_X1 U6940 ( .A(n5946), .ZN(n5947) );
  NOR2_X1 U6941 ( .A1(n5948), .A2(n5947), .ZN(n7959) );
  XNOR2_X1 U6942 ( .A(n5953), .B(n5952), .ZN(n7124) );
  NAND2_X1 U6943 ( .A1(n7124), .A2(n9273), .ZN(n5959) );
  NOR2_X1 U6944 ( .A1(n5932), .A2(n5307), .ZN(n5954) );
  MUX2_X1 U6945 ( .A(n5307), .B(n5954), .S(P1_IR_REG_14__SCAN_IN), .Z(n5957)
         );
  INV_X1 U6946 ( .A(n5955), .ZN(n5956) );
  OR2_X1 U6947 ( .A1(n5957), .A2(n5956), .ZN(n10177) );
  AOI22_X1 U6948 ( .A1(n6032), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6031), .B2(
        n9637), .ZN(n5958) );
  NAND2_X1 U6949 ( .A1(n9986), .A2(n9169), .ZN(n5968) );
  NAND2_X1 U6950 ( .A1(n4916), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5966) );
  INV_X1 U6951 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U6952 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  AND2_X1 U6953 ( .A1(n5976), .A2(n5962), .ZN(n8051) );
  NAND2_X1 U6954 ( .A1(n9184), .A2(n8051), .ZN(n5965) );
  NAND2_X1 U6955 ( .A1(n5786), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U6956 ( .A1(n4918), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5963) );
  OR2_X1 U6957 ( .A1(n8004), .A2(n9170), .ZN(n5967) );
  NAND2_X1 U6958 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  AOI22_X1 U6959 ( .A1(n9986), .A2(n6214), .B1(n6185), .B2(n9561), .ZN(n8049)
         );
  XNOR2_X1 U6960 ( .A(n5971), .B(n5970), .ZN(n7191) );
  NAND2_X1 U6961 ( .A1(n7191), .A2(n9273), .ZN(n5974) );
  NAND2_X1 U6962 ( .A1(n5955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U6963 ( .A(n5972), .B(n5588), .ZN(n9639) );
  INV_X1 U6964 ( .A(n9639), .ZN(n10190) );
  AOI22_X1 U6965 ( .A1(n6032), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6031), .B2(
        n10190), .ZN(n5973) );
  NAND2_X1 U6966 ( .A1(n9980), .A2(n9169), .ZN(n5983) );
  NAND2_X1 U6967 ( .A1(n4916), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5981) );
  INV_X1 U6968 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U6969 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  AND2_X1 U6970 ( .A1(n5997), .A2(n5977), .ZN(n8061) );
  NAND2_X1 U6971 ( .A1(n9184), .A2(n8061), .ZN(n5980) );
  NAND2_X1 U6972 ( .A1(n4918), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U6973 ( .A1(n5786), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5978) );
  NAND4_X1 U6974 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n9560)
         );
  NAND2_X1 U6975 ( .A1(n9560), .A2(n6214), .ZN(n5982) );
  NAND2_X1 U6976 ( .A1(n5983), .A2(n5982), .ZN(n5984) );
  XNOR2_X1 U6977 ( .A(n5984), .B(n9173), .ZN(n8058) );
  AND2_X1 U6978 ( .A1(n9560), .A2(n6185), .ZN(n5985) );
  AOI21_X1 U6979 ( .B1(n9980), .B2(n6214), .A(n5985), .ZN(n5986) );
  NAND2_X1 U6980 ( .A1(n8058), .A2(n5986), .ZN(n5988) );
  INV_X1 U6981 ( .A(n8058), .ZN(n5987) );
  INV_X1 U6982 ( .A(n5986), .ZN(n8057) );
  XNOR2_X1 U6983 ( .A(n5990), .B(n5989), .ZN(n7316) );
  NAND2_X1 U6984 ( .A1(n7316), .A2(n9273), .ZN(n5995) );
  NAND2_X1 U6985 ( .A1(n5991), .A2(n5992), .ZN(n6009) );
  OR2_X1 U6986 ( .A1(n5991), .A2(n5992), .ZN(n5993) );
  AOI22_X1 U6987 ( .A1(n6032), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6031), .B2(
        n9656), .ZN(n5994) );
  NAND2_X1 U6988 ( .A1(n5995), .A2(n5994), .ZN(n9975) );
  NAND2_X1 U6989 ( .A1(n4916), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U6990 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  AND2_X1 U6991 ( .A1(n6014), .A2(n5998), .ZN(n8100) );
  NAND2_X1 U6992 ( .A1(n9184), .A2(n8100), .ZN(n6001) );
  NAND2_X1 U6993 ( .A1(n5786), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U6994 ( .A1(n4918), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5999) );
  OAI22_X1 U6995 ( .A1(n8130), .A2(n6183), .B1(n8108), .B2(n9170), .ZN(n6003)
         );
  XNOR2_X1 U6996 ( .A(n6003), .B(n6216), .ZN(n6005) );
  OAI22_X1 U6997 ( .A1(n8130), .A2(n9170), .B1(n8108), .B2(n9176), .ZN(n6004)
         );
  NOR2_X1 U6998 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  AOI21_X1 U6999 ( .B1(n6005), .B2(n6004), .A(n6006), .ZN(n8123) );
  XNOR2_X1 U7000 ( .A(n6008), .B(n6007), .ZN(n7374) );
  NAND2_X1 U7001 ( .A1(n7374), .A2(n9273), .ZN(n6012) );
  NAND2_X1 U7002 ( .A1(n6009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7003 ( .A(n6010), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U7004 ( .A1(n6032), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6031), .B2(
        n10201), .ZN(n6011) );
  NAND2_X1 U7005 ( .A1(n4916), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6019) );
  INV_X1 U7006 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7007 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  AND2_X1 U7008 ( .A1(n6037), .A2(n6015), .ZN(n9219) );
  NAND2_X1 U7009 ( .A1(n9184), .A2(n9219), .ZN(n6018) );
  NAND2_X1 U7010 ( .A1(n5786), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7011 ( .A1(n4918), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6016) );
  NOR2_X1 U7012 ( .A1(n9674), .A2(n9170), .ZN(n6020) );
  AOI21_X1 U7013 ( .B1(n9970), .B2(n9169), .A(n6020), .ZN(n6021) );
  XNOR2_X1 U7014 ( .A(n6021), .B(n6216), .ZN(n6024) );
  NOR2_X1 U7015 ( .A1(n9674), .A2(n9176), .ZN(n6022) );
  AOI21_X1 U7016 ( .B1(n9970), .B2(n6214), .A(n6022), .ZN(n6023) );
  OR2_X1 U7017 ( .A1(n6024), .A2(n6023), .ZN(n9216) );
  OAI22_X1 U7018 ( .A1(n9880), .A2(n6183), .B1(n9866), .B2(n9170), .ZN(n6025)
         );
  XNOR2_X1 U7019 ( .A(n6025), .B(n6216), .ZN(n6026) );
  NAND2_X1 U7020 ( .A1(n6027), .A2(n6026), .ZN(n9257) );
  AOI21_X2 U7021 ( .B1(n9259), .B2(n9257), .A(n9256), .ZN(n9163) );
  XNOR2_X1 U7022 ( .A(n6029), .B(n6028), .ZN(n7610) );
  NAND2_X1 U7023 ( .A1(n7610), .A2(n9273), .ZN(n6034) );
  AOI22_X1 U7024 ( .A1(n6032), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6031), .B2(
        n9778), .ZN(n6033) );
  NAND2_X1 U7025 ( .A1(n9960), .A2(n9169), .ZN(n6044) );
  INV_X1 U7026 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6036) );
  INV_X1 U7027 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6035) );
  OAI21_X1 U7028 ( .B1(n6037), .B2(n6036), .A(n6035), .ZN(n6038) );
  NAND2_X1 U7029 ( .A1(n6038), .A2(n6053), .ZN(n9860) );
  NAND2_X1 U7030 ( .A1(n4916), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7031 ( .A1(n5786), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6039) );
  AND2_X1 U7032 ( .A1(n6040), .A2(n6039), .ZN(n6042) );
  NAND2_X1 U7033 ( .A1(n4918), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6041) );
  OAI211_X1 U7034 ( .C1(n9860), .C2(n6207), .A(n6042), .B(n6041), .ZN(n9888)
         );
  NAND2_X1 U7035 ( .A1(n9888), .A2(n6214), .ZN(n6043) );
  NAND2_X1 U7036 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  XNOR2_X1 U7037 ( .A(n6045), .B(n6216), .ZN(n6048) );
  INV_X1 U7038 ( .A(n9960), .ZN(n9859) );
  INV_X1 U7039 ( .A(n9888), .ZN(n9678) );
  OAI22_X1 U7040 ( .A1(n9859), .A2(n9170), .B1(n9678), .B2(n9176), .ZN(n6047)
         );
  XNOR2_X1 U7041 ( .A(n6048), .B(n6047), .ZN(n9164) );
  XNOR2_X1 U7042 ( .A(n6050), .B(n6049), .ZN(n7649) );
  NAND2_X1 U7043 ( .A1(n7649), .A2(n9273), .ZN(n6052) );
  OR2_X1 U7044 ( .A1(n5778), .A2(n7650), .ZN(n6051) );
  INV_X1 U7045 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6058) );
  INV_X1 U7046 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U7047 ( .A1(n6053), .A2(n9238), .ZN(n6054) );
  NAND2_X1 U7048 ( .A1(n6055), .A2(n6054), .ZN(n9846) );
  OR2_X1 U7049 ( .A1(n9846), .A2(n6207), .ZN(n6057) );
  AOI22_X1 U7050 ( .A1(n4916), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n4918), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6056) );
  OAI211_X1 U7051 ( .C1(n6257), .C2(n6058), .A(n6057), .B(n6056), .ZN(n9679)
         );
  INV_X1 U7052 ( .A(n9679), .ZN(n9867) );
  OAI22_X1 U7053 ( .A1(n9849), .A2(n9170), .B1(n9867), .B2(n9176), .ZN(n6061)
         );
  OAI22_X1 U7054 ( .A1(n9849), .A2(n6183), .B1(n9867), .B2(n9170), .ZN(n6059)
         );
  XNOR2_X1 U7055 ( .A(n6059), .B(n6216), .ZN(n6060) );
  XOR2_X1 U7056 ( .A(n6061), .B(n6060), .Z(n9234) );
  INV_X1 U7057 ( .A(n6060), .ZN(n6063) );
  INV_X1 U7058 ( .A(n6061), .ZN(n6062) );
  XNOR2_X1 U7059 ( .A(n6065), .B(n6064), .ZN(n9202) );
  NAND2_X1 U7060 ( .A1(n6067), .A2(SI_21_), .ZN(n6092) );
  NAND2_X1 U7061 ( .A1(n6068), .A2(n6092), .ZN(n6069) );
  MUX2_X1 U7062 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n6656), .Z(n6083) );
  XNOR2_X1 U7063 ( .A(n6083), .B(SI_22_), .ZN(n6084) );
  NAND2_X1 U7064 ( .A1(n7819), .A2(n9273), .ZN(n6071) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7832) );
  OR2_X1 U7066 ( .A1(n5778), .A2(n7832), .ZN(n6070) );
  INV_X1 U7067 ( .A(n6073), .ZN(n6072) );
  NAND2_X1 U7068 ( .A1(n6072), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6108) );
  INV_X1 U7069 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U7070 ( .A1(n6073), .A2(n9249), .ZN(n6074) );
  NAND2_X1 U7071 ( .A1(n6108), .A2(n6074), .ZN(n9820) );
  OR2_X1 U7072 ( .A1(n9820), .A2(n6207), .ZN(n6079) );
  INV_X1 U7073 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U7074 ( .A1(n4916), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7075 ( .A1(n4918), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6075) );
  OAI211_X1 U7076 ( .C1(n9821), .C2(n6257), .A(n6076), .B(n6075), .ZN(n6077)
         );
  INV_X1 U7077 ( .A(n6077), .ZN(n6078) );
  AOI22_X1 U7078 ( .A1(n9943), .A2(n9169), .B1(n6214), .B2(n9680), .ZN(n6080)
         );
  XOR2_X1 U7079 ( .A(n6216), .B(n6080), .Z(n6081) );
  INV_X1 U7080 ( .A(n9943), .ZN(n9819) );
  OAI22_X1 U7081 ( .A1(n9819), .A2(n9170), .B1(n9834), .B2(n9176), .ZN(n9247)
         );
  AOI21_X2 U7082 ( .B1(n9244), .B2(n9247), .A(n9245), .ZN(n9156) );
  NAND2_X1 U7083 ( .A1(n6083), .A2(SI_22_), .ZN(n6091) );
  INV_X1 U7084 ( .A(n6091), .ZN(n6086) );
  INV_X1 U7085 ( .A(n6084), .ZN(n6085) );
  INV_X1 U7086 ( .A(n6090), .ZN(n6094) );
  AND2_X1 U7087 ( .A1(n6092), .A2(n6091), .ZN(n6093) );
  MUX2_X1 U7088 ( .A(n7752), .B(n7757), .S(n8141), .Z(n6095) );
  INV_X1 U7089 ( .A(SI_23_), .ZN(n9005) );
  NAND2_X1 U7090 ( .A1(n6095), .A2(n9005), .ZN(n6121) );
  INV_X1 U7091 ( .A(n6095), .ZN(n6096) );
  NAND2_X1 U7092 ( .A1(n6096), .A2(SI_23_), .ZN(n6097) );
  NAND2_X1 U7093 ( .A1(n6121), .A2(n6097), .ZN(n6102) );
  INV_X1 U7094 ( .A(n6102), .ZN(n6098) );
  NAND2_X1 U7095 ( .A1(n6101), .A2(n6100), .ZN(n6103) );
  NAND2_X1 U7096 ( .A1(n6103), .A2(n6102), .ZN(n6104) );
  NAND2_X1 U7097 ( .A1(n6122), .A2(n6104), .ZN(n7755) );
  NAND2_X1 U7098 ( .A1(n7755), .A2(n9273), .ZN(n6106) );
  OR2_X1 U7099 ( .A1(n5778), .A2(n7757), .ZN(n6105) );
  NAND2_X1 U7100 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  AND2_X1 U7101 ( .A1(n6129), .A2(n6109), .ZN(n9800) );
  NAND2_X1 U7102 ( .A1(n9800), .A2(n9184), .ZN(n6115) );
  INV_X1 U7103 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7104 ( .A1(n4916), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7105 ( .A1(n4918), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6110) );
  OAI211_X1 U7106 ( .C1(n6112), .C2(n6257), .A(n6111), .B(n6110), .ZN(n6113)
         );
  INV_X1 U7107 ( .A(n6113), .ZN(n6114) );
  AOI22_X1 U7108 ( .A1(n9939), .A2(n9169), .B1(n6214), .B2(n9783), .ZN(n6116)
         );
  XNOR2_X1 U7109 ( .A(n6116), .B(n6216), .ZN(n6117) );
  OAI22_X1 U7110 ( .A1(n5168), .A2(n9170), .B1(n9809), .B2(n9176), .ZN(n6118)
         );
  XNOR2_X1 U7111 ( .A(n6117), .B(n6118), .ZN(n9157) );
  INV_X1 U7112 ( .A(n6118), .ZN(n6119) );
  NAND2_X1 U7113 ( .A1(n9155), .A2(n6120), .ZN(n9224) );
  INV_X1 U7114 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7921) );
  INV_X1 U7115 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7862) );
  MUX2_X1 U7116 ( .A(n7921), .B(n7862), .S(n6656), .Z(n6123) );
  NAND2_X1 U7117 ( .A1(n6123), .A2(n9017), .ZN(n6149) );
  INV_X1 U7118 ( .A(n6123), .ZN(n6124) );
  NAND2_X1 U7119 ( .A1(n6124), .A2(SI_24_), .ZN(n6125) );
  XNOR2_X1 U7120 ( .A(n6148), .B(n6147), .ZN(n7861) );
  NAND2_X1 U7121 ( .A1(n7861), .A2(n9273), .ZN(n6127) );
  OR2_X1 U7122 ( .A1(n5778), .A2(n7862), .ZN(n6126) );
  NAND2_X1 U7123 ( .A1(n9934), .A2(n9169), .ZN(n6138) );
  INV_X1 U7124 ( .A(n6129), .ZN(n6128) );
  NAND2_X1 U7125 ( .A1(n6128), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6154) );
  INV_X1 U7126 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U7127 ( .A1(n6129), .A2(n9228), .ZN(n6130) );
  NAND2_X1 U7128 ( .A1(n6154), .A2(n6130), .ZN(n9777) );
  INV_X1 U7129 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7130 ( .A1(n4916), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7131 ( .A1(n4918), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6131) );
  OAI211_X1 U7132 ( .C1(n6257), .C2(n6133), .A(n6132), .B(n6131), .ZN(n6134)
         );
  INV_X1 U7133 ( .A(n6134), .ZN(n6135) );
  NAND2_X1 U7134 ( .A1(n9681), .A2(n6214), .ZN(n6137) );
  NAND2_X1 U7135 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  XNOR2_X1 U7136 ( .A(n6139), .B(n6216), .ZN(n6142) );
  NAND2_X1 U7137 ( .A1(n9934), .A2(n6214), .ZN(n6141) );
  NAND2_X1 U7138 ( .A1(n9681), .A2(n6185), .ZN(n6140) );
  NAND2_X1 U7139 ( .A1(n6141), .A2(n6140), .ZN(n6143) );
  NAND2_X1 U7140 ( .A1(n6142), .A2(n6143), .ZN(n9225) );
  NAND2_X1 U7141 ( .A1(n9224), .A2(n9225), .ZN(n6146) );
  INV_X1 U7142 ( .A(n6142), .ZN(n6145) );
  INV_X1 U7143 ( .A(n6143), .ZN(n6144) );
  NAND2_X1 U7144 ( .A1(n6145), .A2(n6144), .ZN(n9226) );
  NAND2_X1 U7145 ( .A1(n6146), .A2(n9226), .ZN(n9208) );
  NAND2_X1 U7146 ( .A1(n6148), .A2(n6147), .ZN(n6150) );
  MUX2_X1 U7147 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n8141), .Z(n6167) );
  INV_X1 U7148 ( .A(SI_25_), .ZN(n9008) );
  XNOR2_X1 U7149 ( .A(n6167), .B(n9008), .ZN(n6164) );
  XNOR2_X1 U7150 ( .A(n6166), .B(n6164), .ZN(n7894) );
  NAND2_X1 U7151 ( .A1(n7894), .A2(n9273), .ZN(n6152) );
  INV_X1 U7152 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7895) );
  OR2_X1 U7153 ( .A1(n5778), .A2(n7895), .ZN(n6151) );
  INV_X1 U7154 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7155 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U7156 ( .A1(n6175), .A2(n6155), .ZN(n9768) );
  INV_X1 U7157 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U7158 ( .A1(n4916), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7159 ( .A1(n4918), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6156) );
  OAI211_X1 U7160 ( .C1(n6257), .C2(n9767), .A(n6157), .B(n6156), .ZN(n6158)
         );
  INV_X1 U7161 ( .A(n6158), .ZN(n6159) );
  OAI22_X1 U7162 ( .A1(n5164), .A2(n9170), .B1(n9786), .B2(n9176), .ZN(n6189)
         );
  NAND2_X1 U7163 ( .A1(n9929), .A2(n9169), .ZN(n6162) );
  INV_X1 U7164 ( .A(n9786), .ZN(n9558) );
  NAND2_X1 U7165 ( .A1(n9558), .A2(n6214), .ZN(n6161) );
  NAND2_X1 U7166 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  XNOR2_X1 U7167 ( .A(n6163), .B(n6216), .ZN(n6188) );
  XOR2_X1 U7168 ( .A(n6189), .B(n6188), .Z(n9209) );
  INV_X1 U7169 ( .A(n6164), .ZN(n6165) );
  NAND2_X1 U7170 ( .A1(n6167), .A2(SI_25_), .ZN(n6168) );
  INV_X1 U7171 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8020) );
  INV_X1 U7172 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8017) );
  MUX2_X1 U7173 ( .A(n8020), .B(n8017), .S(n6656), .Z(n6170) );
  INV_X1 U7174 ( .A(SI_26_), .ZN(n6169) );
  NAND2_X1 U7175 ( .A1(n6170), .A2(n6169), .ZN(n6196) );
  INV_X1 U7176 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7177 ( .A1(n6171), .A2(SI_26_), .ZN(n6172) );
  NAND2_X1 U7178 ( .A1(n6196), .A2(n6172), .ZN(n6197) );
  NAND2_X1 U7179 ( .A1(n8015), .A2(n9273), .ZN(n6174) );
  OR2_X1 U7180 ( .A1(n5778), .A2(n8017), .ZN(n6173) );
  NAND2_X1 U7181 ( .A1(n6175), .A2(n6275), .ZN(n6176) );
  NAND2_X1 U7182 ( .A1(n9754), .A2(n9184), .ZN(n6182) );
  INV_X1 U7183 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7184 ( .A1(n4916), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7185 ( .A1(n4918), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6177) );
  OAI211_X1 U7186 ( .C1(n6179), .C2(n6257), .A(n6178), .B(n6177), .ZN(n6180)
         );
  INV_X1 U7187 ( .A(n6180), .ZN(n6181) );
  OAI22_X1 U7188 ( .A1(n9757), .A2(n6183), .B1(n9763), .B2(n9170), .ZN(n6184)
         );
  XNOR2_X1 U7189 ( .A(n6184), .B(n9173), .ZN(n6193) );
  OR2_X1 U7190 ( .A1(n9757), .A2(n9170), .ZN(n6187) );
  NAND2_X1 U7191 ( .A1(n9684), .A2(n6185), .ZN(n6186) );
  NAND2_X1 U7192 ( .A1(n6187), .A2(n6186), .ZN(n6194) );
  XNOR2_X1 U7193 ( .A(n6193), .B(n6194), .ZN(n6272) );
  INV_X1 U7194 ( .A(n6188), .ZN(n6191) );
  INV_X1 U7195 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7196 ( .A1(n6191), .A2(n6190), .ZN(n6271) );
  INV_X1 U7197 ( .A(n6193), .ZN(n6195) );
  NAND2_X1 U7198 ( .A1(n6195), .A2(n6194), .ZN(n6219) );
  INV_X1 U7199 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6640) );
  INV_X1 U7200 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8001) );
  MUX2_X1 U7201 ( .A(n6640), .B(n8001), .S(n8141), .Z(n6199) );
  INV_X1 U7202 ( .A(SI_27_), .ZN(n8912) );
  NAND2_X1 U7203 ( .A1(n6199), .A2(n8912), .ZN(n6654) );
  INV_X1 U7204 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7205 ( .A1(n6200), .A2(SI_27_), .ZN(n6201) );
  XNOR2_X1 U7206 ( .A(n6653), .B(n6652), .ZN(n7983) );
  NAND2_X1 U7207 ( .A1(n7983), .A2(n9273), .ZN(n6203) );
  OR2_X1 U7208 ( .A1(n5778), .A2(n8001), .ZN(n6202) );
  INV_X1 U7209 ( .A(n6205), .ZN(n6204) );
  NAND2_X1 U7210 ( .A1(n6204), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9183) );
  INV_X1 U7211 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7212 ( .A1(n6205), .A2(n6254), .ZN(n6206) );
  NAND2_X1 U7213 ( .A1(n9183), .A2(n6206), .ZN(n9734) );
  INV_X1 U7214 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7215 ( .A1(n4916), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7216 ( .A1(n4918), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6208) );
  OAI211_X1 U7217 ( .C1(n6210), .C2(n6257), .A(n6209), .B(n6208), .ZN(n6211)
         );
  INV_X1 U7218 ( .A(n6211), .ZN(n6212) );
  AOI22_X1 U7219 ( .A1(n9916), .A2(n9169), .B1(n6214), .B2(n9726), .ZN(n6215)
         );
  XOR2_X1 U7220 ( .A(n6216), .B(n6215), .Z(n6218) );
  INV_X1 U7221 ( .A(n9916), .ZN(n9737) );
  OAI22_X1 U7222 ( .A1(n9737), .A2(n9170), .B1(n9750), .B2(n9176), .ZN(n6217)
         );
  NOR2_X1 U7223 ( .A1(n6218), .A2(n6217), .ZN(n9196) );
  AOI21_X1 U7224 ( .B1(n6218), .B2(n6217), .A(n9196), .ZN(n6220) );
  AOI21_X1 U7225 ( .B1(n6274), .B2(n6219), .A(n6220), .ZN(n6241) );
  NAND2_X1 U7226 ( .A1(n7896), .A2(P1_B_REG_SCAN_IN), .ZN(n6222) );
  INV_X1 U7227 ( .A(n7863), .ZN(n6221) );
  MUX2_X1 U7228 ( .A(n6222), .B(P1_B_REG_SCAN_IN), .S(n6221), .Z(n6223) );
  INV_X1 U7229 ( .A(n6224), .ZN(n8016) );
  NAND2_X1 U7230 ( .A1(n8016), .A2(n7896), .ZN(n10010) );
  OAI21_X1 U7231 ( .B1(n6823), .B2(P1_D_REG_1__SCAN_IN), .A(n10010), .ZN(n7254) );
  INV_X1 U7232 ( .A(n7254), .ZN(n7397) );
  INV_X1 U7233 ( .A(n6823), .ZN(n6233) );
  INV_X1 U7234 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6827) );
  AND2_X1 U7235 ( .A1(n8016), .A2(n7863), .ZN(n6826) );
  NOR4_X1 U7236 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6228) );
  NOR4_X1 U7237 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6227) );
  NOR4_X1 U7238 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6226) );
  NOR4_X1 U7239 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6225) );
  NAND4_X1 U7240 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n6235)
         );
  NOR2_X1 U7241 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6232) );
  NOR4_X1 U7242 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6231) );
  NOR4_X1 U7243 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6230) );
  NOR4_X1 U7244 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6229) );
  NAND4_X1 U7245 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n6234)
         );
  OAI21_X1 U7246 ( .B1(n6235), .B2(n6234), .A(n6233), .ZN(n7251) );
  NAND3_X1 U7247 ( .A1(n7397), .A2(n7320), .A3(n7251), .ZN(n6250) );
  INV_X1 U7248 ( .A(n10444), .ZN(n10451) );
  NAND2_X1 U7249 ( .A1(n6236), .A2(n9550), .ZN(n6251) );
  NOR2_X1 U7250 ( .A1(n10490), .A2(n9471), .ZN(n6246) );
  NAND2_X1 U7251 ( .A1(n6246), .A2(n6824), .ZN(n6240) );
  INV_X1 U7252 ( .A(n6824), .ZN(n9549) );
  OR2_X1 U7253 ( .A1(n10444), .A2(n9544), .ZN(n7405) );
  OR2_X1 U7254 ( .A1(n9549), .A2(n7405), .ZN(n6242) );
  OR2_X1 U7255 ( .A1(n6250), .A2(n6242), .ZN(n6244) );
  OR2_X1 U7256 ( .A1(n9549), .A2(n10450), .ZN(n6248) );
  OR2_X1 U7257 ( .A1(n6250), .A2(n6248), .ZN(n6262) );
  NOR2_X2 U7258 ( .A1(n6262), .A2(n4908), .ZN(n9261) );
  INV_X1 U7259 ( .A(n6246), .ZN(n6247) );
  NAND3_X1 U7260 ( .A1(n6248), .A2(n7405), .A3(n6247), .ZN(n6249) );
  NAND2_X1 U7261 ( .A1(n6250), .A2(n6249), .ZN(n6253) );
  INV_X1 U7262 ( .A(n7237), .ZN(n9545) );
  OAI211_X1 U7263 ( .C1(n9545), .C2(n6251), .A(n5680), .B(n6821), .ZN(n7250)
         );
  INV_X1 U7264 ( .A(n7250), .ZN(n6252) );
  NAND2_X1 U7265 ( .A1(n6253), .A2(n6252), .ZN(n7081) );
  OAI22_X1 U7266 ( .A1(n9734), .A2(n9251), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6254), .ZN(n6265) );
  XNOR2_X1 U7267 ( .A(n9183), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U7268 ( .A1(n9720), .A2(n9184), .ZN(n6261) );
  INV_X1 U7269 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7270 ( .A1(n4916), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7271 ( .A1(n4918), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6255) );
  OAI211_X1 U7272 ( .C1(n6258), .C2(n6257), .A(n6256), .B(n6255), .ZN(n6259)
         );
  INV_X1 U7273 ( .A(n6259), .ZN(n6260) );
  INV_X1 U7274 ( .A(n6262), .ZN(n6263) );
  NOR2_X1 U7275 ( .A1(n9741), .A2(n9264), .ZN(n6264) );
  AOI211_X1 U7276 ( .C1(n9261), .C2(n9684), .A(n6265), .B(n6264), .ZN(n6266)
         );
  OAI21_X1 U7277 ( .B1(n9737), .B2(n9243), .A(n6266), .ZN(n6267) );
  INV_X1 U7278 ( .A(n6267), .ZN(n6268) );
  AND2_X1 U7279 ( .A1(n6270), .A2(n6271), .ZN(n6273) );
  NAND2_X1 U7280 ( .A1(n6274), .A2(n9235), .ZN(n6281) );
  OAI22_X1 U7281 ( .A1(n9786), .A2(n9250), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6275), .ZN(n6277) );
  NOR2_X1 U7282 ( .A1(n9750), .A2(n9264), .ZN(n6276) );
  AOI211_X1 U7283 ( .C1(n9262), .C2(n9754), .A(n6277), .B(n6276), .ZN(n6278)
         );
  INV_X1 U7284 ( .A(n6279), .ZN(n6280) );
  OAI21_X1 U7285 ( .B1(n6282), .B2(n6281), .A(n6280), .ZN(P1_U3240) );
  NOR2_X1 U7286 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6288) );
  NAND2_X1 U7287 ( .A1(n6364), .A2(n6289), .ZN(n6324) );
  INV_X1 U7288 ( .A(n6309), .ZN(n6301) );
  XNOR2_X2 U7289 ( .A(n6295), .B(n6308), .ZN(n6845) );
  NAND2_X1 U7290 ( .A1(n6296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7291 ( .A1(n6297), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6300) );
  NAND2_X4 U7292 ( .A1(n6302), .A2(n6301), .ZN(n8619) );
  NAND2_X1 U7293 ( .A1(n7610), .A2(n8296), .ZN(n6305) );
  NAND2_X1 U7294 ( .A1(n6303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7295 ( .A1(n6565), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6367), .B2(
        n8633), .ZN(n6304) );
  NOR2_X1 U7296 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6306) );
  NAND2_X1 U7297 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  NAND2_X2 U7298 ( .A1(n8204), .A2(n9146), .ZN(n6378) );
  NAND2_X1 U7299 ( .A1(n8306), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6317) );
  INV_X1 U7300 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8852) );
  OR2_X1 U7301 ( .A1(n6677), .A2(n8852), .ZN(n6316) );
  NOR2_X1 U7302 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6413) );
  INV_X1 U7303 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U7304 ( .A1(n6413), .A2(n6414), .ZN(n6428) );
  NAND2_X1 U7305 ( .A1(n6475), .A2(n6474), .ZN(n6489) );
  NOR2_X2 U7306 ( .A1(n6513), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U7307 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  NOR2_X2 U7308 ( .A1(n6343), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U7309 ( .A1(n8604), .A2(n6568), .ZN(n6570) );
  NOR2_X2 U7310 ( .A1(n6570), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6578) );
  AOI21_X1 U7311 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n6570), .A(n6578), .ZN(
        n8775) );
  OR2_X1 U7312 ( .A1(n6376), .A2(n8775), .ZN(n6315) );
  INV_X1 U7313 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8776) );
  OR2_X1 U7314 ( .A1(n6374), .A2(n8776), .ZN(n6314) );
  NAND2_X1 U7315 ( .A1(n8306), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6323) );
  INV_X1 U7316 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6318) );
  OR2_X1 U7317 ( .A1(n6677), .A2(n6318), .ZN(n6322) );
  AND2_X1 U7318 ( .A1(n6343), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6319) );
  NOR2_X1 U7319 ( .A1(n6546), .A2(n6319), .ZN(n7991) );
  OR2_X1 U7320 ( .A1(n6376), .A2(n7991), .ZN(n6321) );
  INV_X1 U7321 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7968) );
  OR2_X1 U7322 ( .A1(n6374), .A2(n7968), .ZN(n6320) );
  NAND4_X1 U7323 ( .A1(n6323), .A2(n6322), .A3(n6321), .A4(n6320), .ZN(n8527)
         );
  NAND2_X1 U7324 ( .A1(n7191), .A2(n8296), .ZN(n6338) );
  NAND4_X1 U7325 ( .A1(n6325), .A2(n6435), .A3(n6420), .A4(n6451), .ZN(n6326)
         );
  INV_X1 U7326 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7327 ( .A1(n6484), .A2(n6327), .ZN(n6328) );
  NAND2_X1 U7328 ( .A1(n6328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6496) );
  INV_X1 U7329 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7330 ( .A1(n6496), .A2(n6329), .ZN(n6330) );
  NAND2_X1 U7331 ( .A1(n6330), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6509) );
  INV_X1 U7332 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7333 ( .A1(n6509), .A2(n6331), .ZN(n6332) );
  NAND2_X1 U7334 ( .A1(n6332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U7335 ( .A1(n6521), .A2(n6333), .ZN(n6334) );
  NAND2_X1 U7336 ( .A1(n6334), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6339) );
  INV_X1 U7337 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7338 ( .A1(n6339), .A2(n6335), .ZN(n6336) );
  NAND2_X1 U7339 ( .A1(n6336), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6539) );
  XNOR2_X1 U7340 ( .A(n6539), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U7341 ( .A1(n6565), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10372), 
        .B2(n6367), .ZN(n6337) );
  NAND2_X1 U7342 ( .A1(n7124), .A2(n8296), .ZN(n6341) );
  XNOR2_X1 U7343 ( .A(n6339), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U7344 ( .A1(n6565), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6367), .B2(
        n10356), .ZN(n6340) );
  NAND2_X1 U7345 ( .A1(n6341), .A2(n6340), .ZN(n7934) );
  INV_X1 U7346 ( .A(n7934), .ZN(n7933) );
  NAND2_X1 U7347 ( .A1(n8306), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6348) );
  INV_X1 U7348 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8550) );
  OR2_X1 U7349 ( .A1(n6677), .A2(n8550), .ZN(n6347) );
  NAND2_X1 U7350 ( .A1(n6527), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6342) );
  AND2_X1 U7351 ( .A1(n6343), .A2(n6342), .ZN(n7904) );
  OR2_X1 U7352 ( .A1(n6376), .A2(n7904), .ZN(n6346) );
  INV_X1 U7353 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6344) );
  OR2_X1 U7354 ( .A1(n6374), .A2(n6344), .ZN(n6345) );
  INV_X1 U7355 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6349) );
  INV_X1 U7356 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6839) );
  INV_X1 U7357 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7011) );
  OR2_X1 U7358 ( .A1(n6374), .A2(n7011), .ZN(n6350) );
  INV_X1 U7359 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6997) );
  NAND2_X1 U7360 ( .A1(n8286), .A2(SI_0_), .ZN(n6354) );
  INV_X1 U7361 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7362 ( .A1(n6354), .A2(n6353), .ZN(n6356) );
  AND2_X1 U7363 ( .A1(n6356), .A2(n6355), .ZN(n9154) );
  MUX2_X1 U7364 ( .A(n4996), .B(n9154), .S(n6357), .Z(n7051) );
  NAND2_X1 U7365 ( .A1(n7132), .A2(n7051), .ZN(n7131) );
  INV_X1 U7366 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7093) );
  INV_X1 U7367 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6358) );
  INV_X1 U7368 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6359) );
  OR2_X1 U7369 ( .A1(n6378), .A2(n6359), .ZN(n6360) );
  OR2_X1 U7370 ( .A1(n6383), .A2(n6362), .ZN(n6370) );
  NAND2_X1 U7371 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6363) );
  MUX2_X1 U7372 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6363), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6366) );
  INV_X1 U7373 ( .A(n6860), .ZN(n6365) );
  NAND2_X1 U7374 ( .A1(n6367), .A2(n6878), .ZN(n6368) );
  INV_X1 U7375 ( .A(n7310), .ZN(n6372) );
  NAND2_X1 U7376 ( .A1(n6371), .A2(n7310), .ZN(n8343) );
  NAND2_X1 U7377 ( .A1(n7131), .A2(n7128), .ZN(n7130) );
  NAND2_X1 U7378 ( .A1(n6371), .A2(n6372), .ZN(n6373) );
  NAND2_X1 U7379 ( .A1(n7130), .A2(n6373), .ZN(n7101) );
  INV_X1 U7380 ( .A(n6374), .ZN(n6375) );
  NAND2_X1 U7381 ( .A1(n6375), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6382) );
  INV_X1 U7382 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10467) );
  OR2_X1 U7383 ( .A1(n6376), .A2(n10467), .ZN(n6381) );
  INV_X1 U7384 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6377) );
  OR2_X1 U7385 ( .A1(n6378), .A2(n6377), .ZN(n6379) );
  OR2_X1 U7386 ( .A1(n6383), .A2(n6793), .ZN(n6388) );
  INV_X1 U7387 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6789) );
  OR2_X1 U7388 ( .A1(n6384), .A2(n6789), .ZN(n6387) );
  NOR2_X1 U7389 ( .A1(n6860), .A2(n9139), .ZN(n6385) );
  OR2_X1 U7390 ( .A1(n6357), .A2(n6863), .ZN(n6386) );
  XNOR2_X1 U7391 ( .A(n8539), .B(n10470), .ZN(n8338) );
  NAND2_X1 U7392 ( .A1(n7101), .A2(n8338), .ZN(n7100) );
  INV_X1 U7393 ( .A(n8539), .ZN(n7109) );
  NAND2_X1 U7394 ( .A1(n7109), .A2(n10470), .ZN(n6389) );
  NAND2_X1 U7395 ( .A1(n7100), .A2(n6389), .ZN(n7107) );
  NAND2_X1 U7396 ( .A1(n8300), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6395) );
  OR2_X1 U7397 ( .A1(n6376), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6394) );
  INV_X1 U7398 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6390) );
  INV_X1 U7399 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6391) );
  OR2_X1 U7400 ( .A1(n6378), .A2(n6391), .ZN(n6392) );
  NAND2_X1 U7401 ( .A1(n6324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6396) );
  MUX2_X1 U7402 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6396), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6397) );
  NAND2_X1 U7403 ( .A1(n6397), .A2(n6408), .ZN(n6949) );
  OR2_X1 U7404 ( .A1(n6383), .A2(n6799), .ZN(n6399) );
  INV_X1 U7405 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6788) );
  OAI211_X1 U7406 ( .C1(n8643), .C2(n6949), .A(n6399), .B(n6398), .ZN(n7073)
         );
  NAND2_X1 U7407 ( .A1(n8538), .A2(n7073), .ZN(n6400) );
  NAND2_X1 U7408 ( .A1(n7107), .A2(n6400), .ZN(n6402) );
  NAND2_X1 U7409 ( .A1(n7140), .A2(n7273), .ZN(n6401) );
  NAND2_X1 U7410 ( .A1(n6402), .A2(n6401), .ZN(n7138) );
  NAND2_X1 U7411 ( .A1(n8306), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6407) );
  INV_X1 U7412 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6953) );
  OR2_X1 U7413 ( .A1(n6677), .A2(n6953), .ZN(n6406) );
  AND2_X1 U7414 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6403) );
  NOR2_X1 U7415 ( .A1(n6413), .A2(n6403), .ZN(n7279) );
  OR2_X1 U7416 ( .A1(n6376), .A2(n7279), .ZN(n6405) );
  INV_X1 U7417 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6956) );
  OR2_X1 U7418 ( .A1(n6374), .A2(n6956), .ZN(n6404) );
  NAND4_X1 U7419 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(n8537)
         );
  NAND2_X1 U7420 ( .A1(n6408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6421) );
  OR2_X1 U7421 ( .A1(n6383), .A2(n6795), .ZN(n6410) );
  OR2_X1 U7422 ( .A1(n8297), .A2(n4993), .ZN(n6409) );
  OAI211_X1 U7423 ( .C1(n8643), .C2(n10270), .A(n6410), .B(n6409), .ZN(n7115)
         );
  NOR2_X1 U7424 ( .A1(n8537), .A2(n7115), .ZN(n6412) );
  NAND2_X1 U7425 ( .A1(n8537), .A2(n7115), .ZN(n6411) );
  NAND2_X1 U7426 ( .A1(n8306), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6419) );
  INV_X1 U7427 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7027) );
  OR2_X1 U7428 ( .A1(n6677), .A2(n7027), .ZN(n6418) );
  OR2_X1 U7429 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  AND2_X1 U7430 ( .A1(n6428), .A2(n6415), .ZN(n7186) );
  OR2_X1 U7431 ( .A1(n6376), .A2(n7186), .ZN(n6417) );
  OR2_X1 U7432 ( .A1(n6374), .A2(n5364), .ZN(n6416) );
  NAND4_X1 U7433 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n8536)
         );
  NAND2_X1 U7434 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  NAND2_X1 U7435 ( .A1(n6422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6436) );
  XNOR2_X1 U7436 ( .A(n6436), .B(n6435), .ZN(n6961) );
  NAND2_X1 U7437 ( .A1(n6423), .A2(n8296), .ZN(n6425) );
  INV_X1 U7438 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6791) );
  OR2_X1 U7439 ( .A1(n8297), .A2(n6791), .ZN(n6424) );
  OAI211_X1 U7440 ( .C1(n8643), .C2(n6961), .A(n6425), .B(n6424), .ZN(n7188)
         );
  AND2_X1 U7441 ( .A1(n8536), .A2(n7188), .ZN(n6426) );
  INV_X1 U7442 ( .A(n7188), .ZN(n7170) );
  NAND2_X1 U7443 ( .A1(n7289), .A2(n7170), .ZN(n6427) );
  NAND2_X1 U7444 ( .A1(n8306), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6433) );
  INV_X1 U7445 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7023) );
  OR2_X1 U7446 ( .A1(n6677), .A2(n7023), .ZN(n6432) );
  NAND2_X1 U7447 ( .A1(n6428), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6429) );
  AND2_X1 U7448 ( .A1(n6442), .A2(n6429), .ZN(n7294) );
  OR2_X1 U7449 ( .A1(n6376), .A2(n7294), .ZN(n6431) );
  INV_X1 U7450 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7144) );
  OR2_X1 U7451 ( .A1(n6374), .A2(n7144), .ZN(n6430) );
  NAND4_X1 U7452 ( .A1(n6433), .A2(n6432), .A3(n6431), .A4(n6430), .ZN(n8535)
         );
  NAND2_X1 U7453 ( .A1(n6434), .A2(n8296), .ZN(n6439) );
  NAND2_X1 U7454 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  NAND2_X1 U7455 ( .A1(n6437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6449) );
  XNOR2_X1 U7456 ( .A(n6449), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8131) );
  AOI22_X1 U7457 ( .A1(n6565), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6367), .B2(
        n8131), .ZN(n6438) );
  NAND2_X1 U7458 ( .A1(n6439), .A2(n6438), .ZN(n7199) );
  AOI21_X2 U7459 ( .B1(n6440), .B2(n5481), .A(n5480), .ZN(n7593) );
  NAND2_X1 U7460 ( .A1(n8300), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6447) );
  INV_X1 U7461 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6441) );
  OR2_X1 U7462 ( .A1(n6378), .A2(n6441), .ZN(n6446) );
  AND2_X1 U7463 ( .A1(n6442), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6443) );
  NOR2_X1 U7464 ( .A1(n6461), .A2(n6443), .ZN(n10566) );
  OR2_X1 U7465 ( .A1(n6376), .A2(n10566), .ZN(n6445) );
  OR2_X1 U7466 ( .A1(n6374), .A2(n5374), .ZN(n6444) );
  NAND2_X1 U7467 ( .A1(n6803), .A2(n8296), .ZN(n6455) );
  INV_X1 U7468 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U7469 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  NAND2_X1 U7470 ( .A1(n6450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6452) );
  NAND2_X1 U7471 ( .A1(n6452), .A2(n6451), .ZN(n6456) );
  OR2_X1 U7472 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  AOI22_X1 U7473 ( .A1(n6565), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6367), .B2(
        n7150), .ZN(n6454) );
  NAND2_X1 U7474 ( .A1(n6455), .A2(n6454), .ZN(n10569) );
  OR2_X1 U7475 ( .A1(n7554), .A2(n10569), .ZN(n7443) );
  NAND2_X1 U7476 ( .A1(n10569), .A2(n7554), .ZN(n8379) );
  NAND2_X1 U7477 ( .A1(n7443), .A2(n8379), .ZN(n8488) );
  NAND2_X1 U7478 ( .A1(n7593), .A2(n8488), .ZN(n7594) );
  OR2_X1 U7479 ( .A1(n8534), .A2(n10569), .ZN(n7438) );
  NAND2_X1 U7480 ( .A1(n7594), .A2(n7438), .ZN(n6467) );
  NAND2_X1 U7481 ( .A1(n6813), .A2(n8296), .ZN(n6459) );
  NAND2_X1 U7482 ( .A1(n6456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6457) );
  XNOR2_X1 U7483 ( .A(n6457), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7459) );
  AOI22_X1 U7484 ( .A1(n6565), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6367), .B2(
        n7459), .ZN(n6458) );
  NAND2_X1 U7485 ( .A1(n6459), .A2(n6458), .ZN(n7615) );
  NAND2_X1 U7486 ( .A1(n8306), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6466) );
  INV_X1 U7487 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6460) );
  OR2_X1 U7488 ( .A1(n6677), .A2(n6460), .ZN(n6465) );
  NOR2_X1 U7489 ( .A1(n6461), .A2(n9078), .ZN(n6462) );
  OR2_X1 U7490 ( .A1(n6376), .A2(n5467), .ZN(n6464) );
  INV_X1 U7491 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7447) );
  OR2_X1 U7492 ( .A1(n6374), .A2(n7447), .ZN(n6463) );
  OR2_X1 U7493 ( .A1(n7615), .A2(n7598), .ZN(n8368) );
  NAND2_X1 U7494 ( .A1(n7615), .A2(n7598), .ZN(n8380) );
  NAND2_X1 U7495 ( .A1(n8368), .A2(n8380), .ZN(n8487) );
  NAND2_X1 U7496 ( .A1(n6467), .A2(n8487), .ZN(n7437) );
  OR2_X1 U7497 ( .A1(n7615), .A2(n8533), .ZN(n7583) );
  NAND2_X1 U7498 ( .A1(n6828), .A2(n8296), .ZN(n6473) );
  NAND2_X1 U7499 ( .A1(n6468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6469) );
  MUX2_X1 U7500 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6469), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n6470) );
  INV_X1 U7501 ( .A(n6470), .ZN(n6471) );
  NOR2_X1 U7502 ( .A1(n6471), .A2(n6484), .ZN(n8541) );
  AOI22_X1 U7503 ( .A1(n6565), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6367), .B2(
        n8541), .ZN(n6472) );
  NAND2_X1 U7504 ( .A1(n8306), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6480) );
  INV_X1 U7505 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7460) );
  OR2_X1 U7506 ( .A1(n6677), .A2(n7460), .ZN(n6479) );
  OR2_X1 U7507 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  AND2_X1 U7508 ( .A1(n6489), .A2(n6476), .ZN(n7696) );
  OR2_X1 U7509 ( .A1(n6376), .A2(n7696), .ZN(n6478) );
  INV_X1 U7510 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7461) );
  OR2_X1 U7511 ( .A1(n6374), .A2(n7461), .ZN(n6477) );
  OR2_X1 U7512 ( .A1(n7703), .A2(n5136), .ZN(n6481) );
  AND2_X1 U7513 ( .A1(n7583), .A2(n6481), .ZN(n6483) );
  INV_X1 U7514 ( .A(n6481), .ZN(n6482) );
  NAND2_X1 U7515 ( .A1(n8369), .A2(n8382), .ZN(n7581) );
  NAND2_X1 U7516 ( .A1(n6833), .A2(n8296), .ZN(n6487) );
  OR2_X1 U7517 ( .A1(n6484), .A2(n9139), .ZN(n6485) );
  XNOR2_X1 U7518 ( .A(n6485), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U7519 ( .A1(n6565), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6367), .B2(
        n10290), .ZN(n6486) );
  NAND2_X1 U7520 ( .A1(n6487), .A2(n6486), .ZN(n7795) );
  NAND2_X1 U7521 ( .A1(n8300), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6494) );
  INV_X1 U7522 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6488) );
  OR2_X1 U7523 ( .A1(n6378), .A2(n6488), .ZN(n6493) );
  NAND2_X1 U7524 ( .A1(n6489), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6490) );
  AND2_X1 U7525 ( .A1(n6500), .A2(n6490), .ZN(n7793) );
  OR2_X1 U7526 ( .A1(n6376), .A2(n7793), .ZN(n6492) );
  INV_X1 U7527 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8565) );
  OR2_X1 U7528 ( .A1(n6374), .A2(n8565), .ZN(n6491) );
  NAND4_X1 U7529 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n8532)
         );
  NAND2_X1 U7530 ( .A1(n7795), .A2(n8532), .ZN(n7622) );
  OR2_X1 U7531 ( .A1(n7795), .A2(n8532), .ZN(n7623) );
  NAND2_X1 U7532 ( .A1(n6915), .A2(n8296), .ZN(n6498) );
  XNOR2_X1 U7533 ( .A(n6496), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U7534 ( .A1(n6565), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6367), .B2(
        n10309), .ZN(n6497) );
  NAND2_X1 U7535 ( .A1(n6498), .A2(n6497), .ZN(n7720) );
  NAND2_X1 U7536 ( .A1(n8306), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6506) );
  INV_X1 U7537 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6499) );
  OR2_X1 U7538 ( .A1(n6677), .A2(n6499), .ZN(n6505) );
  NAND2_X1 U7539 ( .A1(n6500), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6501) );
  AND2_X1 U7540 ( .A1(n6513), .A2(n6501), .ZN(n7850) );
  OR2_X1 U7541 ( .A1(n6376), .A2(n7850), .ZN(n6504) );
  INV_X1 U7542 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6502) );
  OR2_X1 U7543 ( .A1(n6374), .A2(n6502), .ZN(n6503) );
  NAND4_X1 U7544 ( .A1(n6506), .A2(n6505), .A3(n6504), .A4(n6503), .ZN(n8531)
         );
  NOR2_X1 U7545 ( .A1(n7720), .A2(n8531), .ZN(n6508) );
  NAND2_X1 U7546 ( .A1(n7720), .A2(n8531), .ZN(n6507) );
  NAND2_X1 U7547 ( .A1(n7064), .A2(n8296), .ZN(n6511) );
  XNOR2_X1 U7548 ( .A(n6509), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U7549 ( .A1(n6565), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6367), .B2(
        n10324), .ZN(n6510) );
  NAND2_X1 U7550 ( .A1(n6511), .A2(n6510), .ZN(n8870) );
  NAND2_X1 U7551 ( .A1(n8306), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6519) );
  INV_X1 U7552 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6512) );
  OR2_X1 U7553 ( .A1(n6677), .A2(n6512), .ZN(n6518) );
  AND2_X1 U7554 ( .A1(n6513), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6514) );
  NOR2_X1 U7555 ( .A1(n6526), .A2(n6514), .ZN(n7825) );
  OR2_X1 U7556 ( .A1(n6376), .A2(n7825), .ZN(n6517) );
  INV_X1 U7557 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6515) );
  OR2_X1 U7558 ( .A1(n6374), .A2(n6515), .ZN(n6516) );
  NAND4_X1 U7559 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n8530)
         );
  AND2_X1 U7560 ( .A1(n8870), .A2(n8530), .ZN(n6520) );
  NAND2_X1 U7561 ( .A1(n7084), .A2(n8296), .ZN(n6523) );
  XNOR2_X1 U7562 ( .A(n6521), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U7563 ( .A1(n6565), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6367), .B2(
        n10341), .ZN(n6522) );
  NAND2_X1 U7564 ( .A1(n8306), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6533) );
  INV_X1 U7565 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6524) );
  OR2_X1 U7566 ( .A1(n6677), .A2(n6524), .ZN(n6532) );
  OR2_X1 U7567 ( .A1(n6526), .A2(n6525), .ZN(n6528) );
  AND2_X1 U7568 ( .A1(n6528), .A2(n6527), .ZN(n7875) );
  OR2_X1 U7569 ( .A1(n6376), .A2(n7875), .ZN(n6531) );
  INV_X1 U7570 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6529) );
  OR2_X1 U7571 ( .A1(n6374), .A2(n6529), .ZN(n6530) );
  NAND4_X1 U7572 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n8529)
         );
  NAND2_X1 U7573 ( .A1(n6534), .A2(n8529), .ZN(n6537) );
  INV_X1 U7574 ( .A(n7834), .ZN(n6535) );
  NAND2_X1 U7575 ( .A1(n6535), .A2(n7877), .ZN(n6536) );
  OR2_X1 U7576 ( .A1(n7934), .A2(n7994), .ZN(n8413) );
  NAND2_X1 U7577 ( .A1(n7934), .A2(n7994), .ZN(n8412) );
  INV_X1 U7578 ( .A(n8866), .ZN(n7999) );
  INV_X1 U7579 ( .A(n8527), .ZN(n8044) );
  NAND2_X1 U7580 ( .A1(n7316), .A2(n8296), .ZN(n6545) );
  INV_X1 U7581 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7582 ( .A1(n6539), .A2(n6538), .ZN(n6540) );
  NAND2_X1 U7583 ( .A1(n6540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6542) );
  INV_X1 U7584 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6541) );
  NAND2_X1 U7585 ( .A1(n6542), .A2(n6541), .ZN(n6553) );
  OR2_X1 U7586 ( .A1(n6542), .A2(n6541), .ZN(n6543) );
  AOI22_X1 U7587 ( .A1(n10387), .A2(n6367), .B1(n6565), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6544) );
  INV_X1 U7588 ( .A(n6376), .ZN(n6548) );
  OR2_X1 U7589 ( .A1(n6546), .A2(n8999), .ZN(n6547) );
  NAND2_X1 U7590 ( .A1(n6547), .A2(n6557), .ZN(n8071) );
  NAND2_X1 U7591 ( .A1(n6548), .A2(n8071), .ZN(n6552) );
  INV_X1 U7592 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9132) );
  OR2_X1 U7593 ( .A1(n6378), .A2(n9132), .ZN(n6551) );
  INV_X1 U7594 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8863) );
  OR2_X1 U7595 ( .A1(n6677), .A2(n8863), .ZN(n6550) );
  INV_X1 U7596 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8073) );
  OR2_X1 U7597 ( .A1(n6374), .A2(n8073), .ZN(n6549) );
  NAND2_X1 U7598 ( .A1(n8862), .A2(n8802), .ZN(n8421) );
  NAND2_X1 U7599 ( .A1(n8331), .A2(n8421), .ZN(n8067) );
  INV_X1 U7600 ( .A(n8862), .ZN(n8074) );
  NAND2_X1 U7601 ( .A1(n8066), .A2(n5474), .ZN(n8796) );
  NAND2_X1 U7602 ( .A1(n7374), .A2(n8296), .ZN(n6556) );
  NAND2_X1 U7603 ( .A1(n6553), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6554) );
  XNOR2_X1 U7604 ( .A(n6554), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U7605 ( .A1(n10405), .A2(n6367), .B1(n6565), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7606 ( .A1(n8306), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6561) );
  INV_X1 U7607 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8859) );
  OR2_X1 U7608 ( .A1(n6677), .A2(n8859), .ZN(n6560) );
  INV_X1 U7609 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10416) );
  OR2_X1 U7610 ( .A1(n6374), .A2(n10416), .ZN(n6559) );
  AOI21_X1 U7611 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n6557), .A(n6568), .ZN(
        n8803) );
  OR2_X1 U7612 ( .A1(n6376), .A2(n8803), .ZN(n6558) );
  NAND2_X1 U7613 ( .A1(n8858), .A2(n10643), .ZN(n8426) );
  NAND2_X1 U7614 ( .A1(n8425), .A2(n8426), .ZN(n8795) );
  NAND2_X1 U7615 ( .A1(n8796), .A2(n8795), .ZN(n8794) );
  INV_X1 U7616 ( .A(n8858), .ZN(n6562) );
  NAND2_X1 U7617 ( .A1(n8794), .A2(n5482), .ZN(n8783) );
  NAND2_X1 U7618 ( .A1(n7388), .A2(n8296), .ZN(n6567) );
  NAND2_X1 U7619 ( .A1(n6563), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6564) );
  XNOR2_X1 U7620 ( .A(n6564), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8617) );
  AOI22_X1 U7621 ( .A1(n6565), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6367), .B2(
        n8617), .ZN(n6566) );
  NAND2_X1 U7622 ( .A1(n8306), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6575) );
  INV_X1 U7623 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8855) );
  OR2_X1 U7624 ( .A1(n6677), .A2(n8855), .ZN(n6574) );
  INV_X1 U7625 ( .A(n6568), .ZN(n6569) );
  NAND2_X1 U7626 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n6569), .ZN(n6571) );
  AND2_X1 U7627 ( .A1(n6571), .A2(n6570), .ZN(n10654) );
  OR2_X1 U7628 ( .A1(n6376), .A2(n10654), .ZN(n6573) );
  INV_X1 U7629 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8787) );
  OR2_X1 U7630 ( .A1(n6374), .A2(n8787), .ZN(n6572) );
  NAND2_X1 U7631 ( .A1(n10649), .A2(n8222), .ZN(n8429) );
  NAND2_X1 U7632 ( .A1(n8428), .A2(n8429), .ZN(n8782) );
  NAND2_X1 U7633 ( .A1(n8783), .A2(n8782), .ZN(n8766) );
  NAND2_X1 U7634 ( .A1(n10649), .A2(n8798), .ZN(n8767) );
  NAND2_X1 U7635 ( .A1(n8851), .A2(n10642), .ZN(n8433) );
  NAND2_X1 U7636 ( .A1(n7649), .A2(n8296), .ZN(n6577) );
  OR2_X1 U7637 ( .A1(n8297), .A2(n7692), .ZN(n6576) );
  NAND2_X1 U7638 ( .A1(n8306), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6584) );
  INV_X1 U7639 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8848) );
  OR2_X1 U7640 ( .A1(n6677), .A2(n8848), .ZN(n6583) );
  NOR2_X2 U7641 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n6579), .ZN(n6588) );
  AND2_X1 U7642 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n6579), .ZN(n6580) );
  NOR2_X1 U7643 ( .A1(n6588), .A2(n6580), .ZN(n10658) );
  OR2_X1 U7644 ( .A1(n6376), .A2(n10658), .ZN(n6582) );
  INV_X1 U7645 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8757) );
  OR2_X1 U7646 ( .A1(n6374), .A2(n8757), .ZN(n6581) );
  NAND4_X1 U7647 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(n8770)
         );
  NAND2_X1 U7648 ( .A1(n8171), .A2(n8770), .ZN(n8437) );
  INV_X1 U7649 ( .A(n8770), .ZN(n8233) );
  NAND2_X1 U7650 ( .A1(n10668), .A2(n8233), .ZN(n8435) );
  NAND2_X1 U7651 ( .A1(n8437), .A2(n8435), .ZN(n8758) );
  INV_X1 U7652 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7754) );
  OR2_X1 U7653 ( .A1(n8297), .A2(n7754), .ZN(n6585) );
  NAND2_X1 U7654 ( .A1(n8306), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6593) );
  INV_X1 U7655 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6587) );
  OR2_X1 U7656 ( .A1(n6677), .A2(n6587), .ZN(n6592) );
  NOR2_X1 U7657 ( .A1(n6588), .A2(n8974), .ZN(n6589) );
  NOR2_X1 U7658 ( .A1(n6599), .A2(n6589), .ZN(n8746) );
  OR2_X1 U7659 ( .A1(n6376), .A2(n8746), .ZN(n6591) );
  INV_X1 U7660 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8747) );
  OR2_X1 U7661 ( .A1(n6374), .A2(n8747), .ZN(n6590) );
  NAND2_X1 U7662 ( .A1(n8749), .A2(n8259), .ZN(n8441) );
  NAND2_X1 U7663 ( .A1(n8438), .A2(n8441), .ZN(n8742) );
  INV_X1 U7664 ( .A(n8749), .ZN(n8845) );
  NAND2_X1 U7665 ( .A1(n7819), .A2(n8296), .ZN(n6597) );
  INV_X1 U7666 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7821) );
  OR2_X1 U7667 ( .A1(n8297), .A2(n7821), .ZN(n6596) );
  NAND2_X1 U7668 ( .A1(n8300), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6604) );
  INV_X1 U7669 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6598) );
  OR2_X1 U7670 ( .A1(n6378), .A2(n6598), .ZN(n6603) );
  NOR2_X1 U7671 ( .A1(n6599), .A2(n8258), .ZN(n6600) );
  NOR2_X1 U7672 ( .A1(n6607), .A2(n6600), .ZN(n8734) );
  OR2_X1 U7673 ( .A1(n6376), .A2(n8734), .ZN(n6602) );
  INV_X1 U7674 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8735) );
  OR2_X1 U7675 ( .A1(n6374), .A2(n8735), .ZN(n6601) );
  NAND2_X1 U7676 ( .A1(n8835), .A2(n8724), .ZN(n8439) );
  NAND2_X1 U7677 ( .A1(n7755), .A2(n8296), .ZN(n6606) );
  OR2_X1 U7678 ( .A1(n8297), .A2(n7752), .ZN(n6605) );
  NAND2_X1 U7679 ( .A1(n8306), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6612) );
  INV_X1 U7680 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8833) );
  OR2_X1 U7681 ( .A1(n6677), .A2(n8833), .ZN(n6611) );
  OR2_X1 U7682 ( .A1(n6607), .A2(n9075), .ZN(n6608) );
  AND2_X1 U7683 ( .A1(n6608), .A2(n6616), .ZN(n8726) );
  OR2_X1 U7684 ( .A1(n6376), .A2(n8726), .ZN(n6610) );
  INV_X1 U7685 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8727) );
  OR2_X1 U7686 ( .A1(n6374), .A2(n8727), .ZN(n6609) );
  NAND4_X1 U7687 ( .A1(n6612), .A2(n6611), .A3(n6610), .A4(n6609), .ZN(n8732)
         );
  NOR2_X1 U7688 ( .A1(n8832), .A2(n8732), .ZN(n6613) );
  INV_X1 U7689 ( .A(n8832), .ZN(n8218) );
  NAND2_X1 U7690 ( .A1(n7861), .A2(n8296), .ZN(n6615) );
  OR2_X1 U7691 ( .A1(n8297), .A2(n7921), .ZN(n6614) );
  NAND2_X1 U7692 ( .A1(n8300), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6621) );
  INV_X1 U7693 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8890) );
  OR2_X1 U7694 ( .A1(n6378), .A2(n8890), .ZN(n6620) );
  NOR2_X2 U7695 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n6616), .ZN(n6624) );
  AOI21_X1 U7696 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n6616), .A(n6624), .ZN(
        n8714) );
  OR2_X1 U7697 ( .A1(n6376), .A2(n8714), .ZN(n6619) );
  INV_X1 U7698 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6617) );
  OR2_X1 U7699 ( .A1(n6374), .A2(n6617), .ZN(n6618) );
  INV_X1 U7700 ( .A(n8725), .ZN(n8524) );
  NAND2_X1 U7701 ( .A1(n8715), .A2(n8725), .ZN(n8445) );
  NAND2_X1 U7702 ( .A1(n7894), .A2(n8296), .ZN(n6623) );
  INV_X1 U7703 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7908) );
  OR2_X1 U7704 ( .A1(n8297), .A2(n7908), .ZN(n6622) );
  NAND2_X1 U7705 ( .A1(n8306), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6630) );
  INV_X1 U7706 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8825) );
  OR2_X1 U7707 ( .A1(n6677), .A2(n8825), .ZN(n6629) );
  INV_X1 U7708 ( .A(n6624), .ZN(n6626) );
  NAND2_X1 U7709 ( .A1(n6624), .A2(n9092), .ZN(n6633) );
  INV_X1 U7710 ( .A(n6633), .ZN(n6625) );
  AOI21_X1 U7711 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n6626), .A(n6625), .ZN(
        n8700) );
  OR2_X1 U7712 ( .A1(n6376), .A2(n8700), .ZN(n6628) );
  INV_X1 U7713 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8707) );
  OR2_X1 U7714 ( .A1(n6374), .A2(n8707), .ZN(n6627) );
  OR2_X1 U7715 ( .A1(n8824), .A2(n8712), .ZN(n8460) );
  NAND2_X1 U7716 ( .A1(n8824), .A2(n8712), .ZN(n8459) );
  NAND2_X1 U7717 ( .A1(n8460), .A2(n8459), .ZN(n8703) );
  INV_X1 U7718 ( .A(n8824), .ZN(n8701) );
  NAND2_X1 U7719 ( .A1(n8015), .A2(n8296), .ZN(n6632) );
  OR2_X1 U7720 ( .A1(n8297), .A2(n8020), .ZN(n6631) );
  NAND2_X1 U7721 ( .A1(n8300), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6637) );
  INV_X1 U7722 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8882) );
  OR2_X1 U7723 ( .A1(n6378), .A2(n8882), .ZN(n6636) );
  NOR2_X2 U7724 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n6633), .ZN(n6644) );
  AOI21_X1 U7725 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n6633), .A(n6644), .ZN(
        n8691) );
  OR2_X1 U7726 ( .A1(n6376), .A2(n8691), .ZN(n6635) );
  INV_X1 U7727 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8692) );
  OR2_X1 U7728 ( .A1(n6374), .A2(n8692), .ZN(n6634) );
  NAND2_X1 U7729 ( .A1(n8820), .A2(n8522), .ZN(n6639) );
  OR2_X1 U7730 ( .A1(n8820), .A2(n8522), .ZN(n6638) );
  NAND2_X1 U7731 ( .A1(n8687), .A2(n8686), .ZN(n8685) );
  NAND2_X1 U7732 ( .A1(n8685), .A2(n6639), .ZN(n6761) );
  INV_X1 U7733 ( .A(n6761), .ZN(n6651) );
  NAND2_X1 U7734 ( .A1(n7983), .A2(n8296), .ZN(n6642) );
  OR2_X1 U7735 ( .A1(n8297), .A2(n6640), .ZN(n6641) );
  NAND2_X1 U7736 ( .A1(n8300), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6650) );
  INV_X1 U7737 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6643) );
  OR2_X1 U7738 ( .A1(n6378), .A2(n6643), .ZN(n6649) );
  NOR2_X2 U7739 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n6645), .ZN(n6661) );
  AND2_X1 U7740 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n6645), .ZN(n6646) );
  NOR2_X1 U7741 ( .A1(n6661), .A2(n6646), .ZN(n8675) );
  OR2_X1 U7742 ( .A1(n6376), .A2(n8675), .ZN(n6648) );
  INV_X1 U7743 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8676) );
  OR2_X1 U7744 ( .A1(n6374), .A2(n8676), .ZN(n6647) );
  NAND4_X1 U7745 ( .A1(n6650), .A2(n6649), .A3(n6648), .A4(n6647), .ZN(n8688)
         );
  NAND2_X1 U7746 ( .A1(n6653), .A2(n6652), .ZN(n6655) );
  NAND2_X1 U7747 ( .A1(n6655), .A2(n6654), .ZN(n8135) );
  MUX2_X1 U7748 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6656), .Z(n8136) );
  XNOR2_X1 U7749 ( .A(n8136), .B(n8137), .ZN(n8134) );
  XNOR2_X1 U7750 ( .A(n8135), .B(n8134), .ZN(n9149) );
  NAND2_X1 U7751 ( .A1(n9149), .A2(n8296), .ZN(n6658) );
  INV_X1 U7752 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9152) );
  OR2_X1 U7753 ( .A1(n8297), .A2(n9152), .ZN(n6657) );
  NAND2_X1 U7754 ( .A1(n8300), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6666) );
  INV_X1 U7755 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6659) );
  OR2_X1 U7756 ( .A1(n6378), .A2(n6659), .ZN(n6665) );
  INV_X1 U7757 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U7758 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  NOR2_X1 U7759 ( .A1(n8642), .A2(n6662), .ZN(n8667) );
  OR2_X1 U7760 ( .A1(n6376), .A2(n8667), .ZN(n6664) );
  INV_X1 U7761 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8668) );
  OR2_X1 U7762 ( .A1(n6374), .A2(n8668), .ZN(n6663) );
  AND4_X2 U7763 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n8326)
         );
  INV_X1 U7764 ( .A(n8653), .ZN(n8503) );
  XNOR2_X1 U7765 ( .A(n8654), .B(n8503), .ZN(n6683) );
  NAND2_X1 U7766 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  NAND2_X1 U7767 ( .A1(n6673), .A2(n6670), .ZN(n6671) );
  NAND2_X1 U7768 ( .A1(n6684), .A2(n8507), .ZN(n8320) );
  NAND2_X1 U7769 ( .A1(n6685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U7770 ( .A1(n8518), .A2(n8633), .ZN(n6749) );
  INV_X1 U7771 ( .A(n6845), .ZN(n8515) );
  NAND2_X1 U7772 ( .A1(n8515), .A2(n6859), .ZN(n6675) );
  NAND2_X1 U7773 ( .A1(n8643), .A2(n6675), .ZN(n7059) );
  INV_X1 U7774 ( .A(n7059), .ZN(n6990) );
  INV_X1 U7775 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6676) );
  OR2_X1 U7776 ( .A1(n6677), .A2(n6676), .ZN(n6681) );
  INV_X1 U7777 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8663) );
  OR2_X1 U7778 ( .A1(n6374), .A2(n8663), .ZN(n6680) );
  INV_X1 U7779 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6678) );
  OR2_X1 U7780 ( .A1(n6378), .A2(n6678), .ZN(n6679) );
  OAI22_X1 U7781 ( .A1(n8272), .A2(n8801), .B1(n8317), .B2(n8786), .ZN(n6682)
         );
  INV_X1 U7782 ( .A(n8672), .ZN(n8325) );
  INV_X1 U7783 ( .A(n8518), .ZN(n7820) );
  NAND2_X1 U7784 ( .A1(n8674), .A2(n5485), .ZN(n6757) );
  NAND2_X1 U7785 ( .A1(n6718), .A2(n6719), .ZN(n6688) );
  NAND2_X1 U7786 ( .A1(n6690), .A2(n6689), .ZN(n6695) );
  NAND2_X1 U7787 ( .A1(n6692), .A2(n4929), .ZN(n6693) );
  NAND2_X1 U7788 ( .A1(n7920), .A2(n8018), .ZN(n7043) );
  XNOR2_X2 U7789 ( .A(n6697), .B(n6696), .ZN(n6704) );
  XNOR2_X1 U7790 ( .A(n6698), .B(P2_B_REG_SCAN_IN), .ZN(n6699) );
  OR2_X1 U7791 ( .A1(n6703), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U7792 ( .A1(n6704), .A2(n8018), .ZN(n6705) );
  OR2_X1 U7793 ( .A1(n7002), .A2(n7000), .ZN(n6747) );
  NOR2_X1 U7794 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6710) );
  NOR4_X1 U7795 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6709) );
  NOR4_X1 U7796 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6708) );
  NOR4_X1 U7797 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6707) );
  NAND4_X1 U7798 ( .A1(n6710), .A2(n6709), .A3(n6708), .A4(n6707), .ZN(n6716)
         );
  NOR4_X1 U7799 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6714) );
  NOR4_X1 U7800 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6713) );
  NOR4_X1 U7801 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6712) );
  NOR4_X1 U7802 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6711) );
  NAND4_X1 U7803 ( .A1(n6714), .A2(n6713), .A3(n6712), .A4(n6711), .ZN(n6715)
         );
  NOR2_X1 U7804 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  OR2_X1 U7805 ( .A1(n6703), .A2(n6717), .ZN(n6751) );
  AND2_X1 U7806 ( .A1(n6973), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6720) );
  AND2_X1 U7807 ( .A1(n6751), .A2(n7008), .ZN(n6721) );
  NAND2_X1 U7808 ( .A1(n8518), .A2(n7611), .ZN(n6742) );
  OR2_X1 U7809 ( .A1(n6742), .A2(n8322), .ZN(n6722) );
  NAND2_X1 U7810 ( .A1(n8477), .A2(n6722), .ZN(n6999) );
  NAND2_X1 U7811 ( .A1(n7000), .A2(n6999), .ZN(n6725) );
  INV_X1 U7812 ( .A(n7047), .ZN(n6723) );
  OR2_X1 U7813 ( .A1(n8477), .A2(n6723), .ZN(n6974) );
  NAND2_X1 U7814 ( .A1(n6974), .A2(n6999), .ZN(n7001) );
  NAND2_X1 U7815 ( .A1(n7002), .A2(n7001), .ZN(n6724) );
  NAND2_X1 U7816 ( .A1(n8322), .A2(n8633), .ZN(n6992) );
  NAND3_X1 U7817 ( .A1(n6725), .A2(n6724), .A3(n7006), .ZN(n6726) );
  MUX2_X1 U7818 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n6757), .S(n8876), .Z(n6727)
         );
  INV_X1 U7819 ( .A(n6727), .ZN(n6746) );
  INV_X1 U7820 ( .A(n8338), .ZN(n8482) );
  NAND2_X1 U7821 ( .A1(n7099), .A2(n8482), .ZN(n6729) );
  INV_X1 U7822 ( .A(n10470), .ZN(n6728) );
  NAND2_X1 U7823 ( .A1(n7109), .A2(n6728), .ZN(n8346) );
  NAND2_X1 U7824 ( .A1(n7140), .A2(n7073), .ZN(n8351) );
  NAND2_X1 U7825 ( .A1(n8538), .A2(n7273), .ZN(n8356) );
  NAND2_X1 U7826 ( .A1(n7106), .A2(n8479), .ZN(n6730) );
  NAND2_X1 U7827 ( .A1(n6730), .A2(n8351), .ZN(n7137) );
  INV_X1 U7828 ( .A(n7115), .ZN(n7280) );
  NAND2_X1 U7829 ( .A1(n8537), .A2(n7280), .ZN(n8352) );
  NAND2_X1 U7830 ( .A1(n7137), .A2(n8352), .ZN(n6731) );
  INV_X1 U7831 ( .A(n8537), .ZN(n7182) );
  NAND2_X1 U7832 ( .A1(n7182), .A2(n7115), .ZN(n8357) );
  NOR2_X1 U7833 ( .A1(n8536), .A2(n7170), .ZN(n8354) );
  NAND2_X1 U7834 ( .A1(n8536), .A2(n7170), .ZN(n8361) );
  NAND2_X1 U7835 ( .A1(n7599), .A2(n7199), .ZN(n8362) );
  INV_X1 U7836 ( .A(n7199), .ZN(n7293) );
  NAND2_X1 U7837 ( .A1(n7293), .A2(n8535), .ZN(n8370) );
  NAND2_X1 U7838 ( .A1(n8362), .A2(n8370), .ZN(n8486) );
  AND2_X1 U7839 ( .A1(n8368), .A2(n7443), .ZN(n8376) );
  OR2_X1 U7840 ( .A1(n7795), .A2(n7841), .ZN(n8387) );
  AND2_X1 U7841 ( .A1(n8387), .A2(n8369), .ZN(n8375) );
  NAND2_X1 U7842 ( .A1(n7720), .A2(n7843), .ZN(n8389) );
  NAND2_X1 U7843 ( .A1(n7795), .A2(n7841), .ZN(n8381) );
  AND2_X1 U7844 ( .A1(n8389), .A2(n8381), .ZN(n8393) );
  OR2_X1 U7845 ( .A1(n7720), .A2(n7843), .ZN(n8391) );
  OR2_X1 U7846 ( .A1(n8870), .A2(n7868), .ZN(n8401) );
  NAND2_X1 U7847 ( .A1(n8870), .A2(n7868), .ZN(n8400) );
  NAND2_X1 U7848 ( .A1(n7822), .A2(n8398), .ZN(n6734) );
  INV_X1 U7849 ( .A(n8529), .ZN(n8405) );
  NAND2_X1 U7850 ( .A1(n7877), .A2(n8405), .ZN(n6735) );
  NAND2_X1 U7851 ( .A1(n8866), .A2(n8044), .ZN(n8417) );
  OR2_X1 U7852 ( .A1(n8866), .A2(n8044), .ZN(n8414) );
  NAND2_X1 U7853 ( .A1(n8072), .A2(n8499), .ZN(n6736) );
  NAND2_X1 U7854 ( .A1(n6736), .A2(n8331), .ZN(n8791) );
  NAND2_X1 U7855 ( .A1(n8791), .A2(n8792), .ZN(n6737) );
  NAND2_X1 U7856 ( .A1(n6737), .A2(n8425), .ZN(n8780) );
  NAND2_X1 U7857 ( .A1(n8780), .A2(n8781), .ZN(n6738) );
  NOR2_X1 U7858 ( .A1(n8832), .A2(n8713), .ZN(n8448) );
  NAND2_X1 U7859 ( .A1(n8832), .A2(n8713), .ZN(n8450) );
  OR2_X1 U7860 ( .A1(n8828), .A2(n8725), .ZN(n8456) );
  NAND2_X1 U7861 ( .A1(n8708), .A2(n8456), .ZN(n6739) );
  NAND2_X1 U7862 ( .A1(n8828), .A2(n8725), .ZN(n8455) );
  INV_X1 U7863 ( .A(n8703), .ZN(n8696) );
  OR2_X1 U7864 ( .A1(n8820), .A2(n8699), .ZN(n6740) );
  INV_X1 U7865 ( .A(n6740), .ZN(n6741) );
  NAND2_X1 U7866 ( .A1(n8680), .A2(n8272), .ZN(n8467) );
  XNOR2_X1 U7867 ( .A(n8294), .B(n8653), .ZN(n8669) );
  NAND2_X1 U7868 ( .A1(n7047), .A2(n6742), .ZN(n6743) );
  AND2_X1 U7869 ( .A1(n8844), .A2(n6743), .ZN(n6744) );
  OR2_X1 U7870 ( .A1(n6992), .A2(n8518), .ZN(n8814) );
  NAND2_X1 U7871 ( .A1(n6746), .A2(n6745), .ZN(P2_U3487) );
  INV_X1 U7872 ( .A(n6747), .ZN(n6748) );
  NAND2_X1 U7873 ( .A1(n6748), .A2(n6751), .ZN(n6993) );
  AND2_X1 U7874 ( .A1(n8477), .A2(n8844), .ZN(n6982) );
  INV_X1 U7875 ( .A(n6992), .ZN(n7179) );
  OR2_X1 U7876 ( .A1(n8844), .A2(n7179), .ZN(n10469) );
  INV_X1 U7877 ( .A(n10469), .ZN(n6750) );
  AOI21_X1 U7878 ( .B1(n6982), .B2(n6983), .A(n6750), .ZN(n6971) );
  NAND3_X1 U7879 ( .A1(n7002), .A2(n7000), .A3(n6751), .ZN(n6988) );
  OAI22_X1 U7880 ( .A1(n6993), .A2(n6983), .B1(n6971), .B2(n6988), .ZN(n6752)
         );
  NAND2_X1 U7881 ( .A1(n6752), .A2(n7008), .ZN(n6756) );
  INV_X1 U7882 ( .A(n6993), .ZN(n6754) );
  INV_X1 U7883 ( .A(n6753), .ZN(n7005) );
  AND2_X1 U7884 ( .A1(n7008), .A2(n7005), .ZN(n8516) );
  NAND2_X1 U7885 ( .A1(n6754), .A2(n8516), .ZN(n6755) );
  NAND2_X1 U7886 ( .A1(n6757), .A2(n10640), .ZN(n6759) );
  NAND2_X1 U7887 ( .A1(n10637), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6758) );
  INV_X1 U7888 ( .A(n8872), .ZN(n8839) );
  NAND2_X1 U7889 ( .A1(n5469), .A2(n6760), .ZN(P2_U3455) );
  OAI21_X1 U7890 ( .B1(n8211), .B2(n8844), .A(n8682), .ZN(n6771) );
  MUX2_X1 U7891 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n6771), .S(n8876), .Z(n6766)
         );
  INV_X1 U7892 ( .A(n6766), .ZN(n6770) );
  OAI21_X1 U7893 ( .B1(n6768), .B2(n8505), .A(n6767), .ZN(n6769) );
  INV_X1 U7894 ( .A(n6769), .ZN(n8677) );
  NAND2_X1 U7895 ( .A1(n6770), .A2(n5486), .ZN(P2_U3486) );
  MUX2_X1 U7896 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n6771), .S(n10640), .Z(n6772) );
  INV_X1 U7897 ( .A(n6772), .ZN(n6773) );
  NAND2_X1 U7898 ( .A1(n6773), .A2(n5475), .ZN(P2_U3454) );
  INV_X1 U7899 ( .A(n5680), .ZN(n6774) );
  INV_X4 U7900 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X4 U7901 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7902 ( .A1(n6775), .A2(n6776), .ZN(n6779) );
  INV_X1 U7903 ( .A(n6777), .ZN(n6778) );
  AOI211_X1 U7904 ( .C1(n6780), .C2(n6779), .A(n9268), .B(n6778), .ZN(n6784)
         );
  NOR2_X1 U7905 ( .A1(n9251), .A2(n7407), .ZN(n6783) );
  INV_X1 U7906 ( .A(n9572), .ZN(n7395) );
  INV_X1 U7907 ( .A(n9570), .ZN(n7562) );
  OAI22_X1 U7908 ( .A1(n9250), .A2(n7395), .B1(n7562), .B2(n9264), .ZN(n6782)
         );
  NAND2_X1 U7909 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10442) );
  OAI21_X1 U7910 ( .B1(n9243), .B2(n7430), .A(n10442), .ZN(n6781) );
  OR4_X1 U7911 ( .A1(n6784), .A2(n6783), .A3(n6782), .A4(n6781), .ZN(P1_U3230)
         );
  INV_X1 U7912 ( .A(n6847), .ZN(n6786) );
  NAND2_X1 U7913 ( .A1(n8473), .A2(n6973), .ZN(n6785) );
  NAND2_X1 U7914 ( .A1(n6786), .A2(n6785), .ZN(n6858) );
  OR2_X1 U7915 ( .A1(n6858), .A2(n6367), .ZN(n6787) );
  NAND2_X1 U7916 ( .A1(n6787), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X2 U7917 ( .A(n9148), .ZN(n9147) );
  OAI222_X1 U7918 ( .A1(n9153), .A2(n6788), .B1(n9147), .B2(n6799), .C1(
        P2_U3151), .C2(n6949), .ZN(P2_U3292) );
  OAI222_X1 U7919 ( .A1(n9153), .A2(n4993), .B1(n9147), .B2(n6795), .C1(
        P2_U3151), .C2(n10270), .ZN(P2_U3291) );
  INV_X1 U7920 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6838) );
  OAI222_X1 U7921 ( .A1(P2_U3151), .A2(n6878), .B1(n9147), .B2(n6792), .C1(
        n9153), .C2(n6838), .ZN(P2_U3294) );
  OAI222_X1 U7922 ( .A1(n9153), .A2(n6789), .B1(n9147), .B2(n6793), .C1(
        P2_U3151), .C2(n6863), .ZN(P2_U3293) );
  INV_X1 U7923 ( .A(n7008), .ZN(n6807) );
  NAND2_X1 U7924 ( .A1(n6807), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6790) );
  OAI21_X1 U7925 ( .B1(n7000), .B2(n6807), .A(n6790), .ZN(P2_U3377) );
  OAI222_X1 U7926 ( .A1(n9153), .A2(n6791), .B1(n9147), .B2(n6797), .C1(
        P2_U3151), .C2(n6961), .ZN(P2_U3290) );
  INV_X1 U7927 ( .A(n10025), .ZN(n7389) );
  INV_X1 U7928 ( .A(n7389), .ZN(n10018) );
  INV_X2 U7929 ( .A(n10015), .ZN(n8202) );
  OAI222_X1 U7930 ( .A1(n10018), .A2(n5497), .B1(n8202), .B2(n6792), .C1(
        P1_U3086), .C2(n7344), .ZN(P1_U3354) );
  OAI222_X1 U7931 ( .A1(n10018), .A2(n6794), .B1(n8202), .B2(n6793), .C1(
        P1_U3086), .C2(n9596), .ZN(P1_U3353) );
  OAI222_X1 U7932 ( .A1(n10018), .A2(n6796), .B1(n8202), .B2(n6795), .C1(
        P1_U3086), .C2(n10436), .ZN(P1_U3351) );
  OAI222_X1 U7933 ( .A1(n10018), .A2(n6798), .B1(n8202), .B2(n6797), .C1(
        P1_U3086), .C2(n10101), .ZN(P1_U3350) );
  OAI222_X1 U7934 ( .A1(n10018), .A2(n6800), .B1(n8202), .B2(n6799), .C1(
        P1_U3086), .C2(n7348), .ZN(P1_U3352) );
  NAND2_X1 U7935 ( .A1(n7132), .A2(P2_U3893), .ZN(n6801) );
  OAI21_X1 U7936 ( .B1(P2_U3893), .B2(n5676), .A(n6801), .ZN(P2_U3491) );
  OAI222_X1 U7937 ( .A1(n10018), .A2(n6802), .B1(n8202), .B2(n8133), .C1(
        P1_U3086), .C2(n10116), .ZN(P1_U3349) );
  INV_X1 U7938 ( .A(n6803), .ZN(n6805) );
  OAI222_X1 U7939 ( .A1(n10018), .A2(n6804), .B1(n8202), .B2(n6805), .C1(
        P1_U3086), .C2(n10131), .ZN(P1_U3348) );
  INV_X1 U7940 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6806) );
  OAI222_X1 U7941 ( .A1(n9153), .A2(n6806), .B1(n9147), .B2(n6805), .C1(
        P2_U3151), .C2(n7209), .ZN(P2_U3288) );
  INV_X1 U7942 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6808) );
  NOR2_X1 U7943 ( .A1(n6917), .A2(n6808), .ZN(P2_U3260) );
  INV_X1 U7944 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6809) );
  NOR2_X1 U7945 ( .A1(n6917), .A2(n6809), .ZN(P2_U3249) );
  INV_X1 U7946 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6810) );
  NOR2_X1 U7947 ( .A1(n6917), .A2(n6810), .ZN(P2_U3258) );
  INV_X1 U7948 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6811) );
  NOR2_X1 U7949 ( .A1(n6917), .A2(n6811), .ZN(P2_U3259) );
  INV_X1 U7950 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6812) );
  NOR2_X1 U7951 ( .A1(n6917), .A2(n6812), .ZN(P2_U3247) );
  INV_X1 U7952 ( .A(n6813), .ZN(n6815) );
  INV_X1 U7953 ( .A(n7361), .ZN(n10146) );
  OAI222_X1 U7954 ( .A1(n10018), .A2(n6814), .B1(n8202), .B2(n6815), .C1(
        P1_U3086), .C2(n10146), .ZN(P1_U3347) );
  INV_X1 U7955 ( .A(n7459), .ZN(n7452) );
  OAI222_X1 U7956 ( .A1(n9153), .A2(n6816), .B1(n9147), .B2(n6815), .C1(
        P2_U3151), .C2(n7452), .ZN(P2_U3287) );
  NAND4_X1 U7957 ( .A1(n8018), .A2(P2_STATE_REG_SCAN_IN), .A3(n7920), .A4(
        n6973), .ZN(n6817) );
  OAI21_X1 U7958 ( .B1(n6917), .B2(P2_D_REG_0__SCAN_IN), .A(n6817), .ZN(n6818)
         );
  INV_X1 U7959 ( .A(n6818), .ZN(P2_U3376) );
  NAND2_X1 U7960 ( .A1(n9471), .A2(n6821), .ZN(n6819) );
  INV_X1 U7961 ( .A(n7340), .ZN(n6822) );
  OR2_X1 U7962 ( .A1(n6821), .A2(P1_U3086), .ZN(n9551) );
  OR2_X1 U7963 ( .A1(n6824), .A2(n9546), .ZN(n7341) );
  NOR2_X1 U7964 ( .A1(n10439), .A2(P1_U3973), .ZN(P1_U3085) );
  AOI22_X1 U7965 ( .A1(n10027), .A2(n6827), .B1(n6826), .B2(n6825), .ZN(
        P1_U3439) );
  INV_X1 U7966 ( .A(n6828), .ZN(n6830) );
  INV_X1 U7967 ( .A(n7362), .ZN(n10259) );
  OAI222_X1 U7968 ( .A1(n10025), .A2(n6829), .B1(n8202), .B2(n6830), .C1(
        n10259), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U7969 ( .A(n8541), .ZN(n8584) );
  OAI222_X1 U7970 ( .A1(n9153), .A2(n6831), .B1(n9147), .B2(n6830), .C1(n8584), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X2 U7971 ( .A(P1_U3973), .ZN(n9590) );
  NAND2_X1 U7972 ( .A1(n9590), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n6832) );
  OAI21_X1 U7973 ( .B1(n9866), .B2(n9590), .A(n6832), .ZN(P1_U3572) );
  INV_X1 U7974 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6834) );
  INV_X1 U7975 ( .A(n6833), .ZN(n6835) );
  OAI222_X1 U7976 ( .A1(n9153), .A2(n6834), .B1(n9147), .B2(n6835), .C1(n8586), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U7977 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6836) );
  INV_X1 U7978 ( .A(n7363), .ZN(n10244) );
  OAI222_X1 U7979 ( .A1(n10025), .A2(n6836), .B1(n8202), .B2(n6835), .C1(
        n10244), .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U7980 ( .A1(n5284), .A2(P1_U3973), .ZN(n6837) );
  OAI21_X1 U7981 ( .B1(P1_U3973), .B2(n6838), .A(n6837), .ZN(P1_U3555) );
  INV_X1 U7982 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6876) );
  NOR2_X2 U7983 ( .A1(P2_U3150), .A2(n6847), .ZN(n10403) );
  INV_X1 U7984 ( .A(n10403), .ZN(n10288) );
  MUX2_X1 U7985 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8619), .Z(n6840) );
  XOR2_X1 U7986 ( .A(n6878), .B(n6840), .Z(n6877) );
  MUX2_X1 U7987 ( .A(n7011), .B(n6839), .S(n8619), .Z(n6890) );
  NAND2_X1 U7988 ( .A1(n6890), .A2(n4996), .ZN(n6889) );
  AOI22_X1 U7989 ( .A1(n6877), .A2(n6889), .B1(n6840), .B2(n6878), .ZN(n6898)
         );
  MUX2_X1 U7990 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8619), .Z(n6841) );
  XNOR2_X1 U7991 ( .A(n6841), .B(n6863), .ZN(n6897) );
  INV_X1 U7992 ( .A(n6863), .ZN(n6907) );
  INV_X1 U7993 ( .A(n6841), .ZN(n6842) );
  OAI22_X1 U7994 ( .A1(n6898), .A2(n6897), .B1(n6907), .B2(n6842), .ZN(n6946)
         );
  MUX2_X1 U7995 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8619), .Z(n6944) );
  XNOR2_X1 U7996 ( .A(n6944), .B(n6949), .ZN(n6945) );
  XNOR2_X1 U7997 ( .A(n6946), .B(n6945), .ZN(n6843) );
  NAND2_X1 U7998 ( .A1(n6843), .A2(n10412), .ZN(n6875) );
  INV_X1 U7999 ( .A(n6949), .ZN(n6873) );
  NOR2_X1 U8000 ( .A1(n8619), .A2(P2_U3151), .ZN(n7984) );
  NAND2_X1 U8001 ( .A1(n7984), .A2(n6845), .ZN(n6844) );
  OR2_X1 U8002 ( .A1(n6858), .A2(n6844), .ZN(n6849) );
  OR2_X1 U8003 ( .A1(n6845), .A2(P2_U3151), .ZN(n9150) );
  INV_X1 U8004 ( .A(n9150), .ZN(n6846) );
  NAND2_X1 U8005 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  INV_X1 U8006 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9077) );
  NOR2_X1 U8007 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9077), .ZN(n7072) );
  INV_X1 U8008 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6850) );
  MUX2_X1 U8009 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6850), .S(n6863), .Z(n6901)
         );
  NAND2_X1 U8010 ( .A1(n6860), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8011 ( .A1(n6878), .A2(n6855), .ZN(n6854) );
  INV_X1 U8012 ( .A(n4996), .ZN(n6851) );
  NAND2_X1 U8013 ( .A1(n6851), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6852) );
  OR2_X1 U8014 ( .A1(n6852), .A2(n6860), .ZN(n6853) );
  NAND2_X1 U8015 ( .A1(n6854), .A2(n6853), .ZN(n6882) );
  NAND2_X1 U8016 ( .A1(n6882), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8017 ( .A1(n6856), .A2(n6855), .ZN(n6900) );
  NAND2_X1 U8018 ( .A1(n6901), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U8019 ( .A1(n6863), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8020 ( .A1(n6899), .A2(n6857), .ZN(n6950) );
  XNOR2_X1 U8021 ( .A(n6950), .B(n6873), .ZN(n6948) );
  XOR2_X1 U8022 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6948), .Z(n6871) );
  NOR2_X1 U8023 ( .A1(n6858), .A2(n9150), .ZN(n6892) );
  NAND2_X1 U8024 ( .A1(n6892), .A2(n8619), .ZN(n8639) );
  INV_X1 U8025 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10476) );
  NOR2_X1 U8026 ( .A1(n7011), .A2(n4996), .ZN(n6861) );
  NAND2_X1 U8027 ( .A1(n6860), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6862) );
  OAI21_X1 U8028 ( .B1(n6878), .B2(n6861), .A(n6862), .ZN(n6881) );
  OR2_X1 U8029 ( .A1(n6881), .A2(n6358), .ZN(n6879) );
  NAND2_X1 U8030 ( .A1(n6879), .A2(n6862), .ZN(n6903) );
  NAND2_X1 U8031 ( .A1(n6863), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U8032 ( .A1(n6902), .A2(n6864), .ZN(n6865) );
  AND2_X1 U8033 ( .A1(n10273), .A2(n6866), .ZN(n6867) );
  INV_X1 U8034 ( .A(n6867), .ZN(n6869) );
  INV_X1 U8035 ( .A(n10275), .ZN(n6868) );
  AOI21_X1 U8036 ( .B1(n6390), .B2(n6869), .A(n6868), .ZN(n6870) );
  OAI22_X1 U8037 ( .A1(n6871), .A2(n8639), .B1(n10418), .B2(n6870), .ZN(n6872)
         );
  AOI211_X1 U8038 ( .C1(n6873), .C2(n10404), .A(n7072), .B(n6872), .ZN(n6874)
         );
  OAI211_X1 U8039 ( .C1(n6876), .C2(n10288), .A(n6875), .B(n6874), .ZN(
        P2_U3185) );
  XNOR2_X1 U8040 ( .A(n6877), .B(n6889), .ZN(n6888) );
  INV_X1 U8041 ( .A(n10404), .ZN(n10271) );
  OAI22_X1 U8042 ( .A1(n10271), .A2(n6878), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7093), .ZN(n6886) );
  INV_X1 U8043 ( .A(n6879), .ZN(n6880) );
  AOI21_X1 U8044 ( .B1(n6358), .B2(n6881), .A(n6880), .ZN(n6884) );
  XOR2_X1 U8045 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6882), .Z(n6883) );
  OAI22_X1 U8046 ( .A1(n6884), .A2(n10418), .B1(n8639), .B2(n6883), .ZN(n6885)
         );
  AOI211_X1 U8047 ( .C1(n10403), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6886), .B(
        n6885), .ZN(n6887) );
  OAI21_X1 U8048 ( .B1(n10282), .B2(n6888), .A(n6887), .ZN(P2_U3183) );
  INV_X1 U8049 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6896) );
  OAI21_X1 U8050 ( .B1(n4996), .B2(n6890), .A(n6889), .ZN(n6891) );
  OAI21_X1 U8051 ( .B1(n10412), .B2(n6892), .A(n6891), .ZN(n6893) );
  OAI21_X1 U8052 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6997), .A(n6893), .ZN(n6894) );
  AOI21_X1 U8053 ( .B1(n4996), .B2(n10404), .A(n6894), .ZN(n6895) );
  OAI21_X1 U8054 ( .B1(n10288), .B2(n6896), .A(n6895), .ZN(P2_U3182) );
  XNOR2_X1 U8055 ( .A(n6898), .B(n6897), .ZN(n6912) );
  OAI21_X1 U8056 ( .B1(n6901), .B2(n6900), .A(n6899), .ZN(n6906) );
  INV_X1 U8057 ( .A(n10418), .ZN(n8607) );
  OAI21_X1 U8058 ( .B1(n6904), .B2(n6903), .A(n6902), .ZN(n6905) );
  AOI22_X1 U8059 ( .A1(n10413), .A2(n6906), .B1(n8607), .B2(n6905), .ZN(n6909)
         );
  AOI22_X1 U8060 ( .A1(n10404), .A2(n6907), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6908) );
  NAND2_X1 U8061 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  AOI21_X1 U8062 ( .B1(n10403), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n6910), .ZN(
        n6911) );
  OAI21_X1 U8063 ( .B1(n10282), .B2(n6912), .A(n6911), .ZN(P2_U3184) );
  INV_X1 U8064 ( .A(n7051), .ZN(n7015) );
  NAND2_X1 U8065 ( .A1(n7132), .A2(n7015), .ZN(n8334) );
  NAND2_X1 U8066 ( .A1(n8340), .A2(n8334), .ZN(n8480) );
  OAI21_X1 U8067 ( .B1(n8793), .B2(n8872), .A(n8480), .ZN(n6913) );
  OR2_X1 U8068 ( .A1(n6371), .A2(n8786), .ZN(n7012) );
  OAI211_X1 U8069 ( .C1(n8844), .C2(n7015), .A(n6913), .B(n7012), .ZN(n8877)
         );
  NAND2_X1 U8070 ( .A1(n8877), .A2(n10640), .ZN(n6914) );
  OAI21_X1 U8071 ( .B1(n6349), .B2(n10640), .A(n6914), .ZN(P2_U3390) );
  INV_X1 U8072 ( .A(n6915), .ZN(n6969) );
  AOI22_X1 U8073 ( .A1(n10151), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7389), .ZN(n6916) );
  OAI21_X1 U8074 ( .B1(n6969), .B2(n8202), .A(n6916), .ZN(P1_U3344) );
  INV_X1 U8075 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U8076 ( .A1(n6943), .A2(n6918), .ZN(P2_U3253) );
  INV_X1 U8077 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6919) );
  NOR2_X1 U8078 ( .A1(n6943), .A2(n6919), .ZN(P2_U3235) );
  INV_X1 U8079 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6920) );
  NOR2_X1 U8080 ( .A1(n6943), .A2(n6920), .ZN(P2_U3254) );
  INV_X1 U8081 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U8082 ( .A1(n6943), .A2(n6921), .ZN(P2_U3248) );
  INV_X1 U8083 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6922) );
  NOR2_X1 U8084 ( .A1(n6943), .A2(n6922), .ZN(P2_U3236) );
  INV_X1 U8085 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8086 ( .A1(n6943), .A2(n6923), .ZN(P2_U3251) );
  INV_X1 U8087 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8088 ( .A1(n6943), .A2(n6924), .ZN(P2_U3250) );
  INV_X1 U8089 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U8090 ( .A1(n6943), .A2(n6925), .ZN(P2_U3262) );
  INV_X1 U8091 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U8092 ( .A1(n6943), .A2(n6926), .ZN(P2_U3243) );
  INV_X1 U8093 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6927) );
  NOR2_X1 U8094 ( .A1(n6943), .A2(n6927), .ZN(P2_U3242) );
  INV_X1 U8095 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6928) );
  NOR2_X1 U8096 ( .A1(n6943), .A2(n6928), .ZN(P2_U3252) );
  INV_X1 U8097 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6929) );
  NOR2_X1 U8098 ( .A1(n6943), .A2(n6929), .ZN(P2_U3240) );
  INV_X1 U8099 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6930) );
  NOR2_X1 U8100 ( .A1(n6943), .A2(n6930), .ZN(P2_U3255) );
  INV_X1 U8101 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6931) );
  NOR2_X1 U8102 ( .A1(n6943), .A2(n6931), .ZN(P2_U3241) );
  INV_X1 U8103 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6932) );
  NOR2_X1 U8104 ( .A1(n6943), .A2(n6932), .ZN(P2_U3261) );
  INV_X1 U8105 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6933) );
  NOR2_X1 U8106 ( .A1(n6943), .A2(n6933), .ZN(P2_U3239) );
  INV_X1 U8107 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6934) );
  NOR2_X1 U8108 ( .A1(n6943), .A2(n6934), .ZN(P2_U3238) );
  INV_X1 U8109 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6935) );
  NOR2_X1 U8110 ( .A1(n6943), .A2(n6935), .ZN(P2_U3263) );
  INV_X1 U8111 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6936) );
  NOR2_X1 U8112 ( .A1(n6943), .A2(n6936), .ZN(P2_U3237) );
  INV_X1 U8113 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6937) );
  NOR2_X1 U8114 ( .A1(n6943), .A2(n6937), .ZN(P2_U3257) );
  INV_X1 U8115 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6938) );
  NOR2_X1 U8116 ( .A1(n6943), .A2(n6938), .ZN(P2_U3256) );
  INV_X1 U8117 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6939) );
  NOR2_X1 U8118 ( .A1(n6943), .A2(n6939), .ZN(P2_U3244) );
  INV_X1 U8119 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6940) );
  NOR2_X1 U8120 ( .A1(n6943), .A2(n6940), .ZN(P2_U3234) );
  INV_X1 U8121 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6941) );
  NOR2_X1 U8122 ( .A1(n6943), .A2(n6941), .ZN(P2_U3246) );
  INV_X1 U8123 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6942) );
  NOR2_X1 U8124 ( .A1(n6943), .A2(n6942), .ZN(P2_U3245) );
  MUX2_X1 U8125 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8619), .Z(n7016) );
  XNOR2_X1 U8126 ( .A(n7016), .B(n6961), .ZN(n7018) );
  MUX2_X1 U8127 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8619), .Z(n6947) );
  OAI22_X1 U8128 ( .A1(n6946), .A2(n6945), .B1(n6944), .B2(n6949), .ZN(n10283)
         );
  XNOR2_X1 U8129 ( .A(n6947), .B(n10270), .ZN(n10284) );
  NOR2_X1 U8130 ( .A1(n10283), .A2(n10284), .ZN(n10281) );
  AOI21_X1 U8131 ( .B1(n6947), .B2(n10270), .A(n10281), .ZN(n7019) );
  XOR2_X1 U8132 ( .A(n7018), .B(n7019), .Z(n6967) );
  NAND2_X1 U8133 ( .A1(n6948), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8134 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  NAND2_X1 U8135 ( .A1(n6952), .A2(n6951), .ZN(n10266) );
  MUX2_X1 U8136 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6953), .S(n10270), .Z(n10267) );
  NAND2_X1 U8137 ( .A1(n10266), .A2(n10267), .ZN(n10265) );
  NAND2_X1 U8138 ( .A1(n10270), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8139 ( .A1(n10265), .A2(n6954), .ZN(n7024) );
  XNOR2_X1 U8140 ( .A(n7024), .B(n6961), .ZN(n7028) );
  XNOR2_X1 U8141 ( .A(n7028), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6955) );
  NOR2_X1 U8142 ( .A1(n8639), .A2(n6955), .ZN(n6966) );
  NAND2_X1 U8143 ( .A1(n10403), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6964) );
  XNOR2_X1 U8144 ( .A(n10270), .B(n6956), .ZN(n10272) );
  NAND2_X1 U8145 ( .A1(n10270), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8146 ( .A1(n6958), .A2(n6961), .ZN(n7032) );
  OAI21_X1 U8147 ( .B1(n4982), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7033), .ZN(
        n6960) );
  NAND2_X1 U8148 ( .A1(n8607), .A2(n6960), .ZN(n6963) );
  INV_X1 U8149 ( .A(n6961), .ZN(n7026) );
  AND2_X1 U8150 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7171) );
  AOI21_X1 U8151 ( .B1(n10404), .B2(n7026), .A(n7171), .ZN(n6962) );
  NAND3_X1 U8152 ( .A1(n6964), .A2(n6963), .A3(n6962), .ZN(n6965) );
  AOI211_X1 U8153 ( .C1(n6967), .C2(n10412), .A(n6966), .B(n6965), .ZN(n6968)
         );
  INV_X1 U8154 ( .A(n6968), .ZN(P2_U3187) );
  INV_X1 U8155 ( .A(n10309), .ZN(n8562) );
  OAI222_X1 U8156 ( .A1(n9153), .A2(n6970), .B1(n9147), .B2(n6969), .C1(
        P2_U3151), .C2(n8562), .ZN(P2_U3284) );
  INV_X1 U8157 ( .A(n6971), .ZN(n6972) );
  NAND2_X1 U8158 ( .A1(n6993), .A2(n6972), .ZN(n6978) );
  AND2_X1 U8159 ( .A1(n6974), .A2(n6973), .ZN(n6977) );
  INV_X1 U8160 ( .A(n6983), .ZN(n6975) );
  NAND2_X1 U8161 ( .A1(n6988), .A2(n6975), .ZN(n6985) );
  NAND4_X1 U8162 ( .A1(n6978), .A2(n6977), .A3(n6976), .A4(n6985), .ZN(n6979)
         );
  NAND2_X1 U8163 ( .A1(n6979), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6981) );
  NAND2_X1 U8164 ( .A1(n6988), .A2(n8516), .ZN(n6980) );
  INV_X1 U8165 ( .A(n10653), .ZN(n10670) );
  NOR2_X1 U8166 ( .A1(n10670), .A2(P2_U3151), .ZN(n7094) );
  INV_X1 U8167 ( .A(n6982), .ZN(n6984) );
  OAI21_X1 U8168 ( .B1(n6993), .B2(n6984), .A(n6983), .ZN(n6987) );
  AND2_X1 U8169 ( .A1(n6985), .A2(n7008), .ZN(n6986) );
  INV_X1 U8170 ( .A(n8516), .ZN(n6989) );
  OR2_X1 U8171 ( .A1(n6989), .A2(n6988), .ZN(n7060) );
  AOI22_X1 U8172 ( .A1(n10665), .A2(n8480), .B1(n10657), .B2(n6991), .ZN(n6996) );
  NAND2_X1 U8173 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  NAND2_X1 U8174 ( .A1(n10667), .A2(n7051), .ZN(n6995) );
  OAI211_X1 U8175 ( .C1(n7094), .C2(n6997), .A(n6996), .B(n6995), .ZN(P2_U3172) );
  INV_X1 U8176 ( .A(n6998), .ZN(n7004) );
  OAI22_X1 U8177 ( .A1(n7002), .A2(n7001), .B1(n7000), .B2(n6999), .ZN(n7003)
         );
  NAND2_X1 U8178 ( .A1(n7004), .A2(n7003), .ZN(n7010) );
  NOR3_X1 U8179 ( .A1(n7010), .A2(n8871), .A3(n7005), .ZN(n7009) );
  INV_X1 U8180 ( .A(n7006), .ZN(n7007) );
  AOI22_X1 U8181 ( .A1(n8480), .A2(n7009), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10572), .ZN(n7014) );
  MUX2_X1 U8182 ( .A(n7012), .B(n7011), .S(n10577), .Z(n7013) );
  OAI211_X1 U8183 ( .C1(n8649), .C2(n7015), .A(n7014), .B(n7013), .ZN(P2_U3233) );
  INV_X1 U8184 ( .A(n7016), .ZN(n7017) );
  OAI22_X1 U8185 ( .A1(n7019), .A2(n7018), .B1(n7026), .B2(n7017), .ZN(n7022)
         );
  MUX2_X1 U8186 ( .A(n7144), .B(n7023), .S(n8619), .Z(n7020) );
  NAND2_X1 U8187 ( .A1(n7020), .A2(n8131), .ZN(n7156) );
  OAI21_X1 U8188 ( .B1(n7020), .B2(n8131), .A(n7156), .ZN(n7021) );
  NOR2_X1 U8189 ( .A1(n7021), .A2(n7022), .ZN(n7154) );
  AOI21_X1 U8190 ( .B1(n7022), .B2(n7021), .A(n7154), .ZN(n7042) );
  MUX2_X1 U8191 ( .A(n7023), .B(P2_REG1_REG_6__SCAN_IN), .S(n8131), .Z(n7030)
         );
  INV_X1 U8192 ( .A(n7024), .ZN(n7025) );
  OAI22_X1 U8193 ( .A1(n7028), .A2(n7027), .B1(n7026), .B2(n7025), .ZN(n7029)
         );
  NAND2_X1 U8194 ( .A1(n7029), .A2(n7030), .ZN(n7143) );
  OAI21_X1 U8195 ( .B1(n7030), .B2(n7029), .A(n7143), .ZN(n7040) );
  MUX2_X1 U8196 ( .A(n7144), .B(P2_REG2_REG_6__SCAN_IN), .S(n8131), .Z(n7031)
         );
  NAND3_X1 U8197 ( .A1(n7033), .A2(n5365), .A3(n7032), .ZN(n7034) );
  AOI21_X1 U8198 ( .B1(n7146), .B2(n7034), .A(n10418), .ZN(n7039) );
  INV_X1 U8199 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7037) );
  INV_X1 U8200 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7035) );
  NOR2_X1 U8201 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7035), .ZN(n7202) );
  AOI21_X1 U8202 ( .B1(n10404), .B2(n8131), .A(n7202), .ZN(n7036) );
  OAI21_X1 U8203 ( .B1(n10288), .B2(n7037), .A(n7036), .ZN(n7038) );
  AOI211_X1 U8204 ( .C1(n10413), .C2(n7040), .A(n7039), .B(n7038), .ZN(n7041)
         );
  OAI21_X1 U8205 ( .B1(n7042), .B2(n10282), .A(n7041), .ZN(P2_U3188) );
  XNOR2_X1 U8206 ( .A(n7052), .B(n6371), .ZN(n7090) );
  MUX2_X1 U8207 ( .A(n7050), .B(n7132), .S(n7051), .Z(n7089) );
  NOR2_X1 U8208 ( .A1(n7090), .A2(n7089), .ZN(n7054) );
  INV_X1 U8209 ( .A(n7052), .ZN(n7053) );
  NOR2_X1 U8210 ( .A1(n7053), .A2(n6991), .ZN(n7056) );
  XNOR2_X1 U8211 ( .A(n7069), .B(n7109), .ZN(n7055) );
  OAI21_X2 U8212 ( .B1(n7054), .B2(n7056), .A(n7055), .ZN(n7068) );
  INV_X1 U8213 ( .A(n7068), .ZN(n7058) );
  NOR3_X1 U8214 ( .A1(n7091), .A2(n7056), .A3(n7055), .ZN(n7057) );
  OAI21_X1 U8215 ( .B1(n7058), .B2(n7057), .A(n10665), .ZN(n7063) );
  NOR2_X1 U8216 ( .A1(n10470), .A2(n8844), .ZN(n7104) );
  NOR2_X2 U8217 ( .A1(n7060), .A2(n7059), .ZN(n10655) );
  OAI22_X1 U8218 ( .A1(n10644), .A2(n6371), .B1(n7140), .B2(n10641), .ZN(n7061) );
  AOI21_X1 U8219 ( .B1(n7852), .B2(n7104), .A(n7061), .ZN(n7062) );
  OAI211_X1 U8220 ( .C1(n7094), .C2(n10467), .A(n7063), .B(n7062), .ZN(
        P2_U3177) );
  INV_X1 U8221 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7065) );
  INV_X1 U8222 ( .A(n7064), .ZN(n7066) );
  INV_X1 U8223 ( .A(n9634), .ZN(n7370) );
  OAI222_X1 U8224 ( .A1(n10025), .A2(n7065), .B1(n8202), .B2(n7066), .C1(n7370), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8225 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7067) );
  INV_X1 U8226 ( .A(n10324), .ZN(n8590) );
  OAI222_X1 U8227 ( .A1(n9153), .A2(n7067), .B1(n9147), .B2(n7066), .C1(n8590), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  XNOR2_X1 U8228 ( .A(n7050), .B(n7273), .ZN(n7113) );
  XNOR2_X1 U8229 ( .A(n7113), .B(n8538), .ZN(n7071) );
  AOI211_X1 U8230 ( .C1(n7071), .C2(n7070), .A(n8266), .B(n7114), .ZN(n7077)
         );
  AOI21_X1 U8231 ( .B1(n10657), .B2(n8537), .A(n7072), .ZN(n7075) );
  AND2_X1 U8232 ( .A1(n7073), .A2(n8871), .ZN(n7110) );
  AOI22_X1 U8233 ( .A1(n7852), .A2(n7110), .B1(n10655), .B2(n8539), .ZN(n7074)
         );
  OAI211_X1 U8234 ( .C1(n10653), .C2(P2_REG3_REG_3__SCAN_IN), .A(n7075), .B(
        n7074), .ZN(n7076) );
  OR2_X1 U8235 ( .A1(n7077), .A2(n7076), .ZN(P2_U3158) );
  OAI21_X1 U8236 ( .B1(n7080), .B2(n7079), .A(n7078), .ZN(n9586) );
  OR2_X1 U8237 ( .A1(n7081), .A2(P1_U3086), .ZN(n7267) );
  INV_X1 U8238 ( .A(n9404), .ZN(n10445) );
  OAI22_X1 U8239 ( .A1(n9264), .A2(n10446), .B1(n9243), .B2(n10445), .ZN(n7082) );
  AOI21_X1 U8240 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7267), .A(n7082), .ZN(
        n7083) );
  OAI21_X1 U8241 ( .B1(n9268), .B2(n9586), .A(n7083), .ZN(P1_U3232) );
  INV_X1 U8242 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7086) );
  INV_X1 U8243 ( .A(n7084), .ZN(n7087) );
  OAI222_X1 U8244 ( .A1(n10025), .A2(n7086), .B1(n8202), .B2(n7087), .C1(
        P1_U3086), .C2(n7085), .ZN(P1_U3342) );
  INV_X1 U8245 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7088) );
  INV_X1 U8246 ( .A(n10341), .ZN(n8559) );
  OAI222_X1 U8247 ( .A1(n9153), .A2(n7088), .B1(n9147), .B2(n7087), .C1(
        P2_U3151), .C2(n8559), .ZN(P2_U3282) );
  AOI21_X1 U8248 ( .B1(n7089), .B2(n7090), .A(n7091), .ZN(n7098) );
  NOR2_X1 U8249 ( .A1(n6372), .A2(n8844), .ZN(n7135) );
  OAI22_X1 U8250 ( .A1(n10644), .A2(n7092), .B1(n7109), .B2(n10641), .ZN(n7096) );
  NOR2_X1 U8251 ( .A1(n7094), .A2(n7093), .ZN(n7095) );
  AOI211_X1 U8252 ( .C1(n7852), .C2(n7135), .A(n7096), .B(n7095), .ZN(n7097)
         );
  OAI21_X1 U8253 ( .B1(n7098), .B2(n8266), .A(n7097), .ZN(P2_U3162) );
  XNOR2_X1 U8254 ( .A(n7099), .B(n8482), .ZN(n10473) );
  OAI21_X1 U8255 ( .B1(n8338), .B2(n7101), .A(n7100), .ZN(n7102) );
  AOI222_X1 U8256 ( .A1(n8793), .A2(n7102), .B1(n8538), .B2(n8797), .C1(n6991), 
        .C2(n8771), .ZN(n7103) );
  INV_X1 U8257 ( .A(n7103), .ZN(n10471) );
  AOI211_X1 U8258 ( .C1(n8872), .C2(n10473), .A(n7104), .B(n10471), .ZN(n10466) );
  NAND2_X1 U8259 ( .A1(n7621), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7105) );
  OAI21_X1 U8260 ( .B1(n10466), .B2(n7621), .A(n7105), .ZN(P2_U3461) );
  INV_X1 U8261 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7112) );
  XNOR2_X1 U8262 ( .A(n7106), .B(n8479), .ZN(n7277) );
  XNOR2_X1 U8263 ( .A(n7107), .B(n8479), .ZN(n7108) );
  OAI222_X1 U8264 ( .A1(n8786), .A2(n7182), .B1(n8801), .B2(n7109), .C1(n8723), 
        .C2(n7108), .ZN(n7274) );
  AOI211_X1 U8265 ( .C1(n7277), .C2(n8872), .A(n7110), .B(n7274), .ZN(n10485)
         );
  OR2_X1 U8266 ( .A1(n10485), .A2(n7621), .ZN(n7111) );
  OAI21_X1 U8267 ( .B1(n8876), .B2(n7112), .A(n7111), .ZN(P2_U3462) );
  INV_X4 U8268 ( .A(n7050), .ZN(n8194) );
  XNOR2_X1 U8269 ( .A(n8194), .B(n7115), .ZN(n7167) );
  XNOR2_X1 U8270 ( .A(n7167), .B(n7182), .ZN(n7116) );
  OAI21_X1 U8271 ( .B1(n7117), .B2(n7116), .A(n7169), .ZN(n7118) );
  NAND2_X1 U8272 ( .A1(n7118), .A2(n10665), .ZN(n7123) );
  NOR2_X1 U8273 ( .A1(n7280), .A2(n8844), .ZN(n7141) );
  INV_X1 U8274 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7119) );
  NOR2_X1 U8275 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7119), .ZN(n10268) );
  AOI21_X1 U8276 ( .B1(n10655), .B2(n8538), .A(n10268), .ZN(n7120) );
  OAI21_X1 U8277 ( .B1(n7289), .B2(n10641), .A(n7120), .ZN(n7121) );
  AOI21_X1 U8278 ( .B1(n7852), .B2(n7141), .A(n7121), .ZN(n7122) );
  OAI211_X1 U8279 ( .C1(n7279), .C2(n10653), .A(n7123), .B(n7122), .ZN(
        P2_U3170) );
  INV_X1 U8280 ( .A(n7124), .ZN(n7126) );
  INV_X1 U8281 ( .A(n10356), .ZN(n8594) );
  OAI222_X1 U8282 ( .A1(n9153), .A2(n7125), .B1(n9147), .B2(n7126), .C1(
        P2_U3151), .C2(n8594), .ZN(P2_U3281) );
  OAI222_X1 U8283 ( .A1(n10025), .A2(n7127), .B1(n8202), .B2(n7126), .C1(
        P1_U3086), .C2(n10177), .ZN(P1_U3341) );
  OAI21_X1 U8284 ( .B1(n5023), .B2(n5021), .A(n7129), .ZN(n7313) );
  OAI21_X1 U8285 ( .B1(n7131), .B2(n7128), .A(n7130), .ZN(n7133) );
  AOI222_X1 U8286 ( .A1(n8793), .A2(n7133), .B1(n8539), .B2(n8797), .C1(n7132), 
        .C2(n8771), .ZN(n7315) );
  INV_X1 U8287 ( .A(n7315), .ZN(n7134) );
  AOI211_X1 U8288 ( .C1(n8872), .C2(n7313), .A(n7135), .B(n7134), .ZN(n10463)
         );
  OR2_X1 U8289 ( .A1(n10463), .A2(n7621), .ZN(n7136) );
  OAI21_X1 U8290 ( .B1(n8876), .B2(n5036), .A(n7136), .ZN(P2_U3460) );
  AND2_X1 U8291 ( .A1(n8357), .A2(n8352), .ZN(n8484) );
  XNOR2_X1 U8292 ( .A(n7137), .B(n8484), .ZN(n7284) );
  XNOR2_X1 U8293 ( .A(n7138), .B(n8484), .ZN(n7139) );
  OAI222_X1 U8294 ( .A1(n8801), .A2(n7140), .B1(n8786), .B2(n7289), .C1(n8723), 
        .C2(n7139), .ZN(n7281) );
  AOI211_X1 U8295 ( .C1(n7284), .C2(n8872), .A(n7141), .B(n7281), .ZN(n10487)
         );
  OR2_X1 U8296 ( .A1(n10487), .A2(n7621), .ZN(n7142) );
  OAI21_X1 U8297 ( .B1(n8876), .B2(n6953), .A(n7142), .ZN(P2_U3463) );
  OAI21_X1 U8298 ( .B1(n8131), .B2(n7023), .A(n7143), .ZN(n7208) );
  XNOR2_X1 U8299 ( .A(n7208), .B(n7150), .ZN(n7210) );
  INV_X1 U8300 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7149) );
  XNOR2_X1 U8301 ( .A(n7210), .B(n7149), .ZN(n7166) );
  OR2_X1 U8302 ( .A1(n8131), .A2(n7144), .ZN(n7145) );
  NAND2_X1 U8303 ( .A1(n7147), .A2(n7209), .ZN(n7214) );
  OAI21_X1 U8304 ( .B1(n4980), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7215), .ZN(
        n7164) );
  NAND2_X1 U8305 ( .A1(n10403), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7162) );
  INV_X1 U8306 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9065) );
  NOR2_X1 U8307 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9065), .ZN(n7382) );
  AOI21_X1 U8308 ( .B1(n10404), .B2(n7150), .A(n7382), .ZN(n7161) );
  MUX2_X1 U8309 ( .A(n5374), .B(n7149), .S(n8619), .Z(n7151) );
  NAND2_X1 U8310 ( .A1(n7151), .A2(n7150), .ZN(n7217) );
  INV_X1 U8311 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U8312 ( .A1(n7152), .A2(n7209), .ZN(n7153) );
  AND2_X1 U8313 ( .A1(n7217), .A2(n7153), .ZN(n7158) );
  INV_X1 U8314 ( .A(n7154), .ZN(n7155) );
  NAND2_X1 U8315 ( .A1(n7156), .A2(n7155), .ZN(n7157) );
  NAND2_X1 U8316 ( .A1(n7158), .A2(n7157), .ZN(n7218) );
  OAI21_X1 U8317 ( .B1(n7158), .B2(n7157), .A(n7218), .ZN(n7159) );
  NAND2_X1 U8318 ( .A1(n7159), .A2(n10412), .ZN(n7160) );
  NAND3_X1 U8319 ( .A1(n7162), .A2(n7161), .A3(n7160), .ZN(n7163) );
  AOI21_X1 U8320 ( .B1(n7164), .B2(n8607), .A(n7163), .ZN(n7165) );
  OAI21_X1 U8321 ( .B1(n7166), .B2(n8639), .A(n7165), .ZN(P2_U3189) );
  OR2_X1 U8322 ( .A1(n7167), .A2(n8537), .ZN(n7168) );
  XNOR2_X1 U8323 ( .A(n8194), .B(n7188), .ZN(n7195) );
  XNOR2_X1 U8324 ( .A(n7195), .B(n7289), .ZN(n7197) );
  XOR2_X1 U8325 ( .A(n7198), .B(n7197), .Z(n7176) );
  NOR2_X1 U8326 ( .A1(n7170), .A2(n8844), .ZN(n7230) );
  AOI21_X1 U8327 ( .B1(n10657), .B2(n8535), .A(n7171), .ZN(n7173) );
  NAND2_X1 U8328 ( .A1(n10655), .A2(n8537), .ZN(n7172) );
  OAI211_X1 U8329 ( .C1(n10653), .C2(n7186), .A(n7173), .B(n7172), .ZN(n7174)
         );
  AOI21_X1 U8330 ( .B1(n7852), .B2(n7230), .A(n7174), .ZN(n7175) );
  OAI21_X1 U8331 ( .B1(n7176), .B2(n8266), .A(n7175), .ZN(P2_U3167) );
  INV_X1 U8332 ( .A(n8361), .ZN(n7177) );
  OR2_X1 U8333 ( .A1(n7177), .A2(n8354), .ZN(n7180) );
  XNOR2_X1 U8334 ( .A(n7178), .B(n7180), .ZN(n7228) );
  AND2_X1 U8335 ( .A1(n7179), .A2(n6684), .ZN(n7271) );
  NAND2_X1 U8336 ( .A1(n10575), .A2(n7271), .ZN(n10567) );
  INV_X1 U8337 ( .A(n7180), .ZN(n8483) );
  XNOR2_X1 U8338 ( .A(n7181), .B(n8483), .ZN(n7184) );
  OAI22_X1 U8339 ( .A1(n7182), .A2(n8801), .B1(n7599), .B2(n8786), .ZN(n7183)
         );
  AOI21_X1 U8340 ( .B1(n7184), .B2(n8793), .A(n7183), .ZN(n7185) );
  OAI21_X1 U8341 ( .B1(n7228), .B2(n8661), .A(n7185), .ZN(n7229) );
  NAND2_X1 U8342 ( .A1(n7229), .A2(n10575), .ZN(n7190) );
  OAI22_X1 U8343 ( .A1(n10575), .A2(n5364), .B1(n7186), .B2(n10468), .ZN(n7187) );
  AOI21_X1 U8344 ( .B1(n10568), .B2(n7188), .A(n7187), .ZN(n7189) );
  OAI211_X1 U8345 ( .C1(n7228), .C2(n10567), .A(n7190), .B(n7189), .ZN(
        P2_U3228) );
  INV_X1 U8346 ( .A(n7191), .ZN(n7193) );
  OAI222_X1 U8347 ( .A1(n10018), .A2(n7192), .B1(n8202), .B2(n7193), .C1(n9639), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8348 ( .A(n10372), .ZN(n8556) );
  OAI222_X1 U8349 ( .A1(n9153), .A2(n7194), .B1(n9147), .B2(n7193), .C1(n8556), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  INV_X1 U8350 ( .A(n7195), .ZN(n7196) );
  XNOR2_X1 U8351 ( .A(n8194), .B(n7199), .ZN(n7376) );
  XNOR2_X1 U8352 ( .A(n7376), .B(n7599), .ZN(n7200) );
  NAND2_X1 U8353 ( .A1(n7201), .A2(n7200), .ZN(n7378) );
  OAI211_X1 U8354 ( .C1(n7201), .C2(n7200), .A(n7378), .B(n10665), .ZN(n7207)
         );
  NOR2_X1 U8355 ( .A1(n7293), .A2(n8844), .ZN(n7290) );
  AOI21_X1 U8356 ( .B1(n10657), .B2(n8534), .A(n7202), .ZN(n7204) );
  NAND2_X1 U8357 ( .A1(n10655), .A2(n8536), .ZN(n7203) );
  OAI211_X1 U8358 ( .C1(n10653), .C2(n7294), .A(n7204), .B(n7203), .ZN(n7205)
         );
  AOI21_X1 U8359 ( .B1(n7852), .B2(n7290), .A(n7205), .ZN(n7206) );
  NAND2_X1 U8360 ( .A1(n7207), .A2(n7206), .ZN(P2_U3179) );
  MUX2_X1 U8361 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6460), .S(n7459), .Z(n7212)
         );
  AOI22_X1 U8362 ( .A1(n7210), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n7209), .B2(
        n7208), .ZN(n7211) );
  NOR2_X1 U8363 ( .A1(n7211), .A2(n7212), .ZN(n7451) );
  AOI21_X1 U8364 ( .B1(n7212), .B2(n7211), .A(n7451), .ZN(n7227) );
  MUX2_X1 U8365 ( .A(n7447), .B(P2_REG2_REG_8__SCAN_IN), .S(n7459), .Z(n7213)
         );
  NAND3_X1 U8366 ( .A1(n7215), .A2(n5373), .A3(n7214), .ZN(n7216) );
  AOI21_X1 U8367 ( .B1(n7449), .B2(n7216), .A(n10418), .ZN(n7225) );
  AND2_X1 U8368 ( .A1(n7218), .A2(n7217), .ZN(n7220) );
  MUX2_X1 U8369 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8619), .Z(n7456) );
  XNOR2_X1 U8370 ( .A(n7456), .B(n7452), .ZN(n7219) );
  NOR2_X1 U8371 ( .A1(n7220), .A2(n7219), .ZN(n7457) );
  AOI21_X1 U8372 ( .B1(n7220), .B2(n7219), .A(n7457), .ZN(n7223) );
  NOR2_X1 U8373 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9078), .ZN(n7555) );
  NOR2_X1 U8374 ( .A1(n10271), .A2(n7452), .ZN(n7221) );
  AOI211_X1 U8375 ( .C1(n10403), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7555), .B(
        n7221), .ZN(n7222) );
  OAI21_X1 U8376 ( .B1(n7223), .B2(n10282), .A(n7222), .ZN(n7224) );
  NOR2_X1 U8377 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  OAI21_X1 U8378 ( .B1(n7227), .B2(n8639), .A(n7226), .ZN(P2_U3190) );
  INV_X1 U8379 ( .A(n8814), .ZN(n7232) );
  INV_X1 U8380 ( .A(n7228), .ZN(n7231) );
  AOI211_X1 U8381 ( .C1(n7232), .C2(n7231), .A(n7230), .B(n7229), .ZN(n10500)
         );
  OR2_X1 U8382 ( .A1(n10500), .A2(n7621), .ZN(n7233) );
  OAI21_X1 U8383 ( .B1(n8876), .B2(n7027), .A(n7233), .ZN(P2_U3464) );
  NAND2_X1 U8384 ( .A1(n9404), .A2(n9574), .ZN(n7301) );
  NAND2_X1 U8385 ( .A1(n7415), .A2(n10446), .ZN(n7235) );
  INV_X1 U8386 ( .A(n9279), .ZN(n7480) );
  NAND2_X1 U8387 ( .A1(n7480), .A2(n7535), .ZN(n9485) );
  NAND2_X1 U8388 ( .A1(n9279), .A2(n9573), .ZN(n9289) );
  NAND2_X1 U8389 ( .A1(n9485), .A2(n9289), .ZN(n9399) );
  OAI21_X1 U8390 ( .B1(n7236), .B2(n9399), .A(n7394), .ZN(n7249) );
  INV_X1 U8391 ( .A(n10490), .ZN(n10625) );
  OAI211_X1 U8392 ( .C1(n5163), .C2(n9279), .A(n10527), .B(n7492), .ZN(n7477)
         );
  OAI21_X1 U8393 ( .B1(n9279), .B2(n10625), .A(n7477), .ZN(n7248) );
  INV_X1 U8394 ( .A(n7249), .ZN(n7483) );
  NAND2_X1 U8395 ( .A1(n7238), .A2(n7237), .ZN(n7239) );
  AND2_X1 U8396 ( .A1(n7239), .A2(n10444), .ZN(n7240) );
  INV_X1 U8397 ( .A(n9399), .ZN(n7243) );
  NOR2_X1 U8398 ( .A1(n10445), .A2(n9574), .ZN(n7305) );
  NAND2_X1 U8399 ( .A1(n10446), .A2(n7234), .ZN(n7241) );
  NAND2_X1 U8400 ( .A1(n7304), .A2(n7241), .ZN(n7242) );
  OAI21_X1 U8401 ( .B1(n7243), .B2(n7242), .A(n7400), .ZN(n7246) );
  NAND2_X1 U8402 ( .A1(n6236), .A2(n7244), .ZN(n9396) );
  NAND2_X1 U8403 ( .A1(n9550), .A2(n9778), .ZN(n9435) );
  OAI22_X1 U8404 ( .A1(n7395), .A2(n10531), .B1(n10446), .B2(n10533), .ZN(
        n7245) );
  AOI21_X1 U8405 ( .B1(n7246), .B2(n9892), .A(n7245), .ZN(n7247) );
  OAI21_X1 U8406 ( .B1(n7483), .B2(n8025), .A(n7247), .ZN(n7474) );
  AOI211_X1 U8407 ( .C1(n10609), .C2(n7249), .A(n7248), .B(n7474), .ZN(n7322)
         );
  NOR2_X1 U8408 ( .A1(n7250), .A2(P1_U3086), .ZN(n7252) );
  AND2_X1 U8409 ( .A1(n7254), .A2(n7253), .ZN(n7321) );
  NAND2_X1 U8410 ( .A1(n10630), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7255) );
  OAI21_X1 U8411 ( .B1(n7322), .B2(n10630), .A(n7255), .ZN(P1_U3524) );
  INV_X1 U8412 ( .A(n7256), .ZN(n7261) );
  AOI21_X1 U8413 ( .B1(n7260), .B2(n7258), .A(n7257), .ZN(n7259) );
  AOI21_X1 U8414 ( .B1(n7261), .B2(n7260), .A(n7259), .ZN(n7264) );
  AOI22_X1 U8415 ( .A1(n7234), .A2(n9266), .B1(n9261), .B2(n9574), .ZN(n7263)
         );
  AOI22_X1 U8416 ( .A1(n9213), .A2(n9573), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7267), .ZN(n7262) );
  OAI211_X1 U8417 ( .C1(n7264), .C2(n9268), .A(n7263), .B(n7262), .ZN(P1_U3222) );
  XOR2_X1 U8418 ( .A(n7266), .B(n7265), .Z(n7270) );
  AOI22_X1 U8419 ( .A1(n7480), .A2(n9266), .B1(n9261), .B2(n5284), .ZN(n7269)
         );
  AOI22_X1 U8420 ( .A1(n9213), .A2(n9572), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7267), .ZN(n7268) );
  OAI211_X1 U8421 ( .C1(n7270), .C2(n9268), .A(n7269), .B(n7268), .ZN(P1_U3237) );
  INV_X1 U8422 ( .A(n7271), .ZN(n7272) );
  NAND2_X1 U8423 ( .A1(n8661), .A2(n7272), .ZN(n10474) );
  INV_X1 U8424 ( .A(n8807), .ZN(n8752) );
  OAI22_X1 U8425 ( .A1(n8649), .A2(n7273), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10468), .ZN(n7276) );
  MUX2_X1 U8426 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7274), .S(n10575), .Z(n7275)
         );
  AOI211_X1 U8427 ( .C1(n8752), .C2(n7277), .A(n7276), .B(n7275), .ZN(n7278)
         );
  INV_X1 U8428 ( .A(n7278), .ZN(P2_U3230) );
  OAI22_X1 U8429 ( .A1(n8649), .A2(n7280), .B1(n7279), .B2(n10468), .ZN(n7283)
         );
  MUX2_X1 U8430 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7281), .S(n10575), .Z(n7282)
         );
  AOI211_X1 U8431 ( .C1(n8752), .C2(n7284), .A(n7283), .B(n7282), .ZN(n7285)
         );
  INV_X1 U8432 ( .A(n7285), .ZN(P2_U3229) );
  XNOR2_X1 U8433 ( .A(n7286), .B(n8486), .ZN(n7297) );
  XOR2_X1 U8434 ( .A(n7287), .B(n8486), .Z(n7288) );
  OAI222_X1 U8435 ( .A1(n8786), .A2(n7554), .B1(n8801), .B2(n7289), .C1(n8723), 
        .C2(n7288), .ZN(n7292) );
  AOI211_X1 U8436 ( .C1(n8872), .C2(n7297), .A(n7290), .B(n7292), .ZN(n10510)
         );
  NAND2_X1 U8437 ( .A1(n7621), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7291) );
  OAI21_X1 U8438 ( .B1(n10510), .B2(n7621), .A(n7291), .ZN(P2_U3465) );
  INV_X1 U8439 ( .A(n7292), .ZN(n7299) );
  NOR2_X1 U8440 ( .A1(n8649), .A2(n7293), .ZN(n7296) );
  OAI22_X1 U8441 ( .A1(n10575), .A2(n7144), .B1(n7294), .B2(n10468), .ZN(n7295) );
  AOI211_X1 U8442 ( .C1(n7297), .C2(n8752), .A(n7296), .B(n7295), .ZN(n7298)
         );
  OAI21_X1 U8443 ( .B1(n7299), .B2(n10577), .A(n7298), .ZN(P2_U3227) );
  OAI21_X1 U8444 ( .B1(n7302), .B2(n7301), .A(n7300), .ZN(n7417) );
  NAND2_X1 U8445 ( .A1(n7234), .A2(n9404), .ZN(n7411) );
  NAND3_X1 U8446 ( .A1(n7412), .A2(n10527), .A3(n7411), .ZN(n7303) );
  OAI21_X1 U8447 ( .B1(n7415), .B2(n10625), .A(n7303), .ZN(n7308) );
  OAI21_X1 U8448 ( .B1(n9406), .B2(n7305), .A(n7304), .ZN(n7306) );
  AOI222_X1 U8449 ( .A1(n9892), .A2(n7306), .B1(n9573), .B2(n9887), .C1(n9574), 
        .C2(n9889), .ZN(n7419) );
  INV_X1 U8450 ( .A(n7419), .ZN(n7307) );
  AOI211_X1 U8451 ( .C1(n10628), .C2(n7417), .A(n7308), .B(n7307), .ZN(n10465)
         );
  NAND2_X1 U8452 ( .A1(n10630), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7309) );
  OAI21_X1 U8453 ( .B1(n10465), .B2(n10630), .A(n7309), .ZN(P1_U3523) );
  AOI22_X1 U8454 ( .A1(n10568), .A2(n7310), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10572), .ZN(n7311) );
  OAI21_X1 U8455 ( .B1(n6358), .B2(n10575), .A(n7311), .ZN(n7312) );
  AOI21_X1 U8456 ( .B1(n7313), .B2(n8752), .A(n7312), .ZN(n7314) );
  OAI21_X1 U8457 ( .B1(n7315), .B2(n10577), .A(n7314), .ZN(P2_U3232) );
  INV_X1 U8458 ( .A(n7316), .ZN(n7318) );
  INV_X1 U8459 ( .A(n9656), .ZN(n9632) );
  OAI222_X1 U8460 ( .A1(n10018), .A2(n7317), .B1(n8202), .B2(n7318), .C1(
        P1_U3086), .C2(n9632), .ZN(P1_U3339) );
  INV_X1 U8461 ( .A(n10387), .ZN(n8598) );
  OAI222_X1 U8462 ( .A1(n9153), .A2(n7319), .B1(n9147), .B2(n7318), .C1(
        P2_U3151), .C2(n8598), .ZN(P2_U3279) );
  INV_X1 U8463 ( .A(n7320), .ZN(n7398) );
  INV_X1 U8464 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7324) );
  OR2_X1 U8465 ( .A1(n7322), .A2(n10633), .ZN(n7323) );
  OAI21_X1 U8466 ( .B1(n10636), .B2(n7324), .A(n7323), .ZN(P1_U3459) );
  NAND2_X1 U8467 ( .A1(n9590), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7325) );
  OAI21_X1 U8468 ( .B1(n9741), .B2(n9590), .A(n7325), .ZN(P1_U3582) );
  NOR2_X1 U8469 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9634), .ZN(n7326) );
  AOI21_X1 U8470 ( .B1(n9634), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7326), .ZN(
        n7339) );
  INV_X1 U8471 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7327) );
  AOI22_X1 U8472 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10244), .B1(n7363), .B2(
        n7327), .ZN(n10236) );
  NOR2_X1 U8473 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n7362), .ZN(n7328) );
  AOI21_X1 U8474 ( .B1(n7362), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7328), .ZN(
        n10251) );
  XNOR2_X1 U8475 ( .A(n9596), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9600) );
  XNOR2_X1 U8476 ( .A(n7344), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9577) );
  AND2_X1 U8477 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9576) );
  NAND2_X1 U8478 ( .A1(n9577), .A2(n9576), .ZN(n9575) );
  INV_X1 U8479 ( .A(n7344), .ZN(n9581) );
  NAND2_X1 U8480 ( .A1(n9581), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U8481 ( .A1(n9575), .A2(n7329), .ZN(n9599) );
  NAND2_X1 U8482 ( .A1(n9600), .A2(n9599), .ZN(n9598) );
  INV_X1 U8483 ( .A(n9596), .ZN(n7346) );
  NAND2_X1 U8484 ( .A1(n7346), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7330) );
  NAND2_X1 U8485 ( .A1(n9598), .A2(n7330), .ZN(n9615) );
  XNOR2_X1 U8486 ( .A(n7348), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U8487 ( .A1(n9615), .A2(n9616), .ZN(n9614) );
  INV_X1 U8488 ( .A(n7348), .ZN(n9610) );
  NAND2_X1 U8489 ( .A1(n9610), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7331) );
  NAND2_X1 U8490 ( .A1(n9614), .A2(n7331), .ZN(n10428) );
  INV_X1 U8491 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7332) );
  MUX2_X1 U8492 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7332), .S(n7350), .Z(n10429)
         );
  AND2_X1 U8493 ( .A1(n10428), .A2(n10429), .ZN(n10425) );
  AOI21_X1 U8494 ( .B1(n7350), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10425), .ZN(
        n10092) );
  NAND2_X1 U8495 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7353), .ZN(n7333) );
  OAI21_X1 U8496 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7353), .A(n7333), .ZN(
        n10093) );
  NOR2_X1 U8497 ( .A1(n10092), .A2(n10093), .ZN(n10091) );
  AOI21_X1 U8498 ( .B1(n7353), .B2(P1_REG2_REG_5__SCAN_IN), .A(n10091), .ZN(
        n10107) );
  NAND2_X1 U8499 ( .A1(n7356), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7334) );
  OAI21_X1 U8500 ( .B1(n7356), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7334), .ZN(
        n10108) );
  NOR2_X1 U8501 ( .A1(n10107), .A2(n10108), .ZN(n10106) );
  AOI21_X1 U8502 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7356), .A(n10106), .ZN(
        n10122) );
  NAND2_X1 U8503 ( .A1(n7359), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U8504 ( .B1(n7359), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7335), .ZN(
        n10123) );
  NOR2_X1 U8505 ( .A1(n10122), .A2(n10123), .ZN(n10121) );
  AOI21_X1 U8506 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7359), .A(n10121), .ZN(
        n10137) );
  NAND2_X1 U8507 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7361), .ZN(n7336) );
  OAI21_X1 U8508 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7361), .A(n7336), .ZN(
        n10138) );
  NOR2_X1 U8509 ( .A1(n10137), .A2(n10138), .ZN(n10136) );
  AOI21_X1 U8510 ( .B1(n7361), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10136), .ZN(
        n10250) );
  NAND2_X1 U8511 ( .A1(n10251), .A2(n10250), .ZN(n10249) );
  OAI21_X1 U8512 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7362), .A(n10249), .ZN(
        n10235) );
  NOR2_X1 U8513 ( .A1(n10236), .A2(n10235), .ZN(n10234) );
  AOI21_X1 U8514 ( .B1(n7363), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10234), .ZN(
        n10153) );
  NAND2_X1 U8515 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n10151), .ZN(n7337) );
  OAI21_X1 U8516 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10151), .A(n7337), .ZN(
        n10154) );
  NOR2_X1 U8517 ( .A1(n10153), .A2(n10154), .ZN(n10152) );
  AOI21_X1 U8518 ( .B1(n10151), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10152), .ZN(
        n7338) );
  NAND2_X1 U8519 ( .A1(n7339), .A2(n7338), .ZN(n9633) );
  OAI21_X1 U8520 ( .B1(n7339), .B2(n7338), .A(n9633), .ZN(n7372) );
  NAND2_X1 U8521 ( .A1(n7341), .A2(n7340), .ZN(n10090) );
  OR2_X1 U8522 ( .A1(n4908), .A2(n8162), .ZN(n10085) );
  OR2_X1 U8523 ( .A1(n10090), .A2(n10085), .ZN(n10222) );
  OR2_X1 U8524 ( .A1(n10090), .A2(n9588), .ZN(n10437) );
  INV_X1 U8525 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U8526 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9634), .B1(n7370), .B2(
        n10620), .ZN(n7366) );
  INV_X1 U8527 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7342) );
  MUX2_X1 U8528 ( .A(n7342), .B(P1_REG1_REG_10__SCAN_IN), .S(n7363), .Z(n10240) );
  INV_X1 U8529 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7343) );
  MUX2_X1 U8530 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7343), .S(n7362), .Z(n10255)
         );
  XNOR2_X1 U8531 ( .A(n9596), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9603) );
  XNOR2_X1 U8532 ( .A(n7344), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9580) );
  AND2_X1 U8533 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9579) );
  NAND2_X1 U8534 ( .A1(n9580), .A2(n9579), .ZN(n9578) );
  NAND2_X1 U8535 ( .A1(n9581), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7345) );
  NAND2_X1 U8536 ( .A1(n9578), .A2(n7345), .ZN(n9602) );
  NAND2_X1 U8537 ( .A1(n9603), .A2(n9602), .ZN(n9601) );
  NAND2_X1 U8538 ( .A1(n7346), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U8539 ( .A1(n9601), .A2(n7347), .ZN(n9612) );
  XNOR2_X1 U8540 ( .A(n7348), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U8541 ( .A1(n9612), .A2(n9613), .ZN(n9611) );
  NAND2_X1 U8542 ( .A1(n9610), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7349) );
  NAND2_X1 U8543 ( .A1(n9611), .A2(n7349), .ZN(n10432) );
  INV_X1 U8544 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10496) );
  MUX2_X1 U8545 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10496), .S(n7350), .Z(n10433) );
  NAND2_X1 U8546 ( .A1(n10432), .A2(n10433), .ZN(n10430) );
  NAND2_X1 U8547 ( .A1(n7350), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7351) );
  AND2_X1 U8548 ( .A1(n10430), .A2(n7351), .ZN(n10097) );
  NAND2_X1 U8549 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7353), .ZN(n7352) );
  OAI21_X1 U8550 ( .B1(n7353), .B2(P1_REG1_REG_5__SCAN_IN), .A(n7352), .ZN(
        n10096) );
  NOR2_X1 U8551 ( .A1(n10097), .A2(n10096), .ZN(n10095) );
  AOI21_X1 U8552 ( .B1(n7353), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10095), .ZN(
        n10111) );
  OR2_X1 U8553 ( .A1(n7356), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U8554 ( .A1(n7356), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7354) );
  NAND2_X1 U8555 ( .A1(n7355), .A2(n7354), .ZN(n10112) );
  NOR2_X1 U8556 ( .A1(n10111), .A2(n10112), .ZN(n10110) );
  AOI21_X1 U8557 ( .B1(n7356), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10110), .ZN(
        n10126) );
  OR2_X1 U8558 ( .A1(n7359), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U8559 ( .A1(n7359), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U8560 ( .A1(n7358), .A2(n7357), .ZN(n10127) );
  NOR2_X1 U8561 ( .A1(n10126), .A2(n10127), .ZN(n10125) );
  AOI21_X1 U8562 ( .B1(n7359), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10125), .ZN(
        n10141) );
  INV_X1 U8563 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7360) );
  MUX2_X1 U8564 ( .A(n7360), .B(P1_REG1_REG_8__SCAN_IN), .S(n7361), .Z(n10142)
         );
  NOR2_X1 U8565 ( .A1(n10141), .A2(n10142), .ZN(n10140) );
  AOI21_X1 U8566 ( .B1(n7361), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10140), .ZN(
        n10254) );
  NAND2_X1 U8567 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  OAI21_X1 U8568 ( .B1(n7362), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10253), .ZN(
        n10239) );
  NOR2_X1 U8569 ( .A1(n10240), .A2(n10239), .ZN(n10238) );
  AOI21_X1 U8570 ( .B1(n7363), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10238), .ZN(
        n10157) );
  INV_X1 U8571 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7364) );
  MUX2_X1 U8572 ( .A(n7364), .B(P1_REG1_REG_11__SCAN_IN), .S(n10151), .Z(
        n10158) );
  NOR2_X1 U8573 ( .A1(n10157), .A2(n10158), .ZN(n10156) );
  AOI21_X1 U8574 ( .B1(n10151), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10156), .ZN(
        n7365) );
  NAND2_X1 U8575 ( .A1(n7366), .A2(n7365), .ZN(n9621) );
  OAI21_X1 U8576 ( .B1(n7366), .B2(n7365), .A(n9621), .ZN(n7367) );
  INV_X1 U8577 ( .A(n8162), .ZN(n9587) );
  NAND2_X1 U8578 ( .A1(n7367), .A2(n10431), .ZN(n7369) );
  AND2_X1 U8579 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7916) );
  AOI21_X1 U8580 ( .B1(n10439), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7916), .ZN(
        n7368) );
  OAI211_X1 U8581 ( .C1(n10437), .C2(n7370), .A(n7369), .B(n7368), .ZN(n7371)
         );
  AOI21_X1 U8582 ( .B1(n7372), .B2(n10427), .A(n7371), .ZN(n7373) );
  INV_X1 U8583 ( .A(n7373), .ZN(P1_U3255) );
  INV_X1 U8584 ( .A(n7374), .ZN(n7391) );
  AOI22_X1 U8585 ( .A1(n10201), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7389), .ZN(n7375) );
  OAI21_X1 U8586 ( .B1(n7391), .B2(n8202), .A(n7375), .ZN(P1_U3338) );
  XNOR2_X1 U8587 ( .A(n8194), .B(n10569), .ZN(n7551) );
  XNOR2_X1 U8588 ( .A(n7551), .B(n8534), .ZN(n7380) );
  AOI21_X1 U8589 ( .B1(n7380), .B2(n7379), .A(n7552), .ZN(n7387) );
  INV_X1 U8590 ( .A(n10569), .ZN(n7381) );
  NOR2_X1 U8591 ( .A1(n7381), .A2(n8844), .ZN(n7600) );
  AOI21_X1 U8592 ( .B1(n10657), .B2(n8533), .A(n7382), .ZN(n7384) );
  NAND2_X1 U8593 ( .A1(n10655), .A2(n8535), .ZN(n7383) );
  OAI211_X1 U8594 ( .C1(n10653), .C2(n10566), .A(n7384), .B(n7383), .ZN(n7385)
         );
  AOI21_X1 U8595 ( .B1(n7852), .B2(n7600), .A(n7385), .ZN(n7386) );
  OAI21_X1 U8596 ( .B1(n7387), .B2(n8266), .A(n7386), .ZN(P2_U3153) );
  INV_X1 U8597 ( .A(n7388), .ZN(n7436) );
  AOI22_X1 U8598 ( .A1(n10214), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7389), .ZN(n7390) );
  OAI21_X1 U8599 ( .B1(n7436), .B2(n8202), .A(n7390), .ZN(P1_U3337) );
  INV_X1 U8600 ( .A(n10405), .ZN(n8601) );
  OAI222_X1 U8601 ( .A1(n9153), .A2(n7392), .B1(n9147), .B2(n7391), .C1(n8601), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  NAND2_X1 U8602 ( .A1(n9279), .A2(n7535), .ZN(n7393) );
  NAND2_X1 U8603 ( .A1(n10478), .A2(n9572), .ZN(n9290) );
  INV_X1 U8604 ( .A(n10478), .ZN(n7496) );
  NAND2_X1 U8605 ( .A1(n9290), .A2(n9489), .ZN(n7484) );
  NAND2_X1 U8606 ( .A1(n10478), .A2(n7395), .ZN(n7661) );
  INV_X1 U8607 ( .A(n7665), .ZN(n9571) );
  NAND2_X1 U8608 ( .A1(n7430), .A2(n9571), .ZN(n9491) );
  INV_X1 U8609 ( .A(n7430), .ZN(n10489) );
  NAND2_X1 U8610 ( .A1(n7665), .A2(n10489), .ZN(n9493) );
  XNOR2_X1 U8611 ( .A(n7431), .B(n9400), .ZN(n10493) );
  NAND3_X1 U8612 ( .A1(n7398), .A2(n7397), .A3(n7396), .ZN(n7404) );
  NAND2_X1 U8613 ( .A1(n8025), .A2(n7472), .ZN(n7399) );
  NAND2_X1 U8614 ( .A1(n7400), .A2(n9485), .ZN(n7487) );
  INV_X1 U8615 ( .A(n7484), .ZN(n9401) );
  NAND2_X1 U8616 ( .A1(n7487), .A2(n9401), .ZN(n7486) );
  NAND2_X1 U8617 ( .A1(n7486), .A2(n9489), .ZN(n7420) );
  XNOR2_X1 U8618 ( .A(n7420), .B(n9400), .ZN(n7401) );
  NAND2_X1 U8619 ( .A1(n7401), .A2(n9892), .ZN(n7403) );
  AOI22_X1 U8620 ( .A1(n9889), .A2(n9572), .B1(n9570), .B2(n9887), .ZN(n7402)
         );
  AND2_X1 U8621 ( .A1(n7403), .A2(n7402), .ZN(n10491) );
  INV_X2 U8622 ( .A(n9868), .ZN(n10562) );
  MUX2_X1 U8623 ( .A(n10491), .B(n7332), .S(n10562), .Z(n7410) );
  INV_X1 U8624 ( .A(n7425), .ZN(n7426) );
  AOI211_X1 U8625 ( .C1(n10489), .C2(n4981), .A(n10512), .B(n7426), .ZN(n10488) );
  INV_X1 U8626 ( .A(n7405), .ZN(n7406) );
  OAI22_X1 U8627 ( .A1(n9879), .A2(n7430), .B1(n10448), .B2(n7407), .ZN(n7408)
         );
  AOI21_X1 U8628 ( .B1(n10488), .B2(n10556), .A(n7408), .ZN(n7409) );
  OAI211_X1 U8629 ( .C1(n10493), .C2(n9896), .A(n7410), .B(n7409), .ZN(
        P1_U3289) );
  AOI22_X1 U8630 ( .A1(n10562), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10551), .ZN(n7414) );
  NOR2_X1 U8631 ( .A1(n8103), .A2(n10512), .ZN(n9855) );
  NAND3_X1 U8632 ( .A1(n9855), .A2(n7412), .A3(n7411), .ZN(n7413) );
  OAI211_X1 U8633 ( .C1(n7415), .C2(n9879), .A(n7414), .B(n7413), .ZN(n7416)
         );
  AOI21_X1 U8634 ( .B1(n9815), .B2(n7417), .A(n7416), .ZN(n7418) );
  OAI21_X1 U8635 ( .B1(n7419), .B2(n10562), .A(n7418), .ZN(P1_U3292) );
  NAND2_X1 U8636 ( .A1(n7420), .A2(n9491), .ZN(n7422) );
  NAND2_X1 U8637 ( .A1(n7422), .A2(n9493), .ZN(n7421) );
  NAND2_X1 U8638 ( .A1(n10503), .A2(n9570), .ZN(n9497) );
  NAND2_X1 U8639 ( .A1(n9497), .A2(n9494), .ZN(n7670) );
  INV_X1 U8640 ( .A(n7670), .ZN(n9402) );
  NAND2_X1 U8641 ( .A1(n7421), .A2(n9402), .ZN(n7565) );
  NAND3_X1 U8642 ( .A1(n7422), .A2(n7670), .A3(n9493), .ZN(n7423) );
  NAND2_X1 U8643 ( .A1(n7565), .A2(n7423), .ZN(n7424) );
  AOI222_X1 U8644 ( .A1(n9892), .A2(n7424), .B1(n9569), .B2(n9887), .C1(n9571), 
        .C2(n9889), .ZN(n10502) );
  OR2_X1 U8645 ( .A1(n7425), .A2(n7547), .ZN(n7573) );
  OAI211_X1 U8646 ( .C1(n7426), .C2(n10503), .A(n10527), .B(n7573), .ZN(n10501) );
  INV_X1 U8647 ( .A(n10501), .ZN(n7429) );
  AOI22_X1 U8648 ( .A1(n10562), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7545), .B2(
        n10551), .ZN(n7427) );
  OAI21_X1 U8649 ( .B1(n10503), .B2(n9879), .A(n7427), .ZN(n7428) );
  AOI21_X1 U8650 ( .B1(n7429), .B2(n10556), .A(n7428), .ZN(n7434) );
  NAND2_X1 U8651 ( .A1(n7431), .A2(n7665), .ZN(n7432) );
  NAND2_X1 U8652 ( .A1(n7669), .A2(n7432), .ZN(n7561) );
  XNOR2_X1 U8653 ( .A(n7670), .B(n7561), .ZN(n10505) );
  NAND2_X1 U8654 ( .A1(n10505), .A2(n9815), .ZN(n7433) );
  OAI211_X1 U8655 ( .C1(n10502), .C2(n10562), .A(n7434), .B(n7433), .ZN(
        P1_U3288) );
  INV_X1 U8656 ( .A(n8617), .ZN(n8625) );
  INV_X1 U8657 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7435) );
  OAI222_X1 U8658 ( .A1(P2_U3151), .A2(n8625), .B1(n9147), .B2(n7436), .C1(
        n7435), .C2(n9153), .ZN(P2_U3277) );
  INV_X1 U8659 ( .A(n8487), .ZN(n7439) );
  NAND3_X1 U8660 ( .A1(n7594), .A2(n7439), .A3(n7438), .ZN(n7440) );
  NAND2_X1 U8661 ( .A1(n7437), .A2(n7440), .ZN(n7441) );
  AOI222_X1 U8662 ( .A1(n8793), .A2(n7441), .B1(n5136), .B2(n8797), .C1(n8534), 
        .C2(n8771), .ZN(n7616) );
  OAI22_X1 U8663 ( .A1(n10575), .A2(n7447), .B1(n5467), .B2(n10468), .ZN(n7442) );
  AOI21_X1 U8664 ( .B1(n10568), .B2(n7615), .A(n7442), .ZN(n7446) );
  NAND2_X1 U8665 ( .A1(n7592), .A2(n7443), .ZN(n7444) );
  XNOR2_X1 U8666 ( .A(n7444), .B(n8487), .ZN(n7619) );
  NAND2_X1 U8667 ( .A1(n7619), .A2(n8752), .ZN(n7445) );
  OAI211_X1 U8668 ( .C1(n7616), .C2(n10577), .A(n7446), .B(n7445), .ZN(
        P2_U3225) );
  OR2_X1 U8669 ( .A1(n7459), .A2(n7447), .ZN(n7448) );
  NAND2_X1 U8670 ( .A1(n7449), .A2(n7448), .ZN(n8583) );
  NOR2_X1 U8671 ( .A1(n7450), .A2(n7461), .ZN(n8582) );
  AOI21_X1 U8672 ( .B1(n7461), .B2(n7450), .A(n8582), .ZN(n7471) );
  AOI21_X1 U8673 ( .B1(n7452), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7451), .ZN(
        n8542) );
  XNOR2_X1 U8674 ( .A(n8542), .B(n8584), .ZN(n7453) );
  NAND2_X1 U8675 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7453), .ZN(n8543) );
  OAI21_X1 U8676 ( .B1(n7453), .B2(P2_REG1_REG_9__SCAN_IN), .A(n8543), .ZN(
        n7454) );
  NAND2_X1 U8677 ( .A1(n7454), .A2(n10413), .ZN(n7470) );
  NOR2_X1 U8678 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6474), .ZN(n7693) );
  INV_X1 U8679 ( .A(n7693), .ZN(n7455) );
  OAI21_X1 U8680 ( .B1(n10271), .B2(n8584), .A(n7455), .ZN(n7468) );
  INV_X1 U8681 ( .A(n7456), .ZN(n7458) );
  AOI21_X1 U8682 ( .B1(n7459), .B2(n7458), .A(n7457), .ZN(n7465) );
  MUX2_X1 U8683 ( .A(n7461), .B(n7460), .S(n8619), .Z(n7463) );
  AND2_X1 U8684 ( .A1(n7463), .A2(n8541), .ZN(n8564) );
  INV_X1 U8685 ( .A(n8564), .ZN(n7462) );
  OAI21_X1 U8686 ( .B1(n8541), .B2(n7463), .A(n7462), .ZN(n7464) );
  NOR2_X1 U8687 ( .A1(n7465), .A2(n7464), .ZN(n8563) );
  AOI21_X1 U8688 ( .B1(n7465), .B2(n7464), .A(n8563), .ZN(n7466) );
  NOR2_X1 U8689 ( .A1(n7466), .A2(n10282), .ZN(n7467) );
  AOI211_X1 U8690 ( .C1(n10403), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7468), .B(
        n7467), .ZN(n7469) );
  OAI211_X1 U8691 ( .C1(n7471), .C2(n10418), .A(n7470), .B(n7469), .ZN(
        P2_U3191) );
  INV_X1 U8692 ( .A(n7472), .ZN(n7473) );
  NAND2_X1 U8693 ( .A1(n9868), .A2(n7473), .ZN(n8033) );
  NAND2_X1 U8694 ( .A1(n7474), .A2(n9868), .ZN(n7482) );
  INV_X1 U8695 ( .A(n9879), .ZN(n10552) );
  INV_X1 U8696 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7476) );
  INV_X1 U8697 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7475) );
  OAI22_X1 U8698 ( .A1(n9868), .A2(n7476), .B1(n7475), .B2(n10448), .ZN(n7479)
         );
  NOR2_X1 U8699 ( .A1(n7477), .A2(n8103), .ZN(n7478) );
  AOI211_X1 U8700 ( .C1(n10552), .C2(n7480), .A(n7479), .B(n7478), .ZN(n7481)
         );
  OAI211_X1 U8701 ( .C1(n7483), .C2(n8033), .A(n7482), .B(n7481), .ZN(P1_U3291) );
  OAI21_X1 U8702 ( .B1(n7485), .B2(n7484), .A(n7663), .ZN(n10481) );
  INV_X1 U8703 ( .A(n10481), .ZN(n7499) );
  OAI21_X1 U8704 ( .B1(n9401), .B2(n7487), .A(n7486), .ZN(n7489) );
  OAI22_X1 U8705 ( .A1(n7535), .A2(n10533), .B1(n7665), .B2(n10531), .ZN(n7488) );
  AOI21_X1 U8706 ( .B1(n7489), .B2(n9892), .A(n7488), .ZN(n7490) );
  OAI21_X1 U8707 ( .B1(n7499), .B2(n8025), .A(n7490), .ZN(n10479) );
  NAND2_X1 U8708 ( .A1(n10479), .A2(n9868), .ZN(n7498) );
  INV_X1 U8709 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7491) );
  OAI22_X1 U8710 ( .A1(n9868), .A2(n7491), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10448), .ZN(n7495) );
  INV_X1 U8711 ( .A(n7492), .ZN(n7493) );
  OAI211_X1 U8712 ( .C1(n10478), .C2(n7493), .A(n4981), .B(n10527), .ZN(n10477) );
  NOR2_X1 U8713 ( .A1(n10477), .A2(n8103), .ZN(n7494) );
  AOI211_X1 U8714 ( .C1(n10552), .C2(n7496), .A(n7495), .B(n7494), .ZN(n7497)
         );
  OAI211_X1 U8715 ( .C1(n7499), .C2(n8033), .A(n7498), .B(n7497), .ZN(P1_U3290) );
  NOR2_X1 U8716 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7500) );
  AOI21_X1 U8717 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7500), .ZN(n10083) );
  NOR2_X1 U8718 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7501) );
  AOI21_X1 U8719 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7501), .ZN(n10080) );
  NOR2_X1 U8720 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7502) );
  AOI21_X1 U8721 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7502), .ZN(n10077) );
  NOR2_X1 U8722 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7503) );
  AOI21_X1 U8723 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7503), .ZN(n10074) );
  NOR2_X1 U8724 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7504) );
  AOI21_X1 U8725 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7504), .ZN(n10071) );
  NOR2_X1 U8726 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7505) );
  AOI21_X1 U8727 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7505), .ZN(n10068) );
  NOR2_X1 U8728 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7506) );
  AOI21_X1 U8729 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7506), .ZN(n10065) );
  NOR2_X1 U8730 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7507) );
  AOI21_X1 U8731 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7507), .ZN(n10062) );
  NOR2_X1 U8732 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7508) );
  AOI21_X1 U8733 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7508), .ZN(n10059) );
  NOR2_X1 U8734 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7509) );
  AOI21_X1 U8735 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7509), .ZN(n10056) );
  NOR2_X1 U8736 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7510) );
  AOI21_X1 U8737 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7510), .ZN(n10053) );
  NOR2_X1 U8738 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7511) );
  AOI21_X1 U8739 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7511), .ZN(n10050) );
  NOR2_X1 U8740 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7512) );
  AOI21_X1 U8741 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7512), .ZN(n10047) );
  NOR2_X1 U8742 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7513) );
  AOI21_X1 U8743 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7513), .ZN(n10044) );
  NAND2_X1 U8744 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10030) );
  INV_X1 U8745 ( .A(n10030), .ZN(n7514) );
  INV_X1 U8746 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U8747 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  AOI22_X1 U8748 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7514), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10029), .ZN(n10035) );
  NAND2_X1 U8749 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7515) );
  OAI21_X1 U8750 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7515), .ZN(n10034) );
  NOR2_X1 U8751 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  AOI21_X1 U8752 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10033), .ZN(n10038) );
  NAND2_X1 U8753 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7516) );
  OAI21_X1 U8754 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7516), .ZN(n10037) );
  NOR2_X1 U8755 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  AOI21_X1 U8756 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10036), .ZN(n10041) );
  NOR2_X1 U8757 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7517) );
  AOI21_X1 U8758 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7517), .ZN(n10040) );
  NAND2_X1 U8759 ( .A1(n10041), .A2(n10040), .ZN(n10039) );
  OAI21_X1 U8760 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10039), .ZN(n10043) );
  NAND2_X1 U8761 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  OAI21_X1 U8762 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10042), .ZN(n10046) );
  NAND2_X1 U8763 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  OAI21_X1 U8764 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10045), .ZN(n10049) );
  NAND2_X1 U8765 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  OAI21_X1 U8766 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10048), .ZN(n10052) );
  NAND2_X1 U8767 ( .A1(n10053), .A2(n10052), .ZN(n10051) );
  OAI21_X1 U8768 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10051), .ZN(n10055) );
  NAND2_X1 U8769 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  OAI21_X1 U8770 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10054), .ZN(n10058) );
  NAND2_X1 U8771 ( .A1(n10059), .A2(n10058), .ZN(n10057) );
  OAI21_X1 U8772 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10057), .ZN(n10061) );
  NAND2_X1 U8773 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  OAI21_X1 U8774 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10060), .ZN(n10064) );
  NAND2_X1 U8775 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  OAI21_X1 U8776 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10063), .ZN(n10067) );
  NAND2_X1 U8777 ( .A1(n10068), .A2(n10067), .ZN(n10066) );
  OAI21_X1 U8778 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10066), .ZN(n10070) );
  NAND2_X1 U8779 ( .A1(n10071), .A2(n10070), .ZN(n10069) );
  OAI21_X1 U8780 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10069), .ZN(n10073) );
  NAND2_X1 U8781 ( .A1(n10074), .A2(n10073), .ZN(n10072) );
  OAI21_X1 U8782 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10072), .ZN(n10076) );
  NAND2_X1 U8783 ( .A1(n10077), .A2(n10076), .ZN(n10075) );
  OAI21_X1 U8784 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10075), .ZN(n10079) );
  NAND2_X1 U8785 ( .A1(n10080), .A2(n10079), .ZN(n10078) );
  OAI21_X1 U8786 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10078), .ZN(n10082) );
  NAND2_X1 U8787 ( .A1(n10083), .A2(n10082), .ZN(n10081) );
  OAI21_X1 U8788 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10081), .ZN(n7520) );
  XNOR2_X1 U8789 ( .A(n7518), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7519) );
  XNOR2_X1 U8790 ( .A(n7520), .B(n7519), .ZN(ADD_1068_U4) );
  INV_X1 U8791 ( .A(n7522), .ZN(n7524) );
  NAND2_X1 U8792 ( .A1(n7524), .A2(n7523), .ZN(n7541) );
  NAND2_X1 U8793 ( .A1(n7521), .A2(n7541), .ZN(n7527) );
  NAND2_X1 U8794 ( .A1(n7521), .A2(n7525), .ZN(n7603) );
  INV_X1 U8795 ( .A(n7603), .ZN(n7526) );
  AOI21_X1 U8796 ( .B1(n7528), .B2(n7527), .A(n7526), .ZN(n7532) );
  INV_X1 U8797 ( .A(n9568), .ZN(n7675) );
  AOI22_X1 U8798 ( .A1(n9262), .A2(n7575), .B1(n9261), .B2(n9570), .ZN(n7529)
         );
  NAND2_X1 U8799 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10118) );
  OAI211_X1 U8800 ( .C1(n7675), .C2(n9264), .A(n7529), .B(n10118), .ZN(n7530)
         );
  AOI21_X1 U8801 ( .B1(n7576), .B2(n9266), .A(n7530), .ZN(n7531) );
  OAI21_X1 U8802 ( .B1(n7532), .B2(n9268), .A(n7531), .ZN(P1_U3239) );
  XOR2_X1 U8803 ( .A(n7533), .B(n7534), .Z(n7540) );
  NAND2_X1 U8804 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9607) );
  OAI21_X1 U8805 ( .B1(n9243), .B2(n10478), .A(n9607), .ZN(n7537) );
  OAI22_X1 U8806 ( .A1(n9250), .A2(n7535), .B1(n7665), .B2(n9264), .ZN(n7536)
         );
  AOI211_X1 U8807 ( .C1(n9262), .C2(n7538), .A(n7537), .B(n7536), .ZN(n7539)
         );
  OAI21_X1 U8808 ( .B1(n7540), .B2(n9268), .A(n7539), .ZN(P1_U3218) );
  NAND2_X1 U8809 ( .A1(n7542), .A2(n7541), .ZN(n7543) );
  XOR2_X1 U8810 ( .A(n7544), .B(n7543), .Z(n7550) );
  AOI22_X1 U8811 ( .A1(n9262), .A2(n7545), .B1(n9261), .B2(n9571), .ZN(n7549)
         );
  NAND2_X1 U8812 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10103) );
  OAI21_X1 U8813 ( .B1(n9264), .B2(n10534), .A(n10103), .ZN(n7546) );
  AOI21_X1 U8814 ( .B1(n7547), .B2(n9266), .A(n7546), .ZN(n7548) );
  OAI211_X1 U8815 ( .C1(n7550), .C2(n9268), .A(n7549), .B(n7548), .ZN(P1_U3227) );
  INV_X1 U8816 ( .A(n7551), .ZN(n7553) );
  XNOR2_X1 U8817 ( .A(n7615), .B(n8194), .ZN(n7697) );
  XNOR2_X1 U8818 ( .A(n7697), .B(n8533), .ZN(n7698) );
  XOR2_X1 U8819 ( .A(n4978), .B(n7698), .Z(n7560) );
  AOI21_X1 U8820 ( .B1(n10657), .B2(n5136), .A(n7555), .ZN(n7557) );
  NAND2_X1 U8821 ( .A1(n8534), .A2(n10655), .ZN(n7556) );
  OAI211_X1 U8822 ( .C1(n10653), .C2(n5467), .A(n7557), .B(n7556), .ZN(n7558)
         );
  AOI21_X1 U8823 ( .B1(n10667), .B2(n7615), .A(n7558), .ZN(n7559) );
  OAI21_X1 U8824 ( .B1(n7560), .B2(n8266), .A(n7559), .ZN(P2_U3161) );
  NAND2_X1 U8825 ( .A1(n7561), .A2(n7670), .ZN(n7563) );
  NAND2_X1 U8826 ( .A1(n10503), .A2(n7562), .ZN(n7659) );
  NAND2_X1 U8827 ( .A1(n7563), .A2(n7659), .ZN(n7564) );
  XNOR2_X1 U8828 ( .A(n7564), .B(n9300), .ZN(n10515) );
  INV_X1 U8829 ( .A(n8025), .ZN(n10544) );
  NAND2_X1 U8830 ( .A1(n10515), .A2(n10544), .ZN(n7572) );
  NAND2_X1 U8831 ( .A1(n7565), .A2(n9494), .ZN(n7680) );
  INV_X1 U8832 ( .A(n9300), .ZN(n7566) );
  XNOR2_X1 U8833 ( .A(n7680), .B(n7566), .ZN(n7570) );
  NAND2_X1 U8834 ( .A1(n9570), .A2(n9889), .ZN(n7568) );
  NAND2_X1 U8835 ( .A1(n9568), .A2(n9887), .ZN(n7567) );
  NAND2_X1 U8836 ( .A1(n7568), .A2(n7567), .ZN(n7569) );
  AOI21_X1 U8837 ( .B1(n7570), .B2(n9892), .A(n7569), .ZN(n7571) );
  INV_X1 U8838 ( .A(n8033), .ZN(n10557) );
  AND2_X1 U8839 ( .A1(n7573), .A2(n7576), .ZN(n7574) );
  NOR2_X2 U8840 ( .A1(n7573), .A2(n7576), .ZN(n10529) );
  OR2_X1 U8841 ( .A1(n7574), .A2(n10529), .ZN(n10513) );
  INV_X1 U8842 ( .A(n9855), .ZN(n9673) );
  AOI22_X1 U8843 ( .A1(n10562), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7575), .B2(
        n10551), .ZN(n7578) );
  NAND2_X1 U8844 ( .A1(n10552), .A2(n7576), .ZN(n7577) );
  OAI211_X1 U8845 ( .C1(n10513), .C2(n9673), .A(n7578), .B(n7577), .ZN(n7579)
         );
  AOI21_X1 U8846 ( .B1(n10515), .B2(n10557), .A(n7579), .ZN(n7580) );
  OAI21_X1 U8847 ( .B1(n10517), .B2(n10562), .A(n7580), .ZN(P1_U3287) );
  INV_X1 U8848 ( .A(n7581), .ZN(n8491) );
  OAI21_X1 U8849 ( .B1(n5490), .B2(n8491), .A(n7624), .ZN(n7644) );
  NAND2_X1 U8850 ( .A1(n7437), .A2(n7583), .ZN(n7582) );
  NAND2_X1 U8851 ( .A1(n7582), .A2(n7581), .ZN(n7585) );
  NAND3_X1 U8852 ( .A1(n7437), .A2(n8491), .A3(n7583), .ZN(n7584) );
  AND2_X1 U8853 ( .A1(n7585), .A2(n7584), .ZN(n7586) );
  OAI222_X1 U8854 ( .A1(n8801), .A2(n7598), .B1(n8786), .B2(n7841), .C1(n8723), 
        .C2(n7586), .ZN(n7645) );
  NAND2_X1 U8855 ( .A1(n7645), .A2(n10575), .ZN(n7589) );
  OAI22_X1 U8856 ( .A1(n10575), .A2(n7461), .B1(n7696), .B2(n10468), .ZN(n7587) );
  AOI21_X1 U8857 ( .B1(n7703), .B2(n10568), .A(n7587), .ZN(n7588) );
  OAI211_X1 U8858 ( .C1(n8807), .C2(n7644), .A(n7589), .B(n7588), .ZN(P2_U3224) );
  NAND2_X1 U8859 ( .A1(n7590), .A2(n8488), .ZN(n7591) );
  INV_X1 U8860 ( .A(n7593), .ZN(n7596) );
  INV_X1 U8861 ( .A(n7594), .ZN(n7595) );
  AOI21_X1 U8862 ( .B1(n5242), .B2(n7596), .A(n7595), .ZN(n7597) );
  OAI222_X1 U8863 ( .A1(n8801), .A2(n7599), .B1(n8786), .B2(n7598), .C1(n8723), 
        .C2(n7597), .ZN(n10564) );
  AOI211_X1 U8864 ( .C1(n10571), .C2(n8872), .A(n7600), .B(n10564), .ZN(n10563) );
  OR2_X1 U8865 ( .A1(n10563), .A2(n7621), .ZN(n7601) );
  OAI21_X1 U8866 ( .B1(n8876), .B2(n7149), .A(n7601), .ZN(P2_U3466) );
  NAND2_X1 U8867 ( .A1(n7603), .A2(n7602), .ZN(n7604) );
  XOR2_X1 U8868 ( .A(n7605), .B(n7604), .Z(n7609) );
  INV_X1 U8869 ( .A(n10530), .ZN(n10553) );
  AOI22_X1 U8870 ( .A1(n9262), .A2(n10550), .B1(n9261), .B2(n9569), .ZN(n7606)
         );
  NAND2_X1 U8871 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10133) );
  OAI211_X1 U8872 ( .C1(n10532), .C2(n9264), .A(n7606), .B(n10133), .ZN(n7607)
         );
  AOI21_X1 U8873 ( .B1(n10553), .B2(n9266), .A(n7607), .ZN(n7608) );
  OAI21_X1 U8874 ( .B1(n7609), .B2(n9268), .A(n7608), .ZN(P1_U3213) );
  INV_X1 U8875 ( .A(n7610), .ZN(n7613) );
  OAI222_X1 U8876 ( .A1(n9153), .A2(n7612), .B1(n9147), .B2(n7613), .C1(n7611), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U8877 ( .A1(n10018), .A2(n7614), .B1(n8202), .B2(n7613), .C1(
        P1_U3086), .C2(n6030), .ZN(P1_U3336) );
  INV_X1 U8878 ( .A(n7615), .ZN(n7617) );
  OAI21_X1 U8879 ( .B1(n7617), .B2(n8844), .A(n7616), .ZN(n7618) );
  AOI21_X1 U8880 ( .B1(n8872), .B2(n7619), .A(n7618), .ZN(n10587) );
  NAND2_X1 U8881 ( .A1(n7621), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7620) );
  OAI21_X1 U8882 ( .B1(n10587), .B2(n7621), .A(n7620), .ZN(P2_U3467) );
  NAND2_X1 U8883 ( .A1(n7623), .A2(n7622), .ZN(n8490) );
  NAND2_X1 U8884 ( .A1(n7624), .A2(n8369), .ZN(n7625) );
  XOR2_X1 U8885 ( .A(n8490), .B(n7625), .Z(n7629) );
  INV_X1 U8886 ( .A(n7629), .ZN(n7758) );
  XNOR2_X1 U8887 ( .A(n7626), .B(n8490), .ZN(n7631) );
  INV_X1 U8888 ( .A(n8661), .ZN(n10565) );
  OAI22_X1 U8889 ( .A1(n7843), .A2(n8786), .B1(n7627), .B2(n8801), .ZN(n7628)
         );
  AOI21_X1 U8890 ( .B1(n7629), .B2(n10565), .A(n7628), .ZN(n7630) );
  OAI21_X1 U8891 ( .B1(n8723), .B2(n7631), .A(n7630), .ZN(n7759) );
  NAND2_X1 U8892 ( .A1(n7759), .A2(n10575), .ZN(n7634) );
  OAI22_X1 U8893 ( .A1(n10575), .A2(n8565), .B1(n7793), .B2(n10468), .ZN(n7632) );
  AOI21_X1 U8894 ( .B1(n7795), .B2(n10568), .A(n7632), .ZN(n7633) );
  OAI211_X1 U8895 ( .C1(n7758), .C2(n10567), .A(n7634), .B(n7633), .ZN(
        P2_U3223) );
  XNOR2_X1 U8896 ( .A(n7635), .B(n8492), .ZN(n7636) );
  OAI222_X1 U8897 ( .A1(n8786), .A2(n7868), .B1(n8801), .B2(n7841), .C1(n8723), 
        .C2(n7636), .ZN(n7799) );
  INV_X1 U8898 ( .A(n7799), .ZN(n7642) );
  NAND2_X1 U8899 ( .A1(n7637), .A2(n8381), .ZN(n7638) );
  XNOR2_X1 U8900 ( .A(n7638), .B(n8492), .ZN(n7800) );
  INV_X1 U8901 ( .A(n7720), .ZN(n7798) );
  NOR2_X1 U8902 ( .A1(n7798), .A2(n8649), .ZN(n7640) );
  OAI22_X1 U8903 ( .A1(n10575), .A2(n6502), .B1(n7850), .B2(n10468), .ZN(n7639) );
  AOI211_X1 U8904 ( .C1(n7800), .C2(n8752), .A(n7640), .B(n7639), .ZN(n7641)
         );
  OAI21_X1 U8905 ( .B1(n7642), .B2(n10577), .A(n7641), .ZN(P2_U3222) );
  NAND2_X1 U8906 ( .A1(n8580), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7643) );
  OAI21_X1 U8907 ( .B1(n8317), .B2(n8580), .A(n7643), .ZN(P2_U3520) );
  NOR2_X1 U8908 ( .A1(n7644), .A2(n8839), .ZN(n7646) );
  AOI211_X1 U8909 ( .C1(n8871), .C2(n7703), .A(n7646), .B(n7645), .ZN(n10596)
         );
  INV_X1 U8910 ( .A(n10596), .ZN(n7647) );
  NAND2_X1 U8911 ( .A1(n7647), .A2(n8876), .ZN(n7648) );
  OAI21_X1 U8912 ( .B1(n8876), .B2(n7460), .A(n7648), .ZN(P2_U3468) );
  INV_X1 U8913 ( .A(n7649), .ZN(n7691) );
  OAI222_X1 U8914 ( .A1(P1_U3086), .A2(n9544), .B1(n8202), .B2(n7691), .C1(
        n7650), .C2(n10018), .ZN(P1_U3335) );
  XNOR2_X1 U8915 ( .A(n7653), .B(n7652), .ZN(n7654) );
  XNOR2_X1 U8916 ( .A(n7651), .B(n7654), .ZN(n7658) );
  INV_X1 U8917 ( .A(n10532), .ZN(n9567) );
  AOI22_X1 U8918 ( .A1(n9262), .A2(n7740), .B1(n9261), .B2(n9567), .ZN(n7655)
         );
  NAND2_X1 U8919 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10261) );
  OAI211_X1 U8920 ( .C1(n7776), .C2(n9264), .A(n7655), .B(n10261), .ZN(n7656)
         );
  AOI21_X1 U8921 ( .B1(n7775), .B2(n9266), .A(n7656), .ZN(n7657) );
  OAI21_X1 U8922 ( .B1(n7658), .B2(n9268), .A(n7657), .ZN(P1_U3231) );
  INV_X1 U8923 ( .A(n7659), .ZN(n7660) );
  AND2_X1 U8924 ( .A1(n7661), .A2(n7664), .ZN(n7662) );
  NAND2_X1 U8925 ( .A1(n7663), .A2(n7662), .ZN(n7667) );
  INV_X1 U8926 ( .A(n7664), .ZN(n7672) );
  NAND2_X1 U8927 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  NAND2_X1 U8928 ( .A1(n7669), .A2(n7668), .ZN(n10521) );
  AND2_X1 U8929 ( .A1(n7670), .A2(n9300), .ZN(n7671) );
  NAND2_X1 U8930 ( .A1(n10530), .A2(n9568), .ZN(n9302) );
  NAND2_X1 U8931 ( .A1(n7675), .A2(n10553), .ZN(n9308) );
  NAND2_X1 U8932 ( .A1(n9302), .A2(n9308), .ZN(n10536) );
  AND2_X1 U8933 ( .A1(n10522), .A2(n10536), .ZN(n7673) );
  NAND2_X1 U8934 ( .A1(n10521), .A2(n7673), .ZN(n7679) );
  NAND2_X1 U8935 ( .A1(n10511), .A2(n10534), .ZN(n10523) );
  INV_X1 U8936 ( .A(n10523), .ZN(n7674) );
  NAND2_X1 U8937 ( .A1(n10530), .A2(n7675), .ZN(n7676) );
  AND2_X1 U8938 ( .A1(n7677), .A2(n7676), .ZN(n7678) );
  NAND2_X1 U8939 ( .A1(n7679), .A2(n7678), .ZN(n7745) );
  OR2_X1 U8940 ( .A1(n7746), .A2(n10532), .ZN(n9326) );
  NAND2_X1 U8941 ( .A1(n7746), .A2(n10532), .ZN(n9309) );
  NAND2_X1 U8942 ( .A1(n9326), .A2(n9309), .ZN(n7744) );
  XNOR2_X1 U8943 ( .A(n7745), .B(n7744), .ZN(n10581) );
  INV_X1 U8944 ( .A(n9405), .ZN(n9496) );
  INV_X1 U8945 ( .A(n9303), .ZN(n10537) );
  NOR2_X1 U8946 ( .A1(n10536), .A2(n10537), .ZN(n7681) );
  NAND2_X1 U8947 ( .A1(n10535), .A2(n7681), .ZN(n10540) );
  NAND2_X1 U8948 ( .A1(n10540), .A2(n9308), .ZN(n7682) );
  INV_X1 U8949 ( .A(n7744), .ZN(n9307) );
  XNOR2_X1 U8950 ( .A(n7682), .B(n9307), .ZN(n7683) );
  NAND2_X1 U8951 ( .A1(n7683), .A2(n9892), .ZN(n7685) );
  AOI22_X1 U8952 ( .A1(n9566), .A2(n9887), .B1(n9889), .B2(n9568), .ZN(n7684)
         );
  NAND2_X1 U8953 ( .A1(n7685), .A2(n7684), .ZN(n7686) );
  AOI21_X1 U8954 ( .B1(n10581), .B2(n10544), .A(n7686), .ZN(n10583) );
  AND2_X1 U8955 ( .A1(n10529), .A2(n10530), .ZN(n10526) );
  INV_X1 U8956 ( .A(n7746), .ZN(n10579) );
  NAND2_X1 U8957 ( .A1(n10526), .A2(n10579), .ZN(n7738) );
  OAI211_X1 U8958 ( .C1(n10526), .C2(n10579), .A(n10527), .B(n7738), .ZN(
        n10578) );
  AOI22_X1 U8959 ( .A1(n10562), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7712), .B2(
        n10551), .ZN(n7688) );
  NAND2_X1 U8960 ( .A1(n10552), .A2(n7746), .ZN(n7687) );
  OAI211_X1 U8961 ( .C1(n10578), .C2(n8103), .A(n7688), .B(n7687), .ZN(n7689)
         );
  AOI21_X1 U8962 ( .B1(n10581), .B2(n10557), .A(n7689), .ZN(n7690) );
  OAI21_X1 U8963 ( .B1(n10583), .B2(n10562), .A(n7690), .ZN(P1_U3285) );
  OAI222_X1 U8964 ( .A1(n9153), .A2(n7692), .B1(P2_U3151), .B2(n8322), .C1(
        n9147), .C2(n7691), .ZN(P2_U3275) );
  AOI21_X1 U8965 ( .B1(n10657), .B2(n8532), .A(n7693), .ZN(n7695) );
  NAND2_X1 U8966 ( .A1(n8533), .A2(n10655), .ZN(n7694) );
  OAI211_X1 U8967 ( .C1(n10653), .C2(n7696), .A(n7695), .B(n7694), .ZN(n7702)
         );
  XNOR2_X1 U8968 ( .A(n7703), .B(n8194), .ZN(n7719) );
  XNOR2_X1 U8969 ( .A(n7719), .B(n5136), .ZN(n7700) );
  AOI211_X1 U8970 ( .C1(n7700), .C2(n7699), .A(n8266), .B(n7718), .ZN(n7701)
         );
  AOI211_X1 U8971 ( .C1(n10667), .C2(n7703), .A(n7702), .B(n7701), .ZN(n7704)
         );
  INV_X1 U8972 ( .A(n7704), .ZN(P2_U3171) );
  INV_X1 U8973 ( .A(n7707), .ZN(n7711) );
  AOI21_X1 U8974 ( .B1(n7707), .B2(n7706), .A(n7705), .ZN(n7708) );
  NOR2_X1 U8975 ( .A1(n7708), .A2(n9268), .ZN(n7709) );
  OAI21_X1 U8976 ( .B1(n7711), .B2(n7710), .A(n7709), .ZN(n7717) );
  NAND2_X1 U8977 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10148) );
  INV_X1 U8978 ( .A(n10148), .ZN(n7715) );
  INV_X1 U8979 ( .A(n7712), .ZN(n7713) );
  OAI22_X1 U8980 ( .A1(n7734), .A2(n9264), .B1(n9251), .B2(n7713), .ZN(n7714)
         );
  AOI211_X1 U8981 ( .C1(n9261), .C2(n9568), .A(n7715), .B(n7714), .ZN(n7716)
         );
  OAI211_X1 U8982 ( .C1(n10579), .C2(n9243), .A(n7717), .B(n7716), .ZN(
        P1_U3221) );
  XNOR2_X1 U8983 ( .A(n7720), .B(n8194), .ZN(n7844) );
  XNOR2_X1 U8984 ( .A(n7795), .B(n8194), .ZN(n7790) );
  AOI22_X1 U8985 ( .A1(n7844), .A2(n8531), .B1(n7790), .B2(n8532), .ZN(n7724)
         );
  INV_X1 U8986 ( .A(n7790), .ZN(n7839) );
  AOI21_X1 U8987 ( .B1(n7839), .B2(n7841), .A(n7843), .ZN(n7722) );
  NAND2_X1 U8988 ( .A1(n7841), .A2(n7843), .ZN(n7721) );
  OAI22_X1 U8989 ( .A1(n7844), .A2(n7722), .B1(n7790), .B2(n7721), .ZN(n7723)
         );
  XNOR2_X1 U8990 ( .A(n8870), .B(n8194), .ZN(n7867) );
  XNOR2_X1 U8991 ( .A(n7867), .B(n7868), .ZN(n7725) );
  XNOR2_X1 U8992 ( .A(n7866), .B(n7725), .ZN(n7731) );
  NAND2_X1 U8993 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10338) );
  INV_X1 U8994 ( .A(n10338), .ZN(n7727) );
  NOR2_X1 U8995 ( .A1(n10641), .A2(n8405), .ZN(n7726) );
  AOI211_X1 U8996 ( .C1(n10655), .C2(n8531), .A(n7727), .B(n7726), .ZN(n7728)
         );
  OAI21_X1 U8997 ( .B1(n7825), .B2(n10653), .A(n7728), .ZN(n7729) );
  AOI21_X1 U8998 ( .B1(n8870), .B2(n10667), .A(n7729), .ZN(n7730) );
  OAI21_X1 U8999 ( .B1(n7731), .B2(n8266), .A(n7730), .ZN(P2_U3164) );
  INV_X1 U9000 ( .A(n7732), .ZN(n7753) );
  OAI222_X1 U9001 ( .A1(P1_U3086), .A2(n9395), .B1(n8202), .B2(n7753), .C1(
        n7733), .C2(n10018), .ZN(P1_U3334) );
  OR2_X1 U9002 ( .A1(n7775), .A2(n7734), .ZN(n9315) );
  NAND2_X1 U9003 ( .A1(n7775), .A2(n7734), .ZN(n9409) );
  NAND2_X1 U9004 ( .A1(n9315), .A2(n9409), .ZN(n7773) );
  AND2_X1 U9005 ( .A1(n9309), .A2(n9308), .ZN(n9411) );
  INV_X1 U9006 ( .A(n9326), .ZN(n7735) );
  AOI21_X1 U9007 ( .B1(n10540), .B2(n9411), .A(n7735), .ZN(n7736) );
  XOR2_X1 U9008 ( .A(n7773), .B(n7736), .Z(n7737) );
  AOI22_X1 U9009 ( .A1(n7737), .A2(n9892), .B1(n9889), .B2(n9567), .ZN(n10589)
         );
  OR2_X1 U9010 ( .A1(n7738), .A2(n7775), .ZN(n7777) );
  INV_X1 U9011 ( .A(n7777), .ZN(n7779) );
  AOI211_X1 U9012 ( .C1(n7775), .C2(n7738), .A(n10512), .B(n7779), .ZN(n7739)
         );
  AOI21_X1 U9013 ( .B1(n9887), .B2(n9565), .A(n7739), .ZN(n10588) );
  INV_X1 U9014 ( .A(n10588), .ZN(n7743) );
  INV_X1 U9015 ( .A(n7775), .ZN(n10590) );
  AOI22_X1 U9016 ( .A1(n10562), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7740), .B2(
        n10551), .ZN(n7741) );
  OAI21_X1 U9017 ( .B1(n10590), .B2(n9879), .A(n7741), .ZN(n7742) );
  AOI21_X1 U9018 ( .B1(n7743), .B2(n10556), .A(n7742), .ZN(n7749) );
  OR2_X1 U9019 ( .A1(n9567), .A2(n7746), .ZN(n7747) );
  XNOR2_X1 U9020 ( .A(n7774), .B(n7773), .ZN(n10592) );
  NAND2_X1 U9021 ( .A1(n10592), .A2(n9815), .ZN(n7748) );
  OAI211_X1 U9022 ( .C1(n10562), .C2(n10589), .A(n7749), .B(n7748), .ZN(
        P1_U3284) );
  NAND2_X1 U9023 ( .A1(n7755), .A2(n9148), .ZN(n7751) );
  NAND2_X1 U9024 ( .A1(n7750), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8520) );
  OAI211_X1 U9025 ( .C1(n7752), .C2(n9153), .A(n7751), .B(n8520), .ZN(P2_U3272) );
  OAI222_X1 U9026 ( .A1(n9153), .A2(n7754), .B1(P2_U3151), .B2(n8339), .C1(
        n9147), .C2(n7753), .ZN(P2_U3274) );
  NAND2_X1 U9027 ( .A1(n7755), .A2(n10015), .ZN(n7756) );
  OAI211_X1 U9028 ( .C1(n7757), .C2(n10018), .A(n7756), .B(n9551), .ZN(
        P1_U3332) );
  INV_X1 U9029 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8540) );
  NOR2_X1 U9030 ( .A1(n7758), .A2(n8814), .ZN(n7760) );
  AOI211_X1 U9031 ( .C1(n8871), .C2(n7795), .A(n7760), .B(n7759), .ZN(n10603)
         );
  INV_X1 U9032 ( .A(n10603), .ZN(n7761) );
  NAND2_X1 U9033 ( .A1(n7761), .A2(n8876), .ZN(n7762) );
  OAI21_X1 U9034 ( .B1(n8876), .B2(n8540), .A(n7762), .ZN(P2_U3469) );
  XOR2_X1 U9035 ( .A(n7765), .B(n7764), .Z(n7766) );
  XNOR2_X1 U9036 ( .A(n7763), .B(n7766), .ZN(n7772) );
  NAND2_X1 U9037 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10246) );
  INV_X1 U9038 ( .A(n10246), .ZN(n7769) );
  INV_X1 U9039 ( .A(n7784), .ZN(n7767) );
  OAI22_X1 U9040 ( .A1(n7914), .A2(n9264), .B1(n9251), .B2(n7767), .ZN(n7768)
         );
  AOI211_X1 U9041 ( .C1(n9261), .C2(n9566), .A(n7769), .B(n7768), .ZN(n7771)
         );
  NAND2_X1 U9042 ( .A1(n7803), .A2(n9266), .ZN(n7770) );
  OAI211_X1 U9043 ( .C1(n7772), .C2(n9268), .A(n7771), .B(n7770), .ZN(P1_U3217) );
  OR2_X1 U9044 ( .A1(n7803), .A2(n7776), .ZN(n9503) );
  NAND2_X1 U9045 ( .A1(n9503), .A2(n9317), .ZN(n9412) );
  XNOR2_X1 U9046 ( .A(n7805), .B(n9412), .ZN(n10600) );
  INV_X1 U9047 ( .A(n10600), .ZN(n7789) );
  INV_X1 U9048 ( .A(n7813), .ZN(n7778) );
  OAI211_X1 U9049 ( .C1(n5154), .C2(n7779), .A(n7778), .B(n10527), .ZN(n10597)
         );
  NAND2_X1 U9050 ( .A1(n9315), .A2(n9326), .ZN(n7781) );
  NAND2_X1 U9051 ( .A1(n9302), .A2(n9303), .ZN(n7780) );
  NOR2_X1 U9052 ( .A1(n7781), .A2(n7780), .ZN(n9499) );
  OR2_X1 U9053 ( .A1(n7781), .A2(n9411), .ZN(n7782) );
  AND2_X1 U9054 ( .A1(n7782), .A2(n9409), .ZN(n9500) );
  INV_X1 U9055 ( .A(n9412), .ZN(n7806) );
  XNOR2_X1 U9056 ( .A(n7807), .B(n7806), .ZN(n7783) );
  AOI222_X1 U9057 ( .A1(n9892), .A2(n7783), .B1(n9564), .B2(n9887), .C1(n9566), 
        .C2(n9889), .ZN(n10598) );
  OAI21_X1 U9058 ( .B1(n9778), .B2(n10597), .A(n10598), .ZN(n7787) );
  AOI22_X1 U9059 ( .A1(n10562), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7784), .B2(
        n10551), .ZN(n7785) );
  OAI21_X1 U9060 ( .B1(n5154), .B2(n9879), .A(n7785), .ZN(n7786) );
  AOI21_X1 U9061 ( .B1(n7787), .B2(n9868), .A(n7786), .ZN(n7788) );
  OAI21_X1 U9062 ( .B1(n7789), .B2(n9896), .A(n7788), .ZN(P1_U3283) );
  XNOR2_X1 U9063 ( .A(n7840), .B(n7790), .ZN(n7842) );
  XNOR2_X1 U9064 ( .A(n7842), .B(n8532), .ZN(n7797) );
  AOI22_X1 U9065 ( .A1(n5136), .A2(n10655), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3151), .ZN(n7792) );
  NAND2_X1 U9066 ( .A1(n10657), .A2(n8531), .ZN(n7791) );
  OAI211_X1 U9067 ( .C1(n10653), .C2(n7793), .A(n7792), .B(n7791), .ZN(n7794)
         );
  AOI21_X1 U9068 ( .B1(n7795), .B2(n10667), .A(n7794), .ZN(n7796) );
  OAI21_X1 U9069 ( .B1(n7797), .B2(n8266), .A(n7796), .ZN(P2_U3157) );
  NOR2_X1 U9070 ( .A1(n7798), .A2(n8844), .ZN(n7853) );
  AOI211_X1 U9071 ( .C1(n7800), .C2(n8872), .A(n7853), .B(n7799), .ZN(n10605)
         );
  INV_X1 U9072 ( .A(n10605), .ZN(n7801) );
  NAND2_X1 U9073 ( .A1(n7801), .A2(n8876), .ZN(n7802) );
  OAI21_X1 U9074 ( .B1(n8876), .B2(n6499), .A(n7802), .ZN(P2_U3470) );
  NOR2_X1 U9075 ( .A1(n7803), .A2(n9565), .ZN(n7804) );
  AND2_X1 U9076 ( .A1(n7981), .A2(n7914), .ZN(n9319) );
  INV_X1 U9077 ( .A(n9319), .ZN(n9325) );
  OR2_X1 U9078 ( .A1(n7981), .A2(n7914), .ZN(n9327) );
  XNOR2_X1 U9079 ( .A(n4977), .B(n9415), .ZN(n10610) );
  NAND2_X1 U9080 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U9081 ( .A1(n7808), .A2(n9317), .ZN(n7880) );
  XNOR2_X1 U9082 ( .A(n7880), .B(n9415), .ZN(n7809) );
  NAND2_X1 U9083 ( .A1(n7809), .A2(n9892), .ZN(n7811) );
  AOI22_X1 U9084 ( .A1(n9565), .A2(n9889), .B1(n9887), .B2(n9563), .ZN(n7810)
         );
  NAND2_X1 U9085 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  AOI21_X1 U9086 ( .B1(n10610), .B2(n10544), .A(n7812), .ZN(n10612) );
  INV_X1 U9087 ( .A(n7981), .ZN(n10607) );
  OAI21_X1 U9088 ( .B1(n7813), .B2(n10607), .A(n10527), .ZN(n7814) );
  OR2_X1 U9089 ( .A1(n7814), .A2(n7889), .ZN(n10606) );
  AOI22_X1 U9090 ( .A1(n10562), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7972), .B2(
        n10551), .ZN(n7816) );
  NAND2_X1 U9091 ( .A1(n7981), .A2(n10552), .ZN(n7815) );
  OAI211_X1 U9092 ( .C1(n10606), .C2(n8103), .A(n7816), .B(n7815), .ZN(n7817)
         );
  AOI21_X1 U9093 ( .B1(n10610), .B2(n10557), .A(n7817), .ZN(n7818) );
  OAI21_X1 U9094 ( .B1(n10612), .B2(n10562), .A(n7818), .ZN(P1_U3282) );
  INV_X1 U9095 ( .A(n7819), .ZN(n7830) );
  OAI222_X1 U9096 ( .A1(n9153), .A2(n7821), .B1(n9147), .B2(n7830), .C1(
        P2_U3151), .C2(n7820), .ZN(P2_U3273) );
  INV_X1 U9097 ( .A(n8398), .ZN(n8495) );
  XNOR2_X1 U9098 ( .A(n7822), .B(n8495), .ZN(n8873) );
  INV_X1 U9099 ( .A(n8873), .ZN(n7829) );
  XNOR2_X1 U9100 ( .A(n7823), .B(n8398), .ZN(n7824) );
  AOI222_X1 U9101 ( .A1(n8793), .A2(n7824), .B1(n8529), .B2(n8797), .C1(n8531), 
        .C2(n8771), .ZN(n8875) );
  OAI21_X1 U9102 ( .B1(n7825), .B2(n10468), .A(n8875), .ZN(n7826) );
  NAND2_X1 U9103 ( .A1(n7826), .A2(n10575), .ZN(n7828) );
  AOI22_X1 U9104 ( .A1(n8870), .A2(n10568), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n10577), .ZN(n7827) );
  OAI211_X1 U9105 ( .C1(n7829), .C2(n8807), .A(n7828), .B(n7827), .ZN(P2_U3221) );
  OAI222_X1 U9106 ( .A1(n7832), .A2(n10018), .B1(P1_U3086), .B2(n7831), .C1(
        n8202), .C2(n7830), .ZN(P1_U3333) );
  XNOR2_X1 U9107 ( .A(n8406), .B(n8529), .ZN(n8496) );
  XNOR2_X1 U9108 ( .A(n7833), .B(n8403), .ZN(n7856) );
  XNOR2_X1 U9109 ( .A(n7834), .B(n8403), .ZN(n7835) );
  OAI222_X1 U9110 ( .A1(n8786), .A2(n7994), .B1(n8801), .B2(n7868), .C1(n7835), 
        .C2(n8723), .ZN(n7858) );
  OAI22_X1 U9111 ( .A1(n8406), .A2(n10469), .B1(n7875), .B2(n10468), .ZN(n7836) );
  OAI21_X1 U9112 ( .B1(n7858), .B2(n7836), .A(n10575), .ZN(n7838) );
  NAND2_X1 U9113 ( .A1(n10577), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7837) );
  OAI211_X1 U9114 ( .C1(n7856), .C2(n8807), .A(n7838), .B(n7837), .ZN(P2_U3220) );
  AOI22_X1 U9115 ( .A1(n7842), .A2(n7841), .B1(n7840), .B2(n7839), .ZN(n7846)
         );
  XNOR2_X1 U9116 ( .A(n7844), .B(n7843), .ZN(n7845) );
  XNOR2_X1 U9117 ( .A(n7846), .B(n7845), .ZN(n7855) );
  NAND2_X1 U9118 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10321) );
  INV_X1 U9119 ( .A(n10321), .ZN(n7848) );
  NOR2_X1 U9120 ( .A1(n10641), .A2(n7868), .ZN(n7847) );
  AOI211_X1 U9121 ( .C1(n10655), .C2(n8532), .A(n7848), .B(n7847), .ZN(n7849)
         );
  OAI21_X1 U9122 ( .B1(n7850), .B2(n10653), .A(n7849), .ZN(n7851) );
  AOI21_X1 U9123 ( .B1(n7853), .B2(n7852), .A(n7851), .ZN(n7854) );
  OAI21_X1 U9124 ( .B1(n7855), .B2(n8266), .A(n7854), .ZN(P2_U3176) );
  OAI22_X1 U9125 ( .A1(n7856), .A2(n8839), .B1(n8406), .B2(n8844), .ZN(n7857)
         );
  NOR2_X1 U9126 ( .A1(n7858), .A2(n7857), .ZN(n10639) );
  INV_X1 U9127 ( .A(n10639), .ZN(n7859) );
  NAND2_X1 U9128 ( .A1(n7859), .A2(n8876), .ZN(n7860) );
  OAI21_X1 U9129 ( .B1(n8876), .B2(n6524), .A(n7860), .ZN(P2_U3472) );
  INV_X1 U9130 ( .A(n7861), .ZN(n7919) );
  OAI222_X1 U9131 ( .A1(P1_U3086), .A2(n7863), .B1(n8202), .B2(n7919), .C1(
        n7862), .C2(n10018), .ZN(P1_U3331) );
  XNOR2_X1 U9132 ( .A(n8406), .B(n8194), .ZN(n7864) );
  NAND2_X1 U9133 ( .A1(n7864), .A2(n8405), .ZN(n7922) );
  OAI21_X1 U9134 ( .B1(n7864), .B2(n8405), .A(n7922), .ZN(n7871) );
  INV_X1 U9135 ( .A(n7867), .ZN(n7869) );
  AOI21_X1 U9136 ( .B1(n7871), .B2(n4995), .A(n7925), .ZN(n7879) );
  NAND2_X1 U9137 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10353) );
  INV_X1 U9138 ( .A(n10353), .ZN(n7873) );
  NOR2_X1 U9139 ( .A1(n10641), .A2(n7994), .ZN(n7872) );
  AOI211_X1 U9140 ( .C1(n10655), .C2(n8530), .A(n7873), .B(n7872), .ZN(n7874)
         );
  OAI21_X1 U9141 ( .B1(n7875), .B2(n10653), .A(n7874), .ZN(n7876) );
  AOI21_X1 U9142 ( .B1(n7877), .B2(n10667), .A(n7876), .ZN(n7878) );
  OAI21_X1 U9143 ( .B1(n7879), .B2(n8266), .A(n7878), .ZN(P2_U3174) );
  NAND2_X1 U9144 ( .A1(n7880), .A2(n9327), .ZN(n7883) );
  INV_X1 U9145 ( .A(n9563), .ZN(n7974) );
  OR2_X1 U9146 ( .A1(n7948), .A2(n7974), .ZN(n9333) );
  NAND2_X1 U9147 ( .A1(n7948), .A2(n7974), .ZN(n9335) );
  NAND2_X1 U9148 ( .A1(n9333), .A2(n9335), .ZN(n7882) );
  NOR2_X1 U9149 ( .A1(n7882), .A2(n9319), .ZN(n7881) );
  NAND2_X1 U9150 ( .A1(n7883), .A2(n7881), .ZN(n7945) );
  INV_X1 U9151 ( .A(n7945), .ZN(n7942) );
  INV_X1 U9152 ( .A(n7882), .ZN(n9416) );
  AOI21_X1 U9153 ( .B1(n7883), .B2(n9325), .A(n9416), .ZN(n7884) );
  NOR3_X1 U9154 ( .A1(n7942), .A2(n7884), .A3(n10539), .ZN(n7886) );
  OAI22_X1 U9155 ( .A1(n7914), .A2(n10533), .B1(n8053), .B2(n10531), .ZN(n7885) );
  NOR2_X1 U9156 ( .A1(n7886), .A2(n7885), .ZN(n10616) );
  XNOR2_X1 U9157 ( .A(n7950), .B(n9416), .ZN(n10619) );
  NAND2_X1 U9158 ( .A1(n10619), .A2(n9815), .ZN(n7893) );
  INV_X1 U9159 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7888) );
  INV_X1 U9160 ( .A(n7887), .ZN(n7913) );
  OAI22_X1 U9161 ( .A1(n9868), .A2(n7888), .B1(n7913), .B2(n10448), .ZN(n7891)
         );
  OAI211_X1 U9162 ( .C1(n7889), .C2(n10617), .A(n10527), .B(n7953), .ZN(n10615) );
  NOR2_X1 U9163 ( .A1(n10615), .A2(n8103), .ZN(n7890) );
  AOI211_X1 U9164 ( .C1(n10552), .C2(n7948), .A(n7891), .B(n7890), .ZN(n7892)
         );
  OAI211_X1 U9165 ( .C1(n10562), .C2(n10616), .A(n7893), .B(n7892), .ZN(
        P1_U3281) );
  INV_X1 U9166 ( .A(n7894), .ZN(n7907) );
  OAI222_X1 U9167 ( .A1(P1_U3086), .A2(n7896), .B1(n8202), .B2(n7907), .C1(
        n7895), .C2(n10018), .ZN(P1_U3330) );
  OAI21_X1 U9168 ( .B1(n4979), .B2(n8478), .A(n7897), .ZN(n7941) );
  AND2_X1 U9169 ( .A1(n7898), .A2(n8478), .ZN(n7899) );
  OAI21_X1 U9170 ( .B1(n7900), .B2(n7899), .A(n8793), .ZN(n7902) );
  AOI22_X1 U9171 ( .A1(n8771), .A2(n8529), .B1(n8527), .B2(n8797), .ZN(n7901)
         );
  AND2_X1 U9172 ( .A1(n7902), .A2(n7901), .ZN(n7936) );
  OAI21_X1 U9173 ( .B1(n7933), .B2(n10469), .A(n7936), .ZN(n7903) );
  NAND2_X1 U9174 ( .A1(n7903), .A2(n10575), .ZN(n7906) );
  INV_X1 U9175 ( .A(n7904), .ZN(n7930) );
  AOI22_X1 U9176 ( .A1(n10577), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10572), 
        .B2(n7930), .ZN(n7905) );
  OAI211_X1 U9177 ( .C1(n7941), .C2(n8807), .A(n7906), .B(n7905), .ZN(P2_U3219) );
  OAI222_X1 U9178 ( .A1(n9153), .A2(n7908), .B1(P2_U3151), .B2(n6704), .C1(
        n9147), .C2(n7907), .ZN(P2_U3270) );
  AOI21_X1 U9179 ( .B1(n7909), .B2(n7978), .A(n7910), .ZN(n7912) );
  OAI21_X1 U9180 ( .B1(n7912), .B2(n7911), .A(n9235), .ZN(n7918) );
  OAI22_X1 U9181 ( .A1(n9250), .A2(n7914), .B1(n7913), .B2(n9251), .ZN(n7915)
         );
  AOI211_X1 U9182 ( .C1(n9213), .C2(n9562), .A(n7916), .B(n7915), .ZN(n7917)
         );
  OAI211_X1 U9183 ( .C1(n10617), .C2(n9243), .A(n7918), .B(n7917), .ZN(
        P1_U3224) );
  OAI222_X1 U9184 ( .A1(n9153), .A2(n7921), .B1(P2_U3151), .B2(n7920), .C1(
        n9147), .C2(n7919), .ZN(P2_U3271) );
  INV_X1 U9185 ( .A(n7922), .ZN(n7924) );
  XNOR2_X1 U9186 ( .A(n7934), .B(n8194), .ZN(n7986) );
  XNOR2_X1 U9187 ( .A(n7986), .B(n7994), .ZN(n7923) );
  NOR3_X1 U9188 ( .A1(n7925), .A2(n7924), .A3(n7923), .ZN(n7926) );
  OAI21_X1 U9189 ( .B1(n5408), .B2(n7926), .A(n10665), .ZN(n7932) );
  NAND2_X1 U9190 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n10369) );
  INV_X1 U9191 ( .A(n10369), .ZN(n7927) );
  AOI21_X1 U9192 ( .B1(n10655), .B2(n8529), .A(n7927), .ZN(n7928) );
  OAI21_X1 U9193 ( .B1(n8044), .B2(n10641), .A(n7928), .ZN(n7929) );
  AOI21_X1 U9194 ( .B1(n10670), .B2(n7930), .A(n7929), .ZN(n7931) );
  OAI211_X1 U9195 ( .C1(n7933), .C2(n8277), .A(n7932), .B(n7931), .ZN(P2_U3155) );
  INV_X1 U9196 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U9197 ( .A1(n7934), .A2(n8871), .ZN(n7935) );
  AND2_X1 U9198 ( .A1(n7936), .A2(n7935), .ZN(n7939) );
  MUX2_X1 U9199 ( .A(n7937), .B(n7939), .S(n10640), .Z(n7938) );
  OAI21_X1 U9200 ( .B1(n7941), .B2(n9134), .A(n7938), .ZN(P2_U3432) );
  MUX2_X1 U9201 ( .A(n8550), .B(n7939), .S(n8876), .Z(n7940) );
  OAI21_X1 U9202 ( .B1(n8865), .B2(n7941), .A(n7940), .ZN(P2_U3473) );
  INV_X1 U9203 ( .A(n9333), .ZN(n7943) );
  OR2_X1 U9204 ( .A1(n8002), .A2(n8053), .ZN(n9510) );
  NAND2_X1 U9205 ( .A1(n8002), .A2(n8053), .ZN(n9336) );
  NAND2_X1 U9206 ( .A1(n9510), .A2(n9336), .ZN(n9418) );
  OAI21_X1 U9207 ( .B1(n7942), .B2(n7943), .A(n9418), .ZN(n7946) );
  NOR2_X1 U9208 ( .A1(n9418), .A2(n7943), .ZN(n7944) );
  NAND2_X1 U9209 ( .A1(n7945), .A2(n7944), .ZN(n8021) );
  NAND2_X1 U9210 ( .A1(n7946), .A2(n8021), .ZN(n7947) );
  AOI222_X1 U9211 ( .A1(n9892), .A2(n7947), .B1(n9561), .B2(n9887), .C1(n9563), 
        .C2(n9889), .ZN(n10624) );
  AND2_X1 U9212 ( .A1(n7948), .A2(n9563), .ZN(n7949) );
  XOR2_X1 U9213 ( .A(n9418), .B(n4928), .Z(n10629) );
  NAND2_X1 U9214 ( .A1(n10629), .A2(n9815), .ZN(n7957) );
  INV_X1 U9215 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7952) );
  INV_X1 U9216 ( .A(n7951), .ZN(n7962) );
  OAI22_X1 U9217 ( .A1(n9868), .A2(n7952), .B1(n7962), .B2(n10448), .ZN(n7955)
         );
  INV_X1 U9218 ( .A(n8006), .ZN(n8031) );
  OAI211_X1 U9219 ( .C1(n5151), .C2(n10626), .A(n10527), .B(n8031), .ZN(n10623) );
  NOR2_X1 U9220 ( .A1(n10623), .A2(n8103), .ZN(n7954) );
  AOI211_X1 U9221 ( .C1(n10552), .C2(n8002), .A(n7955), .B(n7954), .ZN(n7956)
         );
  OAI211_X1 U9222 ( .C1(n10562), .C2(n10624), .A(n7957), .B(n7956), .ZN(
        P1_U3280) );
  OAI21_X1 U9223 ( .B1(n7911), .B2(n7959), .A(n7958), .ZN(n7960) );
  NAND3_X1 U9224 ( .A1(n4971), .A2(n9235), .A3(n7960), .ZN(n7965) );
  NOR2_X1 U9225 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7961), .ZN(n10230) );
  OAI22_X1 U9226 ( .A1(n8004), .A2(n9264), .B1(n9251), .B2(n7962), .ZN(n7963)
         );
  AOI211_X1 U9227 ( .C1(n9261), .C2(n9563), .A(n10230), .B(n7963), .ZN(n7964)
         );
  OAI211_X1 U9228 ( .C1(n10626), .C2(n9243), .A(n7965), .B(n7964), .ZN(
        P1_U3234) );
  XNOR2_X1 U9229 ( .A(n8866), .B(n8527), .ZN(n8497) );
  XNOR2_X1 U9230 ( .A(n4974), .B(n8497), .ZN(n7966) );
  INV_X1 U9231 ( .A(n7994), .ZN(n8528) );
  INV_X1 U9232 ( .A(n8802), .ZN(n8526) );
  AOI222_X1 U9233 ( .A1(n8793), .A2(n7966), .B1(n8528), .B2(n8771), .C1(n8526), 
        .C2(n8797), .ZN(n8869) );
  XOR2_X1 U9234 ( .A(n7967), .B(n8497), .Z(n8867) );
  NOR2_X1 U9235 ( .A1(n7999), .A2(n8649), .ZN(n7970) );
  OAI22_X1 U9236 ( .A1(n10575), .A2(n7968), .B1(n7991), .B2(n10468), .ZN(n7969) );
  AOI211_X1 U9237 ( .C1(n8867), .C2(n8752), .A(n7970), .B(n7969), .ZN(n7971)
         );
  OAI21_X1 U9238 ( .B1(n8869), .B2(n10577), .A(n7971), .ZN(P2_U3218) );
  AOI22_X1 U9239 ( .A1(n9262), .A2(n7972), .B1(n9261), .B2(n9565), .ZN(n7973)
         );
  NAND2_X1 U9240 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10164) );
  OAI211_X1 U9241 ( .C1(n7974), .C2(n9264), .A(n7973), .B(n10164), .ZN(n7980)
         );
  AOI21_X1 U9242 ( .B1(n7976), .B2(n7978), .A(n7975), .ZN(n7977) );
  AOI211_X1 U9243 ( .C1(n5186), .C2(n7978), .A(n9268), .B(n7977), .ZN(n7979)
         );
  AOI211_X1 U9244 ( .C1(n7981), .C2(n9266), .A(n7980), .B(n7979), .ZN(n7982)
         );
  INV_X1 U9245 ( .A(n7982), .ZN(P1_U3236) );
  INV_X1 U9246 ( .A(n7983), .ZN(n8000) );
  AOI21_X1 U9247 ( .B1(n9141), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7984), .ZN(
        n7985) );
  OAI21_X1 U9248 ( .B1(n8000), .B2(n9147), .A(n7985), .ZN(P2_U3268) );
  XNOR2_X1 U9249 ( .A(n8866), .B(n8194), .ZN(n8037) );
  XNOR2_X1 U9250 ( .A(n8037), .B(n8527), .ZN(n7988) );
  AOI21_X1 U9251 ( .B1(n7989), .B2(n7988), .A(n8266), .ZN(n7990) );
  NAND2_X1 U9252 ( .A1(n7990), .A2(n8039), .ZN(n7998) );
  INV_X1 U9253 ( .A(n7991), .ZN(n7996) );
  NAND2_X1 U9254 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10384) );
  INV_X1 U9255 ( .A(n10384), .ZN(n7992) );
  AOI21_X1 U9256 ( .B1(n10657), .B2(n8526), .A(n7992), .ZN(n7993) );
  OAI21_X1 U9257 ( .B1(n7994), .B2(n10644), .A(n7993), .ZN(n7995) );
  AOI21_X1 U9258 ( .B1(n7996), .B2(n10670), .A(n7995), .ZN(n7997) );
  OAI211_X1 U9259 ( .C1(n7999), .C2(n8277), .A(n7998), .B(n7997), .ZN(P2_U3181) );
  OAI222_X1 U9260 ( .A1(n10025), .A2(n8001), .B1(n8202), .B2(n8000), .C1(n8162), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI21_X1 U9261 ( .B1(n8002), .B2(n9562), .A(n4928), .ZN(n8003) );
  OAI21_X1 U9262 ( .B1(n10626), .B2(n8053), .A(n8003), .ZN(n8024) );
  NAND2_X1 U9263 ( .A1(n9986), .A2(n8004), .ZN(n9340) );
  NAND2_X1 U9264 ( .A1(n9511), .A2(n9340), .ZN(n8023) );
  INV_X1 U9265 ( .A(n9980), .ZN(n8096) );
  AND2_X1 U9266 ( .A1(n8096), .A2(n9560), .ZN(n9514) );
  INV_X1 U9267 ( .A(n9560), .ZN(n8126) );
  NAND2_X1 U9268 ( .A1(n9980), .A2(n8126), .ZN(n9346) );
  NOR2_X1 U9269 ( .A1(n9514), .A2(n5300), .ZN(n9420) );
  XNOR2_X1 U9270 ( .A(n8097), .B(n9420), .ZN(n9984) );
  AOI21_X1 U9271 ( .B1(n9980), .B2(n8029), .A(n8102), .ZN(n9981) );
  AOI22_X1 U9272 ( .A1(n10562), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8061), .B2(
        n10551), .ZN(n8007) );
  OAI21_X1 U9273 ( .B1(n8096), .B2(n9879), .A(n8007), .ZN(n8013) );
  INV_X1 U9274 ( .A(n9336), .ZN(n8008) );
  NOR2_X1 U9275 ( .A1(n8023), .A2(n8008), .ZN(n8009) );
  NAND2_X1 U9276 ( .A1(n8021), .A2(n8009), .ZN(n8010) );
  XOR2_X1 U9277 ( .A(n8094), .B(n9420), .Z(n8011) );
  INV_X1 U9278 ( .A(n8108), .ZN(n9559) );
  AOI222_X1 U9279 ( .A1(n9892), .A2(n8011), .B1(n9559), .B2(n9887), .C1(n9561), 
        .C2(n9889), .ZN(n9983) );
  NOR2_X1 U9280 ( .A1(n9983), .A2(n10562), .ZN(n8012) );
  AOI211_X1 U9281 ( .C1(n9981), .C2(n9855), .A(n8013), .B(n8012), .ZN(n8014)
         );
  OAI21_X1 U9282 ( .B1(n9984), .B2(n9896), .A(n8014), .ZN(P1_U3278) );
  INV_X1 U9283 ( .A(n8015), .ZN(n8019) );
  OAI222_X1 U9284 ( .A1(n10025), .A2(n8017), .B1(n8202), .B2(n8019), .C1(
        P1_U3086), .C2(n8016), .ZN(P1_U3329) );
  OAI222_X1 U9285 ( .A1(n9153), .A2(n8020), .B1(n9147), .B2(n8019), .C1(n8018), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  NAND2_X1 U9286 ( .A1(n8021), .A2(n9336), .ZN(n8022) );
  INV_X1 U9287 ( .A(n8023), .ZN(n9421) );
  XNOR2_X1 U9288 ( .A(n8022), .B(n9421), .ZN(n8028) );
  OAI22_X1 U9289 ( .A1(n8053), .A2(n10533), .B1(n8126), .B2(n10531), .ZN(n8027) );
  XNOR2_X1 U9290 ( .A(n8024), .B(n8023), .ZN(n9989) );
  NOR2_X1 U9291 ( .A1(n9989), .A2(n8025), .ZN(n8026) );
  AOI211_X1 U9292 ( .C1(n8028), .C2(n9892), .A(n8027), .B(n8026), .ZN(n9988)
         );
  INV_X1 U9293 ( .A(n8029), .ZN(n8030) );
  AOI211_X1 U9294 ( .C1(n9986), .C2(n8031), .A(n10512), .B(n8030), .ZN(n9985)
         );
  AOI22_X1 U9295 ( .A1(n10562), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8051), .B2(
        n10551), .ZN(n8032) );
  OAI21_X1 U9296 ( .B1(n8005), .B2(n9879), .A(n8032), .ZN(n8035) );
  NOR2_X1 U9297 ( .A1(n9989), .A2(n8033), .ZN(n8034) );
  AOI211_X1 U9298 ( .C1(n9985), .C2(n10556), .A(n8035), .B(n8034), .ZN(n8036)
         );
  OAI21_X1 U9299 ( .B1(n9988), .B2(n10562), .A(n8036), .ZN(P1_U3279) );
  NAND2_X1 U9300 ( .A1(n8037), .A2(n8527), .ZN(n8038) );
  NAND2_X1 U9301 ( .A1(n8039), .A2(n8038), .ZN(n8079) );
  XNOR2_X1 U9302 ( .A(n8862), .B(n8194), .ZN(n8081) );
  XNOR2_X1 U9303 ( .A(n8081), .B(n8802), .ZN(n8080) );
  XNOR2_X1 U9304 ( .A(n8040), .B(n8080), .ZN(n8047) );
  NAND2_X1 U9305 ( .A1(n10670), .A2(n8071), .ZN(n8043) );
  NAND2_X1 U9306 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10400) );
  INV_X1 U9307 ( .A(n10400), .ZN(n8041) );
  AOI21_X1 U9308 ( .B1(n10657), .B2(n8525), .A(n8041), .ZN(n8042) );
  OAI211_X1 U9309 ( .C1(n8044), .C2(n10644), .A(n8043), .B(n8042), .ZN(n8045)
         );
  AOI21_X1 U9310 ( .B1(n8862), .B2(n10667), .A(n8045), .ZN(n8046) );
  OAI21_X1 U9311 ( .B1(n8047), .B2(n8266), .A(n8046), .ZN(P2_U3166) );
  NAND2_X1 U9312 ( .A1(n4973), .A2(n8048), .ZN(n8050) );
  XNOR2_X1 U9313 ( .A(n8050), .B(n8049), .ZN(n8056) );
  AOI22_X1 U9314 ( .A1(n9213), .A2(n9560), .B1(n9262), .B2(n8051), .ZN(n8052)
         );
  NAND2_X1 U9315 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10179) );
  OAI211_X1 U9316 ( .C1(n8053), .C2(n9250), .A(n8052), .B(n10179), .ZN(n8054)
         );
  AOI21_X1 U9317 ( .B1(n9986), .B2(n9266), .A(n8054), .ZN(n8055) );
  OAI21_X1 U9318 ( .B1(n8056), .B2(n9268), .A(n8055), .ZN(P1_U3215) );
  XNOR2_X1 U9319 ( .A(n8058), .B(n8057), .ZN(n8059) );
  XNOR2_X1 U9320 ( .A(n8060), .B(n8059), .ZN(n8065) );
  AOI22_X1 U9321 ( .A1(n9262), .A2(n8061), .B1(n9261), .B2(n9561), .ZN(n8062)
         );
  NAND2_X1 U9322 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10191) );
  OAI211_X1 U9323 ( .C1(n8108), .C2(n9264), .A(n8062), .B(n10191), .ZN(n8063)
         );
  AOI21_X1 U9324 ( .B1(n9980), .B2(n9266), .A(n8063), .ZN(n8064) );
  OAI21_X1 U9325 ( .B1(n8065), .B2(n9268), .A(n8064), .ZN(P1_U3241) );
  OAI211_X1 U9326 ( .C1(n8068), .C2(n8067), .A(n8066), .B(n8793), .ZN(n8070)
         );
  AOI22_X1 U9327 ( .A1(n8525), .A2(n8797), .B1(n8771), .B2(n8527), .ZN(n8069)
         );
  NAND2_X1 U9328 ( .A1(n8070), .A2(n8069), .ZN(n8861) );
  AOI21_X1 U9329 ( .B1(n10572), .B2(n8071), .A(n8861), .ZN(n8078) );
  XNOR2_X1 U9330 ( .A(n8072), .B(n8499), .ZN(n9135) );
  INV_X1 U9331 ( .A(n9135), .ZN(n8076) );
  OAI22_X1 U9332 ( .A1(n8074), .A2(n8649), .B1(n8073), .B2(n10575), .ZN(n8075)
         );
  AOI21_X1 U9333 ( .B1(n8076), .B2(n8752), .A(n8075), .ZN(n8077) );
  OAI21_X1 U9334 ( .B1(n8078), .B2(n10577), .A(n8077), .ZN(P2_U3217) );
  INV_X1 U9335 ( .A(n8079), .ZN(n8084) );
  INV_X1 U9336 ( .A(n8080), .ZN(n8083) );
  INV_X1 U9337 ( .A(n8081), .ZN(n8082) );
  XNOR2_X1 U9338 ( .A(n8858), .B(n8194), .ZN(n8086) );
  NAND2_X1 U9339 ( .A1(n8086), .A2(n8525), .ZN(n8168) );
  NAND2_X1 U9340 ( .A1(n4919), .A2(n8168), .ZN(n8087) );
  XNOR2_X1 U9341 ( .A(n8085), .B(n8087), .ZN(n8093) );
  NAND2_X1 U9342 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10421) );
  INV_X1 U9343 ( .A(n10421), .ZN(n8089) );
  NOR2_X1 U9344 ( .A1(n10641), .A2(n8222), .ZN(n8088) );
  AOI211_X1 U9345 ( .C1(n10655), .C2(n8526), .A(n8089), .B(n8088), .ZN(n8090)
         );
  OAI21_X1 U9346 ( .B1(n8803), .B2(n10653), .A(n8090), .ZN(n8091) );
  AOI21_X1 U9347 ( .B1(n8858), .B2(n10667), .A(n8091), .ZN(n8092) );
  OAI21_X1 U9348 ( .B1(n8093), .B2(n8266), .A(n8092), .ZN(P2_U3168) );
  OR2_X1 U9349 ( .A1(n9975), .A2(n8108), .ZN(n9517) );
  NAND2_X1 U9350 ( .A1(n9975), .A2(n8108), .ZN(n9347) );
  NAND2_X1 U9351 ( .A1(n9517), .A2(n9347), .ZN(n8098) );
  XNOR2_X1 U9352 ( .A(n8110), .B(n5444), .ZN(n8095) );
  INV_X1 U9353 ( .A(n9674), .ZN(n9890) );
  AOI222_X1 U9354 ( .A1(n9892), .A2(n8095), .B1(n9890), .B2(n9887), .C1(n9560), 
        .C2(n9889), .ZN(n9978) );
  OR2_X1 U9355 ( .A1(n8099), .A2(n8098), .ZN(n9974) );
  NAND3_X1 U9356 ( .A1(n9974), .A2(n9973), .A3(n9815), .ZN(n8107) );
  INV_X1 U9357 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8101) );
  INV_X1 U9358 ( .A(n8100), .ZN(n8125) );
  OAI22_X1 U9359 ( .A1(n9868), .A2(n8101), .B1(n8125), .B2(n10448), .ZN(n8105)
         );
  NAND2_X1 U9360 ( .A1(n8102), .A2(n8130), .ZN(n8116) );
  OAI211_X1 U9361 ( .C1(n8102), .C2(n8130), .A(n8116), .B(n10527), .ZN(n9977)
         );
  NOR2_X1 U9362 ( .A1(n9977), .A2(n8103), .ZN(n8104) );
  AOI211_X1 U9363 ( .C1(n10552), .C2(n9975), .A(n8105), .B(n8104), .ZN(n8106)
         );
  OAI211_X1 U9364 ( .C1(n10562), .C2(n9978), .A(n8107), .B(n8106), .ZN(
        P1_U3277) );
  OR2_X1 U9365 ( .A1(n9970), .A2(n9674), .ZN(n9518) );
  NAND2_X1 U9366 ( .A1(n9970), .A2(n9674), .ZN(n9357) );
  NAND2_X1 U9367 ( .A1(n9518), .A2(n9357), .ZN(n9423) );
  OAI21_X1 U9368 ( .B1(n8109), .B2(n9423), .A(n9676), .ZN(n9972) );
  INV_X1 U9369 ( .A(n9347), .ZN(n9519) );
  INV_X1 U9370 ( .A(n9423), .ZN(n9353) );
  NAND3_X1 U9371 ( .A1(n8112), .A2(n9423), .A3(n9517), .ZN(n8113) );
  NAND3_X1 U9372 ( .A1(n9881), .A2(n9892), .A3(n8113), .ZN(n8115) );
  NAND2_X1 U9373 ( .A1(n9559), .A2(n9889), .ZN(n8114) );
  OAI211_X1 U9374 ( .C1(n9866), .C2(n10531), .A(n8115), .B(n8114), .ZN(n9969)
         );
  INV_X1 U9375 ( .A(n9970), .ZN(n9675) );
  NOR2_X2 U9376 ( .A1(n8116), .A2(n9970), .ZN(n9873) );
  AOI211_X1 U9377 ( .C1(n9970), .C2(n8116), .A(n10512), .B(n9873), .ZN(n9968)
         );
  NAND2_X1 U9378 ( .A1(n9968), .A2(n10556), .ZN(n8118) );
  AOI22_X1 U9379 ( .A1(n10562), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9219), .B2(
        n10551), .ZN(n8117) );
  OAI211_X1 U9380 ( .C1(n9675), .C2(n9879), .A(n8118), .B(n8117), .ZN(n8119)
         );
  AOI21_X1 U9381 ( .B1(n9868), .B2(n9969), .A(n8119), .ZN(n8120) );
  OAI21_X1 U9382 ( .B1(n9972), .B2(n9896), .A(n8120), .ZN(P1_U3276) );
  OAI21_X1 U9383 ( .B1(n8123), .B2(n8122), .A(n8121), .ZN(n8124) );
  NAND2_X1 U9384 ( .A1(n8124), .A2(n9235), .ZN(n8129) );
  AND2_X1 U9385 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9630) );
  OAI22_X1 U9386 ( .A1(n9250), .A2(n8126), .B1(n8125), .B2(n9251), .ZN(n8127)
         );
  AOI211_X1 U9387 ( .C1(n9213), .C2(n9890), .A(n9630), .B(n8127), .ZN(n8128)
         );
  OAI211_X1 U9388 ( .C1(n8130), .C2(n9243), .A(n8129), .B(n8128), .ZN(P1_U3226) );
  AOI22_X1 U9389 ( .A1(n8131), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n9141), .ZN(n8132) );
  OAI21_X1 U9390 ( .B1(n8133), .B2(n9147), .A(n8132), .ZN(P2_U3289) );
  NAND2_X1 U9391 ( .A1(n8135), .A2(n8134), .ZN(n8140) );
  INV_X1 U9392 ( .A(n8136), .ZN(n8138) );
  NAND2_X1 U9393 ( .A1(n8138), .A2(n8137), .ZN(n8139) );
  NAND2_X1 U9394 ( .A1(n8140), .A2(n8139), .ZN(n8144) );
  MUX2_X1 U9395 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n8141), .Z(n8142) );
  NAND2_X1 U9396 ( .A1(n8152), .A2(SI_29_), .ZN(n8146) );
  INV_X1 U9397 ( .A(n8142), .ZN(n8143) );
  OR2_X1 U9398 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  NAND2_X1 U9399 ( .A1(n8146), .A2(n8145), .ZN(n8285) );
  INV_X1 U9400 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10019) );
  INV_X1 U9401 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8280) );
  MUX2_X1 U9402 ( .A(n10019), .B(n8280), .S(n8286), .Z(n8147) );
  NAND2_X1 U9403 ( .A1(n8147), .A2(n9010), .ZN(n8283) );
  INV_X1 U9404 ( .A(n8147), .ZN(n8148) );
  NAND2_X1 U9405 ( .A1(n8148), .A2(SI_30_), .ZN(n8149) );
  NAND2_X1 U9406 ( .A1(n8283), .A2(n8149), .ZN(n8284) );
  XNOR2_X1 U9407 ( .A(n8285), .B(n8284), .ZN(n8279) );
  NOR2_X1 U9408 ( .A1(n5778), .A2(n10019), .ZN(n8150) );
  AOI21_X2 U9409 ( .B1(n8279), .B2(n9273), .A(n8150), .ZN(n9667) );
  INV_X1 U9410 ( .A(SI_29_), .ZN(n8151) );
  XNOR2_X1 U9411 ( .A(n8152), .B(n8151), .ZN(n9144) );
  NAND2_X1 U9412 ( .A1(n9144), .A2(n9273), .ZN(n8154) );
  INV_X1 U9413 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10024) );
  OR2_X1 U9414 ( .A1(n5778), .A2(n10024), .ZN(n8153) );
  NAND2_X1 U9415 ( .A1(n9149), .A2(n9273), .ZN(n8156) );
  INV_X1 U9416 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8203) );
  OR2_X1 U9417 ( .A1(n5778), .A2(n8203), .ZN(n8155) );
  INV_X1 U9418 ( .A(n9934), .ZN(n9682) );
  NAND2_X1 U9419 ( .A1(n9873), .A2(n9880), .ZN(n9874) );
  NAND2_X1 U9420 ( .A1(n9858), .A2(n9849), .ZN(n9843) );
  NOR2_X2 U9421 ( .A1(n9843), .A2(n9950), .ZN(n9835) );
  NAND2_X1 U9422 ( .A1(n9757), .A2(n9766), .ZN(n9751) );
  NOR2_X2 U9423 ( .A1(n9751), .A2(n9916), .ZN(n9733) );
  NAND2_X1 U9424 ( .A1(n9722), .A2(n9733), .ZN(n9717) );
  NOR2_X2 U9425 ( .A1(n9907), .A2(n9717), .ZN(n9687) );
  XNOR2_X1 U9426 ( .A(n9667), .B(n9687), .ZN(n8157) );
  NAND2_X1 U9427 ( .A1(n9900), .A2(n10556), .ZN(n8166) );
  NAND2_X1 U9428 ( .A1(n4916), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U9429 ( .A1(n5786), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U9430 ( .A1(n4918), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8158) );
  NAND3_X1 U9431 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(n9556) );
  INV_X1 U9432 ( .A(n9556), .ZN(n9392) );
  INV_X1 U9433 ( .A(P1_B_REG_SCAN_IN), .ZN(n8161) );
  NOR2_X1 U9434 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  OR2_X1 U9435 ( .A1(n10531), .A2(n8163), .ZN(n9707) );
  NOR2_X1 U9436 ( .A1(n9392), .A2(n9707), .ZN(n9901) );
  INV_X1 U9437 ( .A(n9901), .ZN(n8164) );
  NOR2_X1 U9438 ( .A1(n10562), .A2(n8164), .ZN(n9671) );
  AOI21_X1 U9439 ( .B1(n10562), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9671), .ZN(
        n8165) );
  OAI211_X1 U9440 ( .C1(n9667), .C2(n9879), .A(n8166), .B(n8165), .ZN(P1_U3264) );
  XNOR2_X1 U9441 ( .A(n10649), .B(n8194), .ZN(n8170) );
  XNOR2_X1 U9442 ( .A(n8170), .B(n8798), .ZN(n10647) );
  XNOR2_X1 U9443 ( .A(n8768), .B(n8194), .ZN(n8219) );
  XNOR2_X1 U9444 ( .A(n8171), .B(n8194), .ZN(n8172) );
  NOR2_X1 U9445 ( .A1(n8172), .A2(n8233), .ZN(n10660) );
  NAND2_X1 U9446 ( .A1(n8172), .A2(n8233), .ZN(n10661) );
  OAI21_X1 U9447 ( .B1(n10659), .B2(n10660), .A(n10661), .ZN(n8232) );
  XNOR2_X1 U9448 ( .A(n8749), .B(n8194), .ZN(n8173) );
  NOR2_X1 U9449 ( .A1(n8173), .A2(n6594), .ZN(n8228) );
  NAND2_X1 U9450 ( .A1(n8173), .A2(n6594), .ZN(n8229) );
  XNOR2_X1 U9451 ( .A(n8835), .B(n8194), .ZN(n8175) );
  XNOR2_X1 U9452 ( .A(n8175), .B(n8724), .ZN(n8256) );
  NAND2_X1 U9453 ( .A1(n8175), .A2(n8744), .ZN(n8176) );
  NAND2_X1 U9454 ( .A1(n8255), .A2(n8176), .ZN(n8179) );
  XNOR2_X1 U9455 ( .A(n8832), .B(n7050), .ZN(n8177) );
  XNOR2_X1 U9456 ( .A(n8179), .B(n8177), .ZN(n8213) );
  NAND2_X1 U9457 ( .A1(n8213), .A2(n8732), .ZN(n8212) );
  INV_X1 U9458 ( .A(n8177), .ZN(n8178) );
  NAND2_X1 U9459 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  XNOR2_X1 U9460 ( .A(n8715), .B(n8194), .ZN(n8182) );
  XNOR2_X1 U9461 ( .A(n8182), .B(n8725), .ZN(n8249) );
  NAND2_X1 U9462 ( .A1(n8182), .A2(n8725), .ZN(n8183) );
  XNOR2_X1 U9463 ( .A(n8824), .B(n8194), .ZN(n8184) );
  XNOR2_X1 U9464 ( .A(n8184), .B(n8712), .ZN(n8240) );
  INV_X1 U9465 ( .A(n8184), .ZN(n8185) );
  NAND2_X1 U9466 ( .A1(n8185), .A2(n8712), .ZN(n8186) );
  NAND2_X1 U9467 ( .A1(n8187), .A2(n8186), .ZN(n8265) );
  INV_X1 U9468 ( .A(n8265), .ZN(n8189) );
  XNOR2_X1 U9469 ( .A(n8820), .B(n8194), .ZN(n8190) );
  XNOR2_X1 U9470 ( .A(n8190), .B(n8522), .ZN(n8267) );
  NAND2_X1 U9471 ( .A1(n8189), .A2(n8188), .ZN(n8268) );
  NAND2_X1 U9472 ( .A1(n8190), .A2(n8522), .ZN(n8191) );
  XNOR2_X1 U9473 ( .A(n8680), .B(n7050), .ZN(n8192) );
  NOR2_X1 U9474 ( .A1(n8192), .A2(n8272), .ZN(n8193) );
  AOI21_X1 U9475 ( .B1(n8272), .B2(n8192), .A(n8193), .ZN(n8206) );
  XNOR2_X1 U9476 ( .A(n8653), .B(n8194), .ZN(n8195) );
  NOR2_X1 U9477 ( .A1(n10653), .A2(n8667), .ZN(n8198) );
  AOI22_X1 U9478 ( .A1(n10655), .A2(n8688), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8196) );
  OAI21_X1 U9479 ( .B1(n8317), .B2(n10641), .A(n8196), .ZN(n8197) );
  AOI211_X1 U9480 ( .C1(n8672), .C2(n10667), .A(n8198), .B(n8197), .ZN(n8199)
         );
  OAI21_X1 U9481 ( .B1(n8200), .B2(n8266), .A(n8199), .ZN(P2_U3160) );
  INV_X1 U9482 ( .A(n9149), .ZN(n8201) );
  OAI222_X1 U9483 ( .A1(n10025), .A2(n8203), .B1(n8202), .B2(n8201), .C1(n4908), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U9484 ( .A(n8279), .ZN(n10020) );
  OAI222_X1 U9485 ( .A1(n9153), .A2(n8280), .B1(n9147), .B2(n10020), .C1(n8204), .C2(P2_U3151), .ZN(P2_U3265) );
  INV_X1 U9486 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9068) );
  OAI22_X1 U9487 ( .A1(n10641), .A2(n8326), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9068), .ZN(n8209) );
  NOR2_X1 U9488 ( .A1(n10653), .A2(n8675), .ZN(n8208) );
  AOI211_X1 U9489 ( .C1(n10655), .C2(n8522), .A(n8209), .B(n8208), .ZN(n8210)
         );
  OAI211_X1 U9490 ( .C1(n8213), .C2(n8732), .A(n8212), .B(n10665), .ZN(n8217)
         );
  OAI22_X1 U9491 ( .A1(n10644), .A2(n8724), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9075), .ZN(n8215) );
  NOR2_X1 U9492 ( .A1(n10653), .A2(n8726), .ZN(n8214) );
  AOI211_X1 U9493 ( .C1(n10657), .C2(n8524), .A(n8215), .B(n8214), .ZN(n8216)
         );
  OAI211_X1 U9494 ( .C1(n8218), .C2(n8277), .A(n8217), .B(n8216), .ZN(P2_U3156) );
  INV_X1 U9495 ( .A(n8851), .ZN(n8227) );
  OAI211_X1 U9496 ( .C1(n4972), .C2(n5423), .A(n10665), .B(n8220), .ZN(n8226)
         );
  INV_X1 U9497 ( .A(n8775), .ZN(n8224) );
  AND2_X1 U9498 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8632) );
  AOI21_X1 U9499 ( .B1(n10657), .B2(n8770), .A(n8632), .ZN(n8221) );
  OAI21_X1 U9500 ( .B1(n8222), .B2(n10644), .A(n8221), .ZN(n8223) );
  AOI21_X1 U9501 ( .B1(n8224), .B2(n10670), .A(n8223), .ZN(n8225) );
  OAI211_X1 U9502 ( .C1(n8227), .C2(n8277), .A(n8226), .B(n8225), .ZN(P2_U3159) );
  INV_X1 U9503 ( .A(n8228), .ZN(n8230) );
  NAND2_X1 U9504 ( .A1(n8230), .A2(n8229), .ZN(n8231) );
  XNOR2_X1 U9505 ( .A(n8232), .B(n8231), .ZN(n8238) );
  OAI22_X1 U9506 ( .A1(n10644), .A2(n8233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8974), .ZN(n8234) );
  AOI21_X1 U9507 ( .B1(n10657), .B2(n8744), .A(n8234), .ZN(n8235) );
  OAI21_X1 U9508 ( .B1(n8746), .B2(n10653), .A(n8235), .ZN(n8236) );
  AOI21_X1 U9509 ( .B1(n8749), .B2(n10667), .A(n8236), .ZN(n8237) );
  OAI21_X1 U9510 ( .B1(n8238), .B2(n8266), .A(n8237), .ZN(P2_U3163) );
  XOR2_X1 U9511 ( .A(n8240), .B(n8239), .Z(n8245) );
  OAI22_X1 U9512 ( .A1(n10641), .A2(n8699), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9092), .ZN(n8241) );
  AOI21_X1 U9513 ( .B1(n10655), .B2(n8524), .A(n8241), .ZN(n8242) );
  OAI21_X1 U9514 ( .B1(n8700), .B2(n10653), .A(n8242), .ZN(n8243) );
  AOI21_X1 U9515 ( .B1(n8824), .B2(n10667), .A(n8243), .ZN(n8244) );
  OAI21_X1 U9516 ( .B1(n8245), .B2(n8266), .A(n8244), .ZN(P2_U3165) );
  INV_X1 U9517 ( .A(n8247), .ZN(n8248) );
  AOI21_X1 U9518 ( .B1(n8249), .B2(n8246), .A(n8248), .ZN(n8254) );
  INV_X1 U9519 ( .A(n8712), .ZN(n8523) );
  AOI22_X1 U9520 ( .A1(n10657), .A2(n8523), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8251) );
  NAND2_X1 U9521 ( .A1(n10655), .A2(n8732), .ZN(n8250) );
  OAI211_X1 U9522 ( .C1(n10653), .C2(n8714), .A(n8251), .B(n8250), .ZN(n8252)
         );
  AOI21_X1 U9523 ( .B1(n8828), .B2(n10667), .A(n8252), .ZN(n8253) );
  OAI21_X1 U9524 ( .B1(n8254), .B2(n8266), .A(n8253), .ZN(P2_U3169) );
  INV_X1 U9525 ( .A(n8835), .ZN(n8264) );
  OAI211_X1 U9526 ( .C1(n8257), .C2(n8256), .A(n8255), .B(n10665), .ZN(n8263)
         );
  OAI22_X1 U9527 ( .A1(n10644), .A2(n8259), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8258), .ZN(n8261) );
  NOR2_X1 U9528 ( .A1(n10653), .A2(n8734), .ZN(n8260) );
  AOI211_X1 U9529 ( .C1(n10657), .C2(n8732), .A(n8261), .B(n8260), .ZN(n8262)
         );
  OAI211_X1 U9530 ( .C1(n8264), .C2(n8277), .A(n8263), .B(n8262), .ZN(P2_U3175) );
  INV_X1 U9531 ( .A(n8820), .ZN(n8278) );
  AOI21_X1 U9532 ( .B1(n8265), .B2(n8267), .A(n8266), .ZN(n8270) );
  NAND2_X1 U9534 ( .A1(n8270), .A2(n8269), .ZN(n8276) );
  INV_X1 U9535 ( .A(n8691), .ZN(n8274) );
  AOI22_X1 U9536 ( .A1(n8523), .A2(n10655), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8271) );
  OAI21_X1 U9537 ( .B1(n8272), .B2(n10641), .A(n8271), .ZN(n8273) );
  AOI21_X1 U9538 ( .B1(n8274), .B2(n10670), .A(n8273), .ZN(n8275) );
  OAI211_X1 U9539 ( .C1(n8278), .C2(n8277), .A(n8276), .B(n8275), .ZN(P2_U3180) );
  NAND2_X1 U9540 ( .A1(n8279), .A2(n8296), .ZN(n8282) );
  OR2_X1 U9541 ( .A1(n8297), .A2(n8280), .ZN(n8281) );
  NAND2_X1 U9542 ( .A1(n8282), .A2(n8281), .ZN(n8314) );
  OAI21_X1 U9543 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n8290) );
  MUX2_X1 U9544 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8286), .Z(n8288) );
  INV_X1 U9545 ( .A(SI_31_), .ZN(n8287) );
  XNOR2_X1 U9546 ( .A(n8288), .B(n8287), .ZN(n8289) );
  NAND2_X1 U9547 ( .A1(n10016), .A2(n8296), .ZN(n8293) );
  INV_X1 U9548 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8291) );
  OR2_X1 U9549 ( .A1(n8297), .A2(n8291), .ZN(n8292) );
  NAND2_X1 U9550 ( .A1(n8293), .A2(n8292), .ZN(n8641) );
  NAND2_X1 U9551 ( .A1(n8672), .A2(n8326), .ZN(n8295) );
  NAND2_X1 U9552 ( .A1(n9144), .A2(n8296), .ZN(n8299) );
  INV_X1 U9553 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9145) );
  OR2_X1 U9554 ( .A1(n8297), .A2(n9145), .ZN(n8298) );
  NAND2_X1 U9555 ( .A1(n8299), .A2(n8298), .ZN(n8812) );
  OR2_X1 U9556 ( .A1(n8812), .A2(n8317), .ZN(n8651) );
  NAND2_X1 U9557 ( .A1(n8652), .A2(n8651), .ZN(n8319) );
  NAND2_X1 U9558 ( .A1(n8300), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8305) );
  INV_X1 U9559 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8301) );
  OR2_X1 U9560 ( .A1(n6378), .A2(n8301), .ZN(n8304) );
  INV_X1 U9561 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8302) );
  OR2_X1 U9562 ( .A1(n6374), .A2(n8302), .ZN(n8303) );
  NAND4_X1 U9563 ( .A1(n8312), .A2(n8305), .A3(n8304), .A4(n8303), .ZN(n8644)
         );
  INV_X1 U9564 ( .A(n8644), .ZN(n8511) );
  OR2_X1 U9565 ( .A1(n8641), .A2(n8511), .ZN(n8316) );
  NAND2_X1 U9566 ( .A1(n8306), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8311) );
  INV_X1 U9567 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8307) );
  OR2_X1 U9568 ( .A1(n6677), .A2(n8307), .ZN(n8310) );
  INV_X1 U9569 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8308) );
  OR2_X1 U9570 ( .A1(n6374), .A2(n8308), .ZN(n8309) );
  NAND4_X1 U9571 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), .ZN(n8658)
         );
  INV_X1 U9572 ( .A(n8658), .ZN(n8313) );
  NAND2_X1 U9573 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U9574 ( .A1(n8316), .A2(n8315), .ZN(n8321) );
  NAND2_X1 U9575 ( .A1(n8812), .A2(n8317), .ZN(n8650) );
  INV_X1 U9576 ( .A(n8650), .ZN(n8318) );
  NOR2_X1 U9577 ( .A1(n8321), .A2(n8318), .ZN(n8506) );
  OAI211_X1 U9578 ( .C1(n8810), .C2(n8641), .A(n8319), .B(n8506), .ZN(n8324)
         );
  AND2_X1 U9579 ( .A1(n8810), .A2(n8658), .ZN(n8509) );
  AOI21_X1 U9580 ( .B1(n8509), .B2(n8641), .A(n8320), .ZN(n8323) );
  AOI22_X1 U9581 ( .A1(n8324), .A2(n8323), .B1(n8322), .B2(n8321), .ZN(n8513)
         );
  MUX2_X1 U9582 ( .A(n8657), .B(n8672), .S(n8477), .Z(n8472) );
  INV_X1 U9583 ( .A(n8472), .ZN(n8476) );
  MUX2_X1 U9584 ( .A(n8326), .B(n8325), .S(n8473), .Z(n8471) );
  INV_X1 U9585 ( .A(n8471), .ZN(n8475) );
  INV_X1 U9586 ( .A(n8437), .ZN(n8329) );
  INV_X1 U9587 ( .A(n8327), .ZN(n8328) );
  OAI21_X1 U9588 ( .B1(n8329), .B2(n8328), .A(n8477), .ZN(n8432) );
  NAND2_X1 U9589 ( .A1(n8331), .A2(n8414), .ZN(n8330) );
  NAND2_X1 U9590 ( .A1(n8330), .A2(n8477), .ZN(n8418) );
  INV_X1 U9591 ( .A(n8418), .ZN(n8424) );
  INV_X1 U9592 ( .A(n8417), .ZN(n8333) );
  INV_X1 U9593 ( .A(n8331), .ZN(n8332) );
  AOI21_X1 U9594 ( .B1(n8333), .B2(n8477), .A(n8332), .ZN(n8423) );
  NAND2_X1 U9595 ( .A1(n8335), .A2(n8334), .ZN(n8336) );
  NAND2_X1 U9596 ( .A1(n8343), .A2(n8336), .ZN(n8342) );
  NAND2_X1 U9597 ( .A1(n8539), .A2(n10470), .ZN(n8337) );
  OAI211_X1 U9598 ( .C1(n8342), .C2(n8338), .A(n8356), .B(n8337), .ZN(n8349)
         );
  NAND2_X1 U9599 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  NAND2_X1 U9600 ( .A1(n8342), .A2(n8341), .ZN(n8344) );
  NAND2_X1 U9601 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  NAND2_X1 U9602 ( .A1(n8345), .A2(n8482), .ZN(n8347) );
  NAND3_X1 U9603 ( .A1(n8347), .A2(n8351), .A3(n8346), .ZN(n8348) );
  MUX2_X1 U9604 ( .A(n8349), .B(n8348), .S(n8477), .Z(n8350) );
  NAND2_X1 U9605 ( .A1(n8350), .A2(n8484), .ZN(n8360) );
  INV_X1 U9606 ( .A(n8351), .ZN(n8353) );
  OAI211_X1 U9607 ( .C1(n8360), .C2(n8353), .A(n8361), .B(n8352), .ZN(n8355)
         );
  INV_X1 U9608 ( .A(n8354), .ZN(n8358) );
  NAND3_X1 U9609 ( .A1(n8355), .A2(n8362), .A3(n8358), .ZN(n8367) );
  INV_X1 U9610 ( .A(n8356), .ZN(n8359) );
  OAI211_X1 U9611 ( .C1(n8360), .C2(n8359), .A(n8358), .B(n8357), .ZN(n8365)
         );
  AND2_X1 U9612 ( .A1(n8370), .A2(n8361), .ZN(n8364) );
  INV_X1 U9613 ( .A(n8362), .ZN(n8363) );
  AOI21_X1 U9614 ( .B1(n8365), .B2(n8364), .A(n8363), .ZN(n8366) );
  MUX2_X1 U9615 ( .A(n8367), .B(n8366), .S(n8477), .Z(n8373) );
  INV_X1 U9616 ( .A(n8370), .ZN(n8371) );
  NAND2_X1 U9617 ( .A1(n8371), .A2(n8473), .ZN(n8372) );
  NAND4_X1 U9618 ( .A1(n8373), .A2(n8374), .A3(n5242), .A4(n8372), .ZN(n8386)
         );
  INV_X1 U9619 ( .A(n8374), .ZN(n8377) );
  INV_X1 U9620 ( .A(n8378), .ZN(n8384) );
  AND2_X1 U9621 ( .A1(n8380), .A2(n8379), .ZN(n8383) );
  OAI211_X1 U9622 ( .C1(n8384), .C2(n8383), .A(n8382), .B(n8381), .ZN(n8385)
         );
  INV_X1 U9623 ( .A(n8387), .ZN(n8388) );
  NAND2_X1 U9624 ( .A1(n8389), .A2(n8388), .ZN(n8390) );
  NAND2_X1 U9625 ( .A1(n8390), .A2(n8391), .ZN(n8395) );
  INV_X1 U9626 ( .A(n8391), .ZN(n8392) );
  NOR2_X1 U9627 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  MUX2_X1 U9628 ( .A(n8395), .B(n8394), .S(n8477), .Z(n8396) );
  INV_X1 U9629 ( .A(n8396), .ZN(n8397) );
  NAND3_X1 U9630 ( .A1(n8399), .A2(n8398), .A3(n8397), .ZN(n8404) );
  MUX2_X1 U9631 ( .A(n8401), .B(n8400), .S(n8473), .Z(n8402) );
  NAND3_X1 U9632 ( .A1(n8404), .A2(n8403), .A3(n8402), .ZN(n8410) );
  NAND2_X1 U9633 ( .A1(n8405), .A2(n8477), .ZN(n8408) );
  NAND2_X1 U9634 ( .A1(n8529), .A2(n8473), .ZN(n8407) );
  MUX2_X1 U9635 ( .A(n8408), .B(n8407), .S(n8406), .Z(n8409) );
  NAND2_X1 U9636 ( .A1(n8410), .A2(n8409), .ZN(n8411) );
  AND2_X1 U9637 ( .A1(n8411), .A2(n8478), .ZN(n8420) );
  INV_X1 U9638 ( .A(n8412), .ZN(n8416) );
  NAND2_X1 U9639 ( .A1(n8414), .A2(n8413), .ZN(n8415) );
  MUX2_X1 U9640 ( .A(n8416), .B(n8415), .S(n8473), .Z(n8419) );
  OAI211_X1 U9641 ( .C1(n8420), .C2(n8419), .A(n8418), .B(n8417), .ZN(n8422)
         );
  MUX2_X1 U9642 ( .A(n8426), .B(n8425), .S(n8477), .Z(n8427) );
  MUX2_X1 U9643 ( .A(n8429), .B(n8428), .S(n8473), .Z(n8430) );
  NAND2_X1 U9644 ( .A1(n8432), .A2(n8431), .ZN(n8436) );
  AOI21_X1 U9645 ( .B1(n8435), .B2(n8433), .A(n8477), .ZN(n8434) );
  INV_X1 U9646 ( .A(n8438), .ZN(n8440) );
  INV_X1 U9647 ( .A(n8441), .ZN(n8443) );
  INV_X1 U9648 ( .A(n8450), .ZN(n8444) );
  NOR2_X1 U9649 ( .A1(n8448), .A2(n8444), .ZN(n8721) );
  INV_X1 U9650 ( .A(n8721), .ZN(n8453) );
  INV_X1 U9651 ( .A(n8445), .ZN(n8447) );
  INV_X1 U9652 ( .A(n8709), .ZN(n8452) );
  INV_X1 U9653 ( .A(n8448), .ZN(n8449) );
  MUX2_X1 U9654 ( .A(n8450), .B(n8449), .S(n8477), .Z(n8451) );
  OAI211_X1 U9655 ( .C1(n8454), .C2(n8453), .A(n8452), .B(n8451), .ZN(n8458)
         );
  MUX2_X1 U9656 ( .A(n8456), .B(n8455), .S(n8477), .Z(n8457) );
  NAND3_X1 U9657 ( .A1(n8458), .A2(n8696), .A3(n8457), .ZN(n8462) );
  MUX2_X1 U9658 ( .A(n8460), .B(n8459), .S(n8473), .Z(n8461) );
  NAND2_X1 U9659 ( .A1(n8462), .A2(n8461), .ZN(n8465) );
  MUX2_X1 U9660 ( .A(n8820), .B(n8522), .S(n8477), .Z(n8464) );
  NAND2_X1 U9661 ( .A1(n8465), .A2(n8464), .ZN(n8466) );
  NAND2_X1 U9662 ( .A1(n8466), .A2(n8820), .ZN(n8463) );
  AOI22_X1 U9663 ( .A1(n8463), .A2(n8505), .B1(n8473), .B2(n8474), .ZN(n8470)
         );
  OAI22_X1 U9664 ( .A1(n8465), .A2(n8464), .B1(n8699), .B2(n8477), .ZN(n8468)
         );
  AND3_X1 U9665 ( .A1(n8468), .A2(n8467), .A3(n8466), .ZN(n8469) );
  INV_X1 U9666 ( .A(n8479), .ZN(n8481) );
  NOR4_X1 U9667 ( .A1(n8481), .A2(n8480), .A3(n7128), .A4(n6684), .ZN(n8485)
         );
  NAND4_X1 U9668 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n8489)
         );
  NOR4_X1 U9669 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n8493)
         );
  NAND4_X1 U9670 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n8490), .ZN(n8494)
         );
  NOR4_X1 U9671 ( .A1(n5040), .A2(n8496), .A3(n8495), .A4(n8494), .ZN(n8498)
         );
  NAND4_X1 U9672 ( .A1(n8792), .A2(n8499), .A3(n8498), .A4(n8497), .ZN(n8500)
         );
  NOR4_X1 U9673 ( .A1(n8758), .A2(n5064), .A3(n8782), .A4(n8500), .ZN(n8501)
         );
  NAND4_X1 U9674 ( .A1(n8721), .A2(n8737), .A3(n8750), .A4(n8501), .ZN(n8502)
         );
  NOR4_X1 U9675 ( .A1(n8686), .A2(n8709), .A3(n8703), .A4(n8502), .ZN(n8504)
         );
  AND4_X1 U9676 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(n8508)
         );
  INV_X1 U9677 ( .A(n8509), .ZN(n8510) );
  AOI22_X1 U9678 ( .A1(n8513), .A2(n8512), .B1(n8511), .B2(n8641), .ZN(n8514)
         );
  XNOR2_X1 U9679 ( .A(n8514), .B(n8633), .ZN(n8521) );
  NAND3_X1 U9680 ( .A1(n8516), .A2(n8515), .A3(n8619), .ZN(n8517) );
  OAI211_X1 U9681 ( .C1(n8518), .C2(n8520), .A(n8517), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8519) );
  OAI21_X1 U9682 ( .B1(n8521), .B2(n8520), .A(n8519), .ZN(P2_U3296) );
  MUX2_X1 U9683 ( .A(n8644), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8580), .Z(
        P2_U3522) );
  MUX2_X1 U9684 ( .A(n8658), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8580), .Z(
        P2_U3521) );
  MUX2_X1 U9685 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8657), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9686 ( .A(n8688), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8580), .Z(
        P2_U3518) );
  MUX2_X1 U9687 ( .A(n8522), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8580), .Z(
        P2_U3517) );
  MUX2_X1 U9688 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8523), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9689 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8524), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9690 ( .A(n8732), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8580), .Z(
        P2_U3514) );
  MUX2_X1 U9691 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8744), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9692 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n6594), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9693 ( .A(n8770), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8580), .Z(
        P2_U3511) );
  MUX2_X1 U9694 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n10656), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9695 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8798), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9696 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8525), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9697 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8526), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9698 ( .A(n8527), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8580), .Z(
        P2_U3506) );
  MUX2_X1 U9699 ( .A(n8528), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8580), .Z(
        P2_U3505) );
  MUX2_X1 U9700 ( .A(n8529), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8580), .Z(
        P2_U3504) );
  MUX2_X1 U9701 ( .A(n8530), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8580), .Z(
        P2_U3503) );
  MUX2_X1 U9702 ( .A(n8531), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8580), .Z(
        P2_U3502) );
  MUX2_X1 U9703 ( .A(n8532), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8580), .Z(
        P2_U3501) );
  MUX2_X1 U9704 ( .A(n5136), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8580), .Z(
        P2_U3500) );
  MUX2_X1 U9705 ( .A(n8533), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8580), .Z(
        P2_U3499) );
  MUX2_X1 U9706 ( .A(n8534), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8580), .Z(
        P2_U3498) );
  MUX2_X1 U9707 ( .A(n8535), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8580), .Z(
        P2_U3497) );
  MUX2_X1 U9708 ( .A(n8536), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8580), .Z(
        P2_U3496) );
  MUX2_X1 U9709 ( .A(n8537), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8580), .Z(
        P2_U3495) );
  MUX2_X1 U9710 ( .A(n8538), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8580), .Z(
        P2_U3494) );
  MUX2_X1 U9711 ( .A(n8539), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8580), .Z(
        P2_U3493) );
  MUX2_X1 U9712 ( .A(n6991), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8580), .Z(
        P2_U3492) );
  XNOR2_X1 U9713 ( .A(n8617), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8612) );
  AOI22_X1 U9714 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8598), .B1(n10387), .B2(
        n8863), .ZN(n10390) );
  AOI22_X1 U9715 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8594), .B1(n10356), .B2(
        n8550), .ZN(n10359) );
  AOI22_X1 U9716 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8590), .B1(n10324), .B2(
        n6512), .ZN(n10327) );
  NAND2_X1 U9717 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8586), .ZN(n8545) );
  AOI22_X1 U9718 ( .A1(n10290), .A2(n8540), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n8586), .ZN(n10298) );
  OR2_X1 U9719 ( .A1(n8542), .A2(n8541), .ZN(n8544) );
  NAND2_X1 U9720 ( .A1(n8544), .A2(n8543), .ZN(n10297) );
  NAND2_X1 U9721 ( .A1(n10298), .A2(n10297), .ZN(n10296) );
  NAND2_X1 U9722 ( .A1(n8545), .A2(n10296), .ZN(n8546) );
  NAND2_X1 U9723 ( .A1(n8562), .A2(n8546), .ZN(n8547) );
  XNOR2_X1 U9724 ( .A(n10309), .B(n8546), .ZN(n10314) );
  NAND2_X1 U9725 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10314), .ZN(n10313) );
  NAND2_X1 U9726 ( .A1(n8547), .A2(n10313), .ZN(n10326) );
  NAND2_X1 U9727 ( .A1(n10327), .A2(n10326), .ZN(n10325) );
  OAI21_X1 U9728 ( .B1(n10324), .B2(n6512), .A(n10325), .ZN(n8548) );
  NAND2_X1 U9729 ( .A1(n8559), .A2(n8548), .ZN(n8549) );
  XNOR2_X1 U9730 ( .A(n10341), .B(n8548), .ZN(n10343) );
  NAND2_X1 U9731 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n10343), .ZN(n10342) );
  NAND2_X1 U9732 ( .A1(n8549), .A2(n10342), .ZN(n10358) );
  NAND2_X1 U9733 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  OAI21_X1 U9734 ( .B1(n10356), .B2(n8550), .A(n10357), .ZN(n8551) );
  NAND2_X1 U9735 ( .A1(n8556), .A2(n8551), .ZN(n8552) );
  XNOR2_X1 U9736 ( .A(n10372), .B(n8551), .ZN(n10374) );
  NAND2_X1 U9737 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10374), .ZN(n10373) );
  NAND2_X1 U9738 ( .A1(n8552), .A2(n10373), .ZN(n10389) );
  NAND2_X1 U9739 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  OAI21_X1 U9740 ( .B1(n10387), .B2(n8863), .A(n10388), .ZN(n8553) );
  NAND2_X1 U9741 ( .A1(n8601), .A2(n8553), .ZN(n8554) );
  XNOR2_X1 U9742 ( .A(n10405), .B(n8553), .ZN(n10407) );
  NAND2_X1 U9743 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10407), .ZN(n10406) );
  NAND2_X1 U9744 ( .A1(n8554), .A2(n10406), .ZN(n8613) );
  XOR2_X1 U9745 ( .A(n8612), .B(n8613), .Z(n8611) );
  MUX2_X1 U9746 ( .A(n10416), .B(n8859), .S(n8619), .Z(n8576) );
  XNOR2_X1 U9747 ( .A(n8601), .B(n8576), .ZN(n10410) );
  MUX2_X1 U9748 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8619), .Z(n8555) );
  OR2_X1 U9749 ( .A1(n8555), .A2(n8598), .ZN(n8574) );
  XNOR2_X1 U9750 ( .A(n10387), .B(n8555), .ZN(n10393) );
  MUX2_X1 U9751 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8619), .Z(n8557) );
  OR2_X1 U9752 ( .A1(n8557), .A2(n8556), .ZN(n8573) );
  XNOR2_X1 U9753 ( .A(n10372), .B(n8557), .ZN(n10377) );
  MUX2_X1 U9754 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8619), .Z(n8558) );
  OR2_X1 U9755 ( .A1(n8558), .A2(n8594), .ZN(n8572) );
  XNOR2_X1 U9756 ( .A(n8558), .B(n10356), .ZN(n10362) );
  MUX2_X1 U9757 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8619), .Z(n8560) );
  OR2_X1 U9758 ( .A1(n8560), .A2(n8559), .ZN(n8571) );
  XNOR2_X1 U9759 ( .A(n8560), .B(n10341), .ZN(n10346) );
  MUX2_X1 U9760 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8619), .Z(n8561) );
  OR2_X1 U9761 ( .A1(n8561), .A2(n8590), .ZN(n8570) );
  XNOR2_X1 U9762 ( .A(n8561), .B(n10324), .ZN(n10330) );
  MUX2_X1 U9763 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8619), .Z(n8568) );
  OR2_X1 U9764 ( .A1(n8568), .A2(n8562), .ZN(n8569) );
  NOR2_X1 U9765 ( .A1(n8564), .A2(n8563), .ZN(n10295) );
  MUX2_X1 U9766 ( .A(n8565), .B(n8540), .S(n8619), .Z(n8566) );
  NAND2_X1 U9767 ( .A1(n8566), .A2(n10290), .ZN(n10292) );
  MUX2_X1 U9768 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8619), .Z(n8567) );
  AND2_X1 U9769 ( .A1(n8567), .A2(n8586), .ZN(n10291) );
  AOI21_X1 U9770 ( .B1(n10295), .B2(n10292), .A(n10291), .ZN(n10312) );
  XNOR2_X1 U9771 ( .A(n8568), .B(n10309), .ZN(n10311) );
  NAND2_X1 U9772 ( .A1(n10312), .A2(n10311), .ZN(n10310) );
  NAND2_X1 U9773 ( .A1(n8569), .A2(n10310), .ZN(n10329) );
  NAND2_X1 U9774 ( .A1(n10330), .A2(n10329), .ZN(n10328) );
  NAND2_X1 U9775 ( .A1(n8570), .A2(n10328), .ZN(n10345) );
  NAND2_X1 U9776 ( .A1(n10346), .A2(n10345), .ZN(n10344) );
  NAND2_X1 U9777 ( .A1(n8571), .A2(n10344), .ZN(n10361) );
  NAND2_X1 U9778 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  NAND2_X1 U9779 ( .A1(n8572), .A2(n10360), .ZN(n10376) );
  NAND2_X1 U9780 ( .A1(n10377), .A2(n10376), .ZN(n10375) );
  NAND2_X1 U9781 ( .A1(n8573), .A2(n10375), .ZN(n10392) );
  NAND2_X1 U9782 ( .A1(n10393), .A2(n10392), .ZN(n10391) );
  NAND2_X1 U9783 ( .A1(n8574), .A2(n10391), .ZN(n10409) );
  NAND2_X1 U9784 ( .A1(n10410), .A2(n10409), .ZN(n10408) );
  INV_X1 U9785 ( .A(n10408), .ZN(n8575) );
  AOI21_X1 U9786 ( .B1(n10405), .B2(n8576), .A(n8575), .ZN(n8578) );
  MUX2_X1 U9787 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8619), .Z(n8577) );
  NOR2_X1 U9788 ( .A1(n8578), .A2(n8577), .ZN(n8615) );
  INV_X1 U9789 ( .A(n8615), .ZN(n8579) );
  NAND2_X1 U9790 ( .A1(n8578), .A2(n8577), .ZN(n8616) );
  NAND2_X1 U9791 ( .A1(n8579), .A2(n8616), .ZN(n8581) );
  OAI21_X1 U9792 ( .B1(n8581), .B2(n8580), .A(n10271), .ZN(n8610) );
  INV_X1 U9793 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8609) );
  NAND3_X1 U9794 ( .A1(n8581), .A2(n10412), .A3(n8625), .ZN(n8608) );
  NAND2_X1 U9795 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8586), .ZN(n8585) );
  OAI21_X1 U9796 ( .B1(n8586), .B2(P2_REG2_REG_10__SCAN_IN), .A(n8585), .ZN(
        n10302) );
  NOR2_X1 U9797 ( .A1(n10309), .A2(n8587), .ZN(n8588) );
  NOR2_X1 U9798 ( .A1(n6502), .A2(n10318), .ZN(n10317) );
  MUX2_X1 U9799 ( .A(n6515), .B(P2_REG2_REG_12__SCAN_IN), .S(n10324), .Z(n8589) );
  INV_X1 U9800 ( .A(n8589), .ZN(n10334) );
  NOR2_X1 U9801 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  NOR2_X1 U9802 ( .A1(n10341), .A2(n8591), .ZN(n8592) );
  MUX2_X1 U9803 ( .A(n6344), .B(P2_REG2_REG_14__SCAN_IN), .S(n10356), .Z(n8593) );
  INV_X1 U9804 ( .A(n8593), .ZN(n10366) );
  NOR2_X1 U9805 ( .A1(n10372), .A2(n8595), .ZN(n8596) );
  MUX2_X1 U9806 ( .A(n8073), .B(P2_REG2_REG_16__SCAN_IN), .S(n10387), .Z(n8597) );
  INV_X1 U9807 ( .A(n8597), .ZN(n10397) );
  INV_X1 U9808 ( .A(n8624), .ZN(n8627) );
  INV_X1 U9809 ( .A(n8599), .ZN(n8600) );
  OAI21_X1 U9810 ( .B1(n8601), .B2(n8600), .A(n8624), .ZN(n10417) );
  NOR2_X1 U9811 ( .A1(n8627), .A2(n10415), .ZN(n8603) );
  NOR2_X1 U9812 ( .A1(n8617), .A2(n8787), .ZN(n8602) );
  AOI21_X1 U9813 ( .B1(n8787), .B2(n8617), .A(n8602), .ZN(n8623) );
  XOR2_X1 U9814 ( .A(n8603), .B(n8623), .Z(n8606) );
  NOR2_X1 U9815 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8604), .ZN(n8605) );
  AOI22_X1 U9816 ( .A1(n8613), .A2(n8612), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8625), .ZN(n8614) );
  XNOR2_X1 U9817 ( .A(n8633), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8618) );
  XNOR2_X1 U9818 ( .A(n8614), .B(n8618), .ZN(n8640) );
  AOI21_X1 U9819 ( .B1(n8617), .B2(n8616), .A(n8615), .ZN(n8622) );
  INV_X1 U9820 ( .A(n8618), .ZN(n8620) );
  MUX2_X1 U9821 ( .A(n5489), .B(n8620), .S(n8619), .Z(n8621) );
  XNOR2_X1 U9822 ( .A(n8622), .B(n8621), .ZN(n8638) );
  NAND2_X1 U9823 ( .A1(n10415), .A2(n8623), .ZN(n8630) );
  NAND2_X1 U9824 ( .A1(n8624), .A2(n8787), .ZN(n8626) );
  NAND2_X1 U9825 ( .A1(n8626), .A2(n8625), .ZN(n8629) );
  NAND2_X1 U9826 ( .A1(n8627), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U9827 ( .A1(n8630), .A2(n5478), .ZN(n8631) );
  XNOR2_X1 U9828 ( .A(n8631), .B(n5489), .ZN(n8636) );
  AOI21_X1 U9829 ( .B1(n10404), .B2(n8633), .A(n8632), .ZN(n8635) );
  NAND2_X1 U9830 ( .A1(n10403), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8634) );
  OAI211_X1 U9831 ( .C1(n8636), .C2(n10418), .A(n8635), .B(n8634), .ZN(n8637)
         );
  INV_X1 U9832 ( .A(n8641), .ZN(n8808) );
  AOI21_X1 U9833 ( .B1(n10572), .B2(n8642), .A(n10577), .ZN(n8645) );
  AOI21_X1 U9834 ( .B1(P2_B_REG_SCAN_IN), .B2(n8643), .A(n8786), .ZN(n8659) );
  NAND2_X1 U9835 ( .A1(n8644), .A2(n8659), .ZN(n8809) );
  NAND2_X1 U9836 ( .A1(n8645), .A2(n8809), .ZN(n8647) );
  OAI21_X1 U9837 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n10575), .A(n8647), .ZN(
        n8646) );
  OAI21_X1 U9838 ( .B1(n8808), .B2(n8649), .A(n8646), .ZN(P2_U3202) );
  OAI21_X1 U9839 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(n10575), .A(n8647), .ZN(
        n8648) );
  OAI21_X1 U9840 ( .B1(n8810), .B2(n8649), .A(n8648), .ZN(P2_U3203) );
  NAND2_X1 U9841 ( .A1(n8651), .A2(n8650), .ZN(n8655) );
  INV_X1 U9842 ( .A(n8655), .ZN(n8656) );
  AOI22_X1 U9843 ( .A1(n8659), .A2(n8658), .B1(n8657), .B2(n8771), .ZN(n8660)
         );
  NAND2_X1 U9844 ( .A1(n8811), .A2(n10575), .ZN(n8666) );
  OAI22_X1 U9845 ( .A1(n10575), .A2(n8663), .B1(n8662), .B2(n10468), .ZN(n8664) );
  AOI21_X1 U9846 ( .B1(n8812), .B2(n10568), .A(n8664), .ZN(n8665) );
  OAI211_X1 U9847 ( .C1(n8815), .C2(n10567), .A(n8666), .B(n8665), .ZN(
        P2_U3204) );
  OAI22_X1 U9848 ( .A1(n10575), .A2(n8668), .B1(n8667), .B2(n10468), .ZN(n8671) );
  NOR2_X1 U9849 ( .A1(n8669), .A2(n8807), .ZN(n8670) );
  AOI211_X1 U9850 ( .C1(n10568), .C2(n8672), .A(n8671), .B(n8670), .ZN(n8673)
         );
  OAI21_X1 U9851 ( .B1(n8674), .B2(n10577), .A(n8673), .ZN(P2_U3205) );
  OAI22_X1 U9852 ( .A1(n10575), .A2(n8676), .B1(n8675), .B2(n10468), .ZN(n8679) );
  NOR2_X1 U9853 ( .A1(n8677), .A2(n8807), .ZN(n8678) );
  AOI211_X1 U9854 ( .C1(n10568), .C2(n8680), .A(n8679), .B(n8678), .ZN(n8681)
         );
  OAI21_X1 U9855 ( .B1(n8682), .B2(n10577), .A(n8681), .ZN(P2_U3206) );
  NAND2_X1 U9856 ( .A1(n8683), .A2(n8686), .ZN(n8684) );
  NAND2_X1 U9857 ( .A1(n4954), .A2(n8684), .ZN(n8884) );
  OAI211_X1 U9858 ( .C1(n8687), .C2(n8686), .A(n8685), .B(n8793), .ZN(n8690)
         );
  NAND2_X1 U9859 ( .A1(n8688), .A2(n8797), .ZN(n8689) );
  OAI211_X1 U9860 ( .C1(n8712), .C2(n8801), .A(n8690), .B(n8689), .ZN(n8819)
         );
  NAND2_X1 U9861 ( .A1(n8819), .A2(n10575), .ZN(n8695) );
  OAI22_X1 U9862 ( .A1(n10575), .A2(n8692), .B1(n8691), .B2(n10468), .ZN(n8693) );
  AOI21_X1 U9863 ( .B1(n8820), .B2(n10568), .A(n8693), .ZN(n8694) );
  OAI211_X1 U9864 ( .C1(n8884), .C2(n8807), .A(n8695), .B(n8694), .ZN(P2_U3207) );
  XNOR2_X1 U9865 ( .A(n8697), .B(n8696), .ZN(n8698) );
  OAI222_X1 U9866 ( .A1(n8786), .A2(n8699), .B1(n8801), .B2(n8725), .C1(n8723), 
        .C2(n8698), .ZN(n8823) );
  OAI22_X1 U9867 ( .A1(n8701), .A2(n10469), .B1(n8700), .B2(n10468), .ZN(n8702) );
  OAI21_X1 U9868 ( .B1(n8823), .B2(n8702), .A(n10575), .ZN(n8706) );
  XNOR2_X1 U9869 ( .A(n8704), .B(n8703), .ZN(n8888) );
  OR2_X1 U9870 ( .A1(n8888), .A2(n8807), .ZN(n8705) );
  OAI211_X1 U9871 ( .C1(n10575), .C2(n8707), .A(n8706), .B(n8705), .ZN(
        P2_U3208) );
  XNOR2_X1 U9872 ( .A(n8708), .B(n8709), .ZN(n8892) );
  XNOR2_X1 U9873 ( .A(n8710), .B(n8709), .ZN(n8711) );
  OAI222_X1 U9874 ( .A1(n8801), .A2(n8713), .B1(n8786), .B2(n8712), .C1(n8723), 
        .C2(n8711), .ZN(n8827) );
  OAI22_X1 U9875 ( .A1(n8715), .A2(n10469), .B1(n8714), .B2(n10468), .ZN(n8716) );
  OAI21_X1 U9876 ( .B1(n8827), .B2(n8716), .A(n10575), .ZN(n8718) );
  NAND2_X1 U9877 ( .A1(n10577), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8717) );
  OAI211_X1 U9878 ( .C1(n8892), .C2(n8807), .A(n8718), .B(n8717), .ZN(P2_U3209) );
  XNOR2_X1 U9879 ( .A(n8719), .B(n8721), .ZN(n8896) );
  XNOR2_X1 U9880 ( .A(n8720), .B(n8721), .ZN(n8722) );
  OAI222_X1 U9881 ( .A1(n8786), .A2(n8725), .B1(n8801), .B2(n8724), .C1(n8723), 
        .C2(n8722), .ZN(n8831) );
  NAND2_X1 U9882 ( .A1(n8831), .A2(n10575), .ZN(n8730) );
  OAI22_X1 U9883 ( .A1(n10575), .A2(n8727), .B1(n8726), .B2(n10468), .ZN(n8728) );
  AOI21_X1 U9884 ( .B1(n8832), .B2(n10568), .A(n8728), .ZN(n8729) );
  OAI211_X1 U9885 ( .C1(n8896), .C2(n8807), .A(n8730), .B(n8729), .ZN(P2_U3210) );
  XNOR2_X1 U9886 ( .A(n8731), .B(n8737), .ZN(n8733) );
  AOI222_X1 U9887 ( .A1(n8793), .A2(n8733), .B1(n6594), .B2(n8771), .C1(n8732), 
        .C2(n8797), .ZN(n8837) );
  OAI22_X1 U9888 ( .A1(n10575), .A2(n8735), .B1(n8734), .B2(n10468), .ZN(n8740) );
  OAI21_X1 U9889 ( .B1(n8738), .B2(n8737), .A(n8736), .ZN(n8838) );
  NOR2_X1 U9890 ( .A1(n8838), .A2(n8807), .ZN(n8739) );
  AOI211_X1 U9891 ( .C1(n10568), .C2(n8835), .A(n8740), .B(n8739), .ZN(n8741)
         );
  OAI21_X1 U9892 ( .B1(n8837), .B2(n10577), .A(n8741), .ZN(P2_U3211) );
  XNOR2_X1 U9893 ( .A(n8743), .B(n8742), .ZN(n8745) );
  AOI222_X1 U9894 ( .A1(n8793), .A2(n8745), .B1(n8770), .B2(n8771), .C1(n8744), 
        .C2(n8797), .ZN(n8843) );
  OAI22_X1 U9895 ( .A1(n10575), .A2(n8747), .B1(n8746), .B2(n10468), .ZN(n8748) );
  AOI21_X1 U9896 ( .B1(n8749), .B2(n10568), .A(n8748), .ZN(n8754) );
  OR2_X1 U9897 ( .A1(n8751), .A2(n8750), .ZN(n8841) );
  NAND3_X1 U9898 ( .A1(n8841), .A2(n8752), .A3(n8840), .ZN(n8753) );
  OAI211_X1 U9899 ( .C1(n8843), .C2(n10577), .A(n8754), .B(n8753), .ZN(
        P2_U3212) );
  OAI21_X1 U9900 ( .B1(n4941), .B2(n8758), .A(n8755), .ZN(n8756) );
  AOI222_X1 U9901 ( .A1(n8793), .A2(n8756), .B1(n6594), .B2(n8797), .C1(n10656), .C2(n8771), .ZN(n8846) );
  OAI22_X1 U9902 ( .A1(n10575), .A2(n8757), .B1(n10658), .B2(n10468), .ZN(
        n8763) );
  NAND2_X1 U9903 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  NAND2_X1 U9904 ( .A1(n8761), .A2(n8760), .ZN(n9118) );
  NOR2_X1 U9905 ( .A1(n9118), .A2(n8807), .ZN(n8762) );
  AOI211_X1 U9906 ( .C1(n10568), .C2(n10668), .A(n8763), .B(n8762), .ZN(n8764)
         );
  OAI21_X1 U9907 ( .B1(n8846), .B2(n10577), .A(n8764), .ZN(P2_U3213) );
  XNOR2_X1 U9908 ( .A(n8765), .B(n8768), .ZN(n9122) );
  NAND3_X1 U9909 ( .A1(n8766), .A2(n8768), .A3(n8767), .ZN(n8769) );
  NAND2_X1 U9910 ( .A1(n8769), .A2(n8793), .ZN(n8773) );
  AOI22_X1 U9911 ( .A1(n8798), .A2(n8771), .B1(n8797), .B2(n8770), .ZN(n8772)
         );
  OAI21_X1 U9912 ( .B1(n8774), .B2(n8773), .A(n8772), .ZN(n8850) );
  NAND2_X1 U9913 ( .A1(n8850), .A2(n10575), .ZN(n8779) );
  OAI22_X1 U9914 ( .A1(n10575), .A2(n8776), .B1(n8775), .B2(n10468), .ZN(n8777) );
  AOI21_X1 U9915 ( .B1(n8851), .B2(n10568), .A(n8777), .ZN(n8778) );
  OAI211_X1 U9916 ( .C1(n9122), .C2(n8807), .A(n8779), .B(n8778), .ZN(P2_U3214) );
  XNOR2_X1 U9917 ( .A(n8780), .B(n8781), .ZN(n9126) );
  OAI211_X1 U9918 ( .C1(n8783), .C2(n8782), .A(n8766), .B(n8793), .ZN(n8785)
         );
  OR2_X1 U9919 ( .A1(n10643), .A2(n8801), .ZN(n8784) );
  OAI211_X1 U9920 ( .C1(n10642), .C2(n8786), .A(n8785), .B(n8784), .ZN(n8854)
         );
  NAND2_X1 U9921 ( .A1(n8854), .A2(n10575), .ZN(n8790) );
  OAI22_X1 U9922 ( .A1(n10575), .A2(n8787), .B1(n10654), .B2(n10468), .ZN(
        n8788) );
  AOI21_X1 U9923 ( .B1(n10649), .B2(n10568), .A(n8788), .ZN(n8789) );
  OAI211_X1 U9924 ( .C1(n9126), .C2(n8807), .A(n8790), .B(n8789), .ZN(P2_U3215) );
  XNOR2_X1 U9925 ( .A(n8791), .B(n8792), .ZN(n9130) );
  OAI211_X1 U9926 ( .C1(n8796), .C2(n8795), .A(n8794), .B(n8793), .ZN(n8800)
         );
  NAND2_X1 U9927 ( .A1(n8798), .A2(n8797), .ZN(n8799) );
  OAI211_X1 U9928 ( .C1(n8802), .C2(n8801), .A(n8800), .B(n8799), .ZN(n8857)
         );
  NAND2_X1 U9929 ( .A1(n8857), .A2(n10575), .ZN(n8806) );
  OAI22_X1 U9930 ( .A1(n10575), .A2(n10416), .B1(n8803), .B2(n10468), .ZN(
        n8804) );
  AOI21_X1 U9931 ( .B1(n8858), .B2(n10568), .A(n8804), .ZN(n8805) );
  OAI211_X1 U9932 ( .C1(n9130), .C2(n8807), .A(n8806), .B(n8805), .ZN(P2_U3216) );
  OAI21_X1 U9933 ( .B1(n8808), .B2(n8844), .A(n8809), .ZN(n8878) );
  MUX2_X1 U9934 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8878), .S(n8876), .Z(
        P2_U3490) );
  OAI21_X1 U9935 ( .B1(n8810), .B2(n8844), .A(n8809), .ZN(n8879) );
  MUX2_X1 U9936 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8879), .S(n8876), .Z(
        P2_U3489) );
  INV_X1 U9937 ( .A(n8811), .ZN(n8818) );
  INV_X1 U9938 ( .A(n8812), .ZN(n8813) );
  OAI22_X1 U9939 ( .A1(n8815), .A2(n8814), .B1(n8813), .B2(n8844), .ZN(n8816)
         );
  INV_X1 U9940 ( .A(n8816), .ZN(n8817) );
  NAND2_X1 U9941 ( .A1(n8818), .A2(n8817), .ZN(n8880) );
  MUX2_X1 U9942 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8880), .S(n8876), .Z(
        P2_U3488) );
  INV_X1 U9943 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8821) );
  AOI21_X1 U9944 ( .B1(n8871), .B2(n8820), .A(n8819), .ZN(n8881) );
  MUX2_X1 U9945 ( .A(n8821), .B(n8881), .S(n8876), .Z(n8822) );
  OAI21_X1 U9946 ( .B1(n8865), .B2(n8884), .A(n8822), .ZN(P2_U3485) );
  AOI21_X1 U9947 ( .B1(n8871), .B2(n8824), .A(n8823), .ZN(n8885) );
  MUX2_X1 U9948 ( .A(n8825), .B(n8885), .S(n8876), .Z(n8826) );
  OAI21_X1 U9949 ( .B1(n8865), .B2(n8888), .A(n8826), .ZN(P2_U3484) );
  INV_X1 U9950 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8829) );
  AOI21_X1 U9951 ( .B1(n8871), .B2(n8828), .A(n8827), .ZN(n8889) );
  MUX2_X1 U9952 ( .A(n8829), .B(n8889), .S(n8876), .Z(n8830) );
  OAI21_X1 U9953 ( .B1(n8892), .B2(n8865), .A(n8830), .ZN(P2_U3483) );
  AOI21_X1 U9954 ( .B1(n8871), .B2(n8832), .A(n8831), .ZN(n8893) );
  MUX2_X1 U9955 ( .A(n8833), .B(n8893), .S(n8876), .Z(n8834) );
  OAI21_X1 U9956 ( .B1(n8896), .B2(n8865), .A(n8834), .ZN(P2_U3482) );
  NAND2_X1 U9957 ( .A1(n8835), .A2(n8871), .ZN(n8836) );
  OAI211_X1 U9958 ( .C1(n8839), .C2(n8838), .A(n8837), .B(n8836), .ZN(n9111)
         );
  MUX2_X1 U9959 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9111), .S(n8876), .Z(
        P2_U3481) );
  NAND3_X1 U9960 ( .A1(n8841), .A2(n8840), .A3(n8872), .ZN(n8842) );
  OAI211_X1 U9961 ( .C1(n8845), .C2(n8844), .A(n8843), .B(n8842), .ZN(n9114)
         );
  MUX2_X1 U9962 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9114), .S(n8876), .Z(
        P2_U3480) );
  INV_X1 U9963 ( .A(n8846), .ZN(n8847) );
  AOI21_X1 U9964 ( .B1(n8871), .B2(n10668), .A(n8847), .ZN(n9115) );
  MUX2_X1 U9965 ( .A(n8848), .B(n9115), .S(n8876), .Z(n8849) );
  OAI21_X1 U9966 ( .B1(n8865), .B2(n9118), .A(n8849), .ZN(P2_U3479) );
  AOI21_X1 U9967 ( .B1(n8871), .B2(n8851), .A(n8850), .ZN(n9119) );
  MUX2_X1 U9968 ( .A(n8852), .B(n9119), .S(n8876), .Z(n8853) );
  OAI21_X1 U9969 ( .B1(n9122), .B2(n8865), .A(n8853), .ZN(P2_U3478) );
  AOI21_X1 U9970 ( .B1(n8871), .B2(n10649), .A(n8854), .ZN(n9123) );
  MUX2_X1 U9971 ( .A(n8855), .B(n9123), .S(n8876), .Z(n8856) );
  OAI21_X1 U9972 ( .B1(n9126), .B2(n8865), .A(n8856), .ZN(P2_U3477) );
  AOI21_X1 U9973 ( .B1(n8871), .B2(n8858), .A(n8857), .ZN(n9127) );
  MUX2_X1 U9974 ( .A(n8859), .B(n9127), .S(n8876), .Z(n8860) );
  OAI21_X1 U9975 ( .B1(n9130), .B2(n8865), .A(n8860), .ZN(P2_U3476) );
  AOI21_X1 U9976 ( .B1(n8871), .B2(n8862), .A(n8861), .ZN(n9131) );
  MUX2_X1 U9977 ( .A(n8863), .B(n9131), .S(n8876), .Z(n8864) );
  OAI21_X1 U9978 ( .B1(n9135), .B2(n8865), .A(n8864), .ZN(P2_U3475) );
  AOI22_X1 U9979 ( .A1(n8867), .A2(n8872), .B1(n8871), .B2(n8866), .ZN(n8868)
         );
  NAND2_X1 U9980 ( .A1(n8869), .A2(n8868), .ZN(n9136) );
  MUX2_X1 U9981 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9136), .S(n8876), .Z(
        P2_U3474) );
  AOI22_X1 U9982 ( .A1(n8873), .A2(n8872), .B1(n8871), .B2(n8870), .ZN(n8874)
         );
  NAND2_X1 U9983 ( .A1(n8875), .A2(n8874), .ZN(n9137) );
  MUX2_X1 U9984 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9137), .S(n8876), .Z(
        P2_U3471) );
  MUX2_X1 U9985 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8877), .S(n8876), .Z(
        P2_U3459) );
  MUX2_X1 U9986 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8878), .S(n10640), .Z(
        P2_U3458) );
  MUX2_X1 U9987 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8879), .S(n10640), .Z(
        P2_U3457) );
  MUX2_X1 U9988 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8880), .S(n10640), .Z(
        P2_U3456) );
  MUX2_X1 U9989 ( .A(n8882), .B(n8881), .S(n10640), .Z(n8883) );
  OAI21_X1 U9990 ( .B1(n8884), .B2(n9134), .A(n8883), .ZN(P2_U3453) );
  INV_X1 U9991 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8886) );
  MUX2_X1 U9992 ( .A(n8886), .B(n8885), .S(n10640), .Z(n8887) );
  OAI21_X1 U9993 ( .B1(n8888), .B2(n9134), .A(n8887), .ZN(P2_U3452) );
  MUX2_X1 U9994 ( .A(n8890), .B(n8889), .S(n10640), .Z(n8891) );
  OAI21_X1 U9995 ( .B1(n8892), .B2(n9134), .A(n8891), .ZN(P2_U3451) );
  INV_X1 U9996 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8894) );
  MUX2_X1 U9997 ( .A(n8894), .B(n8893), .S(n10640), .Z(n8895) );
  OAI21_X1 U9998 ( .B1(n8896), .B2(n9134), .A(n8895), .ZN(P2_U3450) );
  OAI22_X1 U9999 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_124), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .ZN(n8897) );
  AOI221_X1 U10000 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        keyinput_125), .C2(P2_REG3_REG_6__SCAN_IN), .A(n8897), .ZN(n8991) );
  AOI22_X1 U10001 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_118), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .ZN(n8898) );
  OAI221_X1 U10002 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_119), .A(n8898), .ZN(n8982) );
  INV_X1 U10003 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8900) );
  AOI22_X1 U10004 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_113), .B1(n8900), 
        .B2(keyinput_114), .ZN(n8899) );
  OAI221_X1 U10005 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(n8900), .C2(keyinput_114), .A(n8899), .ZN(n8903) );
  AOI22_X1 U10006 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_115), .B1(n8999), .B2(keyinput_112), .ZN(n8901) );
  OAI221_X1 U10007 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        n8999), .C2(keyinput_112), .A(n8901), .ZN(n8902) );
  AOI211_X1 U10008 ( .C1(keyinput_116), .C2(P2_REG3_REG_4__SCAN_IN), .A(n8903), 
        .B(n8902), .ZN(n8904) );
  OAI21_X1 U10009 ( .B1(keyinput_116), .B2(P2_REG3_REG_4__SCAN_IN), .A(n8904), 
        .ZN(n8979) );
  XNOR2_X1 U10010 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_103), .ZN(n8969)
         );
  INV_X1 U10011 ( .A(keyinput_102), .ZN(n8963) );
  INV_X1 U10012 ( .A(keyinput_101), .ZN(n8961) );
  INV_X1 U10013 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9071) );
  INV_X1 U10014 ( .A(keyinput_100), .ZN(n8959) );
  INV_X1 U10015 ( .A(keyinput_99), .ZN(n8957) );
  OAI22_X1 U10016 ( .A1(SI_4_), .A2(keyinput_92), .B1(SI_3_), .B2(keyinput_93), 
        .ZN(n8905) );
  AOI221_X1 U10017 ( .B1(SI_4_), .B2(keyinput_92), .C1(keyinput_93), .C2(SI_3_), .A(n8905), .ZN(n8947) );
  OAI22_X1 U10018 ( .A1(n8907), .A2(keyinput_88), .B1(SI_9_), .B2(keyinput_87), 
        .ZN(n8906) );
  AOI221_X1 U10019 ( .B1(n8907), .B2(keyinput_88), .C1(keyinput_87), .C2(SI_9_), .A(n8906), .ZN(n8938) );
  XNOR2_X1 U10020 ( .A(SI_18_), .B(keyinput_78), .ZN(n8927) );
  INV_X1 U10021 ( .A(keyinput_77), .ZN(n8925) );
  INV_X1 U10022 ( .A(keyinput_72), .ZN(n8918) );
  OAI22_X1 U10023 ( .A1(SI_31_), .A2(keyinput_65), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n8908) );
  AOI221_X1 U10024 ( .B1(SI_31_), .B2(keyinput_65), .C1(keyinput_64), .C2(
        P2_WR_REG_SCAN_IN), .A(n8908), .ZN(n8916) );
  AOI22_X1 U10025 ( .A1(SI_25_), .A2(keyinput_71), .B1(SI_26_), .B2(
        keyinput_70), .ZN(n8909) );
  OAI221_X1 U10026 ( .B1(SI_25_), .B2(keyinput_71), .C1(SI_26_), .C2(
        keyinput_70), .A(n8909), .ZN(n8915) );
  AOI22_X1 U10027 ( .A1(SI_29_), .A2(keyinput_67), .B1(SI_28_), .B2(
        keyinput_68), .ZN(n8910) );
  OAI221_X1 U10028 ( .B1(SI_29_), .B2(keyinput_67), .C1(SI_28_), .C2(
        keyinput_68), .A(n8910), .ZN(n8914) );
  AOI22_X1 U10029 ( .A1(n8912), .A2(keyinput_69), .B1(keyinput_66), .B2(n9010), 
        .ZN(n8911) );
  OAI221_X1 U10030 ( .B1(n8912), .B2(keyinput_69), .C1(n9010), .C2(keyinput_66), .A(n8911), .ZN(n8913) );
  NOR4_X1 U10031 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n8917)
         );
  AOI221_X1 U10032 ( .B1(SI_24_), .B2(n8918), .C1(n9017), .C2(keyinput_72), 
        .A(n8917), .ZN(n8923) );
  AOI22_X1 U10033 ( .A1(SI_22_), .A2(keyinput_74), .B1(SI_23_), .B2(
        keyinput_73), .ZN(n8919) );
  OAI221_X1 U10034 ( .B1(SI_22_), .B2(keyinput_74), .C1(SI_23_), .C2(
        keyinput_73), .A(n8919), .ZN(n8922) );
  OAI22_X1 U10035 ( .A1(SI_21_), .A2(keyinput_75), .B1(keyinput_76), .B2(
        SI_20_), .ZN(n8920) );
  AOI221_X1 U10036 ( .B1(SI_21_), .B2(keyinput_75), .C1(SI_20_), .C2(
        keyinput_76), .A(n8920), .ZN(n8921) );
  OAI21_X1 U10037 ( .B1(n8923), .B2(n8922), .A(n8921), .ZN(n8924) );
  OAI221_X1 U10038 ( .B1(SI_19_), .B2(n8925), .C1(n9025), .C2(keyinput_77), 
        .A(n8924), .ZN(n8926) );
  AOI22_X1 U10039 ( .A1(n8927), .A2(n8926), .B1(SI_16_), .B2(keyinput_80), 
        .ZN(n8928) );
  OAI21_X1 U10040 ( .B1(SI_16_), .B2(keyinput_80), .A(n8928), .ZN(n8936) );
  INV_X1 U10041 ( .A(SI_15_), .ZN(n9032) );
  AOI22_X1 U10042 ( .A1(n9032), .A2(keyinput_81), .B1(n8930), .B2(keyinput_79), 
        .ZN(n8929) );
  OAI221_X1 U10043 ( .B1(n9032), .B2(keyinput_81), .C1(n8930), .C2(keyinput_79), .A(n8929), .ZN(n8935) );
  OAI22_X1 U10044 ( .A1(n9035), .A2(keyinput_85), .B1(keyinput_83), .B2(SI_13_), .ZN(n8931) );
  AOI221_X1 U10045 ( .B1(n9035), .B2(keyinput_85), .C1(SI_13_), .C2(
        keyinput_83), .A(n8931), .ZN(n8934) );
  OAI22_X1 U10046 ( .A1(SI_14_), .A2(keyinput_82), .B1(keyinput_84), .B2(
        SI_12_), .ZN(n8932) );
  AOI221_X1 U10047 ( .B1(SI_14_), .B2(keyinput_82), .C1(SI_12_), .C2(
        keyinput_84), .A(n8932), .ZN(n8933) );
  OAI211_X1 U10048 ( .C1(n8936), .C2(n8935), .A(n8934), .B(n8933), .ZN(n8937)
         );
  OAI211_X1 U10049 ( .C1(n8940), .C2(keyinput_86), .A(n8938), .B(n8937), .ZN(
        n8939) );
  AOI21_X1 U10050 ( .B1(n8940), .B2(keyinput_86), .A(n8939), .ZN(n8944) );
  INV_X1 U10051 ( .A(SI_7_), .ZN(n9048) );
  INV_X1 U10052 ( .A(SI_6_), .ZN(n8942) );
  AOI22_X1 U10053 ( .A1(n9048), .A2(keyinput_89), .B1(keyinput_90), .B2(n8942), 
        .ZN(n8941) );
  OAI221_X1 U10054 ( .B1(n9048), .B2(keyinput_89), .C1(n8942), .C2(keyinput_90), .A(n8941), .ZN(n8943) );
  AOI211_X1 U10055 ( .C1(SI_5_), .C2(keyinput_91), .A(n8944), .B(n8943), .ZN(
        n8945) );
  OAI21_X1 U10056 ( .B1(SI_5_), .B2(keyinput_91), .A(n8945), .ZN(n8946) );
  AOI22_X1 U10057 ( .A1(n8947), .A2(n8946), .B1(keyinput_94), .B2(SI_2_), .ZN(
        n8948) );
  OAI21_X1 U10058 ( .B1(keyinput_94), .B2(SI_2_), .A(n8948), .ZN(n8951) );
  INV_X1 U10059 ( .A(keyinput_95), .ZN(n8949) );
  MUX2_X1 U10060 ( .A(keyinput_95), .B(n8949), .S(SI_1_), .Z(n8950) );
  NAND2_X1 U10061 ( .A1(n8951), .A2(n8950), .ZN(n8954) );
  INV_X1 U10062 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10424) );
  OAI22_X1 U10063 ( .A1(n10424), .A2(keyinput_97), .B1(SI_0_), .B2(keyinput_96), .ZN(n8952) );
  AOI221_X1 U10064 ( .B1(n10424), .B2(keyinput_97), .C1(keyinput_96), .C2(
        SI_0_), .A(n8952), .ZN(n8953) );
  AOI22_X1 U10065 ( .A1(n8954), .A2(n8953), .B1(keyinput_98), .B2(P2_U3151), 
        .ZN(n8955) );
  OAI21_X1 U10066 ( .B1(P2_U3151), .B2(keyinput_98), .A(n8955), .ZN(n8956) );
  OAI221_X1 U10067 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(n8957), .C1(n9065), .C2(
        keyinput_99), .A(n8956), .ZN(n8958) );
  OAI221_X1 U10068 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n8959), .C1(n9068), 
        .C2(keyinput_100), .A(n8958), .ZN(n8960) );
  OAI221_X1 U10069 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(n8961), .C1(n9071), 
        .C2(keyinput_101), .A(n8960), .ZN(n8962) );
  OAI221_X1 U10070 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .C1(
        n9075), .C2(n8963), .A(n8962), .ZN(n8968) );
  AOI22_X1 U10071 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_104), .B1(n9078), 
        .B2(keyinput_107), .ZN(n8964) );
  OAI221_X1 U10072 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .C1(n9078), .C2(keyinput_107), .A(n8964), .ZN(n8967) );
  AOI22_X1 U10073 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .ZN(n8965) );
  OAI221_X1 U10074 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_106), .A(n8965), .ZN(n8966) );
  AOI211_X1 U10075 ( .C1(n8969), .C2(n8968), .A(n8967), .B(n8966), .ZN(n8972)
         );
  INV_X1 U10076 ( .A(keyinput_108), .ZN(n8970) );
  MUX2_X1 U10077 ( .A(keyinput_108), .B(n8970), .S(P2_REG3_REG_1__SCAN_IN), 
        .Z(n8971) );
  NOR2_X1 U10078 ( .A1(n8972), .A2(n8971), .ZN(n8976) );
  AOI22_X1 U10079 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_110), .B1(n8974), .B2(keyinput_109), .ZN(n8973) );
  OAI221_X1 U10080 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        n8974), .C2(keyinput_109), .A(n8973), .ZN(n8975) );
  OAI22_X1 U10081 ( .A1(n8976), .A2(n8975), .B1(keyinput_111), .B2(n9092), 
        .ZN(n8977) );
  AOI21_X1 U10082 ( .B1(keyinput_111), .B2(n9092), .A(n8977), .ZN(n8978) );
  OAI22_X1 U10083 ( .A1(keyinput_117), .A2(n6474), .B1(n8979), .B2(n8978), 
        .ZN(n8980) );
  AOI21_X1 U10084 ( .B1(keyinput_117), .B2(n6474), .A(n8980), .ZN(n8981) );
  OAI22_X1 U10085 ( .A1(keyinput_120), .A2(n6525), .B1(n8982), .B2(n8981), 
        .ZN(n8983) );
  AOI21_X1 U10086 ( .B1(keyinput_120), .B2(n6525), .A(n8983), .ZN(n8988) );
  XOR2_X1 U10087 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_123), .Z(n8987) );
  AND2_X1 U10088 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_121), .ZN(n8986)
         );
  INV_X1 U10089 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8984) );
  XNOR2_X1 U10090 ( .A(keyinput_122), .B(n8984), .ZN(n8985) );
  NOR4_X1 U10091 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n8989)
         );
  OAI21_X1 U10092 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .A(n8989), 
        .ZN(n8990) );
  AOI22_X1 U10093 ( .A1(n8991), .A2(n8990), .B1(keyinput_126), .B2(
        P2_REG3_REG_26__SCAN_IN), .ZN(n8992) );
  OAI21_X1 U10094 ( .B1(keyinput_126), .B2(P2_REG3_REG_26__SCAN_IN), .A(n8992), 
        .ZN(n8994) );
  AOI21_X1 U10095 ( .B1(keyinput_127), .B2(n8994), .A(keyinput_63), .ZN(n8997)
         );
  INV_X1 U10096 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8996) );
  INV_X1 U10097 ( .A(keyinput_127), .ZN(n8993) );
  AOI21_X1 U10098 ( .B1(n8994), .B2(n8993), .A(n8996), .ZN(n8995) );
  AOI22_X1 U10099 ( .A1(n8997), .A2(n8996), .B1(n8995), .B2(keyinput_63), .ZN(
        n9110) );
  AOI22_X1 U10100 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_52), .B1(n8999), 
        .B2(keyinput_48), .ZN(n8998) );
  OAI221_X1 U10101 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(n8999), 
        .C2(keyinput_48), .A(n8998), .ZN(n9002) );
  AOI22_X1 U10102 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_49), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .ZN(n9000) );
  OAI221_X1 U10103 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n9000), .ZN(n9001) );
  AOI211_X1 U10104 ( .C1(keyinput_50), .C2(P2_REG3_REG_17__SCAN_IN), .A(n9002), 
        .B(n9001), .ZN(n9003) );
  OAI21_X1 U10105 ( .B1(keyinput_50), .B2(P2_REG3_REG_17__SCAN_IN), .A(n9003), 
        .ZN(n9094) );
  XNOR2_X1 U10106 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n9083)
         );
  INV_X1 U10107 ( .A(keyinput_38), .ZN(n9074) );
  INV_X1 U10108 ( .A(keyinput_37), .ZN(n9072) );
  INV_X1 U10109 ( .A(keyinput_36), .ZN(n9069) );
  INV_X1 U10110 ( .A(keyinput_35), .ZN(n9066) );
  XNOR2_X1 U10111 ( .A(SI_18_), .B(keyinput_14), .ZN(n9028) );
  INV_X1 U10112 ( .A(keyinput_13), .ZN(n9026) );
  OAI22_X1 U10113 ( .A1(n9005), .A2(keyinput_9), .B1(SI_22_), .B2(keyinput_10), 
        .ZN(n9004) );
  AOI221_X1 U10114 ( .B1(n9005), .B2(keyinput_9), .C1(keyinput_10), .C2(SI_22_), .A(n9004), .ZN(n9023) );
  INV_X1 U10115 ( .A(keyinput_8), .ZN(n9018) );
  OAI22_X1 U10116 ( .A1(SI_26_), .A2(keyinput_6), .B1(keyinput_3), .B2(SI_29_), 
        .ZN(n9006) );
  AOI221_X1 U10117 ( .B1(SI_26_), .B2(keyinput_6), .C1(SI_29_), .C2(keyinput_3), .A(n9006), .ZN(n9015) );
  OAI22_X1 U10118 ( .A1(n9008), .A2(keyinput_7), .B1(keyinput_5), .B2(SI_27_), 
        .ZN(n9007) );
  AOI221_X1 U10119 ( .B1(n9008), .B2(keyinput_7), .C1(SI_27_), .C2(keyinput_5), 
        .A(n9007), .ZN(n9014) );
  OAI22_X1 U10120 ( .A1(n8137), .A2(keyinput_4), .B1(n9010), .B2(keyinput_2), 
        .ZN(n9009) );
  AOI221_X1 U10121 ( .B1(n8137), .B2(keyinput_4), .C1(keyinput_2), .C2(n9010), 
        .A(n9009), .ZN(n9013) );
  AOI22_X1 U10122 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n9011) );
  OAI221_X1 U10123 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n9011), .ZN(n9012) );
  NAND4_X1 U10124 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n9016)
         );
  OAI221_X1 U10125 ( .B1(SI_24_), .B2(n9018), .C1(n9017), .C2(keyinput_8), .A(
        n9016), .ZN(n9022) );
  AOI22_X1 U10126 ( .A1(SI_21_), .A2(keyinput_11), .B1(n9020), .B2(keyinput_12), .ZN(n9019) );
  OAI221_X1 U10127 ( .B1(SI_21_), .B2(keyinput_11), .C1(n9020), .C2(
        keyinput_12), .A(n9019), .ZN(n9021) );
  AOI21_X1 U10128 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(n9024) );
  AOI221_X1 U10129 ( .B1(SI_19_), .B2(n9026), .C1(n9025), .C2(keyinput_13), 
        .A(n9024), .ZN(n9027) );
  OAI22_X1 U10130 ( .A1(n9028), .A2(n9027), .B1(n9030), .B2(keyinput_16), .ZN(
        n9029) );
  AOI21_X1 U10131 ( .B1(n9030), .B2(keyinput_16), .A(n9029), .ZN(n9042) );
  OAI22_X1 U10132 ( .A1(n9032), .A2(keyinput_17), .B1(keyinput_15), .B2(SI_17_), .ZN(n9031) );
  AOI221_X1 U10133 ( .B1(n9032), .B2(keyinput_17), .C1(SI_17_), .C2(
        keyinput_15), .A(n9031), .ZN(n9041) );
  AOI22_X1 U10134 ( .A1(n9035), .A2(keyinput_21), .B1(n9034), .B2(keyinput_18), 
        .ZN(n9033) );
  OAI221_X1 U10135 ( .B1(n9035), .B2(keyinput_21), .C1(n9034), .C2(keyinput_18), .A(n9033), .ZN(n9040) );
  INV_X1 U10136 ( .A(SI_13_), .ZN(n9038) );
  AOI22_X1 U10137 ( .A1(n9038), .A2(keyinput_19), .B1(keyinput_20), .B2(n9037), 
        .ZN(n9036) );
  OAI221_X1 U10138 ( .B1(n9038), .B2(keyinput_19), .C1(n9037), .C2(keyinput_20), .A(n9036), .ZN(n9039) );
  AOI211_X1 U10139 ( .C1(n9042), .C2(n9041), .A(n9040), .B(n9039), .ZN(n9046)
         );
  OAI22_X1 U10140 ( .A1(SI_10_), .A2(keyinput_22), .B1(SI_8_), .B2(keyinput_24), .ZN(n9043) );
  AOI221_X1 U10141 ( .B1(SI_10_), .B2(keyinput_22), .C1(keyinput_24), .C2(
        SI_8_), .A(n9043), .ZN(n9044) );
  OAI21_X1 U10142 ( .B1(keyinput_23), .B2(SI_9_), .A(n9044), .ZN(n9045) );
  AOI211_X1 U10143 ( .C1(keyinput_23), .C2(SI_9_), .A(n9046), .B(n9045), .ZN(
        n9050) );
  AOI22_X1 U10144 ( .A1(SI_5_), .A2(keyinput_27), .B1(n9048), .B2(keyinput_25), 
        .ZN(n9047) );
  OAI221_X1 U10145 ( .B1(SI_5_), .B2(keyinput_27), .C1(n9048), .C2(keyinput_25), .A(n9047), .ZN(n9049) );
  AOI211_X1 U10146 ( .C1(SI_6_), .C2(keyinput_26), .A(n9050), .B(n9049), .ZN(
        n9051) );
  OAI21_X1 U10147 ( .B1(SI_6_), .B2(keyinput_26), .A(n9051), .ZN(n9054) );
  OAI22_X1 U10148 ( .A1(SI_4_), .A2(keyinput_28), .B1(SI_3_), .B2(keyinput_29), 
        .ZN(n9052) );
  AOI221_X1 U10149 ( .B1(SI_4_), .B2(keyinput_28), .C1(keyinput_29), .C2(SI_3_), .A(n9052), .ZN(n9053) );
  AND2_X1 U10150 ( .A1(n9054), .A2(n9053), .ZN(n9059) );
  XNOR2_X1 U10151 ( .A(n9055), .B(keyinput_30), .ZN(n9058) );
  INV_X1 U10152 ( .A(keyinput_31), .ZN(n9056) );
  MUX2_X1 U10153 ( .A(n9056), .B(keyinput_31), .S(SI_1_), .Z(n9057) );
  OAI21_X1 U10154 ( .B1(n9059), .B2(n9058), .A(n9057), .ZN(n9062) );
  OAI22_X1 U10155 ( .A1(n10424), .A2(keyinput_33), .B1(SI_0_), .B2(keyinput_32), .ZN(n9060) );
  AOI221_X1 U10156 ( .B1(n10424), .B2(keyinput_33), .C1(keyinput_32), .C2(
        SI_0_), .A(n9060), .ZN(n9061) );
  AOI22_X1 U10157 ( .A1(n9062), .A2(n9061), .B1(keyinput_34), .B2(P2_U3151), 
        .ZN(n9063) );
  OAI21_X1 U10158 ( .B1(P2_U3151), .B2(keyinput_34), .A(n9063), .ZN(n9064) );
  OAI221_X1 U10159 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(n9066), .C1(n9065), .C2(
        keyinput_35), .A(n9064), .ZN(n9067) );
  OAI221_X1 U10160 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n9069), .C1(n9068), 
        .C2(keyinput_36), .A(n9067), .ZN(n9070) );
  OAI221_X1 U10161 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(n9072), .C1(n9071), 
        .C2(keyinput_37), .A(n9070), .ZN(n9073) );
  OAI221_X1 U10162 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(n9075), .C2(n9074), .A(n9073), .ZN(n9082) );
  AOI22_X1 U10163 ( .A1(n9078), .A2(keyinput_43), .B1(keyinput_40), .B2(n9077), 
        .ZN(n9076) );
  OAI221_X1 U10164 ( .B1(n9078), .B2(keyinput_43), .C1(n9077), .C2(keyinput_40), .A(n9076), .ZN(n9081) );
  AOI22_X1 U10165 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_41), .B1(n6660), 
        .B2(keyinput_42), .ZN(n9079) );
  OAI221_X1 U10166 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .C1(n6660), .C2(keyinput_42), .A(n9079), .ZN(n9080) );
  AOI211_X1 U10167 ( .C1(n9083), .C2(n9082), .A(n9081), .B(n9080), .ZN(n9086)
         );
  INV_X1 U10168 ( .A(keyinput_44), .ZN(n9084) );
  MUX2_X1 U10169 ( .A(keyinput_44), .B(n9084), .S(P2_REG3_REG_1__SCAN_IN), .Z(
        n9085) );
  NOR2_X1 U10170 ( .A1(n9086), .A2(n9085), .ZN(n9090) );
  INV_X1 U10171 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9088) );
  AOI22_X1 U10172 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(n9088), 
        .B2(keyinput_46), .ZN(n9087) );
  OAI221_X1 U10173 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(n9088), .C2(keyinput_46), .A(n9087), .ZN(n9089) );
  OAI22_X1 U10174 ( .A1(n9090), .A2(n9089), .B1(keyinput_47), .B2(n9092), .ZN(
        n9091) );
  AOI21_X1 U10175 ( .B1(keyinput_47), .B2(n9092), .A(n9091), .ZN(n9093) );
  OAI22_X1 U10176 ( .A1(keyinput_53), .A2(n6474), .B1(n9094), .B2(n9093), .ZN(
        n9095) );
  AOI21_X1 U10177 ( .B1(keyinput_53), .B2(n6474), .A(n9095), .ZN(n9099) );
  XNOR2_X1 U10178 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n9097)
         );
  XNOR2_X1 U10179 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n9096) );
  NAND2_X1 U10180 ( .A1(n9097), .A2(n9096), .ZN(n9098) );
  OAI22_X1 U10181 ( .A1(n9099), .A2(n9098), .B1(keyinput_56), .B2(n6525), .ZN(
        n9100) );
  AOI21_X1 U10182 ( .B1(keyinput_56), .B2(n6525), .A(n9100), .ZN(n9103) );
  AOI22_X1 U10183 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .ZN(n9101) );
  OAI221_X1 U10184 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n9101), .ZN(n9102) );
  AOI211_X1 U10185 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n9103), 
        .B(n9102), .ZN(n9104) );
  OAI21_X1 U10186 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .A(n9104), 
        .ZN(n9108) );
  OAI22_X1 U10187 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(
        keyinput_61), .B2(P2_REG3_REG_6__SCAN_IN), .ZN(n9105) );
  AOI221_X1 U10188 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n9105), .ZN(n9107) );
  XNOR2_X1 U10189 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n9106)
         );
  AOI21_X1 U10190 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9109) );
  NOR2_X1 U10191 ( .A1(n9110), .A2(n9109), .ZN(n9113) );
  MUX2_X1 U10192 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9111), .S(n10640), .Z(
        n9112) );
  XOR2_X1 U10193 ( .A(n9113), .B(n9112), .Z(P2_U3449) );
  MUX2_X1 U10194 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9114), .S(n10640), .Z(
        P2_U3448) );
  INV_X1 U10195 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9116) );
  MUX2_X1 U10196 ( .A(n9116), .B(n9115), .S(n10640), .Z(n9117) );
  OAI21_X1 U10197 ( .B1(n9118), .B2(n9134), .A(n9117), .ZN(P2_U3447) );
  INV_X1 U10198 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9120) );
  MUX2_X1 U10199 ( .A(n9120), .B(n9119), .S(n10640), .Z(n9121) );
  OAI21_X1 U10200 ( .B1(n9122), .B2(n9134), .A(n9121), .ZN(P2_U3446) );
  INV_X1 U10201 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9124) );
  MUX2_X1 U10202 ( .A(n9124), .B(n9123), .S(n10640), .Z(n9125) );
  OAI21_X1 U10203 ( .B1(n9126), .B2(n9134), .A(n9125), .ZN(P2_U3444) );
  INV_X1 U10204 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9128) );
  MUX2_X1 U10205 ( .A(n9128), .B(n9127), .S(n10640), .Z(n9129) );
  OAI21_X1 U10206 ( .B1(n9130), .B2(n9134), .A(n9129), .ZN(P2_U3441) );
  MUX2_X1 U10207 ( .A(n9132), .B(n9131), .S(n10640), .Z(n9133) );
  OAI21_X1 U10208 ( .B1(n9135), .B2(n9134), .A(n9133), .ZN(P2_U3438) );
  MUX2_X1 U10209 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9136), .S(n10640), .Z(
        P2_U3435) );
  MUX2_X1 U10210 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9137), .S(n10640), .Z(
        P2_U3426) );
  INV_X1 U10211 ( .A(n10016), .ZN(n9143) );
  NOR4_X1 U10212 ( .A1(n9138), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9139), .A4(
        P2_U3151), .ZN(n9140) );
  AOI21_X1 U10213 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9141), .A(n9140), .ZN(
        n9142) );
  OAI21_X1 U10214 ( .B1(n9143), .B2(n9147), .A(n9142), .ZN(P2_U3264) );
  INV_X1 U10215 ( .A(n9144), .ZN(n10023) );
  OAI222_X1 U10216 ( .A1(n9147), .A2(n10023), .B1(P2_U3151), .B2(n9146), .C1(
        n9145), .C2(n9153), .ZN(P2_U3266) );
  NAND2_X1 U10217 ( .A1(n9149), .A2(n9148), .ZN(n9151) );
  OAI211_X1 U10218 ( .C1(n9153), .C2(n9152), .A(n9151), .B(n9150), .ZN(
        P2_U3267) );
  MUX2_X1 U10219 ( .A(n9154), .B(n4996), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10220 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9161) );
  AOI22_X1 U10221 ( .A1(n9681), .A2(n9213), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9159) );
  AOI22_X1 U10222 ( .A1(n9680), .A2(n9261), .B1(n9262), .B2(n9800), .ZN(n9158)
         );
  OAI211_X1 U10223 ( .C1(n5168), .C2(n9243), .A(n9159), .B(n9158), .ZN(n9160)
         );
  AOI21_X1 U10224 ( .B1(n9161), .B2(n9235), .A(n9160), .ZN(n9162) );
  INV_X1 U10225 ( .A(n9162), .ZN(P1_U3216) );
  XOR2_X1 U10226 ( .A(n9164), .B(n9163), .Z(n9168) );
  NAND2_X1 U10227 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9663) );
  OAI21_X1 U10228 ( .B1(n9264), .B2(n9867), .A(n9663), .ZN(n9166) );
  OAI22_X1 U10229 ( .A1(n9250), .A2(n9866), .B1(n9251), .B2(n9860), .ZN(n9165)
         );
  AOI211_X1 U10230 ( .C1(n9960), .C2(n9266), .A(n9166), .B(n9165), .ZN(n9167)
         );
  OAI21_X1 U10231 ( .B1(n9168), .B2(n9268), .A(n9167), .ZN(P1_U3219) );
  INV_X1 U10232 ( .A(n9196), .ZN(n9180) );
  NAND2_X1 U10233 ( .A1(n9910), .A2(n9169), .ZN(n9172) );
  OR2_X1 U10234 ( .A1(n9741), .A2(n9170), .ZN(n9171) );
  NAND2_X1 U10235 ( .A1(n9172), .A2(n9171), .ZN(n9174) );
  XNOR2_X1 U10236 ( .A(n9174), .B(n9173), .ZN(n9178) );
  NAND2_X1 U10237 ( .A1(n9910), .A2(n6214), .ZN(n9175) );
  OAI21_X1 U10238 ( .B1(n9741), .B2(n9176), .A(n9175), .ZN(n9177) );
  XNOR2_X1 U10239 ( .A(n9178), .B(n9177), .ZN(n9195) );
  INV_X1 U10240 ( .A(n9195), .ZN(n9179) );
  NAND4_X1 U10241 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9235), .ZN(n9200)
         );
  NAND3_X1 U10242 ( .A1(n9182), .A2(n9235), .A3(n9195), .ZN(n9199) );
  INV_X1 U10243 ( .A(n9183), .ZN(n9688) );
  NAND3_X1 U10244 ( .A1(n9688), .A2(n9184), .A3(P1_REG3_REG_28__SCAN_IN), .ZN(
        n9191) );
  INV_X1 U10245 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U10246 ( .A1(n5786), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U10247 ( .A1(n4918), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9185) );
  OAI211_X1 U10248 ( .C1(n9188), .C2(n9187), .A(n9186), .B(n9185), .ZN(n9189)
         );
  INV_X1 U10249 ( .A(n9189), .ZN(n9190) );
  INV_X1 U10250 ( .A(n9276), .ZN(n9727) );
  AOI22_X1 U10251 ( .A1(n9727), .A2(n9213), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9192) );
  OAI21_X1 U10252 ( .B1(n9750), .B2(n9250), .A(n9192), .ZN(n9194) );
  NOR2_X1 U10253 ( .A1(n9722), .A2(n9243), .ZN(n9193) );
  AOI211_X1 U10254 ( .C1(n9262), .C2(n9720), .A(n9194), .B(n9193), .ZN(n9198)
         );
  NAND3_X1 U10255 ( .A1(n9196), .A2(n9235), .A3(n9195), .ZN(n9197) );
  NAND4_X1 U10256 ( .A1(n9200), .A2(n9199), .A3(n9198), .A4(n9197), .ZN(
        P1_U3220) );
  OAI211_X1 U10257 ( .C1(n9203), .C2(n9202), .A(n9201), .B(n9235), .ZN(n9207)
         );
  AOI22_X1 U10258 ( .A1(n9261), .A2(n9679), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9206) );
  AOI22_X1 U10259 ( .A1(n9680), .A2(n9213), .B1(n9262), .B2(n9836), .ZN(n9205)
         );
  NAND2_X1 U10260 ( .A1(n9950), .A2(n9266), .ZN(n9204) );
  NAND4_X1 U10261 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), .ZN(
        P1_U3223) );
  OAI21_X1 U10262 ( .B1(n9209), .B2(n9208), .A(n6270), .ZN(n9210) );
  NAND2_X1 U10263 ( .A1(n9210), .A2(n9235), .ZN(n9215) );
  AOI22_X1 U10264 ( .A1(n9681), .A2(n9261), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9211) );
  OAI21_X1 U10265 ( .B1(n9768), .B2(n9251), .A(n9211), .ZN(n9212) );
  AOI21_X1 U10266 ( .B1(n9684), .B2(n9213), .A(n9212), .ZN(n9214) );
  OAI211_X1 U10267 ( .C1(n5164), .C2(n9243), .A(n9215), .B(n9214), .ZN(
        P1_U3225) );
  NAND2_X1 U10268 ( .A1(n4976), .A2(n9216), .ZN(n9217) );
  XNOR2_X1 U10269 ( .A(n9218), .B(n9217), .ZN(n9223) );
  AOI22_X1 U10270 ( .A1(n9262), .A2(n9219), .B1(n9261), .B2(n9559), .ZN(n9220)
         );
  NAND2_X1 U10271 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10203)
         );
  OAI211_X1 U10272 ( .C1(n9866), .C2(n9264), .A(n9220), .B(n10203), .ZN(n9221)
         );
  AOI21_X1 U10273 ( .B1(n9970), .B2(n9266), .A(n9221), .ZN(n9222) );
  OAI21_X1 U10274 ( .B1(n9223), .B2(n9268), .A(n9222), .ZN(P1_U3228) );
  NAND2_X1 U10275 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  XNOR2_X1 U10276 ( .A(n9224), .B(n9227), .ZN(n9232) );
  OAI22_X1 U10277 ( .A1(n9809), .A2(n9250), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9228), .ZN(n9230) );
  OAI22_X1 U10278 ( .A1(n9786), .A2(n9264), .B1(n9251), .B2(n9777), .ZN(n9229)
         );
  AOI211_X1 U10279 ( .C1(n9934), .C2(n9266), .A(n9230), .B(n9229), .ZN(n9231)
         );
  OAI21_X1 U10280 ( .B1(n9232), .B2(n9268), .A(n9231), .ZN(P1_U3229) );
  XNOR2_X1 U10281 ( .A(n9233), .B(n9234), .ZN(n9236) );
  NAND2_X1 U10282 ( .A1(n9236), .A2(n9235), .ZN(n9242) );
  NAND2_X1 U10283 ( .A1(n9261), .A2(n9888), .ZN(n9237) );
  OAI21_X1 U10284 ( .B1(n9251), .B2(n9846), .A(n9237), .ZN(n9240) );
  OAI22_X1 U10285 ( .A1(n9264), .A2(n9808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9238), .ZN(n9239) );
  NOR2_X1 U10286 ( .A1(n9240), .A2(n9239), .ZN(n9241) );
  OAI211_X1 U10287 ( .C1(n9849), .C2(n9243), .A(n9242), .B(n9241), .ZN(
        P1_U3233) );
  INV_X1 U10288 ( .A(n9244), .ZN(n9246) );
  NOR2_X1 U10289 ( .A1(n9246), .A2(n9245), .ZN(n9248) );
  XNOR2_X1 U10290 ( .A(n9248), .B(n9247), .ZN(n9255) );
  OAI22_X1 U10291 ( .A1(n9250), .A2(n9808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9249), .ZN(n9253) );
  OAI22_X1 U10292 ( .A1(n9809), .A2(n9264), .B1(n9251), .B2(n9820), .ZN(n9252)
         );
  AOI211_X1 U10293 ( .C1(n9943), .C2(n9266), .A(n9253), .B(n9252), .ZN(n9254)
         );
  OAI21_X1 U10294 ( .B1(n9255), .B2(n9268), .A(n9254), .ZN(P1_U3235) );
  INV_X1 U10295 ( .A(n9256), .ZN(n9258) );
  NAND2_X1 U10296 ( .A1(n9258), .A2(n9257), .ZN(n9260) );
  XNOR2_X1 U10297 ( .A(n9260), .B(n9259), .ZN(n9269) );
  AOI22_X1 U10298 ( .A1(n9262), .A2(n9877), .B1(n9261), .B2(n9890), .ZN(n9263)
         );
  NAND2_X1 U10299 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10215)
         );
  OAI211_X1 U10300 ( .C1(n9678), .C2(n9264), .A(n9263), .B(n10215), .ZN(n9265)
         );
  AOI21_X1 U10301 ( .B1(n9964), .B2(n9266), .A(n9265), .ZN(n9267) );
  OAI21_X1 U10302 ( .B1(n9269), .B2(n9268), .A(n9267), .ZN(P1_U3238) );
  INV_X1 U10303 ( .A(n9667), .ZN(n9902) );
  NAND2_X1 U10304 ( .A1(n4916), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U10305 ( .A1(n5786), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U10306 ( .A1(n4918), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9270) );
  AND3_X1 U10307 ( .A1(n9272), .A2(n9271), .A3(n9270), .ZN(n9708) );
  OR2_X1 U10308 ( .A1(n9902), .A2(n9708), .ZN(n9538) );
  INV_X1 U10309 ( .A(n9469), .ZN(n9389) );
  INV_X1 U10310 ( .A(n9708), .ZN(n9557) );
  AOI21_X1 U10311 ( .B1(n9557), .B2(n9556), .A(n9667), .ZN(n9466) );
  INV_X1 U10312 ( .A(n9466), .ZN(n9388) );
  MUX2_X1 U10313 ( .A(n9389), .B(n9388), .S(n9383), .Z(n9391) );
  NAND2_X1 U10314 ( .A1(n10016), .A2(n9273), .ZN(n9275) );
  INV_X1 U10315 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10012) );
  OR2_X1 U10316 ( .A1(n5778), .A2(n10012), .ZN(n9274) );
  NAND2_X1 U10317 ( .A1(n9275), .A2(n9274), .ZN(n9897) );
  INV_X1 U10318 ( .A(n9897), .ZN(n9669) );
  AND2_X1 U10319 ( .A1(n9669), .A2(n9556), .ZN(n9472) );
  INV_X1 U10320 ( .A(n9472), .ZN(n9540) );
  NAND2_X1 U10321 ( .A1(n9907), .A2(n9276), .ZN(n9531) );
  MUX2_X1 U10322 ( .A(n9531), .B(n9458), .S(n9383), .Z(n9387) );
  NAND2_X1 U10323 ( .A1(n9929), .A2(n9786), .ZN(n9699) );
  NAND2_X1 U10324 ( .A1(n9934), .A2(n9798), .ZN(n9446) );
  AND2_X1 U10325 ( .A1(n9699), .A2(n9446), .ZN(n9278) );
  OR2_X1 U10326 ( .A1(n9929), .A2(n9786), .ZN(n9443) );
  NAND2_X1 U10327 ( .A1(n9443), .A2(n9699), .ZN(n9764) );
  NOR2_X1 U10328 ( .A1(n9764), .A2(n5315), .ZN(n9277) );
  MUX2_X1 U10329 ( .A(n9278), .B(n9277), .S(n9394), .Z(n9379) );
  MUX2_X1 U10330 ( .A(n9394), .B(n9573), .S(n9279), .Z(n9281) );
  NAND2_X1 U10331 ( .A1(n9573), .A2(n9394), .ZN(n9280) );
  AND2_X1 U10332 ( .A1(n9281), .A2(n9280), .ZN(n9291) );
  INV_X1 U10333 ( .A(n9291), .ZN(n9282) );
  NAND2_X1 U10334 ( .A1(n7242), .A2(n9282), .ZN(n9283) );
  NAND3_X1 U10335 ( .A1(n9283), .A2(n9489), .A3(n9485), .ZN(n9284) );
  NAND4_X1 U10336 ( .A1(n9284), .A2(n9402), .A3(n9491), .A4(n9290), .ZN(n9288)
         );
  INV_X1 U10337 ( .A(n9493), .ZN(n9286) );
  INV_X1 U10338 ( .A(n9494), .ZN(n9285) );
  AOI21_X1 U10339 ( .B1(n9286), .B2(n9497), .A(n9285), .ZN(n9287) );
  NAND2_X1 U10340 ( .A1(n9288), .A2(n9287), .ZN(n9297) );
  AND2_X1 U10341 ( .A1(n9290), .A2(n9289), .ZN(n9487) );
  OAI21_X1 U10342 ( .B1(n9291), .B2(n7242), .A(n9487), .ZN(n9292) );
  NAND3_X1 U10343 ( .A1(n9292), .A2(n9489), .A3(n9493), .ZN(n9293) );
  NAND2_X1 U10344 ( .A1(n9293), .A2(n9491), .ZN(n9294) );
  NAND2_X1 U10345 ( .A1(n9294), .A2(n9402), .ZN(n9295) );
  NAND2_X1 U10346 ( .A1(n9295), .A2(n9497), .ZN(n9296) );
  MUX2_X1 U10347 ( .A(n9297), .B(n9296), .S(n9394), .Z(n9301) );
  NOR2_X1 U10348 ( .A1(n9405), .A2(n9383), .ZN(n9298) );
  NOR2_X1 U10349 ( .A1(n10536), .A2(n9298), .ZN(n9299) );
  OAI21_X1 U10350 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9306) );
  OR2_X1 U10351 ( .A1(n9302), .A2(n9383), .ZN(n9305) );
  NOR2_X1 U10352 ( .A1(n9303), .A2(n9394), .ZN(n9304) );
  AOI21_X1 U10353 ( .B1(n9306), .B2(n9305), .A(n9304), .ZN(n9314) );
  OAI21_X1 U10354 ( .B1(n9394), .B2(n9308), .A(n9307), .ZN(n9313) );
  NAND3_X1 U10355 ( .A1(n9317), .A2(n9409), .A3(n9309), .ZN(n9311) );
  INV_X1 U10356 ( .A(n9315), .ZN(n9310) );
  AOI21_X1 U10357 ( .B1(n9311), .B2(n9394), .A(n9310), .ZN(n9312) );
  OAI21_X1 U10358 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9324) );
  NAND2_X1 U10359 ( .A1(n9503), .A2(n9315), .ZN(n9316) );
  NAND2_X1 U10360 ( .A1(n9316), .A2(n9317), .ZN(n9323) );
  OR2_X1 U10361 ( .A1(n9319), .A2(n9318), .ZN(n9505) );
  INV_X1 U10362 ( .A(n9409), .ZN(n9320) );
  AND2_X1 U10363 ( .A1(n9503), .A2(n9320), .ZN(n9321) );
  NOR2_X1 U10364 ( .A1(n9505), .A2(n9321), .ZN(n9322) );
  MUX2_X1 U10365 ( .A(n9323), .B(n9322), .S(n9383), .Z(n9329) );
  NAND3_X1 U10366 ( .A1(n9324), .A2(n9329), .A3(n9327), .ZN(n9332) );
  AND2_X1 U10367 ( .A1(n9335), .A2(n9325), .ZN(n9331) );
  NAND2_X1 U10368 ( .A1(n9503), .A2(n9326), .ZN(n9328) );
  NAND2_X1 U10369 ( .A1(n9333), .A2(n9327), .ZN(n9506) );
  AOI21_X1 U10370 ( .B1(n9329), .B2(n9328), .A(n9506), .ZN(n9330) );
  NAND2_X1 U10371 ( .A1(n9346), .A2(n9340), .ZN(n9483) );
  AOI21_X1 U10372 ( .B1(n9334), .B2(n9511), .A(n9483), .ZN(n9343) );
  AND2_X1 U10373 ( .A1(n9336), .A2(n9335), .ZN(n9509) );
  NAND2_X1 U10374 ( .A1(n9337), .A2(n9509), .ZN(n9338) );
  NAND2_X1 U10375 ( .A1(n9338), .A2(n9510), .ZN(n9341) );
  OR2_X1 U10376 ( .A1(n9514), .A2(n5303), .ZN(n9339) );
  AOI21_X1 U10377 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(n9342) );
  MUX2_X1 U10378 ( .A(n9343), .B(n9342), .S(n9383), .Z(n9344) );
  NAND2_X1 U10379 ( .A1(n9344), .A2(n5444), .ZN(n9352) );
  NAND2_X1 U10380 ( .A1(n9347), .A2(n9514), .ZN(n9345) );
  AND2_X1 U10381 ( .A1(n9345), .A2(n9517), .ZN(n9350) );
  NAND2_X1 U10382 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NAND2_X1 U10383 ( .A1(n9348), .A2(n9517), .ZN(n9349) );
  MUX2_X1 U10384 ( .A(n9350), .B(n9349), .S(n9383), .Z(n9351) );
  NAND2_X1 U10385 ( .A1(n9352), .A2(n9351), .ZN(n9354) );
  NAND2_X1 U10386 ( .A1(n9354), .A2(n9353), .ZN(n9358) );
  OR2_X1 U10387 ( .A1(n9964), .A2(n9866), .ZN(n9398) );
  AND2_X1 U10388 ( .A1(n9398), .A2(n9518), .ZN(n9356) );
  NAND2_X1 U10389 ( .A1(n9960), .A2(n9678), .ZN(n9523) );
  NAND2_X1 U10390 ( .A1(n9964), .A2(n9866), .ZN(n9455) );
  NAND2_X1 U10391 ( .A1(n9523), .A2(n9455), .ZN(n9355) );
  AOI21_X1 U10392 ( .B1(n9358), .B2(n9356), .A(n9355), .ZN(n9360) );
  AND2_X1 U10393 ( .A1(n9455), .A2(n9357), .ZN(n9522) );
  OR2_X1 U10394 ( .A1(n9960), .A2(n9678), .ZN(n9361) );
  NAND2_X1 U10395 ( .A1(n9361), .A2(n9398), .ZN(n9482) );
  AOI21_X1 U10396 ( .B1(n9358), .B2(n9522), .A(n9482), .ZN(n9359) );
  NAND2_X1 U10397 ( .A1(n9849), .A2(n9679), .ZN(n9694) );
  NAND2_X1 U10398 ( .A1(n9694), .A2(n9361), .ZN(n9363) );
  NAND2_X1 U10399 ( .A1(n9953), .A2(n9867), .ZN(n9829) );
  NAND2_X1 U10400 ( .A1(n9829), .A2(n9523), .ZN(n9362) );
  MUX2_X1 U10401 ( .A(n9363), .B(n9362), .S(n9383), .Z(n9366) );
  OAI21_X1 U10402 ( .B1(n9394), .B2(n9694), .A(n9451), .ZN(n9364) );
  INV_X1 U10403 ( .A(n9364), .ZN(n9365) );
  NAND2_X1 U10404 ( .A1(n9950), .A2(n9808), .ZN(n9426) );
  NAND2_X1 U10405 ( .A1(n9426), .A2(n9829), .ZN(n9693) );
  OAI21_X1 U10406 ( .B1(n9368), .B2(n9693), .A(n9367), .ZN(n9369) );
  NAND2_X1 U10407 ( .A1(n9943), .A2(n9834), .ZN(n9371) );
  AND2_X1 U10408 ( .A1(n9369), .A2(n9814), .ZN(n9375) );
  OR2_X1 U10409 ( .A1(n9939), .A2(n9809), .ZN(n9397) );
  NAND2_X1 U10410 ( .A1(n9397), .A2(n9370), .ZN(n9439) );
  NAND2_X1 U10411 ( .A1(n9939), .A2(n9809), .ZN(n9696) );
  AND2_X1 U10412 ( .A1(n9696), .A2(n9371), .ZN(n9445) );
  INV_X1 U10413 ( .A(n9445), .ZN(n9372) );
  MUX2_X1 U10414 ( .A(n9439), .B(n9372), .S(n9383), .Z(n9374) );
  MUX2_X1 U10415 ( .A(n9696), .B(n9397), .S(n9383), .Z(n9373) );
  NAND2_X1 U10416 ( .A1(n9922), .A2(n9763), .ZN(n9701) );
  AND2_X1 U10417 ( .A1(n9701), .A2(n9699), .ZN(n9449) );
  INV_X1 U10418 ( .A(n9449), .ZN(n9377) );
  INV_X1 U10419 ( .A(n9443), .ZN(n9376) );
  MUX2_X1 U10420 ( .A(n9377), .B(n9376), .S(n9383), .Z(n9378) );
  NAND2_X1 U10421 ( .A1(n9916), .A2(n9750), .ZN(n9462) );
  INV_X1 U10422 ( .A(n9740), .ZN(n9380) );
  OAI21_X1 U10423 ( .B1(n9394), .B2(n9701), .A(n9380), .ZN(n9382) );
  OR2_X1 U10424 ( .A1(n9910), .A2(n9741), .ZN(n9457) );
  NAND2_X1 U10425 ( .A1(n9910), .A2(n9741), .ZN(n9703) );
  NAND2_X1 U10426 ( .A1(n9457), .A2(n9703), .ZN(n9716) );
  INV_X1 U10427 ( .A(n9716), .ZN(n9725) );
  MUX2_X1 U10428 ( .A(n9462), .B(n9459), .S(n9383), .Z(n9381) );
  MUX2_X1 U10429 ( .A(n9457), .B(n9703), .S(n9383), .Z(n9384) );
  NAND3_X1 U10430 ( .A1(n9704), .A2(n9385), .A3(n9384), .ZN(n9386) );
  NAND4_X1 U10431 ( .A1(n9389), .A2(n9388), .A3(n9387), .A4(n9386), .ZN(n9390)
         );
  NAND3_X1 U10432 ( .A1(n9391), .A2(n9540), .A3(n9390), .ZN(n9393) );
  AND2_X1 U10433 ( .A1(n9897), .A2(n9392), .ZN(n9468) );
  MUX2_X1 U10434 ( .A(n9394), .B(n9393), .S(n9542), .Z(n9479) );
  AOI211_X1 U10435 ( .C1(n9472), .C2(n9778), .A(n9550), .B(n9395), .ZN(n9478)
         );
  INV_X1 U10436 ( .A(n9396), .ZN(n9438) );
  NAND2_X1 U10437 ( .A1(n9460), .A2(n9701), .ZN(n9748) );
  NAND2_X1 U10438 ( .A1(n9397), .A2(n9696), .ZN(n9791) );
  NAND2_X1 U10439 ( .A1(n9398), .A2(n9455), .ZN(n9882) );
  INV_X1 U10440 ( .A(n9882), .ZN(n9425) );
  NOR2_X1 U10441 ( .A1(n9399), .A2(n6236), .ZN(n9403) );
  NAND4_X1 U10442 ( .A1(n9403), .A2(n9402), .A3(n9401), .A4(n9400), .ZN(n9408)
         );
  XNOR2_X1 U10443 ( .A(n9574), .B(n9404), .ZN(n10457) );
  NAND3_X1 U10444 ( .A1(n9406), .A2(n10457), .A3(n9405), .ZN(n9407) );
  NOR2_X1 U10445 ( .A1(n9408), .A2(n9407), .ZN(n9410) );
  NAND4_X1 U10446 ( .A1(n9499), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n9413)
         );
  NOR2_X1 U10447 ( .A1(n9413), .A2(n9412), .ZN(n9414) );
  NAND3_X1 U10448 ( .A1(n9416), .A2(n9415), .A3(n9414), .ZN(n9417) );
  NOR2_X1 U10449 ( .A1(n9418), .A2(n9417), .ZN(n9419) );
  NAND4_X1 U10450 ( .A1(n5444), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n9422)
         );
  NOR2_X1 U10451 ( .A1(n9423), .A2(n9422), .ZN(n9424) );
  XNOR2_X1 U10452 ( .A(n9960), .B(n9888), .ZN(n9863) );
  NAND4_X1 U10453 ( .A1(n9850), .A2(n9425), .A3(n9424), .A4(n9863), .ZN(n9427)
         );
  NAND2_X1 U10454 ( .A1(n9451), .A2(n9426), .ZN(n9832) );
  NOR2_X1 U10455 ( .A1(n9427), .A2(n9832), .ZN(n9428) );
  NAND4_X1 U10456 ( .A1(n9781), .A2(n5325), .A3(n9814), .A4(n9428), .ZN(n9429)
         );
  NOR2_X1 U10457 ( .A1(n9764), .A2(n9429), .ZN(n9430) );
  NAND2_X1 U10458 ( .A1(n5316), .A2(n9430), .ZN(n9431) );
  OR2_X1 U10459 ( .A1(n9740), .A2(n9431), .ZN(n9432) );
  NOR2_X1 U10460 ( .A1(n9716), .A2(n9432), .ZN(n9433) );
  NAND2_X1 U10461 ( .A1(n9902), .A2(n9708), .ZN(n9532) );
  AND4_X1 U10462 ( .A1(n9704), .A2(n9538), .A3(n9433), .A4(n9532), .ZN(n9434)
         );
  NAND3_X1 U10463 ( .A1(n9540), .A2(n9434), .A3(n9542), .ZN(n9474) );
  OAI21_X1 U10464 ( .B1(n6236), .B2(n6030), .A(n9435), .ZN(n9436) );
  AOI21_X1 U10465 ( .B1(n9474), .B2(n9436), .A(n9544), .ZN(n9437) );
  AOI21_X1 U10466 ( .B1(n9479), .B2(n9438), .A(n9437), .ZN(n9477) );
  NAND2_X1 U10467 ( .A1(n9439), .A2(n9696), .ZN(n9440) );
  NAND2_X1 U10468 ( .A1(n9698), .A2(n9440), .ZN(n9441) );
  NAND2_X1 U10469 ( .A1(n9441), .A2(n9446), .ZN(n9442) );
  AND2_X1 U10470 ( .A1(n9443), .A2(n9442), .ZN(n9450) );
  NAND2_X1 U10471 ( .A1(n9693), .A2(n9451), .ZN(n9444) );
  NAND3_X1 U10472 ( .A1(n9446), .A2(n9445), .A3(n9444), .ZN(n9447) );
  NAND2_X1 U10473 ( .A1(n9450), .A2(n9447), .ZN(n9448) );
  AND2_X1 U10474 ( .A1(n9449), .A2(n9448), .ZN(n9480) );
  INV_X1 U10475 ( .A(n9450), .ZN(n9453) );
  NAND2_X1 U10476 ( .A1(n9451), .A2(n9694), .ZN(n9452) );
  NOR2_X1 U10477 ( .A1(n9453), .A2(n9452), .ZN(n9481) );
  INV_X1 U10478 ( .A(n9518), .ZN(n9883) );
  NOR2_X1 U10479 ( .A1(n9882), .A2(n9883), .ZN(n9454) );
  NAND2_X1 U10480 ( .A1(n9881), .A2(n9454), .ZN(n9885) );
  NAND2_X1 U10481 ( .A1(n9885), .A2(n9455), .ZN(n9864) );
  NAND2_X1 U10482 ( .A1(n9864), .A2(n9863), .ZN(n9456) );
  NAND2_X1 U10483 ( .A1(n9481), .A2(n9695), .ZN(n9461) );
  NAND2_X1 U10484 ( .A1(n9458), .A2(n9457), .ZN(n9464) );
  INV_X1 U10485 ( .A(n9459), .ZN(n9702) );
  OR3_X1 U10486 ( .A1(n9464), .A2(n9702), .A3(n5122), .ZN(n9537) );
  AOI21_X1 U10487 ( .B1(n9480), .B2(n9461), .A(n9537), .ZN(n9467) );
  INV_X1 U10488 ( .A(n9531), .ZN(n9465) );
  AND2_X1 U10489 ( .A1(n9703), .A2(n9462), .ZN(n9463) );
  NOR2_X1 U10490 ( .A1(n9464), .A2(n9463), .ZN(n9533) );
  NOR4_X1 U10491 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9533), .ZN(n9470)
         );
  NOR3_X1 U10492 ( .A1(n9470), .A2(n9469), .A3(n9468), .ZN(n9473) );
  OAI21_X1 U10493 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(n9475) );
  AOI21_X1 U10494 ( .B1(n9475), .B2(n9474), .A(n9778), .ZN(n9476) );
  AOI211_X1 U10495 ( .C1(n9479), .C2(n9478), .A(n9477), .B(n9476), .ZN(n9555)
         );
  INV_X1 U10496 ( .A(n9480), .ZN(n9530) );
  INV_X1 U10497 ( .A(n9481), .ZN(n9528) );
  INV_X1 U10498 ( .A(n9482), .ZN(n9526) );
  INV_X1 U10499 ( .A(n9483), .ZN(n9516) );
  NAND2_X1 U10500 ( .A1(n10445), .A2(n9574), .ZN(n9484) );
  OAI211_X1 U10501 ( .C1(n10446), .C2(n7234), .A(n9484), .B(n6236), .ZN(n9486)
         );
  NAND2_X1 U10502 ( .A1(n9486), .A2(n9485), .ZN(n9488) );
  OAI21_X1 U10503 ( .B1(n7242), .B2(n9488), .A(n9487), .ZN(n9490) );
  NAND2_X1 U10504 ( .A1(n9490), .A2(n9489), .ZN(n9492) );
  NAND2_X1 U10505 ( .A1(n9492), .A2(n9491), .ZN(n9495) );
  NAND3_X1 U10506 ( .A1(n9495), .A2(n9494), .A3(n9493), .ZN(n9498) );
  AOI21_X1 U10507 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9502) );
  INV_X1 U10508 ( .A(n9499), .ZN(n9501) );
  OAI21_X1 U10509 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9504) );
  NAND2_X1 U10510 ( .A1(n9504), .A2(n9503), .ZN(n9508) );
  INV_X1 U10511 ( .A(n9505), .ZN(n9507) );
  AOI21_X1 U10512 ( .B1(n9508), .B2(n9507), .A(n9506), .ZN(n9513) );
  INV_X1 U10513 ( .A(n9509), .ZN(n9512) );
  OAI211_X1 U10514 ( .C1(n9513), .C2(n9512), .A(n9511), .B(n9510), .ZN(n9515)
         );
  AOI21_X1 U10515 ( .B1(n9516), .B2(n9515), .A(n9514), .ZN(n9520) );
  OAI211_X1 U10516 ( .C1(n9520), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9521)
         );
  NAND2_X1 U10517 ( .A1(n9522), .A2(n9521), .ZN(n9525) );
  INV_X1 U10518 ( .A(n9523), .ZN(n9524) );
  AOI21_X1 U10519 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9527) );
  NOR2_X1 U10520 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  NOR2_X1 U10521 ( .A1(n9530), .A2(n9529), .ZN(n9536) );
  AND2_X1 U10522 ( .A1(n9532), .A2(n9531), .ZN(n9535) );
  INV_X1 U10523 ( .A(n9533), .ZN(n9534) );
  OAI211_X1 U10524 ( .C1(n9537), .C2(n9536), .A(n9535), .B(n9534), .ZN(n9539)
         );
  NAND2_X1 U10525 ( .A1(n9539), .A2(n9538), .ZN(n9541) );
  NAND2_X1 U10526 ( .A1(n9541), .A2(n9540), .ZN(n9543) );
  NAND2_X1 U10527 ( .A1(n9543), .A2(n9542), .ZN(n9548) );
  NAND2_X1 U10528 ( .A1(n9778), .A2(n9544), .ZN(n10455) );
  NAND2_X1 U10529 ( .A1(n9548), .A2(n9545), .ZN(n9547) );
  OAI211_X1 U10530 ( .C1(n9548), .C2(n10455), .A(n9547), .B(n9546), .ZN(n9554)
         );
  NOR3_X1 U10531 ( .A1(n9549), .A2(n10450), .A3(n10085), .ZN(n9553) );
  OAI21_X1 U10532 ( .B1(n9551), .B2(n9550), .A(P1_B_REG_SCAN_IN), .ZN(n9552)
         );
  OAI22_X1 U10533 ( .A1(n9555), .A2(n9554), .B1(n9553), .B2(n9552), .ZN(
        P1_U3242) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9556), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9557), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10536 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9727), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10537 ( .A(n9726), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9590), .Z(
        P1_U3581) );
  MUX2_X1 U10538 ( .A(n9684), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9590), .Z(
        P1_U3580) );
  MUX2_X1 U10539 ( .A(n9558), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9590), .Z(
        P1_U3579) );
  MUX2_X1 U10540 ( .A(n9681), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9590), .Z(
        P1_U3578) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9783), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9680), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9851), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10544 ( .A(n9679), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9590), .Z(
        P1_U3574) );
  MUX2_X1 U10545 ( .A(n9888), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9590), .Z(
        P1_U3573) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9890), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9559), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10548 ( .A(n9560), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9590), .Z(
        P1_U3569) );
  MUX2_X1 U10549 ( .A(n9561), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9590), .Z(
        P1_U3568) );
  MUX2_X1 U10550 ( .A(n9562), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9590), .Z(
        P1_U3567) );
  MUX2_X1 U10551 ( .A(n9563), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9590), .Z(
        P1_U3566) );
  MUX2_X1 U10552 ( .A(n9564), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9590), .Z(
        P1_U3565) );
  MUX2_X1 U10553 ( .A(n9565), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9590), .Z(
        P1_U3564) );
  MUX2_X1 U10554 ( .A(n9566), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9590), .Z(
        P1_U3563) );
  MUX2_X1 U10555 ( .A(n9567), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9590), .Z(
        P1_U3562) );
  MUX2_X1 U10556 ( .A(n9568), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9590), .Z(
        P1_U3561) );
  MUX2_X1 U10557 ( .A(n9569), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9590), .Z(
        P1_U3560) );
  MUX2_X1 U10558 ( .A(n9570), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9590), .Z(
        P1_U3559) );
  MUX2_X1 U10559 ( .A(n9571), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9590), .Z(
        P1_U3558) );
  MUX2_X1 U10560 ( .A(n9572), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9590), .Z(
        P1_U3557) );
  MUX2_X1 U10561 ( .A(n9573), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9590), .Z(
        P1_U3556) );
  MUX2_X1 U10562 ( .A(n9574), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9590), .Z(
        P1_U3554) );
  OAI211_X1 U10563 ( .C1(n9577), .C2(n9576), .A(n10427), .B(n9575), .ZN(n9585)
         );
  OAI211_X1 U10564 ( .C1(n9580), .C2(n9579), .A(n10431), .B(n9578), .ZN(n9584)
         );
  AOI22_X1 U10565 ( .A1(n10439), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9583) );
  NAND2_X1 U10566 ( .A1(n10229), .A2(n9581), .ZN(n9582) );
  NAND4_X1 U10567 ( .A1(n9585), .A2(n9584), .A3(n9583), .A4(n9582), .ZN(
        P1_U3244) );
  INV_X1 U10568 ( .A(n9586), .ZN(n9593) );
  OR2_X1 U10569 ( .A1(n4908), .A2(n9587), .ZN(n10086) );
  NAND2_X1 U10570 ( .A1(n9588), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9589) );
  XOR2_X1 U10571 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9589), .Z(n9591) );
  AOI21_X1 U10572 ( .B1(n9591), .B2(n10086), .A(n9590), .ZN(n9592) );
  OAI21_X1 U10573 ( .B1(n9593), .B2(n10086), .A(n9592), .ZN(n10441) );
  NAND2_X1 U10574 ( .A1(n10439), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U10575 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9594) );
  OAI211_X1 U10576 ( .C1(n10437), .C2(n9596), .A(n9595), .B(n9594), .ZN(n9597)
         );
  INV_X1 U10577 ( .A(n9597), .ZN(n9606) );
  OAI211_X1 U10578 ( .C1(n9600), .C2(n9599), .A(n10427), .B(n9598), .ZN(n9605)
         );
  OAI211_X1 U10579 ( .C1(n9603), .C2(n9602), .A(n10431), .B(n9601), .ZN(n9604)
         );
  NAND4_X1 U10580 ( .A1(n10441), .A2(n9606), .A3(n9605), .A4(n9604), .ZN(
        P1_U3245) );
  INV_X1 U10581 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9608) );
  OAI21_X1 U10582 ( .B1(n10264), .B2(n9608), .A(n9607), .ZN(n9609) );
  AOI21_X1 U10583 ( .B1(n9610), .B2(n10229), .A(n9609), .ZN(n9619) );
  OAI211_X1 U10584 ( .C1(n9613), .C2(n9612), .A(n10431), .B(n9611), .ZN(n9618)
         );
  OAI211_X1 U10585 ( .C1(n9616), .C2(n9615), .A(n10427), .B(n9614), .ZN(n9617)
         );
  NAND3_X1 U10586 ( .A1(n9619), .A2(n9618), .A3(n9617), .ZN(P1_U3246) );
  INV_X1 U10587 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10631) );
  NOR2_X1 U10588 ( .A1(n10228), .A2(n10631), .ZN(n9620) );
  AOI21_X1 U10589 ( .B1(n10228), .B2(n10631), .A(n9620), .ZN(n10220) );
  OAI21_X1 U10590 ( .B1(n9634), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9621), .ZN(
        n10221) );
  NOR2_X1 U10591 ( .A1(n10220), .A2(n10221), .ZN(n10219) );
  AOI21_X1 U10592 ( .B1(n10228), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10219), 
        .ZN(n10172) );
  INV_X1 U10593 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U10594 ( .A1(n9637), .A2(n9622), .ZN(n9624) );
  NAND2_X1 U10595 ( .A1(n10177), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9623) );
  AND2_X1 U10596 ( .A1(n9624), .A2(n9623), .ZN(n10173) );
  NOR2_X1 U10597 ( .A1(n10172), .A2(n10173), .ZN(n10171) );
  AOI21_X1 U10598 ( .B1(n9637), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10171), .ZN(
        n9625) );
  NOR2_X1 U10599 ( .A1(n9625), .A2(n9639), .ZN(n9626) );
  INV_X1 U10600 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10183) );
  XNOR2_X1 U10601 ( .A(n9639), .B(n9625), .ZN(n10184) );
  NOR2_X1 U10602 ( .A1(n10183), .A2(n10184), .ZN(n10182) );
  NOR2_X1 U10603 ( .A1(n9626), .A2(n10182), .ZN(n9629) );
  INV_X1 U10604 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9627) );
  AOI22_X1 U10605 ( .A1(n9656), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9627), .B2(
        n9632), .ZN(n9628) );
  NAND2_X1 U10606 ( .A1(n9628), .A2(n9629), .ZN(n9655) );
  OAI21_X1 U10607 ( .B1(n9629), .B2(n9628), .A(n9655), .ZN(n9646) );
  AOI21_X1 U10608 ( .B1(n10439), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9630), .ZN(
        n9631) );
  OAI21_X1 U10609 ( .B1(n9632), .B2(n10437), .A(n9631), .ZN(n9645) );
  OAI21_X1 U10610 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9634), .A(n9633), .ZN(
        n10225) );
  NAND2_X1 U10611 ( .A1(n10228), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9635) );
  OAI21_X1 U10612 ( .B1(n10228), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9635), .ZN(
        n10224) );
  NOR2_X1 U10613 ( .A1(n10225), .A2(n10224), .ZN(n10223) );
  AOI21_X1 U10614 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10228), .A(n10223), 
        .ZN(n10168) );
  NAND2_X1 U10615 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9637), .ZN(n9636) );
  OAI21_X1 U10616 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9637), .A(n9636), .ZN(
        n10169) );
  NOR2_X1 U10617 ( .A1(n10168), .A2(n10169), .ZN(n10167) );
  AOI21_X1 U10618 ( .B1(n9637), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10167), .ZN(
        n9638) );
  NOR2_X1 U10619 ( .A1(n9638), .A2(n9639), .ZN(n9640) );
  INV_X1 U10620 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10186) );
  XNOR2_X1 U10621 ( .A(n9639), .B(n9638), .ZN(n10187) );
  NOR2_X1 U10622 ( .A1(n10186), .A2(n10187), .ZN(n10185) );
  NOR2_X1 U10623 ( .A1(n9640), .A2(n10185), .ZN(n9643) );
  NAND2_X1 U10624 ( .A1(n9656), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9641) );
  OAI21_X1 U10625 ( .B1(n9656), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9641), .ZN(
        n9642) );
  NOR2_X1 U10626 ( .A1(n9643), .A2(n9642), .ZN(n9649) );
  AOI211_X1 U10627 ( .C1(n9643), .C2(n9642), .A(n9649), .B(n10222), .ZN(n9644)
         );
  AOI211_X1 U10628 ( .C1(n10431), .C2(n9646), .A(n9645), .B(n9644), .ZN(n9647)
         );
  INV_X1 U10629 ( .A(n9647), .ZN(P1_U3259) );
  NAND2_X1 U10630 ( .A1(n10214), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9650) );
  OAI21_X1 U10631 ( .B1(n10214), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9650), .ZN(
        n10210) );
  NOR2_X1 U10632 ( .A1(n10201), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9648) );
  AOI21_X1 U10633 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10201), .A(n9648), .ZN(
        n10195) );
  AOI21_X1 U10634 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9656), .A(n9649), .ZN(
        n10196) );
  NAND2_X1 U10635 ( .A1(n10195), .A2(n10196), .ZN(n10194) );
  OAI21_X1 U10636 ( .B1(n10201), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10194), 
        .ZN(n10211) );
  NOR2_X1 U10637 ( .A1(n10210), .A2(n10211), .ZN(n10209) );
  INV_X1 U10638 ( .A(n10209), .ZN(n9651) );
  NAND2_X1 U10639 ( .A1(n9651), .A2(n9650), .ZN(n9654) );
  INV_X1 U10640 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9652) );
  MUX2_X1 U10641 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9652), .S(n6030), .Z(n9653) );
  XNOR2_X1 U10642 ( .A(n9654), .B(n9653), .ZN(n9662) );
  XOR2_X1 U10643 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10201), .Z(n10198) );
  OAI21_X1 U10644 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9656), .A(n9655), .ZN(
        n10199) );
  NAND2_X1 U10645 ( .A1(n10198), .A2(n10199), .ZN(n10197) );
  OAI21_X1 U10646 ( .B1(n10201), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10197), 
        .ZN(n10207) );
  NAND2_X1 U10647 ( .A1(n10214), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9657) );
  OAI21_X1 U10648 ( .B1(n10214), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9657), .ZN(
        n10208) );
  NOR2_X1 U10649 ( .A1(n10207), .A2(n10208), .ZN(n10206) );
  INV_X1 U10650 ( .A(n9657), .ZN(n9658) );
  NOR2_X1 U10651 ( .A1(n10206), .A2(n9658), .ZN(n9660) );
  XNOR2_X1 U10652 ( .A(n6030), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9659) );
  XNOR2_X1 U10653 ( .A(n9660), .B(n9659), .ZN(n9661) );
  AOI22_X1 U10654 ( .A1(n10427), .A2(n9662), .B1(n10431), .B2(n9661), .ZN(
        n9666) );
  INV_X1 U10655 ( .A(n9663), .ZN(n9664) );
  AOI21_X1 U10656 ( .B1(n10439), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9664), .ZN(
        n9665) );
  OAI211_X1 U10657 ( .C1(n6030), .C2(n10437), .A(n9666), .B(n9665), .ZN(
        P1_U3262) );
  NAND2_X1 U10658 ( .A1(n9667), .A2(n9687), .ZN(n9668) );
  XNOR2_X1 U10659 ( .A(n9897), .B(n9668), .ZN(n9899) );
  NOR2_X1 U10660 ( .A1(n9669), .A2(n9879), .ZN(n9670) );
  AOI211_X1 U10661 ( .C1(n10562), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9671), .B(
        n9670), .ZN(n9672) );
  OAI21_X1 U10662 ( .B1(n9899), .B2(n9673), .A(n9672), .ZN(P1_U3263) );
  NAND2_X1 U10663 ( .A1(n9872), .A2(n9882), .ZN(n9871) );
  OAI21_X1 U10664 ( .B1(n9939), .B2(n9783), .A(n9790), .ZN(n9774) );
  NAND2_X1 U10665 ( .A1(n9934), .A2(n9681), .ZN(n9683) );
  NAND2_X1 U10666 ( .A1(n9765), .A2(n9764), .ZN(n9925) );
  OAI21_X1 U10667 ( .B1(n9786), .B2(n5164), .A(n9925), .ZN(n9747) );
  NAND2_X1 U10668 ( .A1(n9757), .A2(n9763), .ZN(n9685) );
  XNOR2_X1 U10669 ( .A(n9686), .B(n9704), .ZN(n9905) );
  INV_X1 U10670 ( .A(n9905), .ZN(n9715) );
  AOI211_X1 U10671 ( .C1(n9907), .C2(n9717), .A(n10512), .B(n9687), .ZN(n9906)
         );
  INV_X1 U10672 ( .A(n9907), .ZN(n9691) );
  NAND3_X1 U10673 ( .A1(n9688), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n10551), 
        .ZN(n9690) );
  NAND2_X1 U10674 ( .A1(n10562), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9689) );
  OAI211_X1 U10675 ( .C1(n9691), .C2(n9879), .A(n9690), .B(n9689), .ZN(n9692)
         );
  AOI21_X1 U10676 ( .B1(n9906), .B2(n10556), .A(n9692), .ZN(n9714) );
  INV_X1 U10677 ( .A(n9814), .ZN(n9806) );
  INV_X1 U10678 ( .A(n9696), .ZN(n9697) );
  NAND2_X1 U10679 ( .A1(n9782), .A2(n9781), .ZN(n9780) );
  INV_X1 U10680 ( .A(n9699), .ZN(n9700) );
  NOR2_X1 U10681 ( .A1(n9739), .A2(n9740), .ZN(n9738) );
  NOR2_X1 U10682 ( .A1(n9738), .A2(n9702), .ZN(n9724) );
  NAND2_X1 U10683 ( .A1(n9724), .A2(n9725), .ZN(n9723) );
  NAND2_X1 U10684 ( .A1(n9723), .A2(n9703), .ZN(n9705) );
  XNOR2_X1 U10685 ( .A(n9705), .B(n9704), .ZN(n9706) );
  NAND2_X1 U10686 ( .A1(n9706), .A2(n9892), .ZN(n9712) );
  NOR2_X1 U10687 ( .A1(n9708), .A2(n9707), .ZN(n9709) );
  OAI211_X1 U10688 ( .C1(n9715), .C2(n9896), .A(n9714), .B(n9713), .ZN(
        P1_U3356) );
  INV_X1 U10689 ( .A(n9733), .ZN(n9719) );
  INV_X1 U10690 ( .A(n9717), .ZN(n9718) );
  AOI21_X1 U10691 ( .B1(n9910), .B2(n9719), .A(n9718), .ZN(n9911) );
  AOI22_X1 U10692 ( .A1(n9720), .A2(n10551), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10562), .ZN(n9721) );
  OAI21_X1 U10693 ( .B1(n9722), .B2(n9879), .A(n9721), .ZN(n9730) );
  OAI21_X1 U10694 ( .B1(n9725), .B2(n9724), .A(n9723), .ZN(n9728) );
  AOI222_X1 U10695 ( .A1(n9892), .A2(n9728), .B1(n9727), .B2(n9887), .C1(n9726), .C2(n9889), .ZN(n9913) );
  NOR2_X1 U10696 ( .A1(n9913), .A2(n10562), .ZN(n9729) );
  AOI211_X1 U10697 ( .C1(n9911), .C2(n9855), .A(n9730), .B(n9729), .ZN(n9731)
         );
  OAI21_X1 U10698 ( .B1(n9914), .B2(n9896), .A(n9731), .ZN(P1_U3265) );
  XOR2_X1 U10699 ( .A(n9740), .B(n9732), .Z(n9919) );
  AOI211_X1 U10700 ( .C1(n9916), .C2(n9751), .A(n10512), .B(n9733), .ZN(n9915)
         );
  INV_X1 U10701 ( .A(n9734), .ZN(n9735) );
  AOI22_X1 U10702 ( .A1(n9735), .A2(n10551), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10562), .ZN(n9736) );
  OAI21_X1 U10703 ( .B1(n9737), .B2(n9879), .A(n9736), .ZN(n9745) );
  AOI211_X1 U10704 ( .C1(n9740), .C2(n9739), .A(n10539), .B(n9738), .ZN(n9743)
         );
  OAI22_X1 U10705 ( .A1(n9741), .A2(n10531), .B1(n9763), .B2(n10533), .ZN(
        n9742) );
  NOR2_X1 U10706 ( .A1(n9743), .A2(n9742), .ZN(n9918) );
  NOR2_X1 U10707 ( .A1(n9918), .A2(n10562), .ZN(n9744) );
  AOI211_X1 U10708 ( .C1(n10556), .C2(n9915), .A(n9745), .B(n9744), .ZN(n9746)
         );
  OAI21_X1 U10709 ( .B1(n9919), .B2(n9896), .A(n9746), .ZN(P1_U3266) );
  XNOR2_X1 U10710 ( .A(n9747), .B(n9748), .ZN(n9924) );
  XOR2_X1 U10711 ( .A(n9748), .B(n4924), .Z(n9749) );
  OAI222_X1 U10712 ( .A1(n10531), .A2(n9750), .B1(n10533), .B2(n9786), .C1(
        n9749), .C2(n10539), .ZN(n9920) );
  INV_X1 U10713 ( .A(n9766), .ZN(n9753) );
  INV_X1 U10714 ( .A(n9751), .ZN(n9752) );
  AOI211_X1 U10715 ( .C1(n9922), .C2(n9753), .A(n10512), .B(n9752), .ZN(n9921)
         );
  NAND2_X1 U10716 ( .A1(n9921), .A2(n10556), .ZN(n9756) );
  AOI22_X1 U10717 ( .A1(n9754), .A2(n10551), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10562), .ZN(n9755) );
  OAI211_X1 U10718 ( .C1(n9757), .C2(n9879), .A(n9756), .B(n9755), .ZN(n9758)
         );
  AOI21_X1 U10719 ( .B1(n9920), .B2(n9868), .A(n9758), .ZN(n9759) );
  OAI21_X1 U10720 ( .B1(n9924), .B2(n9896), .A(n9759), .ZN(P1_U3267) );
  AOI21_X1 U10721 ( .B1(n9764), .B2(n9761), .A(n9760), .ZN(n9762) );
  OAI222_X1 U10722 ( .A1(n10533), .A2(n9798), .B1(n10531), .B2(n9763), .C1(
        n10539), .C2(n9762), .ZN(n9927) );
  INV_X1 U10723 ( .A(n9927), .ZN(n9773) );
  OR2_X1 U10724 ( .A1(n9765), .A2(n9764), .ZN(n9926) );
  NAND3_X1 U10725 ( .A1(n9926), .A2(n9925), .A3(n9815), .ZN(n9772) );
  AOI211_X1 U10726 ( .C1(n9929), .C2(n9775), .A(n10512), .B(n9766), .ZN(n9928)
         );
  NOR2_X1 U10727 ( .A1(n5164), .A2(n9879), .ZN(n9770) );
  OAI22_X1 U10728 ( .A1(n9768), .A2(n10448), .B1(n9767), .B2(n9868), .ZN(n9769) );
  AOI211_X1 U10729 ( .C1(n9928), .C2(n10556), .A(n9770), .B(n9769), .ZN(n9771)
         );
  OAI211_X1 U10730 ( .C1(n10562), .C2(n9773), .A(n9772), .B(n9771), .ZN(
        P1_U3268) );
  XNOR2_X1 U10731 ( .A(n9774), .B(n9781), .ZN(n9936) );
  AOI22_X1 U10732 ( .A1(n9934), .A2(n10552), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10562), .ZN(n9789) );
  INV_X1 U10733 ( .A(n9775), .ZN(n9776) );
  AOI211_X1 U10734 ( .C1(n9934), .C2(n5169), .A(n10512), .B(n9776), .ZN(n9933)
         );
  INV_X1 U10735 ( .A(n9933), .ZN(n9779) );
  OAI22_X1 U10736 ( .A1(n9779), .A2(n9778), .B1(n10448), .B2(n9777), .ZN(n9787) );
  OAI211_X1 U10737 ( .C1(n9782), .C2(n9781), .A(n9780), .B(n9892), .ZN(n9785)
         );
  NAND2_X1 U10738 ( .A1(n9783), .A2(n9889), .ZN(n9784) );
  OAI211_X1 U10739 ( .C1(n9786), .C2(n10531), .A(n9785), .B(n9784), .ZN(n9932)
         );
  OAI21_X1 U10740 ( .B1(n9787), .B2(n9932), .A(n9868), .ZN(n9788) );
  OAI211_X1 U10741 ( .C1(n9936), .C2(n9896), .A(n9789), .B(n9788), .ZN(
        P1_U3269) );
  OAI21_X1 U10742 ( .B1(n9792), .B2(n9791), .A(n9790), .ZN(n9793) );
  INV_X1 U10743 ( .A(n9793), .ZN(n9941) );
  INV_X1 U10744 ( .A(n9805), .ZN(n9794) );
  AOI21_X1 U10745 ( .B1(n9794), .B2(n9370), .A(n5325), .ZN(n9795) );
  NOR2_X1 U10746 ( .A1(n9796), .A2(n9795), .ZN(n9797) );
  OAI222_X1 U10747 ( .A1(n10533), .A2(n9834), .B1(n10531), .B2(n9798), .C1(
        n10539), .C2(n9797), .ZN(n9937) );
  AOI211_X1 U10748 ( .C1(n9939), .C2(n9816), .A(n10512), .B(n9799), .ZN(n9938)
         );
  NAND2_X1 U10749 ( .A1(n9938), .A2(n10556), .ZN(n9802) );
  AOI22_X1 U10750 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n10562), .B1(n9800), 
        .B2(n10551), .ZN(n9801) );
  OAI211_X1 U10751 ( .C1(n5168), .C2(n9879), .A(n9802), .B(n9801), .ZN(n9803)
         );
  AOI21_X1 U10752 ( .B1(n9937), .B2(n9868), .A(n9803), .ZN(n9804) );
  OAI21_X1 U10753 ( .B1(n9941), .B2(n9896), .A(n9804), .ZN(P1_U3270) );
  AOI211_X1 U10754 ( .C1(n9807), .C2(n9806), .A(n10539), .B(n9805), .ZN(n9811)
         );
  OAI22_X1 U10755 ( .A1(n9809), .A2(n10531), .B1(n9808), .B2(n10533), .ZN(
        n9810) );
  NOR2_X1 U10756 ( .A1(n9811), .A2(n9810), .ZN(n9946) );
  AOI21_X1 U10757 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9942) );
  NAND2_X1 U10758 ( .A1(n9942), .A2(n9815), .ZN(n9825) );
  INV_X1 U10759 ( .A(n9835), .ZN(n9818) );
  INV_X1 U10760 ( .A(n9816), .ZN(n9817) );
  AOI21_X1 U10761 ( .B1(n9943), .B2(n9818), .A(n9817), .ZN(n9944) );
  NOR2_X1 U10762 ( .A1(n9819), .A2(n9879), .ZN(n9823) );
  OAI22_X1 U10763 ( .A1(n9868), .A2(n9821), .B1(n9820), .B2(n10448), .ZN(n9822) );
  AOI211_X1 U10764 ( .C1(n9944), .C2(n9855), .A(n9823), .B(n9822), .ZN(n9824)
         );
  OAI211_X1 U10765 ( .C1(n10562), .C2(n9946), .A(n9825), .B(n9824), .ZN(
        P1_U3271) );
  OAI21_X1 U10766 ( .B1(n9827), .B2(n9832), .A(n9826), .ZN(n9828) );
  INV_X1 U10767 ( .A(n9828), .ZN(n9952) );
  INV_X1 U10768 ( .A(n9829), .ZN(n9830) );
  AOI21_X1 U10769 ( .B1(n9695), .B2(n9850), .A(n9830), .ZN(n9831) );
  XOR2_X1 U10770 ( .A(n9832), .B(n9831), .Z(n9833) );
  OAI222_X1 U10771 ( .A1(n10531), .A2(n9834), .B1(n10533), .B2(n9867), .C1(
        n9833), .C2(n10539), .ZN(n9948) );
  AOI211_X1 U10772 ( .C1(n9950), .C2(n9843), .A(n10512), .B(n9835), .ZN(n9949)
         );
  NAND2_X1 U10773 ( .A1(n9949), .A2(n10556), .ZN(n9838) );
  AOI22_X1 U10774 ( .A1(n10562), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9836), 
        .B2(n10551), .ZN(n9837) );
  OAI211_X1 U10775 ( .C1(n9839), .C2(n9879), .A(n9838), .B(n9837), .ZN(n9840)
         );
  AOI21_X1 U10776 ( .B1(n9868), .B2(n9948), .A(n9840), .ZN(n9841) );
  OAI21_X1 U10777 ( .B1(n9952), .B2(n9896), .A(n9841), .ZN(P1_U3272) );
  XOR2_X1 U10778 ( .A(n9842), .B(n9850), .Z(n9957) );
  INV_X1 U10779 ( .A(n9858), .ZN(n9845) );
  INV_X1 U10780 ( .A(n9843), .ZN(n9844) );
  AOI21_X1 U10781 ( .B1(n9953), .B2(n9845), .A(n9844), .ZN(n9954) );
  INV_X1 U10782 ( .A(n9846), .ZN(n9847) );
  AOI22_X1 U10783 ( .A1(n10562), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9847), 
        .B2(n10551), .ZN(n9848) );
  OAI21_X1 U10784 ( .B1(n9849), .B2(n9879), .A(n9848), .ZN(n9854) );
  XNOR2_X1 U10785 ( .A(n9695), .B(n9850), .ZN(n9852) );
  AOI222_X1 U10786 ( .A1(n9892), .A2(n9852), .B1(n9851), .B2(n9887), .C1(n9888), .C2(n9889), .ZN(n9956) );
  NOR2_X1 U10787 ( .A1(n9956), .A2(n10562), .ZN(n9853) );
  AOI211_X1 U10788 ( .C1(n9954), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9856)
         );
  OAI21_X1 U10789 ( .B1(n9957), .B2(n9896), .A(n9856), .ZN(P1_U3273) );
  XOR2_X1 U10790 ( .A(n9857), .B(n9863), .Z(n9962) );
  AOI211_X1 U10791 ( .C1(n9960), .C2(n9874), .A(n10512), .B(n9858), .ZN(n9959)
         );
  NOR2_X1 U10792 ( .A1(n9859), .A2(n9879), .ZN(n9862) );
  OAI22_X1 U10793 ( .A1(n9868), .A2(n9652), .B1(n9860), .B2(n10448), .ZN(n9861) );
  AOI211_X1 U10794 ( .C1(n9959), .C2(n10556), .A(n9862), .B(n9861), .ZN(n9870)
         );
  XOR2_X1 U10795 ( .A(n9864), .B(n9863), .Z(n9865) );
  OAI222_X1 U10796 ( .A1(n10531), .A2(n9867), .B1(n10533), .B2(n9866), .C1(
        n10539), .C2(n9865), .ZN(n9958) );
  NAND2_X1 U10797 ( .A1(n9958), .A2(n9868), .ZN(n9869) );
  OAI211_X1 U10798 ( .C1(n9962), .C2(n9896), .A(n9870), .B(n9869), .ZN(
        P1_U3274) );
  OAI21_X1 U10799 ( .B1(n9872), .B2(n9882), .A(n9871), .ZN(n9967) );
  INV_X1 U10800 ( .A(n9873), .ZN(n9876) );
  INV_X1 U10801 ( .A(n9874), .ZN(n9875) );
  AOI211_X1 U10802 ( .C1(n9964), .C2(n9876), .A(n10512), .B(n9875), .ZN(n9963)
         );
  AOI22_X1 U10803 ( .A1(n10562), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9877), 
        .B2(n10551), .ZN(n9878) );
  OAI21_X1 U10804 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(n9894) );
  INV_X1 U10805 ( .A(n9881), .ZN(n9884) );
  OAI21_X1 U10806 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9886) );
  NAND2_X1 U10807 ( .A1(n9886), .A2(n9885), .ZN(n9891) );
  AOI222_X1 U10808 ( .A1(n9892), .A2(n9891), .B1(n9890), .B2(n9889), .C1(n9888), .C2(n9887), .ZN(n9966) );
  NOR2_X1 U10809 ( .A1(n9966), .A2(n10562), .ZN(n9893) );
  AOI211_X1 U10810 ( .C1(n9963), .C2(n10556), .A(n9894), .B(n9893), .ZN(n9895)
         );
  OAI21_X1 U10811 ( .B1(n9967), .B2(n9896), .A(n9895), .ZN(P1_U3275) );
  AOI21_X1 U10812 ( .B1(n9897), .B2(n10490), .A(n9901), .ZN(n9898) );
  OAI21_X1 U10813 ( .B1(n9899), .B2(n10512), .A(n9898), .ZN(n9991) );
  MUX2_X1 U10814 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9991), .S(n10632), .Z(
        P1_U3553) );
  INV_X1 U10815 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9903) );
  MUX2_X1 U10816 ( .A(n9903), .B(n9992), .S(n10632), .Z(n9904) );
  INV_X1 U10817 ( .A(n9904), .ZN(P1_U3552) );
  NAND2_X1 U10818 ( .A1(n9905), .A2(n10628), .ZN(n9909) );
  NAND2_X1 U10819 ( .A1(n9909), .A2(n9908), .ZN(n9994) );
  MUX2_X1 U10820 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9994), .S(n10632), .Z(
        P1_U3551) );
  AOI22_X1 U10821 ( .A1(n9911), .A2(n10527), .B1(n10490), .B2(n9910), .ZN(
        n9912) );
  OAI211_X1 U10822 ( .C1(n9914), .C2(n10494), .A(n9913), .B(n9912), .ZN(n9995)
         );
  MUX2_X1 U10823 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9995), .S(n10632), .Z(
        P1_U3550) );
  AOI21_X1 U10824 ( .B1(n10490), .B2(n9916), .A(n9915), .ZN(n9917) );
  OAI211_X1 U10825 ( .C1(n9919), .C2(n10494), .A(n9918), .B(n9917), .ZN(n9996)
         );
  MUX2_X1 U10826 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9996), .S(n10632), .Z(
        P1_U3549) );
  AOI211_X1 U10827 ( .C1(n10490), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9923)
         );
  OAI21_X1 U10828 ( .B1(n9924), .B2(n10494), .A(n9923), .ZN(n9997) );
  MUX2_X1 U10829 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9997), .S(n10632), .Z(
        P1_U3548) );
  NAND3_X1 U10830 ( .A1(n9926), .A2(n9925), .A3(n10628), .ZN(n9931) );
  AOI211_X1 U10831 ( .C1(n10490), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9930)
         );
  NAND2_X1 U10832 ( .A1(n9931), .A2(n9930), .ZN(n9998) );
  MUX2_X1 U10833 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9998), .S(n10632), .Z(
        P1_U3547) );
  AOI211_X1 U10834 ( .C1(n10490), .C2(n9934), .A(n9933), .B(n9932), .ZN(n9935)
         );
  OAI21_X1 U10835 ( .B1(n9936), .B2(n10494), .A(n9935), .ZN(n9999) );
  MUX2_X1 U10836 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9999), .S(n10632), .Z(
        P1_U3546) );
  AOI211_X1 U10837 ( .C1(n10490), .C2(n9939), .A(n9938), .B(n9937), .ZN(n9940)
         );
  OAI21_X1 U10838 ( .B1(n9941), .B2(n10494), .A(n9940), .ZN(n10000) );
  MUX2_X1 U10839 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10000), .S(n10632), .Z(
        P1_U3545) );
  INV_X1 U10840 ( .A(n9942), .ZN(n9947) );
  AOI22_X1 U10841 ( .A1(n9944), .A2(n10527), .B1(n10490), .B2(n9943), .ZN(
        n9945) );
  OAI211_X1 U10842 ( .C1(n9947), .C2(n10494), .A(n9946), .B(n9945), .ZN(n10001) );
  MUX2_X1 U10843 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10001), .S(n10632), .Z(
        P1_U3544) );
  AOI211_X1 U10844 ( .C1(n10490), .C2(n9950), .A(n9949), .B(n9948), .ZN(n9951)
         );
  OAI21_X1 U10845 ( .B1(n9952), .B2(n10494), .A(n9951), .ZN(n10002) );
  MUX2_X1 U10846 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10002), .S(n10632), .Z(
        P1_U3543) );
  AOI22_X1 U10847 ( .A1(n9954), .A2(n10527), .B1(n10490), .B2(n9953), .ZN(
        n9955) );
  OAI211_X1 U10848 ( .C1(n9957), .C2(n10494), .A(n9956), .B(n9955), .ZN(n10003) );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10003), .S(n10632), .Z(
        P1_U3542) );
  AOI211_X1 U10850 ( .C1(n10490), .C2(n9960), .A(n9959), .B(n9958), .ZN(n9961)
         );
  OAI21_X1 U10851 ( .B1(n9962), .B2(n10494), .A(n9961), .ZN(n10004) );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10004), .S(n10632), .Z(
        P1_U3541) );
  AOI21_X1 U10853 ( .B1(n10490), .B2(n9964), .A(n9963), .ZN(n9965) );
  OAI211_X1 U10854 ( .C1(n9967), .C2(n10494), .A(n9966), .B(n9965), .ZN(n10005) );
  MUX2_X1 U10855 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10005), .S(n10632), .Z(
        P1_U3540) );
  AOI211_X1 U10856 ( .C1(n10490), .C2(n9970), .A(n9969), .B(n9968), .ZN(n9971)
         );
  OAI21_X1 U10857 ( .B1(n9972), .B2(n10494), .A(n9971), .ZN(n10006) );
  MUX2_X1 U10858 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10006), .S(n10632), .Z(
        P1_U3539) );
  NAND3_X1 U10859 ( .A1(n9974), .A2(n9973), .A3(n10628), .ZN(n9979) );
  NAND2_X1 U10860 ( .A1(n9975), .A2(n10490), .ZN(n9976) );
  NAND4_X1 U10861 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n10007) );
  MUX2_X1 U10862 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10007), .S(n10632), .Z(
        P1_U3538) );
  AOI22_X1 U10863 ( .A1(n9981), .A2(n10527), .B1(n10490), .B2(n9980), .ZN(
        n9982) );
  OAI211_X1 U10864 ( .C1(n9984), .C2(n10494), .A(n9983), .B(n9982), .ZN(n10008) );
  MUX2_X1 U10865 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10008), .S(n10632), .Z(
        P1_U3537) );
  AOI21_X1 U10866 ( .B1(n10490), .B2(n9986), .A(n9985), .ZN(n9987) );
  OAI211_X1 U10867 ( .C1(n9990), .C2(n9989), .A(n9988), .B(n9987), .ZN(n10009)
         );
  MUX2_X1 U10868 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10009), .S(n10632), .Z(
        P1_U3536) );
  MUX2_X1 U10869 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9991), .S(n10636), .Z(
        P1_U3521) );
  INV_X1 U10870 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9993) );
  MUX2_X1 U10871 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9994), .S(n10636), .Z(
        P1_U3519) );
  MUX2_X1 U10872 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9995), .S(n10636), .Z(
        P1_U3518) );
  MUX2_X1 U10873 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9996), .S(n10636), .Z(
        P1_U3517) );
  MUX2_X1 U10874 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9997), .S(n10636), .Z(
        P1_U3516) );
  MUX2_X1 U10875 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9998), .S(n10636), .Z(
        P1_U3515) );
  MUX2_X1 U10876 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9999), .S(n10636), .Z(
        P1_U3514) );
  MUX2_X1 U10877 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10000), .S(n10636), .Z(
        P1_U3513) );
  MUX2_X1 U10878 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10001), .S(n10636), .Z(
        P1_U3512) );
  MUX2_X1 U10879 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10002), .S(n10636), .Z(
        P1_U3511) );
  MUX2_X1 U10880 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10003), .S(n10636), .Z(
        P1_U3510) );
  MUX2_X1 U10881 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10004), .S(n10636), .Z(
        P1_U3509) );
  MUX2_X1 U10882 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10005), .S(n10636), .Z(
        P1_U3507) );
  MUX2_X1 U10883 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10006), .S(n10636), .Z(
        P1_U3504) );
  MUX2_X1 U10884 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10007), .S(n10636), .Z(
        P1_U3501) );
  MUX2_X1 U10885 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10008), .S(n10636), .Z(
        P1_U3498) );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10009), .S(n10636), .Z(
        P1_U3495) );
  MUX2_X1 U10887 ( .A(n10010), .B(P1_D_REG_1__SCAN_IN), .S(n10027), .Z(
        P1_U3440) );
  NAND3_X1 U10888 ( .A1(n10011), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10013) );
  OAI22_X1 U10889 ( .A1(n5636), .A2(n10013), .B1(n10012), .B2(n10018), .ZN(
        n10014) );
  AOI21_X1 U10890 ( .B1(n10016), .B2(n10015), .A(n10014), .ZN(n10017) );
  INV_X1 U10891 ( .A(n10017), .ZN(P1_U3324) );
  OAI222_X1 U10892 ( .A1(P1_U3086), .A2(n10021), .B1(n8202), .B2(n10020), .C1(
        n10019), .C2(n10018), .ZN(P1_U3325) );
  OAI222_X1 U10893 ( .A1(n10025), .A2(n10024), .B1(n8202), .B2(n10023), .C1(
        n10022), .C2(P1_U3086), .ZN(P1_U3326) );
  MUX2_X1 U10894 ( .A(n10026), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U10895 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10027), .ZN(P1_U3323) );
  AND2_X1 U10896 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10027), .ZN(P1_U3322) );
  AND2_X1 U10897 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10027), .ZN(P1_U3321) );
  AND2_X1 U10898 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10027), .ZN(P1_U3320) );
  AND2_X1 U10899 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10027), .ZN(P1_U3319) );
  AND2_X1 U10900 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10027), .ZN(P1_U3318) );
  AND2_X1 U10901 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10027), .ZN(P1_U3317) );
  AND2_X1 U10902 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10027), .ZN(P1_U3316) );
  AND2_X1 U10903 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10027), .ZN(P1_U3315) );
  AND2_X1 U10904 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10027), .ZN(P1_U3314) );
  AND2_X1 U10905 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10027), .ZN(P1_U3313) );
  AND2_X1 U10906 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10027), .ZN(P1_U3312) );
  AND2_X1 U10907 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10027), .ZN(P1_U3311) );
  AND2_X1 U10908 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10027), .ZN(P1_U3310) );
  AND2_X1 U10909 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10027), .ZN(P1_U3309) );
  AND2_X1 U10910 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10027), .ZN(P1_U3308) );
  AND2_X1 U10911 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10027), .ZN(P1_U3307) );
  AND2_X1 U10912 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10027), .ZN(P1_U3306) );
  AND2_X1 U10913 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10027), .ZN(P1_U3305) );
  AND2_X1 U10914 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10027), .ZN(P1_U3304) );
  AND2_X1 U10915 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10027), .ZN(P1_U3303) );
  AND2_X1 U10916 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10027), .ZN(P1_U3302) );
  AND2_X1 U10917 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10027), .ZN(P1_U3301) );
  AND2_X1 U10918 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10027), .ZN(P1_U3300) );
  AND2_X1 U10919 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10027), .ZN(P1_U3299) );
  AND2_X1 U10920 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10027), .ZN(P1_U3298) );
  AND2_X1 U10921 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10027), .ZN(P1_U3297) );
  AND2_X1 U10922 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10027), .ZN(P1_U3296) );
  AND2_X1 U10923 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10027), .ZN(P1_U3295) );
  AND2_X1 U10924 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10027), .ZN(P1_U3294) );
  OAI21_X1 U10925 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10030), .ZN(n10028) );
  INV_X1 U10926 ( .A(n10028), .ZN(ADD_1068_U46) );
  OAI21_X1 U10927 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10032) );
  XNOR2_X1 U10928 ( .A(n10032), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  AOI21_X1 U10929 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(ADD_1068_U54) );
  AOI21_X1 U10930 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(ADD_1068_U53) );
  OAI21_X1 U10931 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(ADD_1068_U52) );
  OAI21_X1 U10932 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(ADD_1068_U51) );
  OAI21_X1 U10933 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(ADD_1068_U50) );
  OAI21_X1 U10934 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(ADD_1068_U49) );
  OAI21_X1 U10935 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(ADD_1068_U48) );
  OAI21_X1 U10936 ( .B1(n10056), .B2(n10055), .A(n10054), .ZN(ADD_1068_U47) );
  OAI21_X1 U10937 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(ADD_1068_U63) );
  OAI21_X1 U10938 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(ADD_1068_U62) );
  OAI21_X1 U10939 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(ADD_1068_U61) );
  OAI21_X1 U10940 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(ADD_1068_U60) );
  OAI21_X1 U10941 ( .B1(n10071), .B2(n10070), .A(n10069), .ZN(ADD_1068_U59) );
  OAI21_X1 U10942 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(ADD_1068_U58) );
  OAI21_X1 U10943 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(ADD_1068_U57) );
  OAI21_X1 U10944 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(ADD_1068_U56) );
  OAI21_X1 U10945 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(ADD_1068_U55) );
  INV_X1 U10946 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10084) );
  OAI22_X1 U10947 ( .A1(n5681), .A2(n10086), .B1(n10085), .B2(n10084), .ZN(
        n10087) );
  XNOR2_X1 U10948 ( .A(n10087), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U10949 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10439), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10088) );
  OAI21_X1 U10950 ( .B1(n10090), .B2(n10089), .A(n10088), .ZN(P1_U3243) );
  INV_X1 U10951 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10105) );
  AOI21_X1 U10952 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10094) );
  NAND2_X1 U10953 ( .A1(n10427), .A2(n10094), .ZN(n10100) );
  AOI21_X1 U10954 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10098) );
  NAND2_X1 U10955 ( .A1(n10431), .A2(n10098), .ZN(n10099) );
  OAI211_X1 U10956 ( .C1(n10437), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10102) );
  INV_X1 U10957 ( .A(n10102), .ZN(n10104) );
  OAI211_X1 U10958 ( .C1(n10264), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        P1_U3248) );
  INV_X1 U10959 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10120) );
  AOI21_X1 U10960 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(n10109) );
  NAND2_X1 U10961 ( .A1(n10427), .A2(n10109), .ZN(n10115) );
  AOI21_X1 U10962 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(n10113) );
  NAND2_X1 U10963 ( .A1(n10431), .A2(n10113), .ZN(n10114) );
  OAI211_X1 U10964 ( .C1(n10437), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        n10117) );
  INV_X1 U10965 ( .A(n10117), .ZN(n10119) );
  OAI211_X1 U10966 ( .C1(n10264), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        P1_U3249) );
  INV_X1 U10967 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10135) );
  AOI21_X1 U10968 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(n10124) );
  NAND2_X1 U10969 ( .A1(n10427), .A2(n10124), .ZN(n10130) );
  AOI21_X1 U10970 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(n10128) );
  NAND2_X1 U10971 ( .A1(n10431), .A2(n10128), .ZN(n10129) );
  OAI211_X1 U10972 ( .C1(n10437), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        n10132) );
  INV_X1 U10973 ( .A(n10132), .ZN(n10134) );
  OAI211_X1 U10974 ( .C1(n10264), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        P1_U3250) );
  INV_X1 U10975 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10150) );
  AOI21_X1 U10976 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(n10139) );
  NAND2_X1 U10977 ( .A1(n10427), .A2(n10139), .ZN(n10145) );
  AOI21_X1 U10978 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(n10143) );
  NAND2_X1 U10979 ( .A1(n10431), .A2(n10143), .ZN(n10144) );
  OAI211_X1 U10980 ( .C1(n10437), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        n10147) );
  INV_X1 U10981 ( .A(n10147), .ZN(n10149) );
  OAI211_X1 U10982 ( .C1(n10264), .C2(n10150), .A(n10149), .B(n10148), .ZN(
        P1_U3251) );
  INV_X1 U10983 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10166) );
  INV_X1 U10984 ( .A(n10151), .ZN(n10162) );
  AOI21_X1 U10985 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10155) );
  NAND2_X1 U10986 ( .A1(n10427), .A2(n10155), .ZN(n10161) );
  AOI21_X1 U10987 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10159) );
  NAND2_X1 U10988 ( .A1(n10431), .A2(n10159), .ZN(n10160) );
  OAI211_X1 U10989 ( .C1(n10437), .C2(n10162), .A(n10161), .B(n10160), .ZN(
        n10163) );
  INV_X1 U10990 ( .A(n10163), .ZN(n10165) );
  OAI211_X1 U10991 ( .C1(n10264), .C2(n10166), .A(n10165), .B(n10164), .ZN(
        P1_U3254) );
  INV_X1 U10992 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10181) );
  AOI21_X1 U10993 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(n10170) );
  NAND2_X1 U10994 ( .A1(n10427), .A2(n10170), .ZN(n10176) );
  AOI21_X1 U10995 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(n10174) );
  NAND2_X1 U10996 ( .A1(n10431), .A2(n10174), .ZN(n10175) );
  OAI211_X1 U10997 ( .C1(n10437), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10178) );
  INV_X1 U10998 ( .A(n10178), .ZN(n10180) );
  OAI211_X1 U10999 ( .C1(n10264), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        P1_U3257) );
  INV_X1 U11000 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10193) );
  AOI211_X1 U11001 ( .C1(n10184), .C2(n10183), .A(n10182), .B(n10218), .ZN(
        n10189) );
  AOI211_X1 U11002 ( .C1(n10187), .C2(n10186), .A(n10185), .B(n10222), .ZN(
        n10188) );
  AOI211_X1 U11003 ( .C1(n10229), .C2(n10190), .A(n10189), .B(n10188), .ZN(
        n10192) );
  OAI211_X1 U11004 ( .C1(n10264), .C2(n10193), .A(n10192), .B(n10191), .ZN(
        P1_U3258) );
  INV_X1 U11005 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10205) );
  OAI21_X1 U11006 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10202) );
  OAI21_X1 U11007 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(n10200) );
  AOI222_X1 U11008 ( .A1(n10202), .A2(n10427), .B1(n10201), .B2(n10229), .C1(
        n10200), .C2(n10431), .ZN(n10204) );
  OAI211_X1 U11009 ( .C1(n10264), .C2(n10205), .A(n10204), .B(n10203), .ZN(
        P1_U3260) );
  INV_X1 U11010 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10217) );
  AOI211_X1 U11011 ( .C1(n10208), .C2(n10207), .A(n10206), .B(n10218), .ZN(
        n10213) );
  AOI211_X1 U11012 ( .C1(n10211), .C2(n10210), .A(n10209), .B(n10222), .ZN(
        n10212) );
  AOI211_X1 U11013 ( .C1(n10229), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        n10216) );
  OAI211_X1 U11014 ( .C1(n10264), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        P1_U3261) );
  INV_X1 U11015 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10233) );
  AOI211_X1 U11016 ( .C1(n10221), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10227) );
  AOI211_X1 U11017 ( .C1(n10225), .C2(n10224), .A(n10223), .B(n10222), .ZN(
        n10226) );
  AOI211_X1 U11018 ( .C1(n10229), .C2(n10228), .A(n10227), .B(n10226), .ZN(
        n10232) );
  INV_X1 U11019 ( .A(n10230), .ZN(n10231) );
  OAI211_X1 U11020 ( .C1(n10264), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        P1_U3256) );
  INV_X1 U11021 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10248) );
  AOI21_X1 U11022 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(n10237) );
  NAND2_X1 U11023 ( .A1(n10427), .A2(n10237), .ZN(n10243) );
  AOI21_X1 U11024 ( .B1(n10240), .B2(n10239), .A(n10238), .ZN(n10241) );
  NAND2_X1 U11025 ( .A1(n10431), .A2(n10241), .ZN(n10242) );
  OAI211_X1 U11026 ( .C1(n10437), .C2(n10244), .A(n10243), .B(n10242), .ZN(
        n10245) );
  INV_X1 U11027 ( .A(n10245), .ZN(n10247) );
  OAI211_X1 U11028 ( .C1(n10264), .C2(n10248), .A(n10247), .B(n10246), .ZN(
        P1_U3253) );
  INV_X1 U11029 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10263) );
  OAI21_X1 U11030 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(n10252) );
  NAND2_X1 U11031 ( .A1(n10427), .A2(n10252), .ZN(n10258) );
  OAI21_X1 U11032 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(n10256) );
  NAND2_X1 U11033 ( .A1(n10431), .A2(n10256), .ZN(n10257) );
  OAI211_X1 U11034 ( .C1(n10437), .C2(n10259), .A(n10258), .B(n10257), .ZN(
        n10260) );
  INV_X1 U11035 ( .A(n10260), .ZN(n10262) );
  OAI211_X1 U11036 ( .C1(n10264), .C2(n10263), .A(n10262), .B(n10261), .ZN(
        P1_U3252) );
  INV_X1 U11037 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10289) );
  OAI21_X1 U11038 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(n10280) );
  INV_X1 U11039 ( .A(n10268), .ZN(n10269) );
  OAI21_X1 U11040 ( .B1(n10271), .B2(n10270), .A(n10269), .ZN(n10279) );
  INV_X1 U11041 ( .A(n10272), .ZN(n10274) );
  NAND3_X1 U11042 ( .A1(n10275), .A2(n10274), .A3(n10273), .ZN(n10276) );
  AOI21_X1 U11043 ( .B1(n10277), .B2(n10276), .A(n10418), .ZN(n10278) );
  AOI211_X1 U11044 ( .C1(n10413), .C2(n10280), .A(n10279), .B(n10278), .ZN(
        n10287) );
  AOI211_X1 U11045 ( .C1(n10284), .C2(n10283), .A(n10282), .B(n10281), .ZN(
        n10285) );
  INV_X1 U11046 ( .A(n10285), .ZN(n10286) );
  OAI211_X1 U11047 ( .C1(n10289), .C2(n10288), .A(n10287), .B(n10286), .ZN(
        P2_U3186) );
  AOI22_X1 U11048 ( .A1(n10290), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n10308) );
  INV_X1 U11049 ( .A(n10291), .ZN(n10293) );
  NAND2_X1 U11050 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  XNOR2_X1 U11051 ( .A(n10295), .B(n10294), .ZN(n10300) );
  OAI21_X1 U11052 ( .B1(n10298), .B2(n10297), .A(n10296), .ZN(n10299) );
  AOI22_X1 U11053 ( .A1(n10300), .A2(n10412), .B1(n10413), .B2(n10299), .ZN(
        n10307) );
  NAND2_X1 U11054 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3151), .ZN(n10306)
         );
  AOI21_X1 U11055 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(n10304) );
  OR2_X1 U11056 ( .A1(n10304), .A2(n10418), .ZN(n10305) );
  NAND4_X1 U11057 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        P2_U3192) );
  AOI22_X1 U11058 ( .A1(n10309), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n10323) );
  OAI21_X1 U11059 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(n10316) );
  OAI21_X1 U11060 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n10314), .A(n10313), 
        .ZN(n10315) );
  AOI22_X1 U11061 ( .A1(n10316), .A2(n10412), .B1(n10413), .B2(n10315), .ZN(
        n10322) );
  AOI21_X1 U11062 ( .B1(n10318), .B2(n6502), .A(n10317), .ZN(n10319) );
  OR2_X1 U11063 ( .A1(n10418), .A2(n10319), .ZN(n10320) );
  NAND4_X1 U11064 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        P2_U3193) );
  AOI22_X1 U11065 ( .A1(n10324), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n10340) );
  OAI21_X1 U11066 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10332) );
  OAI21_X1 U11067 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(n10331) );
  AOI22_X1 U11068 ( .A1(n10332), .A2(n10413), .B1(n10412), .B2(n10331), .ZN(
        n10339) );
  AOI21_X1 U11069 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(n10336) );
  OR2_X1 U11070 ( .A1(n10336), .A2(n10418), .ZN(n10337) );
  NAND4_X1 U11071 ( .A1(n10340), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        P2_U3194) );
  AOI22_X1 U11072 ( .A1(n10341), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10355) );
  OAI21_X1 U11073 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10343), .A(n10342), 
        .ZN(n10348) );
  OAI21_X1 U11074 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(n10347) );
  AOI22_X1 U11075 ( .A1(n10348), .A2(n10413), .B1(n10412), .B2(n10347), .ZN(
        n10354) );
  AOI21_X1 U11076 ( .B1(n10350), .B2(n6529), .A(n10349), .ZN(n10351) );
  OR2_X1 U11077 ( .A1(n10418), .A2(n10351), .ZN(n10352) );
  NAND4_X1 U11078 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        P2_U3195) );
  AOI22_X1 U11079 ( .A1(n10356), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10371) );
  OAI21_X1 U11080 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(n10364) );
  OAI21_X1 U11081 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n10363) );
  AOI22_X1 U11082 ( .A1(n10364), .A2(n10413), .B1(n10412), .B2(n10363), .ZN(
        n10370) );
  AOI21_X1 U11083 ( .B1(n4970), .B2(n10366), .A(n10365), .ZN(n10367) );
  OR2_X1 U11084 ( .A1(n10367), .A2(n10418), .ZN(n10368) );
  NAND4_X1 U11085 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        P2_U3196) );
  AOI22_X1 U11086 ( .A1(n10372), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n10386) );
  OAI21_X1 U11087 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10374), .A(n10373), 
        .ZN(n10379) );
  OAI21_X1 U11088 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(n10378) );
  AOI22_X1 U11089 ( .A1(n10379), .A2(n10413), .B1(n10412), .B2(n10378), .ZN(
        n10385) );
  AOI21_X1 U11090 ( .B1(n10381), .B2(n7968), .A(n10380), .ZN(n10382) );
  OR2_X1 U11091 ( .A1(n10418), .A2(n10382), .ZN(n10383) );
  NAND4_X1 U11092 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        P2_U3197) );
  AOI22_X1 U11093 ( .A1(n10387), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10402) );
  OAI21_X1 U11094 ( .B1(n10390), .B2(n10389), .A(n10388), .ZN(n10395) );
  OAI21_X1 U11095 ( .B1(n10393), .B2(n10392), .A(n10391), .ZN(n10394) );
  AOI22_X1 U11096 ( .A1(n10395), .A2(n10413), .B1(n10412), .B2(n10394), .ZN(
        n10401) );
  AOI21_X1 U11097 ( .B1(n4943), .B2(n10397), .A(n10396), .ZN(n10398) );
  OR2_X1 U11098 ( .A1(n10398), .A2(n10418), .ZN(n10399) );
  NAND4_X1 U11099 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        P2_U3198) );
  AOI22_X1 U11100 ( .A1(n10405), .A2(n10404), .B1(n10403), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10423) );
  OAI21_X1 U11101 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10407), .A(n10406), 
        .ZN(n10414) );
  OAI21_X1 U11102 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(n10411) );
  AOI22_X1 U11103 ( .A1(n10414), .A2(n10413), .B1(n10412), .B2(n10411), .ZN(
        n10422) );
  AOI21_X1 U11104 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10419) );
  OR2_X1 U11105 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  NAND4_X1 U11106 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        P2_U3199) );
  XOR2_X1 U11107 ( .A(P1_RD_REG_SCAN_IN), .B(n10424), .Z(U126) );
  INV_X1 U11108 ( .A(n10425), .ZN(n10426) );
  OAI211_X1 U11109 ( .C1(n10429), .C2(n10428), .A(n10427), .B(n10426), .ZN(
        n10435) );
  OAI211_X1 U11110 ( .C1(n10433), .C2(n10432), .A(n10431), .B(n10430), .ZN(
        n10434) );
  OAI211_X1 U11111 ( .C1(n10437), .C2(n10436), .A(n10435), .B(n10434), .ZN(
        n10438) );
  INV_X1 U11112 ( .A(n10438), .ZN(n10443) );
  NAND2_X1 U11113 ( .A1(n10439), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10440) );
  NAND4_X1 U11114 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        P1_U3247) );
  NOR2_X1 U11115 ( .A1(n10445), .A2(n10444), .ZN(n10459) );
  INV_X1 U11116 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10449) );
  NOR2_X1 U11117 ( .A1(n10446), .A2(n10531), .ZN(n10458) );
  INV_X1 U11118 ( .A(n10458), .ZN(n10447) );
  OAI21_X1 U11119 ( .B1(n10449), .B2(n10448), .A(n10447), .ZN(n10454) );
  INV_X1 U11120 ( .A(n10450), .ZN(n10452) );
  NOR3_X1 U11121 ( .A1(n10457), .A2(n10452), .A3(n10451), .ZN(n10453) );
  AOI211_X1 U11122 ( .C1(n10459), .C2(n10455), .A(n10454), .B(n10453), .ZN(
        n10456) );
  AOI22_X1 U11123 ( .A1(n10562), .A2(n10084), .B1(n10456), .B2(n9868), .ZN(
        P1_U3293) );
  AOI21_X1 U11124 ( .B1(n10539), .B2(n10494), .A(n10457), .ZN(n10460) );
  NOR3_X1 U11125 ( .A1(n10460), .A2(n10459), .A3(n10458), .ZN(n10462) );
  AOI22_X1 U11126 ( .A1(n10632), .A2(n10462), .B1(n5681), .B2(n10630), .ZN(
        P1_U3522) );
  INV_X1 U11127 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U11128 ( .A1(n10636), .A2(n10462), .B1(n10461), .B2(n10633), .ZN(
        P1_U3453) );
  AOI22_X1 U11129 ( .A1(n10640), .A2(n10463), .B1(n6359), .B2(n10637), .ZN(
        P2_U3393) );
  INV_X1 U11130 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U11131 ( .A1(n10636), .A2(n10465), .B1(n10464), .B2(n10633), .ZN(
        P1_U3456) );
  AOI22_X1 U11132 ( .A1(n10640), .A2(n10466), .B1(n6377), .B2(n10637), .ZN(
        P2_U3396) );
  OAI22_X1 U11133 ( .A1(n10470), .A2(n10469), .B1(n10468), .B2(n10467), .ZN(
        n10472) );
  AOI211_X1 U11134 ( .C1(n10474), .C2(n10473), .A(n10472), .B(n10471), .ZN(
        n10475) );
  AOI22_X1 U11135 ( .A1(n10577), .A2(n10476), .B1(n10475), .B2(n10575), .ZN(
        P2_U3231) );
  OAI21_X1 U11136 ( .B1(n10478), .B2(n10625), .A(n10477), .ZN(n10480) );
  AOI211_X1 U11137 ( .C1(n10609), .C2(n10481), .A(n10480), .B(n10479), .ZN(
        n10484) );
  INV_X1 U11138 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U11139 ( .A1(n10632), .A2(n10484), .B1(n10482), .B2(n10630), .ZN(
        P1_U3525) );
  INV_X1 U11140 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U11141 ( .A1(n10636), .A2(n10484), .B1(n10483), .B2(n10633), .ZN(
        P1_U3462) );
  AOI22_X1 U11142 ( .A1(n10640), .A2(n10485), .B1(n6391), .B2(n10637), .ZN(
        P2_U3399) );
  INV_X1 U11143 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U11144 ( .A1(n10640), .A2(n10487), .B1(n10486), .B2(n10637), .ZN(
        P2_U3402) );
  AOI21_X1 U11145 ( .B1(n10490), .B2(n10489), .A(n10488), .ZN(n10492) );
  OAI211_X1 U11146 ( .C1(n10494), .C2(n10493), .A(n10492), .B(n10491), .ZN(
        n10495) );
  INV_X1 U11147 ( .A(n10495), .ZN(n10498) );
  AOI22_X1 U11148 ( .A1(n10632), .A2(n10498), .B1(n10496), .B2(n10630), .ZN(
        P1_U3526) );
  INV_X1 U11149 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U11150 ( .A1(n10636), .A2(n10498), .B1(n10497), .B2(n10633), .ZN(
        P1_U3465) );
  INV_X1 U11151 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U11152 ( .A1(n10640), .A2(n10500), .B1(n10499), .B2(n10637), .ZN(
        P2_U3405) );
  OAI211_X1 U11153 ( .C1(n10503), .C2(n10625), .A(n10502), .B(n10501), .ZN(
        n10504) );
  AOI21_X1 U11154 ( .B1(n10628), .B2(n10505), .A(n10504), .ZN(n10508) );
  INV_X1 U11155 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U11156 ( .A1(n10632), .A2(n10508), .B1(n10506), .B2(n10630), .ZN(
        P1_U3527) );
  INV_X1 U11157 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U11158 ( .A1(n10636), .A2(n10508), .B1(n10507), .B2(n10633), .ZN(
        P1_U3468) );
  INV_X1 U11159 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U11160 ( .A1(n10640), .A2(n10510), .B1(n10509), .B2(n10637), .ZN(
        P2_U3408) );
  OAI22_X1 U11161 ( .A1(n10513), .A2(n10512), .B1(n10511), .B2(n10625), .ZN(
        n10514) );
  AOI21_X1 U11162 ( .B1(n10515), .B2(n10609), .A(n10514), .ZN(n10516) );
  INV_X1 U11163 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U11164 ( .A1(n10632), .A2(n10520), .B1(n10518), .B2(n10630), .ZN(
        P1_U3528) );
  INV_X1 U11165 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U11166 ( .A1(n10636), .A2(n10520), .B1(n10519), .B2(n10633), .ZN(
        P1_U3471) );
  NAND2_X1 U11167 ( .A1(n10521), .A2(n10522), .ZN(n10524) );
  NAND2_X1 U11168 ( .A1(n10524), .A2(n10523), .ZN(n10525) );
  XNOR2_X1 U11169 ( .A(n10525), .B(n10536), .ZN(n10558) );
  INV_X1 U11170 ( .A(n10526), .ZN(n10528) );
  OAI211_X1 U11171 ( .C1(n10530), .C2(n10529), .A(n10528), .B(n10527), .ZN(
        n10554) );
  OAI21_X1 U11172 ( .B1(n10530), .B2(n10625), .A(n10554), .ZN(n10546) );
  OAI22_X1 U11173 ( .A1(n10534), .A2(n10533), .B1(n10532), .B2(n10531), .ZN(
        n10543) );
  INV_X1 U11174 ( .A(n10535), .ZN(n10538) );
  OAI21_X1 U11175 ( .B1(n10538), .B2(n10537), .A(n10536), .ZN(n10541) );
  AOI21_X1 U11176 ( .B1(n10541), .B2(n10540), .A(n10539), .ZN(n10542) );
  AOI211_X1 U11177 ( .C1(n10544), .C2(n10558), .A(n10543), .B(n10542), .ZN(
        n10561) );
  INV_X1 U11178 ( .A(n10561), .ZN(n10545) );
  AOI211_X1 U11179 ( .C1(n10609), .C2(n10558), .A(n10546), .B(n10545), .ZN(
        n10549) );
  INV_X1 U11180 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U11181 ( .A1(n10632), .A2(n10549), .B1(n10547), .B2(n10630), .ZN(
        P1_U3529) );
  INV_X1 U11182 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U11183 ( .A1(n10636), .A2(n10549), .B1(n10548), .B2(n10633), .ZN(
        P1_U3474) );
  AOI222_X1 U11184 ( .A1(n10553), .A2(n10552), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n10562), .C1(n10551), .C2(n10550), .ZN(n10560) );
  INV_X1 U11185 ( .A(n10554), .ZN(n10555) );
  AOI22_X1 U11186 ( .A1(n10558), .A2(n10557), .B1(n10556), .B2(n10555), .ZN(
        n10559) );
  OAI211_X1 U11187 ( .C1(n10562), .C2(n10561), .A(n10560), .B(n10559), .ZN(
        P1_U3286) );
  AOI22_X1 U11188 ( .A1(n10640), .A2(n10563), .B1(n6441), .B2(n10637), .ZN(
        P2_U3411) );
  AOI21_X1 U11189 ( .B1(n10565), .B2(n10571), .A(n10564), .ZN(n10576) );
  INV_X1 U11190 ( .A(n10566), .ZN(n10573) );
  INV_X1 U11191 ( .A(n10567), .ZN(n10570) );
  AOI222_X1 U11192 ( .A1(n10573), .A2(n10572), .B1(n10571), .B2(n10570), .C1(
        n10569), .C2(n10568), .ZN(n10574) );
  OAI221_X1 U11193 ( .B1(n10577), .B2(n10576), .C1(n10575), .C2(n5374), .A(
        n10574), .ZN(P2_U3226) );
  OAI21_X1 U11194 ( .B1(n10579), .B2(n10625), .A(n10578), .ZN(n10580) );
  AOI21_X1 U11195 ( .B1(n10581), .B2(n10609), .A(n10580), .ZN(n10582) );
  AND2_X1 U11196 ( .A1(n10583), .A2(n10582), .ZN(n10585) );
  AOI22_X1 U11197 ( .A1(n10632), .A2(n10585), .B1(n7360), .B2(n10630), .ZN(
        P1_U3530) );
  INV_X1 U11198 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U11199 ( .A1(n10636), .A2(n10585), .B1(n10584), .B2(n10633), .ZN(
        P1_U3477) );
  INV_X1 U11200 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U11201 ( .A1(n10640), .A2(n10587), .B1(n10586), .B2(n10637), .ZN(
        P2_U3414) );
  OAI211_X1 U11202 ( .C1(n10590), .C2(n10625), .A(n10589), .B(n10588), .ZN(
        n10591) );
  AOI21_X1 U11203 ( .B1(n10628), .B2(n10592), .A(n10591), .ZN(n10594) );
  AOI22_X1 U11204 ( .A1(n10632), .A2(n10594), .B1(n7343), .B2(n10630), .ZN(
        P1_U3531) );
  INV_X1 U11205 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U11206 ( .A1(n10636), .A2(n10594), .B1(n10593), .B2(n10633), .ZN(
        P1_U3480) );
  INV_X1 U11207 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U11208 ( .A1(n10640), .A2(n10596), .B1(n10595), .B2(n10637), .ZN(
        P2_U3417) );
  OAI211_X1 U11209 ( .C1(n5154), .C2(n10625), .A(n10598), .B(n10597), .ZN(
        n10599) );
  AOI21_X1 U11210 ( .B1(n10628), .B2(n10600), .A(n10599), .ZN(n10602) );
  AOI22_X1 U11211 ( .A1(n10632), .A2(n10602), .B1(n7342), .B2(n10630), .ZN(
        P1_U3532) );
  INV_X1 U11212 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U11213 ( .A1(n10636), .A2(n10602), .B1(n10601), .B2(n10633), .ZN(
        P1_U3483) );
  AOI22_X1 U11214 ( .A1(n10640), .A2(n10603), .B1(n6488), .B2(n10637), .ZN(
        P2_U3420) );
  INV_X1 U11215 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U11216 ( .A1(n10640), .A2(n10605), .B1(n10604), .B2(n10637), .ZN(
        P2_U3423) );
  OAI21_X1 U11217 ( .B1(n10607), .B2(n10625), .A(n10606), .ZN(n10608) );
  AOI21_X1 U11218 ( .B1(n10610), .B2(n10609), .A(n10608), .ZN(n10611) );
  AND2_X1 U11219 ( .A1(n10612), .A2(n10611), .ZN(n10614) );
  AOI22_X1 U11220 ( .A1(n10632), .A2(n10614), .B1(n7364), .B2(n10630), .ZN(
        P1_U3533) );
  INV_X1 U11221 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U11222 ( .A1(n10636), .A2(n10614), .B1(n10613), .B2(n10633), .ZN(
        P1_U3486) );
  OAI211_X1 U11223 ( .C1(n10617), .C2(n10625), .A(n10616), .B(n10615), .ZN(
        n10618) );
  AOI21_X1 U11224 ( .B1(n10619), .B2(n10628), .A(n10618), .ZN(n10622) );
  AOI22_X1 U11225 ( .A1(n10632), .A2(n10622), .B1(n10620), .B2(n10630), .ZN(
        P1_U3534) );
  INV_X1 U11226 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U11227 ( .A1(n10636), .A2(n10622), .B1(n10621), .B2(n10633), .ZN(
        P1_U3489) );
  OAI211_X1 U11228 ( .C1(n10626), .C2(n10625), .A(n10624), .B(n10623), .ZN(
        n10627) );
  AOI21_X1 U11229 ( .B1(n10629), .B2(n10628), .A(n10627), .ZN(n10635) );
  AOI22_X1 U11230 ( .A1(n10632), .A2(n10635), .B1(n10631), .B2(n10630), .ZN(
        P1_U3535) );
  INV_X1 U11231 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U11232 ( .A1(n10636), .A2(n10635), .B1(n10634), .B2(n10633), .ZN(
        P1_U3492) );
  INV_X1 U11233 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U11234 ( .A1(n10640), .A2(n10639), .B1(n10638), .B2(n10637), .ZN(
        P2_U3429) );
  OAI22_X1 U11235 ( .A1(n10644), .A2(n10643), .B1(n10642), .B2(n10641), .ZN(
        n10645) );
  AOI21_X1 U11236 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(P2_U3151), .A(n10645), 
        .ZN(n10652) );
  XNOR2_X1 U11237 ( .A(n10648), .B(n10647), .ZN(n10650) );
  AOI22_X1 U11238 ( .A1(n10650), .A2(n10665), .B1(n10667), .B2(n10649), .ZN(
        n10651) );
  OAI211_X1 U11239 ( .C1(n10654), .C2(n10653), .A(n10652), .B(n10651), .ZN(
        P2_U3178) );
  INV_X1 U11240 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U11241 ( .A1(n10657), .A2(n6594), .B1(n10656), .B2(n10655), .ZN(
        n10672) );
  INV_X1 U11242 ( .A(n10658), .ZN(n10669) );
  INV_X1 U11243 ( .A(n10660), .ZN(n10662) );
  NAND2_X1 U11244 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  XNOR2_X1 U11245 ( .A(n10664), .B(n10663), .ZN(n10666) );
  AOI222_X1 U11246 ( .A1(n10670), .A2(n10669), .B1(n10668), .B2(n10667), .C1(
        n10666), .C2(n10665), .ZN(n10671) );
  OAI211_X1 U11247 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10673), .A(n10672), .B(
        n10671), .ZN(P2_U3173) );
  XNOR2_X1 U11248 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U4981 ( .A(n5708), .Z(n9169) );
  INV_X1 U4991 ( .A(n5708), .ZN(n6183) );
  CLKBUF_X1 U5555 ( .A(n5683), .Z(n9176) );
  CLKBUF_X1 U6677 ( .A(n8268), .Z(n8269) );
  CLKBUF_X1 U9533 ( .A(n6245), .Z(n4908) );
endmodule

