

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175;

  OR2_X1 U34680 ( .A1(n5135), .A2(n3438), .ZN(n3446) );
  CLKBUF_X2 U34690 ( .A(n3829), .Z(n3437) );
  CLKBUF_X2 U34700 ( .A(n3659), .Z(n4374) );
  AND2_X2 U34710 ( .A1(n5115), .A2(n5086), .ZN(n3712) );
  AND4_X1 U34720 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3690)
         );
  AND2_X2 U34730 ( .A1(n5828), .A2(n5086), .ZN(n3706) );
  NAND4_X2 U34740 ( .A1(n3625), .A2(n3622), .A3(n3623), .A4(n3624), .ZN(n3692)
         );
  NAND4_X1 U3475 ( .A1(n3691), .A2(n3688), .A3(n3689), .A4(n3690), .ZN(n4836)
         );
  AND2_X1 U3476 ( .A1(n3828), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4519) );
  NAND2_X1 U3477 ( .A1(n5370), .A2(n5000), .ZN(n4743) );
  NAND2_X1 U3478 ( .A1(n3975), .A2(n3974), .ZN(n4444) );
  INV_X2 U3479 ( .A(n5338), .ZN(n4872) );
  OR2_X1 U3480 ( .A1(n3621), .A2(n3620), .ZN(n4402) );
  AND2_X1 U3481 ( .A1(n3730), .A2(n3849), .ZN(n3555) );
  NOR2_X2 U3482 ( .A1(n3468), .A2(n5454), .ZN(n5444) );
  AND2_X1 U3483 ( .A1(n3847), .A2(n3849), .ZN(n3480) );
  INV_X2 U3484 ( .A(n5629), .ZN(n5704) );
  INV_X1 U3485 ( .A(n3849), .ZN(n3722) );
  INV_X1 U3486 ( .A(n6188), .ZN(n6211) );
  INV_X1 U3487 ( .A(n6526), .ZN(n6510) );
  OR2_X1 U3488 ( .A1(n4562), .A2(n4546), .ZN(n3435) );
  AND2_X4 U3489 ( .A1(n5828), .A2(n3581), .ZN(n3711) );
  AND2_X4 U3490 ( .A1(n3567), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5828)
         );
  NOR2_X4 U3491 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5115) );
  XNOR2_X2 U3492 ( .A(n3814), .B(n3815), .ZN(n3853) );
  NAND2_X2 U3493 ( .A1(n3779), .A2(n3778), .ZN(n3814) );
  OAI21_X1 U3494 ( .B1(n5704), .B2(n3565), .A(n4563), .ZN(n4565) );
  AOI211_X1 U3495 ( .C1(n5409), .C2(n6206), .A(n5332), .B(n5331), .ZN(n5333)
         );
  NAND2_X1 U3496 ( .A1(n5444), .A2(n3521), .ZN(n5329) );
  NAND2_X1 U3497 ( .A1(n5293), .A2(n4076), .ZN(n5299) );
  NAND2_X1 U3498 ( .A1(n3973), .A2(n3972), .ZN(n4961) );
  INV_X2 U3499 ( .A(n5629), .ZN(n5689) );
  NAND2_X1 U3500 ( .A1(n4444), .A2(n4394), .ZN(n4466) );
  CLKBUF_X1 U3501 ( .A(n4941), .Z(n3458) );
  NAND2_X1 U3502 ( .A1(n6162), .A2(n5561), .ZN(n5558) );
  NAND2_X1 U3504 ( .A1(n3864), .A2(n3865), .ZN(n3819) );
  AND2_X2 U3505 ( .A1(n4750), .A2(n4872), .ZN(n4742) );
  INV_X2 U3506 ( .A(n5370), .ZN(n3528) );
  CLKBUF_X2 U3507 ( .A(n3998), .Z(n4345) );
  BUF_X2 U3508 ( .A(n3770), .Z(n4372) );
  CLKBUF_X2 U3509 ( .A(n3641), .Z(n4045) );
  CLKBUF_X2 U3510 ( .A(n3706), .Z(n4371) );
  BUF_X4 U3511 ( .A(n3670), .Z(n3436) );
  NOR2_X1 U3512 ( .A1(n3451), .A2(n5396), .ZN(n5608) );
  OR2_X1 U3513 ( .A1(n5373), .A2(n6188), .ZN(n4545) );
  XNOR2_X1 U3514 ( .A(n4556), .B(n4555), .ZN(n5342) );
  AOI21_X1 U3515 ( .B1(n5415), .B2(n3460), .A(n3461), .ZN(n5618) );
  NAND2_X1 U3516 ( .A1(n6203), .A2(n4469), .ZN(n5703) );
  CLKBUF_X1 U3517 ( .A(n5533), .Z(n5544) );
  OR2_X1 U3518 ( .A1(n3448), .A2(n3449), .ZN(n5533) );
  NAND2_X1 U3519 ( .A1(n5299), .A2(n3513), .ZN(n5304) );
  AOI21_X1 U3520 ( .B1(n3553), .B2(n3547), .A(n3486), .ZN(n3546) );
  OR3_X1 U3521 ( .A1(n5210), .A2(n5227), .A3(n4066), .ZN(n4076) );
  NOR2_X2 U3522 ( .A1(n4961), .A2(n3446), .ZN(n5143) );
  NOR2_X1 U3523 ( .A1(n4961), .A2(n5135), .ZN(n5134) );
  OR2_X1 U3524 ( .A1(n4460), .A2(n4459), .ZN(n3463) );
  NOR2_X1 U3525 ( .A1(n5689), .A2(n3487), .ZN(n4475) );
  NAND2_X1 U3526 ( .A1(n5704), .A2(n5810), .ZN(n3561) );
  AND2_X1 U3527 ( .A1(n3908), .A2(n3447), .ZN(n4912) );
  AND2_X1 U3528 ( .A1(n3951), .A2(n3950), .ZN(n3975) );
  NOR2_X1 U3529 ( .A1(n6718), .A2(n6799), .ZN(n7118) );
  AND2_X1 U3530 ( .A1(n4415), .A2(n4414), .ZN(n6172) );
  OAI21_X1 U3531 ( .B1(n4938), .B2(n4107), .A(n4071), .ZN(n3872) );
  OR2_X1 U3532 ( .A1(n4938), .A2(n4611), .ZN(n4415) );
  NAND2_X1 U3533 ( .A1(n3508), .A2(n3842), .ZN(n3845) );
  XNOR2_X1 U3534 ( .A(n5107), .B(n5105), .ZN(n4941) );
  NAND2_X1 U3535 ( .A1(n3877), .A2(n3879), .ZN(n5107) );
  NAND2_X1 U3536 ( .A1(n4534), .A2(n4533), .ZN(n5365) );
  NAND2_X1 U3537 ( .A1(n3886), .A2(n3885), .ZN(n5105) );
  CLKBUF_X1 U3538 ( .A(n4594), .Z(n5109) );
  AND4_X1 U3539 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3762)
         );
  AND2_X1 U3540 ( .A1(n3813), .A2(n4393), .ZN(n3852) );
  AND3_X1 U3541 ( .A1(n4607), .A2(n6580), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3761) );
  INV_X1 U3542 ( .A(n5160), .ZN(n3438) );
  AND2_X1 U3543 ( .A1(n3757), .A2(n3684), .ZN(n3728) );
  NAND2_X1 U3544 ( .A1(n3793), .A2(n3792), .ZN(n3815) );
  AND2_X1 U3545 ( .A1(n3683), .A2(n5009), .ZN(n3684) );
  OAI211_X1 U3546 ( .C1(n4836), .C2(n3731), .A(n4402), .B(n3635), .ZN(n4581)
         );
  NOR2_X1 U3547 ( .A1(n4398), .A2(n3730), .ZN(n3733) );
  NAND2_X1 U3548 ( .A1(n3847), .A2(n3692), .ZN(n3731) );
  CLKBUF_X1 U3549 ( .A(n3726), .Z(n3727) );
  INV_X2 U3550 ( .A(n4750), .ZN(n5337) );
  AND2_X2 U3551 ( .A1(n3725), .A2(n5370), .ZN(n4396) );
  OR2_X1 U3552 ( .A1(n3805), .A2(n3804), .ZN(n4403) );
  INV_X4 U3553 ( .A(n4593), .ZN(n3725) );
  OR2_X1 U3554 ( .A1(n3776), .A2(n3775), .ZN(n4397) );
  AND2_X2 U3555 ( .A1(n4402), .A2(n4593), .ZN(n4750) );
  OR2_X1 U3556 ( .A1(n3789), .A2(n3788), .ZN(n4462) );
  NAND2_X1 U3557 ( .A1(n5370), .A2(n4593), .ZN(n5338) );
  AND4_X2 U3558 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n5009)
         );
  NAND4_X2 U3559 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(n4593)
         );
  AND2_X1 U3560 ( .A1(n3665), .A2(n3664), .ZN(n3682) );
  AND4_X1 U3561 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(n3622)
         );
  AND4_X1 U3562 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3656)
         );
  AND4_X1 U3563 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3718)
         );
  AND4_X1 U3564 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3559)
         );
  AND4_X1 U3565 ( .A1(n3674), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(n3680)
         );
  AND4_X1 U3566 ( .A1(n3593), .A2(n3592), .A3(n3591), .A4(n3590), .ZN(n3594)
         );
  AND4_X1 U3567 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3624)
         );
  AND4_X1 U3568 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3595)
         );
  AND4_X1 U3569 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3681)
         );
  AND4_X1 U3570 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3657)
         );
  AND4_X1 U3571 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3689)
         );
  NAND2_X2 U3572 ( .A1(n6808), .A2(n4392), .ZN(n6188) );
  AND4_X1 U3573 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3688)
         );
  AND4_X1 U3574 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3623)
         );
  AND4_X1 U3575 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3720)
         );
  AND4_X1 U3576 ( .A1(n3653), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3654)
         );
  AND4_X1 U3577 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3679)
         );
  AND4_X1 U3578 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3717)
         );
  AND4_X1 U3579 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(n3655)
         );
  AND4_X1 U3580 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3719)
         );
  CLKBUF_X2 U3581 ( .A(n3834), .Z(n4350) );
  AND2_X2 U3582 ( .A1(n5827), .A2(n5090), .ZN(n3659) );
  AND2_X2 U3583 ( .A1(n3581), .A2(n4877), .ZN(n3770) );
  BUF_X4 U3584 ( .A(n3663), .Z(n4373) );
  AND2_X2 U3585 ( .A1(n3576), .A2(n5827), .ZN(n3829) );
  AND2_X2 U3586 ( .A1(n4877), .A2(n5090), .ZN(n3663) );
  AND2_X2 U3587 ( .A1(n3880), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3576)
         );
  CLKBUF_X1 U3588 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n6544) );
  AND2_X2 U3589 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4877) );
  AND2_X2 U3590 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5086) );
  AND2_X1 U3591 ( .A1(n3541), .A2(n3439), .ZN(n4476) );
  NOR2_X1 U3592 ( .A1(n3538), .A2(n4475), .ZN(n3439) );
  INV_X2 U3593 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3566) );
  AND2_X1 U3594 ( .A1(n3928), .A2(n6725), .ZN(n5127) );
  NAND2_X1 U3595 ( .A1(n6181), .A2(n3443), .ZN(n3440) );
  AND2_X2 U3596 ( .A1(n3440), .A2(n3441), .ZN(n6192) );
  OR2_X2 U3597 ( .A1(n3442), .A2(n6184), .ZN(n3441) );
  INV_X1 U3598 ( .A(n4442), .ZN(n3442) );
  AND2_X1 U3599 ( .A1(n4433), .A2(n4442), .ZN(n3443) );
  AND2_X2 U3600 ( .A1(n4471), .A2(n3444), .ZN(n4472) );
  AND2_X1 U3601 ( .A1(n3485), .A2(n3561), .ZN(n3444) );
  NOR2_X1 U3602 ( .A1(n4562), .A2(n4546), .ZN(n3445) );
  NOR2_X1 U3603 ( .A1(n4562), .A2(n4546), .ZN(n5599) );
  NOR2_X1 U3604 ( .A1(n4865), .A2(n4931), .ZN(n3447) );
  NAND2_X1 U3605 ( .A1(n5299), .A2(n3513), .ZN(n3448) );
  OR2_X1 U3606 ( .A1(n3450), .A2(n5549), .ZN(n3449) );
  INV_X1 U3607 ( .A(n5542), .ZN(n3450) );
  AND2_X1 U3608 ( .A1(n5397), .A2(n5329), .ZN(n3451) );
  NAND2_X1 U3609 ( .A1(n3541), .A2(n3537), .ZN(n3452) );
  AND2_X1 U3610 ( .A1(n4877), .A2(n5086), .ZN(n3453) );
  AND2_X1 U3611 ( .A1(n4877), .A2(n5086), .ZN(n3454) );
  AND2_X2 U3612 ( .A1(n3576), .A2(n5828), .ZN(n3834) );
  INV_X2 U3613 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3824) );
  NAND2_X1 U3614 ( .A1(n4407), .A2(n4852), .ZN(n6171) );
  NAND2_X1 U3615 ( .A1(n3822), .A2(n3821), .ZN(n3878) );
  NOR2_X1 U3616 ( .A1(n3452), .A2(n5668), .ZN(n5662) );
  AOI21_X1 U3617 ( .B1(n5127), .B2(n4485), .A(n4423), .ZN(n4861) );
  OR2_X1 U3618 ( .A1(n3750), .A2(n3749), .ZN(n4606) );
  AOI22_X1 U3619 ( .A1(n3732), .A2(n4396), .B1(n3693), .B2(n4750), .ZN(n3760)
         );
  AND4_X2 U3620 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3763)
         );
  NAND2_X2 U3621 ( .A1(n3559), .A2(n3470), .ZN(n3849) );
  NAND2_X2 U3622 ( .A1(n3480), .A2(n4836), .ZN(n3751) );
  XNOR2_X1 U3623 ( .A(n3878), .B(n3877), .ZN(n4878) );
  AND2_X1 U3624 ( .A1(n3576), .A2(n4877), .ZN(n3456) );
  AND2_X1 U3625 ( .A1(n3576), .A2(n4877), .ZN(n3701) );
  BUF_X8 U3626 ( .A(n4206), .Z(n3457) );
  AND2_X2 U3627 ( .A1(n5115), .A2(n5090), .ZN(n4206) );
  OAI22_X2 U3628 ( .A1(n5175), .A2(n5174), .B1(n5179), .B2(n5704), .ZN(n5196)
         );
  AOI21_X2 U3629 ( .B1(n5168), .B2(n5169), .A(n3475), .ZN(n5175) );
  OR2_X2 U3630 ( .A1(n5469), .A2(n5514), .ZN(n3468) );
  OAI21_X2 U3631 ( .B1(n3471), .B2(n3522), .A(n3460), .ZN(n5624) );
  AND2_X2 U3632 ( .A1(n3576), .A2(n4877), .ZN(n3459) );
  OAI222_X1 U3633 ( .A1(n6600), .A2(n4942), .B1(n6601), .B2(n5133), .C1(n6793), 
        .C2(n6606), .ZN(U3464) );
  XNOR2_X2 U3634 ( .A(n3818), .B(n3819), .ZN(n4942) );
  OAI21_X1 U3635 ( .B1(n5373), .B2(n6490), .A(n3505), .ZN(n3504) );
  OR3_X1 U3636 ( .A1(n6226), .A2(n5023), .A3(n5022), .ZN(n6402) );
  OR2_X1 U3637 ( .A1(n5295), .A2(n5296), .ZN(n5822) );
  OR2_X1 U3638 ( .A1(n5365), .A2(n4884), .ZN(n4901) );
  AND2_X1 U3639 ( .A1(n3524), .A2(n4391), .ZN(n3523) );
  OAI21_X1 U3640 ( .B1(n5196), .B2(n3548), .A(n3546), .ZN(n6205) );
  NAND2_X1 U3641 ( .A1(n3512), .A2(n4066), .ZN(n4067) );
  NAND2_X1 U3642 ( .A1(n5143), .A2(n3481), .ZN(n3512) );
  AND2_X1 U3643 ( .A1(n5365), .A2(n6572), .ZN(n4777) );
  NAND2_X1 U3644 ( .A1(n5337), .A2(n4743), .ZN(n5339) );
  NAND2_X1 U3645 ( .A1(n4778), .A2(n4766), .ZN(n6226) );
  NAND2_X1 U3646 ( .A1(n3692), .A2(n3763), .ZN(n3726) );
  AND2_X2 U3647 ( .A1(n3824), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3581)
         );
  NAND2_X1 U3648 ( .A1(n3930), .A2(n3929), .ZN(n3949) );
  INV_X1 U3649 ( .A(n3928), .ZN(n3930) );
  AND2_X1 U3650 ( .A1(n3743), .A2(n3742), .ZN(n3745) );
  NAND2_X1 U3651 ( .A1(n3777), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3778) );
  NAND2_X1 U3652 ( .A1(n3729), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3823) );
  OR2_X1 U3653 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  INV_X1 U3654 ( .A(n5397), .ZN(n4343) );
  NAND2_X1 U3655 ( .A1(n5528), .A2(n3519), .ZN(n3518) );
  AND2_X1 U3656 ( .A1(n3520), .A2(n4156), .ZN(n3519) );
  INV_X1 U3657 ( .A(n5483), .ZN(n3520) );
  INV_X1 U3658 ( .A(n5227), .ZN(n3509) );
  AND2_X1 U3659 ( .A1(n3478), .A2(n5211), .ZN(n3510) );
  INV_X1 U3660 ( .A(n4341), .ZN(n4301) );
  NOR2_X1 U3661 ( .A1(n5516), .A2(n5515), .ZN(n3498) );
  OR2_X1 U3662 ( .A1(n3564), .A2(n3540), .ZN(n3539) );
  INV_X1 U3663 ( .A(n3563), .ZN(n3540) );
  NOR2_X1 U3664 ( .A1(n5629), .A2(n4473), .ZN(n3545) );
  NAND2_X1 U3665 ( .A1(n5629), .A2(n3488), .ZN(n3544) );
  INV_X1 U3666 ( .A(n3564), .ZN(n3543) );
  INV_X1 U3667 ( .A(n3545), .ZN(n3542) );
  NOR2_X1 U3668 ( .A1(n5137), .A2(n3502), .ZN(n3501) );
  INV_X1 U3669 ( .A(n5162), .ZN(n3502) );
  INV_X1 U3670 ( .A(n5138), .ZN(n3500) );
  INV_X1 U3671 ( .A(n3532), .ZN(n3531) );
  NAND2_X1 U3672 ( .A1(n5337), .A2(n4872), .ZN(n4729) );
  NAND2_X1 U3673 ( .A1(n4878), .A2(n6594), .ZN(n3508) );
  AND2_X1 U3674 ( .A1(n4943), .A2(n3825), .ZN(n4993) );
  INV_X1 U3675 ( .A(n3878), .ZN(n3879) );
  OR2_X1 U3676 ( .A1(n4880), .A2(n4838), .ZN(n4922) );
  NAND2_X1 U3677 ( .A1(n3528), .A2(n3725), .ZN(n4921) );
  OR2_X1 U3678 ( .A1(n4778), .A2(READY_N), .ZN(n4779) );
  AND2_X1 U3679 ( .A1(n3477), .A2(n5330), .ZN(n3521) );
  INV_X1 U3680 ( .A(n5291), .ZN(n4074) );
  NAND2_X1 U3681 ( .A1(n4038), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4068)
         );
  AND2_X1 U3682 ( .A1(n4011), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4025)
         );
  AND2_X1 U3683 ( .A1(n3966), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3977)
         );
  NAND2_X1 U3684 ( .A1(n5426), .A2(n5411), .ZN(n5413) );
  AND2_X1 U3685 ( .A1(n5552), .A2(n3484), .ZN(n5525) );
  INV_X1 U3686 ( .A(n5485), .ZN(n3494) );
  NAND2_X1 U3687 ( .A1(n5552), .A2(n3495), .ZN(n5538) );
  NAND2_X1 U3688 ( .A1(n5552), .A2(n3476), .ZN(n5547) );
  AND2_X1 U3689 ( .A1(n5552), .A2(n5551), .ZN(n5554) );
  NAND2_X1 U3690 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4470) );
  NAND2_X1 U3691 ( .A1(n3474), .A2(n3462), .ZN(n3551) );
  OR2_X1 U3692 ( .A1(n5147), .A2(n5191), .ZN(n5212) );
  MUX2_X1 U3693 ( .A(n3863), .B(n3862), .S(n3861), .Z(n6780) );
  INV_X1 U3694 ( .A(n6598), .ZN(n6572) );
  AOI21_X1 U3695 ( .B1(n5380), .B2(n5379), .A(n5378), .ZN(n3505) );
  AND2_X1 U3696 ( .A1(n6402), .A2(n5024), .ZN(n6530) );
  XNOR2_X1 U3697 ( .A(n4751), .B(n5336), .ZN(n5377) );
  AND2_X1 U3698 ( .A1(n5564), .A2(n5563), .ZN(n6838) );
  INV_X1 U3699 ( .A(n5564), .ZN(n6837) );
  AND2_X1 U3700 ( .A1(n5564), .A2(n4929), .ZN(n5306) );
  INV_X1 U3701 ( .A(n6209), .ZN(n6210) );
  NAND2_X1 U3702 ( .A1(n6209), .A2(n4541), .ZN(n6216) );
  AOI21_X1 U3703 ( .B1(n3731), .B2(n4402), .A(n4593), .ZN(n3754) );
  NOR2_X1 U3704 ( .A1(n4581), .A2(n3636), .ZN(n3757) );
  NAND2_X1 U3705 ( .A1(n4484), .A2(n4483), .ZN(n4514) );
  NAND2_X1 U3706 ( .A1(n3920), .A2(n3919), .ZN(n3929) );
  INV_X1 U3707 ( .A(n3949), .ZN(n3951) );
  OR2_X1 U3708 ( .A1(n3940), .A2(n3939), .ZN(n4452) );
  NOR2_X1 U3709 ( .A1(n4593), .A2(n4567), .ZN(n3739) );
  OR2_X1 U3710 ( .A1(n3841), .A2(n3840), .ZN(n4408) );
  OR2_X1 U3711 ( .A1(n3757), .A2(n3725), .ZN(n3758) );
  AOI22_X1 U3712 ( .A1(n3770), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U3713 ( .A1(n3712), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3591) );
  AND2_X1 U3714 ( .A1(n4836), .A2(n5370), .ZN(n3828) );
  INV_X1 U3715 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4525) );
  INV_X1 U3716 ( .A(n4524), .ZN(n4518) );
  AOI22_X1 U3717 ( .A1(n3835), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3701), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3634) );
  INV_X1 U3718 ( .A(n3731), .ZN(n4927) );
  AND2_X1 U3719 ( .A1(n4343), .A2(n3525), .ZN(n3524) );
  INV_X1 U3720 ( .A(n5382), .ZN(n3525) );
  INV_X1 U3721 ( .A(n5445), .ZN(n4264) );
  NAND2_X1 U3722 ( .A1(n5318), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4386) );
  INV_X1 U3723 ( .A(n5245), .ZN(n3549) );
  INV_X1 U3724 ( .A(n5189), .ZN(n3511) );
  AND2_X1 U3725 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4547)
         );
  AND2_X1 U3726 ( .A1(n3476), .A2(n3496), .ZN(n3495) );
  INV_X1 U3727 ( .A(n5536), .ZN(n3496) );
  AND2_X1 U3728 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3563)
         );
  OR2_X1 U3729 ( .A1(n3961), .A2(n3960), .ZN(n4451) );
  INV_X1 U3730 ( .A(n5339), .ZN(n4747) );
  INV_X1 U3731 ( .A(n6153), .ZN(n3492) );
  OR2_X1 U3732 ( .A1(n3896), .A2(n3895), .ZN(n4421) );
  AND2_X1 U3733 ( .A1(n3692), .A2(n4593), .ZN(n4485) );
  OR2_X1 U3734 ( .A1(n6252), .A2(n6242), .ZN(n4614) );
  NAND2_X1 U3735 ( .A1(n4395), .A2(n4485), .ZN(n3536) );
  NOR2_X1 U3736 ( .A1(n4402), .A2(n5370), .ZN(n3752) );
  NAND2_X1 U3737 ( .A1(n3735), .A2(n3725), .ZN(n4594) );
  OAI211_X1 U3738 ( .C1(n4905), .C2(n4904), .A(n4903), .B(n4902), .ZN(n5101)
         );
  AND2_X1 U3739 ( .A1(n4938), .A2(n6677), .ZN(n6778) );
  AND4_X1 U3740 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3625)
         );
  OAI21_X1 U3741 ( .B1(n6232), .B2(n6587), .A(n6590), .ZN(n4949) );
  AND2_X1 U3742 ( .A1(n4519), .A2(n4485), .ZN(n4532) );
  NOR2_X1 U3743 ( .A1(n3828), .A2(n6594), .ZN(n4529) );
  OR2_X1 U3745 ( .A1(n3823), .A2(n3880), .ZN(n3886) );
  INV_X1 U3746 ( .A(n5043), .ZN(n5029) );
  INV_X1 U3747 ( .A(n4921), .ZN(n3527) );
  NOR2_X1 U3748 ( .A1(n4917), .A2(n4647), .ZN(n6154) );
  AND2_X1 U3749 ( .A1(n4777), .A2(n4769), .ZN(n6049) );
  AND2_X1 U3750 ( .A1(n4389), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4557)
         );
  INV_X1 U3751 ( .A(n4071), .ZN(n4553) );
  NOR2_X1 U3752 ( .A1(n4337), .A2(n5328), .ZN(n4338) );
  INV_X1 U3753 ( .A(n4319), .ZN(n5330) );
  AND2_X1 U3754 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4283), .ZN(n4284)
         );
  NAND2_X1 U3755 ( .A1(n4279), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4282)
         );
  AND2_X1 U3756 ( .A1(n4259), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4279)
         );
  NOR2_X1 U3757 ( .A1(n4218), .A2(n4217), .ZN(n4219) );
  NOR2_X1 U3758 ( .A1(n3518), .A2(n3516), .ZN(n3515) );
  INV_X1 U3759 ( .A(n5470), .ZN(n3516) );
  AND2_X1 U3760 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4172), .ZN(n4173)
         );
  NAND2_X1 U3761 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4218)
         );
  INV_X1 U3762 ( .A(n3519), .ZN(n3517) );
  NOR2_X1 U3763 ( .A1(n4152), .A2(n5685), .ZN(n4153) );
  NAND2_X1 U3764 ( .A1(n4153), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4171)
         );
  NAND2_X1 U3765 ( .A1(n4124), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4152)
         );
  NOR2_X1 U3766 ( .A1(n4093), .A2(n4092), .ZN(n4110) );
  NOR2_X1 U3767 ( .A1(n5303), .A2(n3514), .ZN(n3513) );
  INV_X1 U3768 ( .A(n5301), .ZN(n3514) );
  NOR2_X1 U3769 ( .A1(n4068), .A2(n5230), .ZN(n4069) );
  AND2_X1 U3770 ( .A1(n4054), .A2(n4053), .ZN(n5227) );
  AND2_X1 U3771 ( .A1(n4025), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4038)
         );
  INV_X1 U3772 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3996) );
  CLKBUF_X1 U3773 ( .A(n5143), .Z(n5144) );
  NAND2_X1 U3774 ( .A1(n3977), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3997)
         );
  INV_X1 U3775 ( .A(n6193), .ZN(n3533) );
  AND2_X1 U3776 ( .A1(n6193), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3535)
         );
  AOI21_X1 U3777 ( .B1(n4443), .B2(n3848), .A(n3971), .ZN(n4962) );
  NOR2_X1 U3778 ( .A1(n3945), .A2(n3944), .ZN(n3966) );
  INV_X1 U3779 ( .A(n4865), .ZN(n3907) );
  NAND2_X1 U3780 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3902) );
  NOR2_X1 U3781 ( .A1(n5459), .A2(n4725), .ZN(n5426) );
  NAND2_X1 U3782 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4477) );
  NAND2_X1 U3783 ( .A1(n3498), .A2(n3497), .ZN(n5459) );
  INV_X1 U3784 ( .A(n5457), .ZN(n3497) );
  INV_X1 U3785 ( .A(n3498), .ZN(n5518) );
  AND2_X1 U3786 ( .A1(n4710), .A2(n4709), .ZN(n5471) );
  AND2_X1 U3787 ( .A1(n5525), .A2(n5524), .ZN(n5527) );
  INV_X1 U3788 ( .A(n3538), .ZN(n3537) );
  OAI21_X1 U3789 ( .B1(n3545), .B2(n3539), .A(n3544), .ZN(n3538) );
  NOR2_X1 U3790 ( .A1(n4472), .A2(n3563), .ZN(n5691) );
  NOR2_X2 U3791 ( .A1(n5822), .A2(n4689), .ZN(n5552) );
  NAND2_X1 U3792 ( .A1(n5689), .A2(n6259), .ZN(n4469) );
  INV_X1 U3793 ( .A(n6345), .ZN(n6252) );
  NOR2_X1 U3794 ( .A1(n5212), .A2(n5213), .ZN(n5232) );
  AND2_X1 U3795 ( .A1(n4673), .A2(n4672), .ZN(n5191) );
  INV_X1 U3796 ( .A(n5149), .ZN(n3499) );
  NAND2_X1 U3797 ( .A1(n3500), .A2(n3501), .ZN(n5165) );
  NOR2_X1 U3798 ( .A1(n5138), .A2(n5137), .ZN(n5163) );
  NAND2_X1 U3799 ( .A1(n4661), .A2(n4660), .ZN(n5138) );
  INV_X1 U3800 ( .A(n4964), .ZN(n4660) );
  INV_X1 U3801 ( .A(n4965), .ZN(n4661) );
  NAND3_X1 U3802 ( .A1(n3490), .A2(n3493), .A3(n3489), .ZN(n4965) );
  INV_X1 U3803 ( .A(n4647), .ZN(n3493) );
  NOR2_X1 U3804 ( .A1(n4914), .A2(n3492), .ZN(n3489) );
  NAND2_X1 U3805 ( .A1(n3490), .A2(n3491), .ZN(n6156) );
  NOR2_X1 U3806 ( .A1(n4647), .A2(n3492), .ZN(n3491) );
  INV_X1 U3807 ( .A(n4614), .ZN(n5051) );
  INV_X1 U3808 ( .A(n4880), .ZN(n3737) );
  AND3_X1 U3809 ( .A1(n3528), .A2(n3725), .A3(n3555), .ZN(n3738) );
  NAND2_X1 U3810 ( .A1(n4591), .A2(n6572), .ZN(n4738) );
  NAND2_X1 U3811 ( .A1(n3821), .A2(n3748), .ZN(n3818) );
  OR2_X1 U3812 ( .A1(n3823), .A2(n3824), .ZN(n3827) );
  NAND2_X1 U3813 ( .A1(n6594), .A2(n4949), .ZN(n5121) );
  AND2_X2 U3814 ( .A1(n3566), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5827)
         );
  OR3_X1 U3815 ( .A1(n6677), .A2(n4938), .A3(n3900), .ZN(n6718) );
  INV_X1 U3816 ( .A(n5121), .ZN(n6680) );
  NOR2_X1 U3817 ( .A1(n4985), .A2(n4939), .ZN(n6654) );
  AND4_X2 U3818 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n5562)
         );
  CLKBUF_X1 U3819 ( .A(n4341), .Z(n5020) );
  AND2_X1 U3820 ( .A1(n6585), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4535) );
  INV_X1 U3821 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6220) );
  AND2_X1 U3822 ( .A1(n6808), .A2(n6585), .ZN(n5229) );
  INV_X2 U3823 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6797) );
  AND2_X1 U3824 ( .A1(n6402), .A2(n5036), .ZN(n6528) );
  INV_X1 U3825 ( .A(n6524), .ZN(n6457) );
  INV_X1 U3826 ( .A(n6521), .ZN(n6434) );
  INV_X1 U3827 ( .A(n6157), .ZN(n6150) );
  NAND2_X1 U3828 ( .A1(n4901), .A2(n4840), .ZN(n4841) );
  NAND2_X1 U3829 ( .A1(n6162), .A2(n3722), .ZN(n6157) );
  OAI21_X1 U3830 ( .B1(n4924), .B2(n4923), .A(n6572), .ZN(n4925) );
  INV_X1 U3831 ( .A(n5306), .ZN(n5255) );
  AND2_X2 U3832 ( .A1(n4779), .A2(n4800), .ZN(n4847) );
  INV_X1 U3833 ( .A(n4800), .ZN(n4848) );
  INV_X1 U3834 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5685) );
  XNOR2_X1 U3835 ( .A(n5341), .B(n5340), .ZN(n5710) );
  OR2_X1 U3836 ( .A1(n5377), .A2(n6339), .ZN(n4756) );
  XNOR2_X1 U3837 ( .A(n5604), .B(n5603), .ZN(n5742) );
  NAND2_X1 U3838 ( .A1(n3435), .A2(n5602), .ZN(n5604) );
  AND2_X1 U3839 ( .A1(n5770), .A2(n4633), .ZN(n6321) );
  OR2_X1 U3840 ( .A1(n4738), .A2(n4884), .ZN(n6288) );
  NAND2_X1 U3841 ( .A1(n3550), .A2(n3551), .ZN(n5247) );
  NAND2_X1 U3842 ( .A1(n5196), .A2(n3552), .ZN(n3550) );
  AND2_X1 U3843 ( .A1(n3554), .A2(n4467), .ZN(n5216) );
  NAND2_X1 U3844 ( .A1(n5196), .A2(n5195), .ZN(n3554) );
  NOR2_X1 U3845 ( .A1(n5051), .A2(n5062), .ZN(n6292) );
  INV_X1 U3846 ( .A(n6339), .ZN(n6326) );
  INV_X1 U3847 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6794) );
  INV_X1 U3848 ( .A(n6780), .ZN(n6799) );
  INV_X1 U3849 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6793) );
  CLKBUF_X1 U3850 ( .A(n4395), .Z(n4939) );
  OR2_X1 U3851 ( .A1(n6800), .A2(n6799), .ZN(n7174) );
  INV_X1 U3852 ( .A(n7174), .ZN(n7158) );
  OAI211_X1 U3853 ( .C1(n6789), .C2(n7149), .A(n6788), .B(n6819), .ZN(n7151)
         );
  INV_X1 U3854 ( .A(n7061), .ZN(n7142) );
  OR2_X1 U3855 ( .A1(n6668), .A2(n6780), .ZN(n7046) );
  NAND2_X1 U3856 ( .A1(n6654), .A2(n6799), .ZN(n7084) );
  INV_X1 U3857 ( .A(n6872), .ZN(n6874) );
  INV_X1 U3858 ( .A(n6880), .ZN(n6913) );
  INV_X1 U3859 ( .A(n6910), .ZN(n6912) );
  INV_X1 U3860 ( .A(n6948), .ZN(n6950) );
  INV_X1 U3861 ( .A(n6986), .ZN(n6988) );
  INV_X1 U3862 ( .A(n7030), .ZN(n7032) );
  INV_X1 U3863 ( .A(n7070), .ZN(n7072) );
  AND2_X1 U3864 ( .A1(n6571), .A2(n6570), .ZN(n6599) );
  NAND2_X1 U3865 ( .A1(n5365), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6590) );
  NOR2_X1 U3866 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6580) );
  INV_X1 U3867 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6594) );
  INV_X1 U3868 ( .A(n6591), .ZN(n6232) );
  INV_X1 U3869 ( .A(n6579), .ZN(n6589) );
  NOR2_X1 U3870 ( .A1(n6220), .A2(STATE_REG_0__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U3871 ( .A1(n3506), .A2(n3503), .ZN(U2797) );
  OR2_X1 U3872 ( .A1(n5377), .A2(n6510), .ZN(n3506) );
  INV_X1 U3873 ( .A(n3504), .ZN(n3503) );
  AND2_X2 U3874 ( .A1(n5115), .A2(n3581), .ZN(n3835) );
  AND2_X2 U3875 ( .A1(n3576), .A2(n5115), .ZN(n3998) );
  NAND2_X1 U3876 ( .A1(n5444), .A2(n3466), .ZN(n3460) );
  AND2_X1 U3877 ( .A1(n5444), .A2(n3477), .ZN(n3461) );
  NOR2_X1 U3878 ( .A1(n5544), .A2(n3517), .ZN(n5482) );
  NAND2_X1 U3879 ( .A1(n5704), .A2(n5250), .ZN(n3462) );
  AND2_X2 U3880 ( .A1(n3581), .A2(n5827), .ZN(n3626) );
  NOR2_X1 U3881 ( .A1(n3518), .A2(n5544), .ZN(n5468) );
  AND2_X1 U3882 ( .A1(n5143), .A2(n3478), .ZN(n5188) );
  OAI21_X1 U3883 ( .B1(n3823), .B2(n3566), .A(n3794), .ZN(n3864) );
  INV_X1 U3884 ( .A(n3553), .ZN(n3552) );
  NAND2_X1 U3885 ( .A1(n3462), .A2(n5195), .ZN(n3553) );
  AND2_X1 U3886 ( .A1(n3501), .A2(n3499), .ZN(n3464) );
  AND2_X1 U3887 ( .A1(n4401), .A2(n5066), .ZN(n3465) );
  INV_X1 U3888 ( .A(n4467), .ZN(n4468) );
  INV_X1 U3889 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3880) );
  AND2_X1 U3890 ( .A1(n4264), .A2(n3522), .ZN(n3466) );
  OR2_X1 U3891 ( .A1(n5413), .A2(n4732), .ZN(n3467) );
  OR2_X1 U3893 ( .A1(n5691), .A2(n3564), .ZN(n3469) );
  OAI211_X1 U3894 ( .C1(n3823), .C2(n3567), .A(n3744), .B(n3745), .ZN(n3821)
         );
  AND4_X1 U3895 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3470)
         );
  NOR2_X1 U3896 ( .A1(n5304), .A2(n5549), .ZN(n5541) );
  NAND2_X1 U3897 ( .A1(n4157), .A2(n4156), .ZN(n5481) );
  XNOR2_X1 U3898 ( .A(n3928), .B(n3929), .ZN(n4426) );
  AND2_X1 U3899 ( .A1(n5444), .A2(n4264), .ZN(n3471) );
  NAND2_X1 U3900 ( .A1(n4429), .A2(n4428), .ZN(n4432) );
  XNOR2_X1 U3901 ( .A(n4432), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6179)
         );
  OR2_X1 U3902 ( .A1(n4403), .A2(n4393), .ZN(n3472) );
  AND2_X1 U3903 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3473)
         );
  INV_X1 U3904 ( .A(n3548), .ZN(n3547) );
  NAND2_X1 U3905 ( .A1(n3551), .A2(n3549), .ZN(n3548) );
  OR2_X1 U3906 ( .A1(n4468), .A2(n3473), .ZN(n3474) );
  NAND2_X1 U3907 ( .A1(n3827), .A2(n3826), .ZN(n3877) );
  AND2_X1 U3908 ( .A1(n4465), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3475)
         );
  NOR2_X4 U3909 ( .A1(n5561), .A2(n6797), .ZN(n3927) );
  NAND2_X1 U3910 ( .A1(n5299), .A2(n5301), .ZN(n5300) );
  INV_X1 U3911 ( .A(n3764), .ZN(n4307) );
  NAND2_X1 U3912 ( .A1(n5143), .A2(n5146), .ZN(n5145) );
  INV_X1 U3913 ( .A(n3730), .ZN(n3847) );
  AND2_X1 U3914 ( .A1(n5545), .A2(n5551), .ZN(n3476) );
  AND2_X1 U3915 ( .A1(n3466), .A2(n5414), .ZN(n3477) );
  NAND2_X1 U3916 ( .A1(n3534), .A2(n3532), .ZN(n6197) );
  AND2_X1 U3917 ( .A1(n3511), .A2(n5146), .ZN(n3478) );
  AND2_X1 U3918 ( .A1(n5704), .A2(n4632), .ZN(n3479) );
  INV_X1 U3919 ( .A(n3900), .ZN(n5126) );
  NAND2_X1 U3920 ( .A1(n3898), .A2(n3897), .ZN(n3900) );
  AND2_X1 U3921 ( .A1(n3510), .A2(n3509), .ZN(n3481) );
  OR2_X1 U3922 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3482)
         );
  OR2_X1 U3923 ( .A1(n5365), .A2(n3527), .ZN(n3483) );
  AND2_X1 U3924 ( .A1(n3495), .A2(n3494), .ZN(n3484) );
  OR2_X1 U3925 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3485)
         );
  BUF_X1 U3926 ( .A(n3712), .Z(n4046) );
  INV_X1 U3927 ( .A(n3507), .ZN(n4569) );
  NAND2_X1 U3928 ( .A1(n3733), .A2(n4585), .ZN(n3507) );
  NAND2_X1 U3929 ( .A1(n4419), .A2(n4418), .ZN(n4860) );
  AND2_X1 U3930 ( .A1(n5704), .A2(n4676), .ZN(n3486) );
  NAND2_X1 U3931 ( .A1(n3875), .A2(n3874), .ZN(n4935) );
  AND4_X1 U3932 ( .A1(n5772), .A2(n5788), .A3(n5754), .A4(n5768), .ZN(n3487)
         );
  NAND3_X1 U3933 ( .A1(n4695), .A2(n5678), .A3(n4474), .ZN(n3488) );
  NOR2_X2 U3934 ( .A1(n5274), .A2(n5009), .ZN(n6911) );
  NAND3_X1 U3935 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6594), .A3(n4949), .ZN(
        n5274) );
  INV_X1 U3936 ( .A(n4917), .ZN(n3490) );
  NAND2_X1 U3937 ( .A1(n3500), .A2(n3464), .ZN(n5147) );
  NAND3_X1 U3938 ( .A1(n3733), .A2(n4585), .A3(n5370), .ZN(n4758) );
  NAND2_X1 U3939 ( .A1(n5143), .A2(n3510), .ZN(n5210) );
  NAND2_X1 U3940 ( .A1(n4157), .A2(n3515), .ZN(n5469) );
  NAND2_X2 U3941 ( .A1(n6724), .A2(n3901), .ZN(n4938) );
  INV_X1 U3942 ( .A(n4281), .ZN(n3522) );
  NAND2_X1 U3943 ( .A1(n4344), .A2(n4343), .ZN(n5395) );
  AND2_X1 U3944 ( .A1(n4344), .A2(n3524), .ZN(n5381) );
  NAND2_X1 U3945 ( .A1(n4344), .A2(n3523), .ZN(n4556) );
  NAND2_X1 U3946 ( .A1(n3526), .A2(n4861), .ZN(n4425) );
  NAND3_X1 U3947 ( .A1(n4419), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n4418), 
        .ZN(n3526) );
  NAND2_X1 U3948 ( .A1(n4860), .A2(n5055), .ZN(n4424) );
  AND2_X1 U3949 ( .A1(n4592), .A2(n3527), .ZN(n4894) );
  NAND2_X1 U3950 ( .A1(n5029), .A2(n3527), .ZN(n5025) );
  NAND2_X1 U3951 ( .A1(n3529), .A2(n3463), .ZN(n5168) );
  NAND2_X1 U3952 ( .A1(n3534), .A2(n3530), .ZN(n3529) );
  NOR2_X1 U3953 ( .A1(n6198), .A2(n3531), .ZN(n3530) );
  NAND2_X1 U3954 ( .A1(n3533), .A2(n6274), .ZN(n3532) );
  OR2_X2 U3955 ( .A1(n6192), .A2(n3535), .ZN(n3534) );
  NAND2_X1 U3956 ( .A1(n3536), .A2(n4401), .ZN(n4406) );
  NAND2_X1 U3957 ( .A1(n3536), .A2(n3465), .ZN(n4851) );
  NAND3_X1 U3958 ( .A1(n4472), .A2(n3543), .A3(n3542), .ZN(n3541) );
  XNOR2_X1 U3959 ( .A(n4565), .B(n4564), .ZN(n5334) );
  AOI22_X1 U3960 ( .A1(n3998), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3633) );
  NAND2_X1 U3961 ( .A1(n3626), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3599)
         );
  AOI22_X1 U3962 ( .A1(n3711), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3626), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3587) );
  AND2_X2 U3963 ( .A1(n5827), .A2(n5086), .ZN(n3670) );
  OAI22_X1 U3964 ( .A1(n5599), .A2(n5588), .B1(n5629), .B2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5592) );
  OAI21_X1 U3965 ( .B1(n5381), .B2(n4391), .A(n4556), .ZN(n5373) );
  INV_X1 U3966 ( .A(n5329), .ZN(n4344) );
  AOI21_X1 U3967 ( .B1(n5342), .B2(n6211), .A(n4560), .ZN(n4561) );
  NAND2_X1 U3968 ( .A1(n3847), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4107) );
  AND2_X1 U3969 ( .A1(n4756), .A2(n4755), .ZN(n3556) );
  AND2_X1 U3970 ( .A1(n3998), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3557) );
  AND2_X1 U3971 ( .A1(n5455), .A2(n5445), .ZN(n3558) );
  AND2_X1 U3972 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3560) );
  OR2_X1 U3973 ( .A1(n3746), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3562)
         );
  NAND2_X1 U3974 ( .A1(n5051), .A2(n6288), .ZN(n5817) );
  INV_X1 U3975 ( .A(n5817), .ZN(n5807) );
  AND2_X1 U3976 ( .A1(n5704), .A2(n5678), .ZN(n3564) );
  NAND2_X1 U3977 ( .A1(n3844), .A2(n3843), .ZN(n6724) );
  INV_X1 U3978 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5132) );
  INV_X1 U3979 ( .A(n5303), .ZN(n4109) );
  INV_X1 U3980 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4517) );
  INV_X1 U3981 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4482) );
  AND2_X1 U3982 ( .A1(n4562), .A2(n5611), .ZN(n3565) );
  OR2_X1 U3983 ( .A1(n3918), .A2(n3917), .ZN(n4435) );
  NOR2_X1 U3984 ( .A1(n4836), .A2(n3722), .ZN(n3724) );
  AND2_X1 U3985 ( .A1(n3723), .A2(n3849), .ZN(n3635) );
  INV_X1 U3986 ( .A(n4532), .ZN(n4520) );
  INV_X1 U3987 ( .A(n4491), .ZN(n4493) );
  AOI22_X1 U3988 ( .A1(n3770), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3706), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3631) );
  INV_X1 U3989 ( .A(n5534), .ZN(n4156) );
  INV_X1 U3990 ( .A(n4962), .ZN(n3972) );
  NAND2_X1 U3991 ( .A1(n3712), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3582)
         );
  INV_X1 U3992 ( .A(n4386), .ZN(n4363) );
  INV_X1 U3993 ( .A(n4485), .ZN(n4611) );
  AND2_X1 U3994 ( .A1(n5089), .A2(n5088), .ZN(n6559) );
  NAND2_X1 U3995 ( .A1(n4528), .A2(n4527), .ZN(n4574) );
  INV_X1 U3996 ( .A(n4742), .ZN(n4728) );
  INV_X1 U3997 ( .A(n3927), .ZN(n4361) );
  INV_X1 U3998 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4217) );
  AOI21_X1 U3999 ( .B1(n3981), .B2(n3848), .A(n3980), .ZN(n5135) );
  AND2_X1 U4000 ( .A1(n4547), .A2(n3560), .ZN(n4548) );
  AND2_X1 U4001 ( .A1(n4694), .A2(n4693), .ZN(n5545) );
  NAND2_X1 U4002 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U4003 ( .A1(n3738), .A2(n3737), .ZN(n4734) );
  NAND2_X1 U4004 ( .A1(n4532), .A2(n4574), .ZN(n4533) );
  INV_X1 U4005 ( .A(n4939), .ZN(n6677) );
  NAND2_X1 U4006 ( .A1(n4518), .A2(n4517), .ZN(n4575) );
  AND2_X1 U4007 ( .A1(n5416), .A2(n5348), .ZN(n5383) );
  INV_X1 U4008 ( .A(n4171), .ZN(n4172) );
  AND2_X1 U4009 ( .A1(n4110), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4124)
         );
  INV_X1 U4010 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5230) );
  OR2_X1 U4011 ( .A1(n6322), .A2(n5021), .ZN(n5022) );
  NAND2_X1 U4012 ( .A1(n6402), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U4013 ( .A1(n5029), .A2(n5028), .ZN(n6521) );
  AND3_X1 U4014 ( .A1(n4024), .A2(n4023), .A3(n4022), .ZN(n5189) );
  NAND2_X1 U4015 ( .A1(n4897), .A2(n4896), .ZN(n4924) );
  NAND2_X1 U4016 ( .A1(n4284), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4337)
         );
  AND2_X1 U4017 ( .A1(n4219), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4259)
         );
  INV_X1 U4018 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4092) );
  NOR2_X1 U4019 ( .A1(n3997), .A2(n3996), .ZN(n4011) );
  INV_X1 U4020 ( .A(n3902), .ZN(n3903) );
  NAND2_X1 U4021 ( .A1(n5629), .A2(n5601), .ZN(n5602) );
  NOR2_X1 U4022 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6252), .ZN(n5062)
         );
  INV_X1 U4023 ( .A(n5101), .ZN(n6555) );
  OR3_X1 U4024 ( .A1(n6726), .A2(n4939), .A3(n6725), .ZN(n6738) );
  NAND2_X1 U4025 ( .A1(n6785), .A2(n6808), .ZN(n6825) );
  AOI21_X1 U4026 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6794), .A(n5121), .ZN(
        n6806) );
  NOR2_X1 U4027 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4341) );
  INV_X1 U4028 ( .A(n5650), .ZN(n6529) );
  NAND2_X1 U4029 ( .A1(n4069), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4093)
         );
  INV_X1 U4030 ( .A(n6455), .ZN(n6499) );
  AND2_X1 U4031 ( .A1(n5350), .A2(n5040), .ZN(n6526) );
  INV_X1 U4032 ( .A(n6162), .ZN(n5531) );
  INV_X1 U4033 ( .A(n4926), .ZN(n4815) );
  INV_X1 U4034 ( .A(n6216), .ZN(n6206) );
  NAND2_X1 U4035 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3903), .ZN(n3945)
         );
  AND2_X1 U4036 ( .A1(n4777), .A2(n6563), .ZN(n6212) );
  OR2_X1 U4037 ( .A1(n4738), .A2(n4737), .ZN(n6339) );
  OAI21_X1 U4038 ( .B1(n6289), .B2(n6288), .A(n6268), .ZN(n6276) );
  INV_X1 U4039 ( .A(n6334), .ZN(n6327) );
  OR2_X1 U4040 ( .A1(n4586), .A2(n3725), .ZN(n6550) );
  INV_X1 U4041 ( .A(n7001), .ZN(n7169) );
  NOR2_X1 U4042 ( .A1(n5127), .A2(n6748), .ZN(n6767) );
  INV_X1 U4043 ( .A(n7141), .ZN(n7129) );
  INV_X1 U4044 ( .A(n6711), .ZN(n7116) );
  INV_X1 U4045 ( .A(n7115), .ZN(n7103) );
  INV_X1 U4046 ( .A(n7102), .ZN(n7043) );
  INV_X1 U4047 ( .A(n7046), .ZN(n7091) );
  INV_X1 U4048 ( .A(n7090), .ZN(n7078) );
  INV_X1 U4049 ( .A(n6811), .ZN(n6828) );
  INV_X1 U4050 ( .A(n7162), .ZN(n7167) );
  AND2_X1 U4051 ( .A1(n6578), .A2(n6577), .ZN(n6579) );
  NAND2_X1 U4052 ( .A1(n4777), .A2(n5361), .ZN(n4778) );
  INV_X1 U4053 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6817) );
  INV_X1 U4054 ( .A(n6506), .ZN(n6533) );
  INV_X1 U4055 ( .A(n6530), .ZN(n6490) );
  INV_X1 U4056 ( .A(n6528), .ZN(n6515) );
  AND2_X2 U4057 ( .A1(n4841), .A2(n6572), .ZN(n6162) );
  INV_X1 U4058 ( .A(n5260), .ZN(n5288) );
  NAND2_X1 U4059 ( .A1(n4926), .A2(n4925), .ZN(n5564) );
  NAND2_X2 U4060 ( .A1(n5564), .A2(n4928), .ZN(n6635) );
  INV_X1 U4061 ( .A(n6049), .ZN(n6078) );
  NAND2_X1 U4062 ( .A1(n4777), .A2(n4776), .ZN(n4800) );
  OR2_X1 U4063 ( .A1(n6212), .A2(n4538), .ZN(n6209) );
  INV_X1 U4064 ( .A(n6212), .ZN(n6535) );
  AND2_X1 U4065 ( .A1(n5769), .A2(n4624), .ZN(n6332) );
  OR2_X1 U4066 ( .A1(n4738), .A2(n4597), .ZN(n6334) );
  OR2_X1 U4067 ( .A1(n4738), .A2(n6550), .ZN(n6345) );
  INV_X1 U4068 ( .A(n3458), .ZN(n6785) );
  INV_X1 U4069 ( .A(n6798), .ZN(n7163) );
  NAND2_X1 U4070 ( .A1(n6767), .A2(n6780), .ZN(n7154) );
  NAND2_X1 U4071 ( .A1(n6767), .A2(n6799), .ZN(n7061) );
  INV_X1 U4072 ( .A(n6740), .ZN(n7135) );
  INV_X1 U4073 ( .A(n7118), .ZN(n7128) );
  INV_X1 U4074 ( .A(n6717), .ZN(n7122) );
  OR2_X1 U4075 ( .A1(n6692), .A2(n6799), .ZN(n7115) );
  INV_X1 U4076 ( .A(n6691), .ZN(n7109) );
  OR2_X1 U4077 ( .A1(n6668), .A2(n6799), .ZN(n7102) );
  NAND2_X1 U4078 ( .A1(n6654), .A2(n6780), .ZN(n7090) );
  AND2_X1 U4079 ( .A1(n4992), .A2(n4991), .ZN(n5287) );
  OR2_X1 U4080 ( .A1(n4950), .A2(n6780), .ZN(n7001) );
  INV_X1 U4081 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6585) );
  INV_X1 U4082 ( .A(n6612), .ZN(n6046) );
  INV_X1 U4083 ( .A(n6119), .ZN(n6115) );
  NAND2_X1 U4084 ( .A1(n3436), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3571)
         );
  INV_X1 U4085 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U4086 ( .A1(n3706), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3570)
         );
  NAND2_X1 U4087 ( .A1(n3835), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3569) );
  NOR2_X4 U4088 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U4089 ( .A1(n3457), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3568) );
  AND4_X2 U4090 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3691)
         );
  AND2_X2 U4091 ( .A1(n5828), .A2(n5090), .ZN(n3641) );
  NAND2_X1 U4092 ( .A1(n3641), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3575) );
  NAND2_X1 U4093 ( .A1(n3829), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4094 ( .A1(n3834), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3573) );
  NAND2_X1 U4095 ( .A1(n3456), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3572) );
  NAND2_X1 U4096 ( .A1(n3998), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4097 ( .A1(n3770), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3579)
         );
  NAND2_X1 U4098 ( .A1(n3659), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3578) );
  NAND2_X1 U4099 ( .A1(n3663), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U4100 ( .A1(n3711), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3585) );
  NAND2_X1 U4101 ( .A1(n3626), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3584)
         );
  AND2_X4 U4102 ( .A1(n4877), .A2(n5086), .ZN(n3765) );
  NAND2_X1 U4103 ( .A1(n3454), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3583)
         );
  AOI22_X1 U4104 ( .A1(n3835), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4206), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4105 ( .A1(n3829), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4106 ( .A1(n3998), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3706), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4107 ( .A1(n3834), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3701), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4108 ( .A1(n3659), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3590) );
  NAND2_X2 U4109 ( .A1(n3595), .A2(n3594), .ZN(n3730) );
  NAND2_X1 U4110 ( .A1(n3711), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3598) );
  NAND2_X1 U4111 ( .A1(n3998), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3597) );
  NAND2_X1 U4112 ( .A1(n3765), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3596)
         );
  NAND2_X1 U4113 ( .A1(n3436), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3603)
         );
  NAND2_X1 U4114 ( .A1(n3706), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3602)
         );
  NAND2_X1 U4115 ( .A1(n3641), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3601) );
  NAND2_X1 U4116 ( .A1(n3835), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3600) );
  NAND2_X1 U4117 ( .A1(n3829), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4118 ( .A1(n3834), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4119 ( .A1(n3701), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4120 ( .A1(n3457), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4121 ( .A1(n3770), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3611)
         );
  NAND2_X1 U4122 ( .A1(n3659), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4123 ( .A1(n3663), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3609) );
  NAND2_X1 U4124 ( .A1(n3712), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3608)
         );
  AOI22_X1 U4125 ( .A1(n3626), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4126 ( .A1(n3770), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4127 ( .A1(n3829), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4128 ( .A1(n3641), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3701), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4129 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3621)
         );
  AOI22_X1 U4130 ( .A1(n3711), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4131 ( .A1(n3834), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4132 ( .A1(n3712), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4133 ( .A1(n3659), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3706), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3616) );
  NAND4_X1 U4134 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3620)
         );
  NAND2_X1 U4135 ( .A1(n5562), .A2(n3730), .ZN(n3723) );
  AOI22_X1 U4136 ( .A1(n3829), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4137 ( .A1(n3436), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3712), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4138 ( .A1(n3711), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3626), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4139 ( .A1(n3834), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4140 ( .A1(n3659), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3632) );
  AND2_X1 U4141 ( .A1(n3731), .A2(n4836), .ZN(n3636) );
  NAND2_X1 U4142 ( .A1(n3706), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3640)
         );
  NAND2_X1 U4143 ( .A1(n3834), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U4144 ( .A1(n3701), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4145 ( .A1(n3457), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4146 ( .A1(n3835), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4147 ( .A1(n3436), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3644)
         );
  NAND2_X1 U4148 ( .A1(n3829), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3643) );
  NAND2_X1 U4149 ( .A1(n3641), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4150 ( .A1(n3998), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3649) );
  NAND2_X1 U4151 ( .A1(n3711), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3648) );
  NAND2_X1 U4152 ( .A1(n3770), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3647)
         );
  NAND2_X1 U4153 ( .A1(n3663), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U4154 ( .A1(n3626), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3653)
         );
  NAND2_X1 U4155 ( .A1(n3659), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4156 ( .A1(n3765), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3651)
         );
  NAND2_X1 U4157 ( .A1(n3712), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3650)
         );
  XNOR2_X1 U4158 ( .A(n6220), .B(STATE_REG_2__SCAN_IN), .ZN(n4567) );
  INV_X1 U4159 ( .A(n3739), .ZN(n3658) );
  NAND2_X1 U4160 ( .A1(n3658), .A2(n5562), .ZN(n3683) );
  NAND2_X1 U4161 ( .A1(n3659), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4162 ( .A1(n3770), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3660)
         );
  NAND2_X1 U4163 ( .A1(n3661), .A2(n3660), .ZN(n3662) );
  NOR2_X1 U4164 ( .A1(n3557), .A2(n3662), .ZN(n3665) );
  NAND2_X1 U4165 ( .A1(n4373), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3664) );
  NAND2_X1 U4166 ( .A1(n3711), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4167 ( .A1(n3626), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3668)
         );
  NAND2_X1 U4168 ( .A1(n3765), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3667)
         );
  NAND2_X1 U4169 ( .A1(n3712), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3666)
         );
  NAND2_X1 U4170 ( .A1(n3436), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3674)
         );
  NAND2_X1 U4171 ( .A1(n3706), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3673)
         );
  NAND2_X1 U4172 ( .A1(n3835), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3672) );
  NAND2_X1 U4173 ( .A1(n3457), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4174 ( .A1(n3641), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4175 ( .A1(n3829), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4176 ( .A1(n3834), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4177 ( .A1(n3701), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3675) );
  INV_X1 U4178 ( .A(n3692), .ZN(n3685) );
  NAND2_X1 U4179 ( .A1(n3685), .A2(n3555), .ZN(n3686) );
  NAND2_X1 U4180 ( .A1(n3751), .A2(n3686), .ZN(n3687) );
  NAND2_X1 U4181 ( .A1(n3687), .A2(n5009), .ZN(n3695) );
  INV_X1 U4182 ( .A(n3726), .ZN(n3693) );
  NAND2_X1 U4183 ( .A1(n3693), .A2(n3555), .ZN(n4536) );
  NOR2_X2 U4184 ( .A1(n4536), .A2(n5009), .ZN(n3734) );
  INV_X1 U4185 ( .A(n3734), .ZN(n3694) );
  NAND2_X1 U4186 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  NAND2_X1 U4187 ( .A1(n3696), .A2(n3754), .ZN(n3721) );
  NAND2_X1 U4188 ( .A1(n3998), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4189 ( .A1(n3770), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3699)
         );
  NAND2_X1 U4190 ( .A1(n3659), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U4191 ( .A1(n3663), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U4192 ( .A1(n3641), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3705) );
  NAND2_X1 U4193 ( .A1(n3829), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U4194 ( .A1(n3834), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4195 ( .A1(n3701), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4196 ( .A1(n3436), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3710)
         );
  NAND2_X1 U4197 ( .A1(n3706), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3709)
         );
  NAND2_X1 U4198 ( .A1(n3835), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U4199 ( .A1(n3457), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U4200 ( .A1(n3626), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3716)
         );
  NAND2_X1 U4201 ( .A1(n3711), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4202 ( .A1(n3765), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3714)
         );
  NAND2_X1 U4203 ( .A1(n3712), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3713)
         );
  NAND4_X4 U4204 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n5370)
         );
  NAND2_X1 U4205 ( .A1(n3721), .A2(n3528), .ZN(n3750) );
  NAND2_X1 U4206 ( .A1(n3724), .A2(n3723), .ZN(n3732) );
  NAND3_X1 U4207 ( .A1(n3728), .A2(n3750), .A3(n3760), .ZN(n3729) );
  NAND2_X1 U4208 ( .A1(n5009), .A2(n4402), .ZN(n4398) );
  NOR2_X2 U4209 ( .A1(n3732), .A2(n4927), .ZN(n4585) );
  NAND2_X1 U4210 ( .A1(n3734), .A2(n3752), .ZN(n4586) );
  INV_X1 U4211 ( .A(n4586), .ZN(n3735) );
  NOR2_X1 U4212 ( .A1(n4402), .A2(n3692), .ZN(n3736) );
  NAND2_X1 U4213 ( .A1(n3736), .A2(n5009), .ZN(n4880) );
  OAI211_X1 U4214 ( .C1(n4758), .C2(n3739), .A(n4594), .B(n4734), .ZN(n3740)
         );
  NAND2_X1 U4215 ( .A1(n3740), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4216 ( .A1(n6580), .A2(n6594), .ZN(n4537) );
  NAND2_X1 U4217 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6766) );
  NOR2_X1 U4218 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6813) );
  INV_X1 U4219 ( .A(n6813), .ZN(n3741) );
  NAND2_X1 U4220 ( .A1(n6766), .A2(n3741), .ZN(n6727) );
  OR2_X1 U4221 ( .A1(n4537), .A2(n6727), .ZN(n3743) );
  INV_X1 U4222 ( .A(n4535), .ZN(n3883) );
  NAND2_X1 U4223 ( .A1(n3883), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3742) );
  INV_X1 U4224 ( .A(n3744), .ZN(n3747) );
  INV_X1 U4225 ( .A(n3745), .ZN(n3746) );
  NAND2_X1 U4226 ( .A1(n3747), .A2(n3562), .ZN(n3748) );
  MUX2_X1 U4227 ( .A(n4535), .B(n4537), .S(n6794), .Z(n3794) );
  NOR2_X1 U4228 ( .A1(n3727), .A2(n3725), .ZN(n3749) );
  INV_X1 U4229 ( .A(n3751), .ZN(n5318) );
  AND2_X1 U4230 ( .A1(n3752), .A2(n5009), .ZN(n3753) );
  NAND2_X1 U4231 ( .A1(n5318), .A2(n3753), .ZN(n4607) );
  INV_X1 U4232 ( .A(n3754), .ZN(n3755) );
  NAND2_X1 U4233 ( .A1(n3755), .A2(n5009), .ZN(n3756) );
  NAND2_X1 U4234 ( .A1(n3756), .A2(n5370), .ZN(n3759) );
  NAND2_X1 U4235 ( .A1(n4606), .A2(n3762), .ZN(n3865) );
  NAND2_X1 U4236 ( .A1(n4942), .A2(n6594), .ZN(n3779) );
  INV_X1 U4237 ( .A(n3626), .ZN(n3764) );
  AOI22_X1 U4238 ( .A1(n4307), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4239 ( .A1(n4366), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4240 ( .A1(n4045), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4241 ( .A1(n4201), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3766) );
  NAND4_X1 U4242 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3776)
         );
  AOI22_X1 U4243 ( .A1(n3437), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4244 ( .A1(n4372), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4245 ( .A1(n3712), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4246 ( .A1(n3706), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4247 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3775)
         );
  NAND2_X1 U4248 ( .A1(n3763), .A2(n4397), .ZN(n3777) );
  NAND2_X1 U4249 ( .A1(n4519), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3793) );
  INV_X1 U4250 ( .A(n4397), .ZN(n3790) );
  AOI22_X1 U4251 ( .A1(n4345), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4252 ( .A1(n4372), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3706), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4253 ( .A1(n3437), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3781) );
  BUF_X1 U4254 ( .A(n3436), .Z(n4366) );
  AOI22_X1 U4255 ( .A1(n4366), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4256 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4257 ( .A1(n3834), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4258 ( .A1(n4307), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3712), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4259 ( .A1(n3795), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4260 ( .A1(n3711), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4261 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  OAI22_X1 U4262 ( .A1(n3790), .A2(n5370), .B1(n4836), .B2(n4462), .ZN(n3791)
         );
  NAND2_X1 U4263 ( .A1(n3791), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3792) );
  AND2_X1 U4264 ( .A1(n3794), .A2(n6594), .ZN(n3859) );
  NOR2_X1 U4265 ( .A1(n4836), .A2(n6594), .ZN(n3806) );
  INV_X1 U4266 ( .A(n4462), .ZN(n3809) );
  AOI22_X1 U4267 ( .A1(n4374), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3706), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4268 ( .A1(n4045), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4269 ( .A1(n4345), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3712), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3797) );
  BUF_X1 U4270 ( .A(n3835), .Z(n3795) );
  AOI22_X1 U4271 ( .A1(n3795), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3796) );
  NAND4_X1 U4272 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3805)
         );
  AOI22_X1 U4273 ( .A1(n3437), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4274 ( .A1(n4372), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4275 ( .A1(n3711), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4276 ( .A1(n4307), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3800) );
  NAND4_X1 U4277 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3804)
         );
  NAND3_X1 U4278 ( .A1(n3806), .A2(n3809), .A3(n4403), .ZN(n3807) );
  NAND2_X1 U4279 ( .A1(n3806), .A2(n4462), .ZN(n4393) );
  NAND2_X1 U4280 ( .A1(n3807), .A2(n3472), .ZN(n3861) );
  NAND2_X1 U4281 ( .A1(n4519), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4282 ( .A1(n3528), .A2(n4403), .ZN(n3808) );
  OAI211_X1 U4283 ( .C1(n3809), .C2(n4836), .A(STATE2_REG_0__SCAN_IN), .B(
        n3808), .ZN(n3810) );
  INV_X1 U4284 ( .A(n3810), .ZN(n3811) );
  NAND2_X1 U4285 ( .A1(n3812), .A2(n3811), .ZN(n3862) );
  OAI21_X1 U4286 ( .B1(n3859), .B2(n3861), .A(n3862), .ZN(n3813) );
  INV_X1 U4287 ( .A(n3814), .ZN(n3816) );
  NOR2_X1 U4288 ( .A1(n3816), .A2(n3815), .ZN(n3817) );
  AOI21_X2 U4289 ( .B1(n3853), .B2(n3852), .A(n3817), .ZN(n3846) );
  INV_X1 U4290 ( .A(n3846), .ZN(n3844) );
  INV_X1 U4291 ( .A(n3818), .ZN(n3820) );
  NAND2_X1 U4292 ( .A1(n3820), .A2(n3819), .ZN(n3822) );
  INV_X1 U4293 ( .A(n6766), .ZN(n3881) );
  NAND2_X1 U4294 ( .A1(n3881), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U4295 ( .A1(n6766), .A2(n4482), .ZN(n3825) );
  INV_X1 U4296 ( .A(n4537), .ZN(n3884) );
  AOI22_X1 U4297 ( .A1(n4993), .A2(n3884), .B1(n3883), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4298 ( .A1(n4201), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4299 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n4366), .B1(n4374), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4300 ( .A1(n3437), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4301 ( .A1(n3712), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4302 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3841)
         );
  AOI22_X1 U4303 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n4372), .B1(n4371), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4304 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n4350), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4305 ( .A1(n4345), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4306 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n3795), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3836) );
  NAND4_X1 U4307 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3840)
         );
  AOI22_X1 U4308 ( .A1(n4529), .A2(n4408), .B1(n4519), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3842) );
  INV_X1 U4309 ( .A(n3845), .ZN(n3843) );
  NAND2_X2 U4310 ( .A1(n3846), .A2(n3845), .ZN(n3901) );
  INV_X1 U4311 ( .A(n4107), .ZN(n3848) );
  NAND2_X1 U4312 ( .A1(n6797), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4071) );
  INV_X1 U4313 ( .A(n3555), .ZN(n4599) );
  OR2_X1 U4314 ( .A1(n4599), .A2(n6797), .ZN(n3923) );
  OAI21_X1 U4315 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3902), .ZN(n6177) );
  AOI22_X1 U4316 ( .A1(n4553), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5020), 
        .B2(n6177), .ZN(n3851) );
  INV_X1 U4317 ( .A(n3722), .ZN(n5561) );
  NAND2_X1 U4318 ( .A1(n3927), .A2(EAX_REG_2__SCAN_IN), .ZN(n3850) );
  OAI211_X1 U4319 ( .C1(n3923), .C2(n3824), .A(n3851), .B(n3850), .ZN(n3873)
         );
  NAND2_X1 U4320 ( .A1(n3872), .A2(n3873), .ZN(n3871) );
  XNOR2_X1 U4321 ( .A(n3853), .B(n3852), .ZN(n4395) );
  NAND2_X1 U4322 ( .A1(n4395), .A2(n3848), .ZN(n3858) );
  NAND2_X1 U4323 ( .A1(n6797), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3855)
         );
  NAND2_X1 U4324 ( .A1(n3927), .A2(EAX_REG_1__SCAN_IN), .ZN(n3854) );
  OAI211_X1 U4325 ( .C1(n3923), .C2(n3567), .A(n3855), .B(n3854), .ZN(n3856)
         );
  INV_X1 U4326 ( .A(n3856), .ZN(n3857) );
  NAND2_X1 U4327 ( .A1(n3858), .A2(n3857), .ZN(n4856) );
  INV_X1 U4328 ( .A(n3859), .ZN(n3860) );
  NAND2_X1 U4329 ( .A1(n3862), .A2(n3860), .ZN(n3863) );
  AOI21_X1 U4330 ( .B1(n6780), .B2(n3480), .A(n6797), .ZN(n4844) );
  OAI21_X1 U4331 ( .B1(n3864), .B2(n3865), .A(n3819), .ZN(n6713) );
  OR2_X1 U4332 ( .A1(n6713), .A2(n4107), .ZN(n3870) );
  NAND2_X1 U4333 ( .A1(n6797), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3867)
         );
  NAND2_X1 U4334 ( .A1(n3927), .A2(EAX_REG_0__SCAN_IN), .ZN(n3866) );
  OAI211_X1 U4335 ( .C1(n3923), .C2(n3566), .A(n3867), .B(n3866), .ZN(n3868)
         );
  INV_X1 U4336 ( .A(n3868), .ZN(n3869) );
  NAND2_X1 U4337 ( .A1(n3870), .A2(n3869), .ZN(n4845) );
  MUX2_X1 U4338 ( .A(n5020), .B(n4844), .S(n4845), .Z(n4855) );
  NAND2_X1 U4339 ( .A1(n4856), .A2(n4855), .ZN(n4936) );
  NAND2_X1 U4340 ( .A1(n3871), .A2(n4936), .ZN(n3876) );
  INV_X1 U4341 ( .A(n3872), .ZN(n3875) );
  INV_X1 U4342 ( .A(n3873), .ZN(n3874) );
  NAND2_X1 U4343 ( .A1(n3876), .A2(n4935), .ZN(n4864) );
  INV_X1 U4344 ( .A(n4864), .ZN(n3908) );
  INV_X1 U4345 ( .A(n3901), .ZN(n3899) );
  NAND2_X1 U4346 ( .A1(n4943), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3882) );
  NOR2_X1 U4347 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4482), .ZN(n6753)
         );
  NAND2_X1 U4348 ( .A1(n3881), .A2(n6753), .ZN(n6714) );
  NAND2_X1 U4349 ( .A1(n3882), .A2(n6714), .ZN(n6750) );
  AOI22_X1 U4350 ( .A1(n6750), .A2(n3884), .B1(n3883), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3885) );
  NAND2_X1 U4351 ( .A1(n4941), .A2(n6594), .ZN(n3898) );
  AOI22_X1 U4352 ( .A1(n4366), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4353 ( .A1(n3437), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4354 ( .A1(n4350), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4355 ( .A1(n3795), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4356 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3896)
         );
  AOI22_X1 U4357 ( .A1(n4372), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4358 ( .A1(n4326), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3712), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4359 ( .A1(n4345), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3892) );
  INV_X1 U4360 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U4361 ( .A1(n4201), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4362 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3895)
         );
  AOI22_X1 U4363 ( .A1(n4529), .A2(n4421), .B1(n4519), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3897) );
  NAND2_X2 U4364 ( .A1(n3899), .A2(n3900), .ZN(n3928) );
  NAND2_X1 U4365 ( .A1(n3901), .A2(n5126), .ZN(n6725) );
  OAI21_X1 U4366 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3903), .A(n3945), 
        .ZN(n5037) );
  AOI22_X1 U4367 ( .A1(n5020), .A2(n5037), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U4368 ( .A1(n3927), .A2(EAX_REG_3__SCAN_IN), .ZN(n3904) );
  OAI211_X1 U4369 ( .C1(n3923), .C2(n3880), .A(n3905), .B(n3904), .ZN(n3906)
         );
  AOI21_X1 U4370 ( .B1(n5127), .B2(n3848), .A(n3906), .ZN(n4865) );
  NAND2_X1 U4371 ( .A1(n3908), .A2(n3907), .ZN(n4863) );
  AOI22_X1 U4372 ( .A1(n4201), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4373 ( .A1(n4374), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4374 ( .A1(n3437), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4375 ( .A1(n4350), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4376 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3918)
         );
  AOI22_X1 U4377 ( .A1(n4372), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4378 ( .A1(n3712), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4379 ( .A1(n4045), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3914) );
  INV_X1 U4380 ( .A(n3764), .ZN(n4326) );
  AOI22_X1 U4381 ( .A1(n4326), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4382 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3917)
         );
  NAND2_X1 U4383 ( .A1(n4529), .A2(n4435), .ZN(n3920) );
  NAND2_X1 U4384 ( .A1(n4519), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3919) );
  NAND2_X1 U4385 ( .A1(n6797), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3922)
         );
  NAND2_X1 U4386 ( .A1(n3927), .A2(EAX_REG_4__SCAN_IN), .ZN(n3921) );
  OAI211_X1 U4387 ( .C1(n3923), .C2(n4517), .A(n3922), .B(n3921), .ZN(n3925)
         );
  INV_X1 U4388 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3924) );
  XNOR2_X1 U4389 ( .A(n3924), .B(n3945), .ZN(n6360) );
  MUX2_X1 U4390 ( .A(n3925), .B(n6360), .S(n5020), .Z(n3926) );
  AOI21_X1 U4391 ( .B1(n4426), .B2(n3848), .A(n3926), .ZN(n4931) );
  INV_X1 U4392 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U4393 ( .A1(n4366), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4394 ( .A1(n3437), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4395 ( .A1(n4350), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4396 ( .A1(n3795), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4397 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3940)
         );
  AOI22_X1 U4398 ( .A1(n4372), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4399 ( .A1(n4326), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3712), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4400 ( .A1(n4345), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3936) );
  INV_X1 U4401 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n7037) );
  AOI22_X1 U4402 ( .A1(n4201), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3935) );
  NAND4_X1 U4403 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3939)
         );
  NAND2_X1 U4404 ( .A1(n4529), .A2(n4452), .ZN(n3942) );
  NAND2_X1 U4405 ( .A1(n4519), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U4406 ( .A1(n3942), .A2(n3941), .ZN(n3950) );
  XNOR2_X1 U4407 ( .A(n3949), .B(n3950), .ZN(n4434) );
  NAND2_X1 U4408 ( .A1(n4434), .A2(n3848), .ZN(n3948) );
  INV_X1 U4409 ( .A(n3945), .ZN(n3943) );
  AOI21_X1 U4410 ( .B1(n3943), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4411 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3944) );
  OR2_X1 U4412 ( .A1(n3946), .A2(n3966), .ZN(n6376) );
  AOI22_X1 U4413 ( .A1(n6376), .A2(n4341), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3947) );
  OAI211_X1 U4414 ( .C1(n4361), .C2(n4788), .A(n3948), .B(n3947), .ZN(n4911)
         );
  NAND2_X1 U4415 ( .A1(n4912), .A2(n4911), .ZN(n4910) );
  INV_X1 U4416 ( .A(n4910), .ZN(n3973) );
  INV_X1 U4417 ( .A(n3975), .ZN(n3965) );
  AOI22_X1 U4418 ( .A1(n3795), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4419 ( .A1(n4350), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4420 ( .A1(n4201), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4421 ( .A1(n4345), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3712), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3952) );
  NAND4_X1 U4422 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3961)
         );
  AOI22_X1 U4423 ( .A1(n4372), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4424 ( .A1(n4366), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4425 ( .A1(n4326), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4426 ( .A1(n3437), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4427 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3960)
         );
  NAND2_X1 U4428 ( .A1(n4529), .A2(n4451), .ZN(n3963) );
  NAND2_X1 U4429 ( .A1(n4519), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3962) );
  NAND2_X1 U4430 ( .A1(n3963), .A2(n3962), .ZN(n3974) );
  INV_X1 U4431 ( .A(n3974), .ZN(n3964) );
  NAND2_X1 U4432 ( .A1(n3965), .A2(n3964), .ZN(n4443) );
  NOR2_X1 U4433 ( .A1(n3966), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3967)
         );
  OR2_X1 U4434 ( .A1(n3977), .A2(n3967), .ZN(n6387) );
  INV_X1 U4435 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3969) );
  INV_X1 U4436 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3968) );
  OAI22_X1 U4437 ( .A1(n4361), .A2(n3969), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3968), .ZN(n3970) );
  MUX2_X1 U4438 ( .A(n6387), .B(n3970), .S(n4301), .Z(n3971) );
  AOI22_X1 U4439 ( .A1(n4529), .A2(n4462), .B1(n4519), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3976) );
  XNOR2_X1 U4440 ( .A(n4444), .B(n3976), .ZN(n4450) );
  INV_X1 U4441 ( .A(n4450), .ZN(n3981) );
  INV_X1 U4442 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4781) );
  OR2_X1 U4443 ( .A1(n3977), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3978) );
  NAND2_X1 U4444 ( .A1(n3978), .A2(n3997), .ZN(n6400) );
  AOI22_X1 U4445 ( .A1(n6400), .A2(n4341), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3979) );
  OAI21_X1 U4446 ( .B1(n4361), .B2(n4781), .A(n3979), .ZN(n3980) );
  AOI22_X1 U4447 ( .A1(n4372), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4448 ( .A1(n4366), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4449 ( .A1(n4350), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4450 ( .A1(n4345), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4451 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3991)
         );
  AOI22_X1 U4452 ( .A1(n3437), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4453 ( .A1(n4326), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4454 ( .A1(n3795), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4455 ( .A1(n4201), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3986) );
  NAND4_X1 U4456 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3990)
         );
  NOR2_X1 U4457 ( .A1(n3991), .A2(n3990), .ZN(n3995) );
  INV_X1 U4458 ( .A(n3997), .ZN(n3992) );
  XNOR2_X1 U4459 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3992), .ZN(n6408) );
  AOI22_X1 U4460 ( .A1(n5020), .A2(n6408), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4461 ( .A1(n3927), .A2(EAX_REG_8__SCAN_IN), .ZN(n3993) );
  OAI211_X1 U4462 ( .C1(n4107), .C2(n3995), .A(n3994), .B(n3993), .ZN(n5160)
         );
  XOR2_X1 U4463 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4011), .Z(n6418) );
  AOI22_X1 U4464 ( .A1(n3927), .A2(EAX_REG_9__SCAN_IN), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4465 ( .A1(n3437), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4466 ( .A1(n4345), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4467 ( .A1(n4046), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4468 ( .A1(n3795), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4469 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4008)
         );
  AOI22_X1 U4470 ( .A1(n4201), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4326), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4471 ( .A1(n4372), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4472 ( .A1(n4045), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4473 ( .A1(n4374), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4003) );
  NAND4_X1 U4474 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(n4007)
         );
  OAI21_X1 U4475 ( .B1(n4008), .B2(n4007), .A(n3848), .ZN(n4009) );
  OAI211_X1 U4476 ( .C1(n6418), .C2(n4301), .A(n4010), .B(n4009), .ZN(n5146)
         );
  XNOR2_X1 U4477 ( .A(n4025), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6426)
         );
  NAND2_X1 U4478 ( .A1(n6426), .A2(n4341), .ZN(n4024) );
  AOI22_X1 U4479 ( .A1(n3927), .A2(EAX_REG_10__SCAN_IN), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4480 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n4371), .B1(n4366), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4481 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n4350), .B1(n4045), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4482 ( .A1(n4201), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4483 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n3437), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U4484 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4021)
         );
  AOI22_X1 U4485 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(n4374), .B1(n4372), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4486 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n3459), .B1(n3795), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4487 ( .A1(n4326), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4488 ( .A1(n4345), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4489 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4020)
         );
  OAI21_X1 U4490 ( .B1(n4021), .B2(n4020), .A(n3848), .ZN(n4022) );
  XOR2_X1 U4491 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4038), .Z(n6445) );
  AOI22_X1 U4492 ( .A1(n3927), .A2(EAX_REG_11__SCAN_IN), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4493 ( .A1(n4345), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4494 ( .A1(n4045), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4495 ( .A1(n4371), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4496 ( .A1(n4326), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U4497 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4035)
         );
  AOI22_X1 U4498 ( .A1(n4201), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4499 ( .A1(n4372), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4500 ( .A1(n3437), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4501 ( .A1(n4350), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4502 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4034)
         );
  OAI21_X1 U4503 ( .B1(n4035), .B2(n4034), .A(n3848), .ZN(n4036) );
  OAI211_X1 U4504 ( .C1(n6445), .C2(n4301), .A(n4037), .B(n4036), .ZN(n5211)
         );
  XNOR2_X1 U4505 ( .A(n4068), .B(n5230), .ZN(n5258) );
  AOI21_X1 U4506 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5230), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4040) );
  AND2_X1 U4507 ( .A1(n3927), .A2(EAX_REG_12__SCAN_IN), .ZN(n4039) );
  OAI22_X1 U4508 ( .A1(n5258), .A2(n4301), .B1(n4040), .B2(n4039), .ZN(n4054)
         );
  AOI22_X1 U4509 ( .A1(n4345), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4510 ( .A1(n3437), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4511 ( .A1(n4366), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4512 ( .A1(n4201), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U4513 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4052)
         );
  AOI22_X1 U4514 ( .A1(n4045), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4515 ( .A1(n4326), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4516 ( .A1(n3795), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4517 ( .A1(n4374), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4047) );
  NAND4_X1 U4518 ( .A1(n4050), .A2(n4049), .A3(n4048), .A4(n4047), .ZN(n4051)
         );
  OAI21_X1 U4519 ( .B1(n4052), .B2(n4051), .A(n3848), .ZN(n4053) );
  AOI22_X1 U4520 ( .A1(n4201), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4521 ( .A1(n4366), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4522 ( .A1(n4350), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U4523 ( .A1(n4045), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U4524 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4064)
         );
  AOI22_X1 U4525 ( .A1(n3437), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4526 ( .A1(n4345), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4527 ( .A1(n4374), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4528 ( .A1(n4326), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U4529 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  OR2_X1 U4530 ( .A1(n4064), .A2(n4063), .ZN(n4065) );
  NAND2_X1 U4531 ( .A1(n3848), .A2(n4065), .ZN(n4066) );
  NAND2_X1 U4532 ( .A1(n4076), .A2(n4067), .ZN(n5290) );
  INV_X1 U4533 ( .A(n5290), .ZN(n4075) );
  INV_X1 U4534 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4072) );
  OAI21_X1 U4535 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4069), .A(n4093), 
        .ZN(n6462) );
  NAND2_X1 U4536 ( .A1(n6462), .A2(n4341), .ZN(n4070) );
  OAI21_X1 U4537 ( .B1(n4072), .B2(n4071), .A(n4070), .ZN(n4073) );
  AOI21_X1 U4538 ( .B1(n3927), .B2(EAX_REG_13__SCAN_IN), .A(n4073), .ZN(n5291)
         );
  NAND2_X1 U4539 ( .A1(n4075), .A2(n4074), .ZN(n5293) );
  XOR2_X1 U4540 ( .A(n4092), .B(n4093), .Z(n6468) );
  NAND2_X1 U4541 ( .A1(n6468), .A2(n5020), .ZN(n4079) );
  INV_X1 U4542 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4799) );
  OAI21_X1 U4543 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6817), .A(n6797), 
        .ZN(n4077) );
  OAI21_X1 U4544 ( .B1(n4361), .B2(n4799), .A(n4077), .ZN(n4078) );
  NAND2_X1 U4545 ( .A1(n4079), .A2(n4078), .ZN(n4091) );
  AOI22_X1 U4546 ( .A1(n4372), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4547 ( .A1(n4350), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U4548 ( .A1(n4345), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U4549 ( .A1(n3835), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U4550 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4089)
         );
  AOI22_X1 U4551 ( .A1(n4374), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4552 ( .A1(n3437), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U4553 ( .A1(n4201), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U4554 ( .A1(n4326), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4084) );
  NAND4_X1 U4555 ( .A1(n4087), .A2(n4086), .A3(n4085), .A4(n4084), .ZN(n4088)
         );
  OAI21_X1 U4556 ( .B1(n4089), .B2(n4088), .A(n3848), .ZN(n4090) );
  NAND2_X1 U4557 ( .A1(n4091), .A2(n4090), .ZN(n5301) );
  XNOR2_X1 U4558 ( .A(n4110), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5698)
         );
  AOI22_X1 U4559 ( .A1(n4372), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U4560 ( .A1(n4371), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U4561 ( .A1(n3437), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U4562 ( .A1(n4345), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4094) );
  NAND4_X1 U4563 ( .A1(n4097), .A2(n4096), .A3(n4095), .A4(n4094), .ZN(n4103)
         );
  AOI22_X1 U4564 ( .A1(n4350), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U4565 ( .A1(n4326), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U4566 ( .A1(n4366), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U4567 ( .A1(n4201), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4098) );
  NAND4_X1 U4568 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4098), .ZN(n4102)
         );
  NOR2_X1 U4569 ( .A1(n4103), .A2(n4102), .ZN(n4106) );
  NAND2_X1 U4570 ( .A1(n3927), .A2(EAX_REG_15__SCAN_IN), .ZN(n4105) );
  NAND2_X1 U4571 ( .A1(n4553), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4104)
         );
  OAI211_X1 U4572 ( .C1(n4107), .C2(n4106), .A(n4105), .B(n4104), .ZN(n4108)
         );
  AOI21_X1 U4573 ( .B1(n5698), .B2(n4341), .A(n4108), .ZN(n5303) );
  XOR2_X1 U4574 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4124), .Z(n6481) );
  INV_X1 U4575 ( .A(n6481), .ZN(n5693) );
  AOI22_X1 U4576 ( .A1(n4326), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U4577 ( .A1(n4372), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4578 ( .A1(n3835), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4579 ( .A1(n4201), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U4580 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4120)
         );
  AOI22_X1 U4581 ( .A1(n4350), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U4582 ( .A1(n3998), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U4583 ( .A1(n3437), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U4584 ( .A1(n4371), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4115) );
  NAND4_X1 U4585 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4119)
         );
  NOR2_X1 U4586 ( .A1(n4120), .A2(n4119), .ZN(n4122) );
  AOI22_X1 U4587 ( .A1(n3927), .A2(EAX_REG_16__SCAN_IN), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4121) );
  OAI21_X1 U4588 ( .B1(n4386), .B2(n4122), .A(n4121), .ZN(n4123) );
  AOI21_X1 U4589 ( .B1(n5693), .B2(n4341), .A(n4123), .ZN(n5549) );
  XNOR2_X1 U4590 ( .A(n4152), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6488)
         );
  AOI21_X1 U4591 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5685), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4125) );
  AOI21_X1 U4592 ( .B1(n3927), .B2(EAX_REG_17__SCAN_IN), .A(n4125), .ZN(n4137)
         );
  AOI22_X1 U4593 ( .A1(n3436), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U4594 ( .A1(n3998), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U4595 ( .A1(n4350), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U4596 ( .A1(n4201), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4126) );
  NAND4_X1 U4597 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4135)
         );
  AOI22_X1 U4598 ( .A1(n4372), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U4599 ( .A1(n3437), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U4600 ( .A1(n4045), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U4601 ( .A1(n4326), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U4602 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4134)
         );
  OAI21_X1 U4603 ( .B1(n4135), .B2(n4134), .A(n4363), .ZN(n4136) );
  AOI22_X1 U4604 ( .A1(n6488), .A2(n4341), .B1(n4137), .B2(n4136), .ZN(n5542)
         );
  INV_X1 U4605 ( .A(n5533), .ZN(n4157) );
  AOI22_X1 U4606 ( .A1(n4372), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U4607 ( .A1(n4366), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U4608 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n3459), .B1(n4045), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U4609 ( .A1(n4307), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4138) );
  NAND4_X1 U4610 ( .A1(n4141), .A2(n4140), .A3(n4139), .A4(n4138), .ZN(n4147)
         );
  AOI22_X1 U4611 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n3437), .B1(n4350), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U4612 ( .A1(n4201), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U4613 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n3795), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U4614 ( .A1(n4345), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4142) );
  NAND4_X1 U4615 ( .A1(n4145), .A2(n4144), .A3(n4143), .A4(n4142), .ZN(n4146)
         );
  NOR2_X1 U4616 ( .A1(n4147), .A2(n4146), .ZN(n4151) );
  OAI21_X1 U4617 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6817), .A(n6797), 
        .ZN(n4148) );
  INV_X1 U4618 ( .A(n4148), .ZN(n4149) );
  AOI21_X1 U4619 ( .B1(n3927), .B2(EAX_REG_18__SCAN_IN), .A(n4149), .ZN(n4150)
         );
  OAI21_X1 U4620 ( .B1(n4386), .B2(n4151), .A(n4150), .ZN(n4155) );
  OAI21_X1 U4621 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4153), .A(n4171), 
        .ZN(n6502) );
  OR2_X1 U4622 ( .A1(n4301), .A2(n6502), .ZN(n4154) );
  NAND2_X1 U4623 ( .A1(n4155), .A2(n4154), .ZN(n5534) );
  XNOR2_X1 U4624 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4171), .ZN(n5674)
         );
  AOI22_X1 U4625 ( .A1(n4372), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U4626 ( .A1(n4371), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U4627 ( .A1(n4350), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U4628 ( .A1(n4345), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4158) );
  NAND4_X1 U4629 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4167)
         );
  AOI22_X1 U4630 ( .A1(n3437), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4631 ( .A1(n3626), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4632 ( .A1(n4366), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U4633 ( .A1(n4201), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4162) );
  NAND4_X1 U4634 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4166)
         );
  OR2_X1 U4635 ( .A1(n4167), .A2(n4166), .ZN(n4169) );
  INV_X1 U4636 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4792) );
  INV_X1 U4637 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5672) );
  OAI22_X1 U4638 ( .A1(n4361), .A2(n4792), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5672), .ZN(n4168) );
  AOI21_X1 U4639 ( .B1(n4363), .B2(n4169), .A(n4168), .ZN(n4170) );
  MUX2_X1 U4640 ( .A(n5674), .B(n4170), .S(n4301), .Z(n5483) );
  OAI21_X1 U4641 ( .B1(n4173), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4218), 
        .ZN(n6516) );
  AOI22_X1 U4642 ( .A1(n3626), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U4643 ( .A1(n4372), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U4644 ( .A1(n4350), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U4645 ( .A1(n4366), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4174) );
  NAND4_X1 U4646 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(n4183)
         );
  AOI22_X1 U4647 ( .A1(n3437), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U4648 ( .A1(n3998), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U4649 ( .A1(n3795), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U4650 ( .A1(n4201), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4178) );
  NAND4_X1 U4651 ( .A1(n4181), .A2(n4180), .A3(n4179), .A4(n4178), .ZN(n4182)
         );
  NOR2_X1 U4652 ( .A1(n4183), .A2(n4182), .ZN(n4185) );
  AOI22_X1 U4653 ( .A1(n3927), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6797), .ZN(n4184) );
  OAI21_X1 U4654 ( .B1(n4386), .B2(n4185), .A(n4184), .ZN(n4186) );
  MUX2_X1 U4655 ( .A(n6516), .B(n4186), .S(n4301), .Z(n5528) );
  XNOR2_X1 U4656 ( .A(n4218), .B(n4217), .ZN(n5657) );
  AOI22_X1 U4657 ( .A1(n4201), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4326), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U4658 ( .A1(n4372), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U4659 ( .A1(n4350), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U4660 ( .A1(n4345), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4187) );
  NAND4_X1 U4661 ( .A1(n4190), .A2(n4189), .A3(n4188), .A4(n4187), .ZN(n4196)
         );
  AOI22_X1 U4662 ( .A1(n4374), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U4663 ( .A1(n3437), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U4664 ( .A1(n4373), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U4665 ( .A1(n3835), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4191) );
  NAND4_X1 U4666 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4195)
         );
  NOR2_X1 U4667 ( .A1(n4196), .A2(n4195), .ZN(n4199) );
  NOR2_X1 U4668 ( .A1(n4217), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4197) );
  AOI21_X1 U4669 ( .B1(n3927), .B2(EAX_REG_21__SCAN_IN), .A(n4197), .ZN(n4198)
         );
  OAI21_X1 U4670 ( .B1(n4386), .B2(n4199), .A(n4198), .ZN(n4200) );
  MUX2_X1 U4671 ( .A(n5657), .B(n4200), .S(n4301), .Z(n5470) );
  AOI22_X1 U4672 ( .A1(n4307), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U4673 ( .A1(n3437), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U4674 ( .A1(n4045), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4675 ( .A1(n4201), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4202) );
  NAND4_X1 U4676 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(n4212)
         );
  AOI22_X1 U4677 ( .A1(n4372), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U4678 ( .A1(n3436), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4679 ( .A1(n4046), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U4680 ( .A1(n4350), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4207) );
  NAND4_X1 U4681 ( .A1(n4210), .A2(n4209), .A3(n4208), .A4(n4207), .ZN(n4211)
         );
  NOR2_X1 U4682 ( .A1(n4212), .A2(n4211), .ZN(n4216) );
  OAI21_X1 U4683 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6817), .A(n6797), 
        .ZN(n4213) );
  INV_X1 U4684 ( .A(n4213), .ZN(n4214) );
  AOI21_X1 U4685 ( .B1(n3927), .B2(EAX_REG_22__SCAN_IN), .A(n4214), .ZN(n4215)
         );
  OAI21_X1 U4686 ( .B1(n4386), .B2(n4216), .A(n4215), .ZN(n4222) );
  NOR2_X1 U4687 ( .A1(n4219), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4220)
         );
  OR2_X1 U4688 ( .A1(n4259), .A2(n4220), .ZN(n5650) );
  NAND2_X1 U4689 ( .A1(n6529), .A2(n4341), .ZN(n4221) );
  NAND2_X1 U4690 ( .A1(n4222), .A2(n4221), .ZN(n5514) );
  AOI22_X1 U4691 ( .A1(n4374), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4226) );
  AOI22_X1 U4692 ( .A1(n4045), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U4693 ( .A1(n3711), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U4694 ( .A1(n4326), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4223) );
  NAND4_X1 U4695 ( .A1(n4226), .A2(n4225), .A3(n4224), .A4(n4223), .ZN(n4232)
         );
  AOI22_X1 U4696 ( .A1(n3437), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U4697 ( .A1(n4372), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U4698 ( .A1(n4345), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U4699 ( .A1(n3795), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4227) );
  NAND4_X1 U4700 ( .A1(n4230), .A2(n4229), .A3(n4228), .A4(n4227), .ZN(n4231)
         );
  NOR2_X1 U4701 ( .A1(n4232), .A2(n4231), .ZN(n4246) );
  AOI22_X1 U4702 ( .A1(n3711), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4326), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U4703 ( .A1(n3437), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4704 ( .A1(n4045), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U4705 ( .A1(n4046), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4233) );
  NAND4_X1 U4706 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), .ZN(n4242)
         );
  AOI22_X1 U4707 ( .A1(n4372), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U4708 ( .A1(n4366), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U4709 ( .A1(n4345), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U4710 ( .A1(n4350), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4237) );
  NAND4_X1 U4711 ( .A1(n4240), .A2(n4239), .A3(n4238), .A4(n4237), .ZN(n4241)
         );
  NOR2_X1 U4712 ( .A1(n4242), .A2(n4241), .ZN(n4247) );
  XOR2_X1 U4713 ( .A(n4246), .B(n4247), .Z(n4244) );
  INV_X1 U4714 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4784) );
  INV_X1 U4715 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5641) );
  OAI22_X1 U4716 ( .A1(n4361), .A2(n4784), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5641), .ZN(n4243) );
  AOI21_X1 U4717 ( .B1(n4363), .B2(n4244), .A(n4243), .ZN(n4245) );
  XNOR2_X1 U4718 ( .A(n4259), .B(n5641), .ZN(n5643) );
  MUX2_X1 U4719 ( .A(n4245), .B(n5643), .S(n5020), .Z(n5454) );
  OR2_X1 U4720 ( .A1(n4247), .A2(n4246), .ZN(n4276) );
  AOI22_X1 U4721 ( .A1(n3437), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4722 ( .A1(n3711), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U4723 ( .A1(n4366), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U4724 ( .A1(n4326), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4248) );
  NAND4_X1 U4725 ( .A1(n4251), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4257)
         );
  AOI22_X1 U4726 ( .A1(n4372), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U4727 ( .A1(n4350), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4254) );
  INV_X1 U4728 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6879) );
  AOI22_X1 U4729 ( .A1(n4045), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U4730 ( .A1(n3459), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4252) );
  NAND4_X1 U4731 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4256)
         );
  NOR2_X1 U4732 ( .A1(n4257), .A2(n4256), .ZN(n4275) );
  INV_X1 U4733 ( .A(n4275), .ZN(n4258) );
  XNOR2_X1 U4734 ( .A(n4276), .B(n4258), .ZN(n4263) );
  INV_X1 U4735 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4790) );
  XNOR2_X1 U4736 ( .A(n4279), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5635)
         );
  NAND2_X1 U4737 ( .A1(n5635), .A2(n5020), .ZN(n4261) );
  NAND2_X1 U4738 ( .A1(n4553), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4260)
         );
  OAI211_X1 U4739 ( .C1(n4361), .C2(n4790), .A(n4261), .B(n4260), .ZN(n4262)
         );
  AOI21_X1 U4740 ( .B1(n4263), .B2(n4363), .A(n4262), .ZN(n5445) );
  AOI22_X1 U4741 ( .A1(n4374), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U4742 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n3437), .B1(n3795), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U4743 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4350), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U4744 ( .A1(n4373), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4265) );
  NAND4_X1 U4745 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(n4274)
         );
  AOI22_X1 U4746 ( .A1(n3711), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4326), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U4747 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n4372), .B1(n3436), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U4748 ( .A1(n4345), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U4749 ( .A1(n4045), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4269) );
  NAND4_X1 U4750 ( .A1(n4272), .A2(n4271), .A3(n4270), .A4(n4269), .ZN(n4273)
         );
  NOR2_X1 U4751 ( .A1(n4274), .A2(n4273), .ZN(n4288) );
  OR2_X1 U4752 ( .A1(n4276), .A2(n4275), .ZN(n4287) );
  XOR2_X1 U4753 ( .A(n4288), .B(n4287), .Z(n4278) );
  INV_X1 U4754 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4797) );
  INV_X1 U4755 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5623) );
  OAI22_X1 U4756 ( .A1(n4361), .A2(n4797), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5623), .ZN(n4277) );
  AOI21_X1 U4757 ( .B1(n4278), .B2(n4363), .A(n4277), .ZN(n4280) );
  XNOR2_X1 U4758 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4282), .ZN(n5627)
         );
  MUX2_X1 U4759 ( .A(n4280), .B(n5627), .S(n5020), .Z(n4281) );
  INV_X1 U4760 ( .A(n4282), .ZN(n4283) );
  INV_X1 U4761 ( .A(n4284), .ZN(n4285) );
  INV_X1 U4762 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U4763 ( .A1(n4285), .A2(n5419), .ZN(n4286) );
  NAND2_X1 U4764 ( .A1(n4337), .A2(n4286), .ZN(n5616) );
  NOR2_X1 U4765 ( .A1(n4288), .A2(n4287), .ZN(n4315) );
  AOI22_X1 U4766 ( .A1(n4366), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U4767 ( .A1(n3437), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4291) );
  AOI22_X1 U4768 ( .A1(n4350), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4290) );
  AOI22_X1 U4769 ( .A1(n3795), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4289) );
  NAND4_X1 U4770 ( .A1(n4292), .A2(n4291), .A3(n4290), .A4(n4289), .ZN(n4298)
         );
  AOI22_X1 U4771 ( .A1(n4372), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U4772 ( .A1(n4326), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4773 ( .A1(n4345), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U4774 ( .A1(n4201), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4293) );
  NAND4_X1 U4775 ( .A1(n4296), .A2(n4295), .A3(n4294), .A4(n4293), .ZN(n4297)
         );
  OR2_X1 U4776 ( .A1(n4298), .A2(n4297), .ZN(n4314) );
  XNOR2_X1 U4777 ( .A(n4315), .B(n4314), .ZN(n4300) );
  AOI22_X1 U4778 ( .A1(n3927), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6797), .ZN(n4299) );
  OAI21_X1 U4779 ( .B1(n4300), .B2(n4386), .A(n4299), .ZN(n4302) );
  MUX2_X1 U4780 ( .A(n5616), .B(n4302), .S(n4301), .Z(n5414) );
  AOI22_X1 U4781 ( .A1(n3437), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4306) );
  AOI22_X1 U4782 ( .A1(n4374), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U4783 ( .A1(n4345), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U4784 ( .A1(n3795), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4303) );
  NAND4_X1 U4785 ( .A1(n4306), .A2(n4305), .A3(n4304), .A4(n4303), .ZN(n4313)
         );
  AOI22_X1 U4786 ( .A1(n4201), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4311) );
  AOI22_X1 U4787 ( .A1(n4372), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U4788 ( .A1(n4045), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4309) );
  AOI22_X1 U4789 ( .A1(n4046), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4308) );
  NAND4_X1 U4790 ( .A1(n4311), .A2(n4310), .A3(n4309), .A4(n4308), .ZN(n4312)
         );
  NOR2_X1 U4791 ( .A1(n4313), .A2(n4312), .ZN(n4321) );
  NAND2_X1 U4792 ( .A1(n4315), .A2(n4314), .ZN(n4320) );
  XOR2_X1 U4793 ( .A(n4321), .B(n4320), .Z(n4317) );
  INV_X1 U4794 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4795) );
  INV_X1 U4795 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5328) );
  OAI22_X1 U4796 ( .A1(n4361), .A2(n4795), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5328), .ZN(n4316) );
  AOI21_X1 U4797 ( .B1(n4317), .B2(n4363), .A(n4316), .ZN(n4318) );
  XNOR2_X1 U4798 ( .A(n4337), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5409)
         );
  MUX2_X1 U4799 ( .A(n4318), .B(n5409), .S(n5020), .Z(n4319) );
  NOR2_X1 U4800 ( .A1(n4321), .A2(n4320), .ZN(n4359) );
  AOI22_X1 U4801 ( .A1(n3436), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U4802 ( .A1(n3437), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U4803 ( .A1(n4350), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U4804 ( .A1(n3795), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4322) );
  NAND4_X1 U4805 ( .A1(n4325), .A2(n4324), .A3(n4323), .A4(n4322), .ZN(n4332)
         );
  AOI22_X1 U4806 ( .A1(n4372), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U4807 ( .A1(n4326), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U4808 ( .A1(n4345), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U4809 ( .A1(n3711), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4327) );
  NAND4_X1 U4810 ( .A1(n4330), .A2(n4329), .A3(n4328), .A4(n4327), .ZN(n4331)
         );
  OR2_X1 U4811 ( .A1(n4332), .A2(n4331), .ZN(n4358) );
  INV_X1 U4812 ( .A(n4358), .ZN(n4333) );
  XNOR2_X1 U4813 ( .A(n4359), .B(n4333), .ZN(n4336) );
  INV_X1 U4814 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4334) );
  INV_X1 U4815 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5605) );
  OAI22_X1 U4816 ( .A1(n4361), .A2(n4334), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5605), .ZN(n4335) );
  AOI21_X1 U4817 ( .B1(n4336), .B2(n4363), .A(n4335), .ZN(n4342) );
  NAND2_X1 U4818 ( .A1(n4338), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4388)
         );
  INV_X1 U4819 ( .A(n4338), .ZN(n4339) );
  NAND2_X1 U4820 ( .A1(n4339), .A2(n5605), .ZN(n4340) );
  AND2_X1 U4821 ( .A1(n4388), .A2(n4340), .ZN(n5607) );
  MUX2_X1 U4822 ( .A(n4342), .B(n5607), .S(n4341), .Z(n5397) );
  AOI22_X1 U4823 ( .A1(n3711), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4326), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4824 ( .A1(n3436), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4825 ( .A1(n4045), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U4826 ( .A1(n4345), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4346) );
  NAND4_X1 U4827 ( .A1(n4349), .A2(n4348), .A3(n4347), .A4(n4346), .ZN(n4357)
         );
  AOI22_X1 U4828 ( .A1(n3437), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4355) );
  AOI22_X1 U4829 ( .A1(n4372), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U4830 ( .A1(n4046), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3765), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U4831 ( .A1(n3835), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4352) );
  NAND4_X1 U4832 ( .A1(n4355), .A2(n4354), .A3(n4353), .A4(n4352), .ZN(n4356)
         );
  NOR2_X1 U4833 ( .A1(n4357), .A2(n4356), .ZN(n4382) );
  NAND2_X1 U4834 ( .A1(n4359), .A2(n4358), .ZN(n4381) );
  XOR2_X1 U4835 ( .A(n4382), .B(n4381), .Z(n4364) );
  INV_X1 U4836 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4360) );
  INV_X1 U4837 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5593) );
  OAI22_X1 U4838 ( .A1(n4361), .A2(n4360), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5593), .ZN(n4362) );
  AOI21_X1 U4839 ( .B1(n4364), .B2(n4363), .A(n4362), .ZN(n4365) );
  XNOR2_X1 U4840 ( .A(n4388), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5595)
         );
  MUX2_X1 U4841 ( .A(n4365), .B(n5595), .S(n5020), .Z(n5382) );
  AOI22_X1 U4842 ( .A1(n4350), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U4843 ( .A1(n4366), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4844 ( .A1(n3835), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U4845 ( .A1(n3711), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4367) );
  NAND4_X1 U4846 ( .A1(n4370), .A2(n4369), .A3(n4368), .A4(n4367), .ZN(n4380)
         );
  AOI22_X1 U4847 ( .A1(n4326), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U4848 ( .A1(n4372), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U4849 ( .A1(n3437), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U4850 ( .A1(n4374), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4375) );
  NAND4_X1 U4851 ( .A1(n4378), .A2(n4377), .A3(n4376), .A4(n4375), .ZN(n4379)
         );
  NOR2_X1 U4852 ( .A1(n4380), .A2(n4379), .ZN(n4384) );
  NOR2_X1 U4853 ( .A1(n4382), .A2(n4381), .ZN(n4383) );
  XOR2_X1 U4854 ( .A(n4384), .B(n4383), .Z(n4387) );
  AOI22_X1 U4855 ( .A1(n3927), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6797), .ZN(n4385) );
  OAI21_X1 U4856 ( .B1(n4387), .B2(n4386), .A(n4385), .ZN(n4390) );
  INV_X1 U4857 ( .A(n4388), .ZN(n4389) );
  XNOR2_X1 U4858 ( .A(n4557), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5374)
         );
  MUX2_X1 U4859 ( .A(n4390), .B(n5374), .S(n5020), .Z(n4391) );
  NOR2_X2 U4860 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6808) );
  NOR2_X1 U4861 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6585), .ZN(n5019) );
  NAND2_X1 U4862 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5019), .ZN(n6224) );
  INV_X1 U4863 ( .A(n6224), .ZN(n4392) );
  NOR2_X1 U4864 ( .A1(n4393), .A2(n4611), .ZN(n4394) );
  INV_X1 U4865 ( .A(n4547), .ZN(n5590) );
  INV_X1 U4866 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U4867 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4752) );
  NOR3_X1 U4868 ( .A1(n5590), .A2(n5611), .A3(n4752), .ZN(n4478) );
  NAND2_X1 U4869 ( .A1(n4403), .A2(n4397), .ZN(n4409) );
  OAI211_X1 U4870 ( .C1(n4397), .C2(n4403), .A(n4396), .B(n4409), .ZN(n4400)
         );
  NOR2_X1 U4871 ( .A1(n4398), .A2(n5562), .ZN(n4399) );
  AND2_X1 U4872 ( .A1(n4400), .A2(n4399), .ZN(n4401) );
  INV_X1 U4873 ( .A(n4396), .ZN(n6229) );
  NAND2_X1 U4874 ( .A1(n3528), .A2(n4402), .ZN(n4411) );
  OAI21_X1 U4875 ( .B1(n6229), .B2(n4403), .A(n4411), .ZN(n4404) );
  INV_X1 U4876 ( .A(n4404), .ZN(n4405) );
  OAI21_X1 U4877 ( .B1(n6780), .B2(n4611), .A(n4405), .ZN(n6163) );
  AND2_X1 U4878 ( .A1(n6163), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6165)
         );
  NAND2_X1 U4879 ( .A1(n4851), .A2(n6165), .ZN(n4407) );
  NAND2_X1 U4880 ( .A1(n4406), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4852)
         );
  NAND2_X1 U4881 ( .A1(n6171), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4416)
         );
  INV_X1 U4882 ( .A(n4408), .ZN(n4410) );
  NAND2_X1 U4883 ( .A1(n4409), .A2(n4410), .ZN(n4420) );
  OAI21_X1 U4884 ( .B1(n4410), .B2(n4409), .A(n4420), .ZN(n4413) );
  INV_X1 U4885 ( .A(n4411), .ZN(n4412) );
  AOI21_X1 U4886 ( .B1(n4413), .B2(n4396), .A(n4412), .ZN(n4414) );
  NAND2_X1 U4887 ( .A1(n6172), .A2(n4416), .ZN(n4419) );
  INV_X1 U4888 ( .A(n6171), .ZN(n4417) );
  INV_X1 U4889 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U4890 ( .A1(n4417), .A2(n6291), .ZN(n4418) );
  INV_X1 U4891 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U4892 ( .A1(n4420), .A2(n4421), .ZN(n4437) );
  OAI211_X1 U4893 ( .C1(n4421), .C2(n4420), .A(n4437), .B(n4396), .ZN(n4422)
         );
  INV_X1 U4894 ( .A(n4422), .ZN(n4423) );
  NAND2_X1 U4895 ( .A1(n4425), .A2(n4424), .ZN(n6178) );
  INV_X1 U4896 ( .A(n6178), .ZN(n4431) );
  NAND2_X1 U4897 ( .A1(n4426), .A2(n4485), .ZN(n4429) );
  XNOR2_X1 U4898 ( .A(n4437), .B(n4435), .ZN(n4427) );
  NAND2_X1 U4899 ( .A1(n4427), .A2(n4396), .ZN(n4428) );
  INV_X1 U4900 ( .A(n6179), .ZN(n4430) );
  NAND2_X1 U4901 ( .A1(n4431), .A2(n4430), .ZN(n6181) );
  NAND2_X1 U4902 ( .A1(n4432), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4433)
         );
  NAND2_X1 U4903 ( .A1(n6181), .A2(n4433), .ZN(n6185) );
  NAND2_X1 U4904 ( .A1(n4434), .A2(n4485), .ZN(n4440) );
  INV_X1 U4905 ( .A(n4435), .ZN(n4436) );
  OR2_X1 U4906 ( .A1(n4437), .A2(n4436), .ZN(n4445) );
  XNOR2_X1 U4907 ( .A(n4445), .B(n4452), .ZN(n4438) );
  NAND2_X1 U4908 ( .A1(n4438), .A2(n4396), .ZN(n4439) );
  NAND2_X1 U4909 ( .A1(n4440), .A2(n4439), .ZN(n4441) );
  INV_X1 U4910 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4652) );
  XNOR2_X1 U4911 ( .A(n4441), .B(n4652), .ZN(n6184) );
  NAND2_X1 U4912 ( .A1(n6185), .A2(n6184), .ZN(n6187) );
  NAND2_X1 U4913 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4442)
         );
  NAND3_X1 U4914 ( .A1(n4444), .A2(n4485), .A3(n4443), .ZN(n4449) );
  INV_X1 U4915 ( .A(n4445), .ZN(n4454) );
  NAND2_X1 U4916 ( .A1(n4454), .A2(n4452), .ZN(n4446) );
  XNOR2_X1 U4917 ( .A(n4446), .B(n4451), .ZN(n4447) );
  NAND2_X1 U4918 ( .A1(n4447), .A2(n4396), .ZN(n4448) );
  NAND2_X1 U4919 ( .A1(n4449), .A2(n4448), .ZN(n6193) );
  OR2_X1 U4920 ( .A1(n4450), .A2(n4611), .ZN(n4457) );
  AND2_X1 U4921 ( .A1(n4452), .A2(n4451), .ZN(n4453) );
  NAND2_X1 U4922 ( .A1(n4454), .A2(n4453), .ZN(n4461) );
  XNOR2_X1 U4923 ( .A(n4461), .B(n4462), .ZN(n4455) );
  NAND2_X1 U4924 ( .A1(n4455), .A2(n4396), .ZN(n4456) );
  NAND2_X1 U4925 ( .A1(n4457), .A2(n4456), .ZN(n4458) );
  XNOR2_X1 U4926 ( .A(n4458), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6198)
         );
  INV_X1 U4927 ( .A(n4458), .ZN(n4460) );
  INV_X1 U4928 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4459) );
  INV_X1 U4929 ( .A(n4461), .ZN(n4463) );
  NAND3_X1 U4930 ( .A1(n4463), .A2(n4396), .A3(n4462), .ZN(n4464) );
  NAND2_X1 U4931 ( .A1(n4466), .A2(n4464), .ZN(n4465) );
  XOR2_X1 U4932 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .B(n4465), .Z(n5169) );
  XOR2_X1 U4933 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .B(n5689), .Z(n5174) );
  INV_X4 U4934 ( .A(n4466), .ZN(n5629) );
  INV_X1 U4935 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5179) );
  XNOR2_X1 U4936 ( .A(n5704), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5195)
         );
  INV_X1 U4937 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5250) );
  INV_X1 U4938 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4676) );
  NOR2_X1 U4939 ( .A1(n5689), .A2(n4676), .ZN(n5245) );
  XNOR2_X1 U4940 ( .A(n5704), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6204)
         );
  NAND2_X1 U4941 ( .A1(n6205), .A2(n6204), .ZN(n6203) );
  INV_X1 U4942 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U4943 ( .A1(n5703), .A2(n4470), .ZN(n4471) );
  NAND2_X1 U4944 ( .A1(n4471), .A2(n3485), .ZN(n5696) );
  INV_X1 U4945 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5810) );
  INV_X1 U4946 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U4947 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4627) );
  INV_X1 U4948 ( .A(n4627), .ZN(n4473) );
  INV_X1 U4949 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4474) );
  NOR2_X1 U4950 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5772) );
  NOR2_X1 U4951 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5788) );
  INV_X1 U4952 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5754) );
  INV_X1 U4953 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5768) );
  AND2_X1 U4954 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5787) );
  AND2_X1 U4955 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5771) );
  AND2_X1 U4956 ( .A1(n5787), .A2(n5771), .ZN(n5752) );
  AND2_X1 U4957 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U4958 ( .A1(n5752), .A2(n4622), .ZN(n4632) );
  NOR2_X2 U4959 ( .A1(n4476), .A2(n3479), .ZN(n5622) );
  XNOR2_X1 U4960 ( .A(n5689), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5621)
         );
  NAND2_X1 U4961 ( .A1(n5622), .A2(n5621), .ZN(n5620) );
  INV_X1 U4962 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6331) );
  NAND2_X2 U4963 ( .A1(n5620), .A2(n4477), .ZN(n5612) );
  NOR2_X1 U4964 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5600) );
  INV_X1 U4965 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5732) );
  AOI21_X1 U4966 ( .B1(n5600), .B2(n5732), .A(n5689), .ZN(n5588) );
  OR2_X1 U4967 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5589)
         );
  NOR3_X2 U4968 ( .A1(n5612), .A2(n5588), .A3(n5589), .ZN(n4549) );
  AOI21_X1 U4969 ( .B1(n4478), .B2(n5612), .A(n4549), .ZN(n4479) );
  XNOR2_X1 U4970 ( .A(n4479), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4741)
         );
  NAND2_X1 U4971 ( .A1(n6794), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4491) );
  XNOR2_X1 U4972 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U4973 ( .A1(n4493), .A2(n4492), .ZN(n4481) );
  NAND2_X1 U4974 ( .A1(n6793), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U4975 ( .A1(n4481), .A2(n4480), .ZN(n4487) );
  MUX2_X1 U4976 ( .A(n4482), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4486) );
  NAND2_X1 U4977 ( .A1(n4487), .A2(n4486), .ZN(n4484) );
  NAND2_X1 U4978 ( .A1(n4482), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4483) );
  MUX2_X1 U4979 ( .A(n5132), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(n6544), 
        .Z(n4513) );
  XNOR2_X1 U4980 ( .A(n4514), .B(n4513), .ZN(n4572) );
  INV_X1 U4981 ( .A(n4519), .ZN(n4511) );
  XNOR2_X1 U4982 ( .A(n4487), .B(n4486), .ZN(n4570) );
  INV_X1 U4983 ( .A(n5562), .ZN(n4494) );
  OAI21_X1 U4984 ( .B1(n3528), .B2(n4494), .A(n3725), .ZN(n4501) );
  INV_X1 U4985 ( .A(n4501), .ZN(n4490) );
  INV_X1 U4986 ( .A(n4570), .ZN(n4488) );
  NAND2_X1 U4987 ( .A1(n4529), .A2(n4488), .ZN(n4502) );
  INV_X1 U4988 ( .A(n4502), .ZN(n4489) );
  AOI211_X1 U4989 ( .C1(n4519), .C2(n4570), .A(n4490), .B(n4489), .ZN(n4510)
         );
  OAI21_X1 U4990 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6794), .A(n4491), 
        .ZN(n4498) );
  INV_X1 U4991 ( .A(n4498), .ZN(n4500) );
  XNOR2_X1 U4992 ( .A(n4493), .B(n4492), .ZN(n4571) );
  INV_X1 U4993 ( .A(n4529), .ZN(n4497) );
  OAI21_X1 U4994 ( .B1(n4497), .B2(n3725), .A(n4494), .ZN(n4495) );
  AOI21_X1 U4995 ( .B1(n4519), .B2(n4571), .A(n4495), .ZN(n4504) );
  INV_X1 U4996 ( .A(n4571), .ZN(n4496) );
  NAND2_X1 U4997 ( .A1(n4496), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4505) );
  AOI211_X1 U4998 ( .C1(n4504), .C2(n4505), .A(n4498), .B(n4497), .ZN(n4499)
         );
  NOR2_X1 U4999 ( .A1(n4499), .A2(n4532), .ZN(n4503) );
  AOI211_X1 U5000 ( .C1(n3727), .C2(n4500), .A(n3528), .B(n4503), .ZN(n4508)
         );
  AOI21_X1 U5001 ( .B1(n4503), .B2(n4502), .A(n4501), .ZN(n4507) );
  AOI21_X1 U5002 ( .B1(n4520), .B2(n4505), .A(n4504), .ZN(n4506) );
  NOR3_X1 U5003 ( .A1(n4508), .A2(n4507), .A3(n4506), .ZN(n4509) );
  AOI211_X1 U5004 ( .C1(n4511), .C2(n4572), .A(n4510), .B(n4509), .ZN(n4512)
         );
  AOI21_X1 U5005 ( .B1(n4572), .B2(n4532), .A(n4512), .ZN(n4522) );
  NAND2_X1 U5006 ( .A1(n4514), .A2(n4513), .ZN(n4516) );
  NAND2_X1 U5007 ( .A1(n5132), .A2(n6544), .ZN(n4515) );
  NAND2_X1 U5008 ( .A1(n4516), .A2(n4515), .ZN(n4526) );
  NOR2_X1 U5009 ( .A1(n4519), .A2(n4575), .ZN(n4521) );
  OAI22_X1 U5010 ( .A1(n4522), .A2(n4521), .B1(n4520), .B2(n4575), .ZN(n4523)
         );
  AOI21_X1 U5011 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6594), .A(n4523), 
        .ZN(n4531) );
  NAND2_X1 U5012 ( .A1(n4524), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5013 ( .A1(n4526), .A2(n4525), .ZN(n4527) );
  NAND2_X1 U5014 ( .A1(n4529), .A2(n4574), .ZN(n4530) );
  NAND2_X1 U5015 ( .A1(n4531), .A2(n4530), .ZN(n4534) );
  NAND2_X1 U5016 ( .A1(n4535), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6598) );
  NAND3_X1 U5017 ( .A1(n5009), .A2(n4402), .A3(n5370), .ZN(n4610) );
  NOR2_X1 U5018 ( .A1(n4536), .A2(n4610), .ZN(n6563) );
  NAND2_X1 U5019 ( .A1(n4741), .A2(n6212), .ZN(n4544) );
  INV_X1 U5020 ( .A(n6808), .ZN(n6768) );
  NAND2_X1 U5021 ( .A1(n6768), .A2(n4537), .ZN(n6227) );
  AND2_X1 U5022 ( .A1(n6227), .A2(n6594), .ZN(n4538) );
  AND2_X2 U5023 ( .A1(n5229), .A2(n6594), .ZN(n6322) );
  INV_X1 U5024 ( .A(n6322), .ZN(n6262) );
  INV_X1 U5025 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6118) );
  NOR2_X1 U5026 ( .A1(n6262), .A2(n6118), .ZN(n4754) );
  NAND2_X1 U5027 ( .A1(n6594), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U5028 ( .A1(n6817), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4539) );
  AND2_X1 U5029 ( .A1(n4540), .A2(n4539), .ZN(n6166) );
  INV_X1 U5030 ( .A(n6166), .ZN(n4541) );
  NOR2_X1 U5031 ( .A1(n6216), .A2(n5374), .ZN(n4542) );
  AOI211_X1 U5032 ( .C1(PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n6210), .A(n4754), 
        .B(n4542), .ZN(n4543) );
  NAND3_X1 U5033 ( .A1(n4545), .A2(n4544), .A3(n4543), .ZN(U2956) );
  NAND2_X2 U5034 ( .A1(n5612), .A2(n3482), .ZN(n4562) );
  NOR2_X1 U5035 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4546)
         );
  NAND2_X1 U5036 ( .A1(n3445), .A2(n4548), .ZN(n4551) );
  INV_X1 U5037 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U5038 ( .A1(n4549), .A2(n5712), .ZN(n4550) );
  NAND2_X1 U5039 ( .A1(n4551), .A2(n4550), .ZN(n4552) );
  XNOR2_X1 U5040 ( .A(n4552), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5720)
         );
  AOI22_X1 U5041 ( .A1(n3927), .A2(EAX_REG_31__SCAN_IN), .B1(n4553), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4554) );
  INV_X1 U5042 ( .A(n4554), .ZN(n4555) );
  NAND2_X1 U5043 ( .A1(n4557), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4558)
         );
  INV_X1 U5044 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5351) );
  XNOR2_X1 U5045 ( .A(n4558), .B(n5351), .ZN(n5035) );
  NAND2_X1 U5046 ( .A1(n6322), .A2(REIP_REG_31__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U5047 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4559)
         );
  OAI211_X1 U5048 ( .C1(n6216), .C2(n5035), .A(n5714), .B(n4559), .ZN(n4560)
         );
  OAI21_X1 U5049 ( .B1(n5720), .B2(n6535), .A(n4561), .ZN(U2955) );
  NAND2_X1 U5050 ( .A1(n4562), .A2(n5689), .ZN(n4563) );
  INV_X1 U5051 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4564) );
  INV_X1 U5052 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U5053 ( .A1(n4567), .A2(n4566), .ZN(n6221) );
  NAND2_X1 U5054 ( .A1(n3725), .A2(n6221), .ZN(n4568) );
  NAND2_X1 U5055 ( .A1(n5365), .A2(n4568), .ZN(n4905) );
  NOR3_X1 U5056 ( .A1(n4572), .A2(n4571), .A3(n4570), .ZN(n4573) );
  OR2_X1 U5057 ( .A1(n4574), .A2(n4573), .ZN(n4576) );
  NAND2_X1 U5058 ( .A1(n4576), .A2(n4575), .ZN(n5368) );
  INV_X1 U5059 ( .A(n5009), .ZN(n4601) );
  NAND2_X1 U5060 ( .A1(n4593), .A2(n6221), .ZN(n5371) );
  NAND3_X1 U5061 ( .A1(n5368), .A2(n4601), .A3(n5371), .ZN(n4577) );
  OAI21_X1 U5062 ( .B1(n4905), .B2(n3507), .A(n4577), .ZN(n4578) );
  INV_X1 U5063 ( .A(READY_N), .ZN(n6619) );
  NAND2_X1 U5064 ( .A1(n4578), .A2(n6619), .ZN(n4590) );
  NOR2_X1 U5065 ( .A1(n3751), .A2(n4611), .ZN(n4580) );
  NAND3_X1 U5066 ( .A1(n5365), .A2(n5370), .A3(n4599), .ZN(n4579) );
  OAI211_X1 U5067 ( .C1(n5365), .C2(n4580), .A(n4579), .B(n5009), .ZN(n4588)
         );
  OR2_X1 U5068 ( .A1(n4581), .A2(n4601), .ZN(n4598) );
  OAI21_X1 U5069 ( .B1(n3751), .B2(n5562), .A(n3528), .ZN(n4582) );
  INV_X1 U5070 ( .A(n4582), .ZN(n4583) );
  NOR2_X1 U5071 ( .A1(n4598), .A2(n4583), .ZN(n4592) );
  AOI21_X1 U5072 ( .B1(n3731), .B2(n5370), .A(n4396), .ZN(n4584) );
  OR2_X1 U5073 ( .A1(n4585), .A2(n4584), .ZN(n4604) );
  NAND2_X1 U5074 ( .A1(n4592), .A2(n4604), .ZN(n4587) );
  NAND2_X1 U5075 ( .A1(n4587), .A2(n4586), .ZN(n4899) );
  AND2_X1 U5076 ( .A1(n4588), .A2(n4899), .ZN(n4589) );
  NAND2_X1 U5077 ( .A1(n4590), .A2(n4589), .ZN(n4591) );
  OR2_X1 U5078 ( .A1(n4894), .A2(n6563), .ZN(n5362) );
  NAND2_X1 U5079 ( .A1(n4569), .A2(n4872), .ZN(n4595) );
  OAI211_X1 U5080 ( .C1(n3763), .C2(n4734), .A(n4595), .B(n5109), .ZN(n4596)
         );
  NOR2_X1 U5081 ( .A1(n5362), .A2(n4596), .ZN(n4597) );
  INV_X1 U5082 ( .A(n4402), .ZN(n5000) );
  NAND2_X1 U5083 ( .A1(n4598), .A2(n5339), .ZN(n4603) );
  OAI21_X1 U5084 ( .B1(n4599), .B2(n5370), .A(n4601), .ZN(n4602) );
  NAND2_X1 U5085 ( .A1(n3528), .A2(n4593), .ZN(n5042) );
  OR2_X1 U5086 ( .A1(n5042), .A2(n4601), .ZN(n4898) );
  AND4_X1 U5087 ( .A1(n4604), .A2(n4603), .A3(n4602), .A4(n4898), .ZN(n4605)
         );
  NAND2_X1 U5088 ( .A1(n4606), .A2(n4605), .ZN(n4879) );
  INV_X1 U5089 ( .A(n4607), .ZN(n4608) );
  NOR2_X1 U5090 ( .A1(n4879), .A2(n4608), .ZN(n4609) );
  NOR2_X1 U5091 ( .A1(n4738), .A2(n4609), .ZN(n6242) );
  NOR2_X1 U5092 ( .A1(n4611), .A2(n4610), .ZN(n4612) );
  NAND2_X1 U5093 ( .A1(n5318), .A2(n4612), .ZN(n4884) );
  AND2_X1 U5094 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U5095 ( .A1(n6262), .A2(n4738), .ZN(n6344) );
  INV_X1 U5096 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U5097 ( .A1(n6242), .A2(n6346), .ZN(n6336) );
  NAND2_X1 U5098 ( .A1(n6344), .A2(n6336), .ZN(n5176) );
  INV_X1 U5099 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5066) );
  NOR2_X1 U5100 ( .A1(n6291), .A2(n5066), .ZN(n5054) );
  INV_X1 U5101 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4648) );
  NOR2_X1 U5102 ( .A1(n4648), .A2(n5055), .ZN(n6277) );
  NAND3_X1 U5103 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6277), .ZN(n5177) );
  INV_X1 U5104 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5204) );
  NOR2_X1 U5105 ( .A1(n5204), .A2(n4459), .ZN(n5203) );
  INV_X1 U5106 ( .A(n5203), .ZN(n5178) );
  NAND2_X1 U5107 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5218) );
  NOR3_X1 U5108 ( .A1(n5177), .A2(n5178), .A3(n5218), .ZN(n5219) );
  NAND2_X1 U5109 ( .A1(n5054), .A2(n5219), .ZN(n6247) );
  NAND3_X1 U5110 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5818) );
  NOR2_X1 U5111 ( .A1(n5819), .A2(n5818), .ZN(n5809) );
  NAND3_X1 U5112 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5809), .ZN(n4615) );
  NOR2_X1 U5113 ( .A1(n6247), .A2(n4615), .ZN(n4628) );
  INV_X1 U5114 ( .A(n4628), .ZN(n4613) );
  NAND2_X1 U5115 ( .A1(n4614), .A2(n4613), .ZN(n4617) );
  INV_X1 U5116 ( .A(n4615), .ZN(n6312) );
  NAND2_X1 U5117 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6312), .ZN(n5799) );
  AOI21_X1 U5118 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6289) );
  INV_X1 U5119 ( .A(n6289), .ZN(n5053) );
  NAND2_X1 U5120 ( .A1(n5219), .A2(n5053), .ZN(n6244) );
  NOR2_X1 U5121 ( .A1(n5799), .A2(n6244), .ZN(n4625) );
  OR2_X1 U5122 ( .A1(n6288), .A2(n4625), .ZN(n4616) );
  NAND2_X1 U5123 ( .A1(n4617), .A2(n4616), .ZN(n4618) );
  NOR2_X1 U5124 ( .A1(n5176), .A2(n4618), .ZN(n6313) );
  NAND2_X1 U5125 ( .A1(n5817), .A2(n4627), .ZN(n4619) );
  NAND2_X1 U5126 ( .A1(n6313), .A2(n4619), .ZN(n6236) );
  INV_X1 U5127 ( .A(n5752), .ZN(n5762) );
  AND2_X1 U5128 ( .A1(n5817), .A2(n5762), .ZN(n4620) );
  NOR2_X1 U5129 ( .A1(n6236), .A2(n4620), .ZN(n5769) );
  INV_X1 U5130 ( .A(n6292), .ZN(n4621) );
  NAND2_X1 U5131 ( .A1(n6288), .A2(n4621), .ZN(n5248) );
  INV_X1 U5132 ( .A(n4622), .ZN(n4623) );
  NAND2_X1 U5133 ( .A1(n5248), .A2(n4623), .ZN(n4624) );
  OAI21_X1 U5134 ( .B1(n5807), .B2(n5743), .A(n6332), .ZN(n5739) );
  NAND2_X1 U5135 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n4625), .ZN(n4626) );
  OR2_X1 U5136 ( .A1(n6288), .A2(n4626), .ZN(n4631) );
  NAND2_X1 U5137 ( .A1(n6292), .A2(n4628), .ZN(n5800) );
  INV_X1 U5138 ( .A(n5800), .ZN(n4629) );
  NAND2_X1 U5139 ( .A1(n4473), .A2(n4629), .ZN(n4630) );
  NAND2_X1 U5140 ( .A1(n4631), .A2(n4630), .ZN(n5770) );
  INV_X1 U5141 ( .A(n4632), .ZN(n4633) );
  NAND2_X1 U5142 ( .A1(n6321), .A2(n5743), .ZN(n5731) );
  NOR2_X1 U5143 ( .A1(n5731), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5738)
         );
  INV_X1 U5144 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5145 ( .A1(n4742), .A2(n4634), .ZN(n4638) );
  NAND2_X1 U5146 ( .A1(n4743), .A2(n5066), .ZN(n4636) );
  NAND2_X1 U5147 ( .A1(n4872), .A2(n4634), .ZN(n4635) );
  NAND3_X1 U5148 ( .A1(n4636), .A2(n5337), .A3(n4635), .ZN(n4637) );
  NAND2_X1 U5149 ( .A1(n4638), .A2(n4637), .ZN(n4640) );
  NAND2_X1 U5150 ( .A1(n4743), .A2(EBX_REG_0__SCAN_IN), .ZN(n4639) );
  OAI21_X1 U5151 ( .B1(n4750), .B2(EBX_REG_0__SCAN_IN), .A(n4639), .ZN(n4842)
         );
  XNOR2_X1 U5152 ( .A(n4640), .B(n4842), .ZN(n5075) );
  NAND2_X1 U5153 ( .A1(n5075), .A2(n4872), .ZN(n4874) );
  NAND2_X1 U5154 ( .A1(n4874), .A2(n4640), .ZN(n4917) );
  MUX2_X1 U5155 ( .A(n4729), .B(n5337), .S(EBX_REG_3__SCAN_IN), .Z(n4642) );
  OR2_X1 U5156 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4641)
         );
  AND2_X1 U5157 ( .A1(n4642), .A2(n4641), .ZN(n4918) );
  INV_X1 U5158 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U5159 ( .A1(n4742), .A2(n6148), .ZN(n4646) );
  NAND2_X1 U5160 ( .A1(n4743), .A2(n6291), .ZN(n4644) );
  NAND2_X1 U5161 ( .A1(n4872), .A2(n6148), .ZN(n4643) );
  NAND3_X1 U5162 ( .A1(n4644), .A2(n5337), .A3(n4643), .ZN(n4645) );
  NAND2_X1 U5163 ( .A1(n4646), .A2(n4645), .ZN(n5151) );
  NAND2_X1 U5164 ( .A1(n4918), .A2(n5151), .ZN(n4647) );
  NAND2_X1 U5165 ( .A1(n4743), .A2(n4648), .ZN(n4650) );
  INV_X1 U5166 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U5167 ( .A1(n4872), .A2(n6161), .ZN(n4649) );
  NAND3_X1 U5168 ( .A1(n4650), .A2(n5337), .A3(n4649), .ZN(n4651) );
  OAI21_X1 U5169 ( .B1(n4728), .B2(EBX_REG_4__SCAN_IN), .A(n4651), .ZN(n6153)
         );
  NAND2_X1 U5170 ( .A1(n4652), .A2(n4747), .ZN(n4654) );
  MUX2_X1 U5171 ( .A(n4729), .B(n5337), .S(EBX_REG_5__SCAN_IN), .Z(n4653) );
  NAND2_X1 U5172 ( .A1(n4654), .A2(n4653), .ZN(n4914) );
  INV_X1 U5173 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U5174 ( .A1(n4742), .A2(n4655), .ZN(n4659) );
  NAND2_X1 U5175 ( .A1(n4743), .A2(n6274), .ZN(n4657) );
  NAND2_X1 U5176 ( .A1(n4872), .A2(n4655), .ZN(n4656) );
  NAND3_X1 U5177 ( .A1(n4657), .A2(n5337), .A3(n4656), .ZN(n4658) );
  AND2_X1 U5178 ( .A1(n4659), .A2(n4658), .ZN(n4964) );
  NAND2_X1 U5179 ( .A1(n4459), .A2(n4747), .ZN(n4663) );
  MUX2_X1 U5180 ( .A(n4729), .B(n5337), .S(EBX_REG_7__SCAN_IN), .Z(n4662) );
  NAND2_X1 U5181 ( .A1(n4663), .A2(n4662), .ZN(n5137) );
  NAND2_X1 U5182 ( .A1(n4743), .A2(n5204), .ZN(n4665) );
  INV_X1 U5183 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U5184 ( .A1(n4872), .A2(n6406), .ZN(n4664) );
  NAND3_X1 U5185 ( .A1(n4665), .A2(n5337), .A3(n4664), .ZN(n4666) );
  OAI21_X1 U5186 ( .B1(n4728), .B2(EBX_REG_8__SCAN_IN), .A(n4666), .ZN(n5162)
         );
  NAND2_X1 U5187 ( .A1(n5179), .A2(n4747), .ZN(n4668) );
  MUX2_X1 U5188 ( .A(n4729), .B(n5337), .S(EBX_REG_9__SCAN_IN), .Z(n4667) );
  NAND2_X1 U5189 ( .A1(n4668), .A2(n4667), .ZN(n5149) );
  INV_X1 U5190 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U5191 ( .A1(n4742), .A2(n6424), .ZN(n4673) );
  INV_X1 U5192 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5193 ( .A1(n4743), .A2(n4669), .ZN(n4671) );
  NAND2_X1 U5194 ( .A1(n4872), .A2(n6424), .ZN(n4670) );
  NAND3_X1 U5195 ( .A1(n4671), .A2(n5337), .A3(n4670), .ZN(n4672) );
  NAND2_X1 U5196 ( .A1(n5250), .A2(n4747), .ZN(n4675) );
  MUX2_X1 U5197 ( .A(n4729), .B(n5337), .S(EBX_REG_11__SCAN_IN), .Z(n4674) );
  NAND2_X1 U5198 ( .A1(n4675), .A2(n4674), .ZN(n5213) );
  OAI21_X1 U5199 ( .B1(n4750), .B2(n4676), .A(n4743), .ZN(n4679) );
  INV_X1 U5200 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4677) );
  NAND2_X1 U5201 ( .A1(n4872), .A2(n4677), .ZN(n4678) );
  NAND2_X1 U5202 ( .A1(n4679), .A2(n4678), .ZN(n4680) );
  OAI21_X1 U5203 ( .B1(EBX_REG_12__SCAN_IN), .B2(n4728), .A(n4680), .ZN(n5231)
         );
  NAND2_X1 U5204 ( .A1(n5232), .A2(n5231), .ZN(n5295) );
  INV_X1 U5205 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U5206 ( .A1(n6259), .A2(n4747), .ZN(n4682) );
  MUX2_X1 U5207 ( .A(n4729), .B(n5337), .S(EBX_REG_13__SCAN_IN), .Z(n4681) );
  NAND2_X1 U5208 ( .A1(n4682), .A2(n4681), .ZN(n5296) );
  MUX2_X1 U5209 ( .A(n4729), .B(n5337), .S(EBX_REG_15__SCAN_IN), .Z(n4684) );
  OR2_X1 U5210 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4683)
         );
  AND2_X1 U5211 ( .A1(n4684), .A2(n4683), .ZN(n5308) );
  INV_X1 U5212 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U5213 ( .A1(n4742), .A2(n6152), .ZN(n4688) );
  NAND2_X1 U5214 ( .A1(n4743), .A2(n5819), .ZN(n4686) );
  NAND2_X1 U5215 ( .A1(n4872), .A2(n6152), .ZN(n4685) );
  NAND3_X1 U5216 ( .A1(n4686), .A2(n5337), .A3(n4685), .ZN(n4687) );
  NAND2_X1 U5217 ( .A1(n4688), .A2(n4687), .ZN(n5821) );
  NAND2_X1 U5218 ( .A1(n5308), .A2(n5821), .ZN(n4689) );
  NAND2_X1 U5219 ( .A1(n4743), .A2(n5678), .ZN(n4691) );
  INV_X1 U5220 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U5221 ( .A1(n4872), .A2(n5555), .ZN(n4690) );
  NAND3_X1 U5222 ( .A1(n4691), .A2(n5337), .A3(n4690), .ZN(n4692) );
  OAI21_X1 U5223 ( .B1(n4728), .B2(EBX_REG_16__SCAN_IN), .A(n4692), .ZN(n5551)
         );
  MUX2_X1 U5224 ( .A(n4729), .B(n5337), .S(EBX_REG_17__SCAN_IN), .Z(n4694) );
  OR2_X1 U5225 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4693)
         );
  INV_X1 U5226 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U5227 ( .A1(n4742), .A2(n6497), .ZN(n4699) );
  INV_X1 U5228 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U5229 ( .A1(n4743), .A2(n4695), .ZN(n4697) );
  NAND2_X1 U5230 ( .A1(n4872), .A2(n6497), .ZN(n4696) );
  NAND3_X1 U5231 ( .A1(n4697), .A2(n5337), .A3(n4696), .ZN(n4698) );
  AND2_X1 U5232 ( .A1(n4699), .A2(n4698), .ZN(n5536) );
  INV_X1 U5233 ( .A(n4729), .ZN(n4706) );
  INV_X1 U5234 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U5235 ( .A1(n4706), .A2(n5498), .ZN(n4702) );
  INV_X1 U5236 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U5237 ( .A1(n4872), .A2(n5498), .ZN(n4700) );
  OAI211_X1 U5238 ( .C1(n4750), .C2(n5661), .A(n4700), .B(n4743), .ZN(n4701)
         );
  NAND2_X1 U5239 ( .A1(n4702), .A2(n4701), .ZN(n5485) );
  INV_X1 U5240 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5794) );
  OAI21_X1 U5241 ( .B1(n4750), .B2(n5794), .A(n4743), .ZN(n4704) );
  INV_X1 U5242 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U5243 ( .A1(n4872), .A2(n5530), .ZN(n4703) );
  NAND2_X1 U5244 ( .A1(n4704), .A2(n4703), .ZN(n4705) );
  OAI21_X1 U5245 ( .B1(EBX_REG_20__SCAN_IN), .B2(n4728), .A(n4705), .ZN(n5524)
         );
  INV_X1 U5246 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U5247 ( .A1(n4706), .A2(n5521), .ZN(n4710) );
  INV_X1 U5248 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U5249 ( .A1(n4872), .A2(n5521), .ZN(n4707) );
  OAI211_X1 U5250 ( .C1(n4750), .C2(n4708), .A(n4707), .B(n4743), .ZN(n4709)
         );
  NAND2_X1 U5251 ( .A1(n5527), .A2(n5471), .ZN(n5516) );
  INV_X1 U5252 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U5253 ( .A1(n4742), .A2(n6534), .ZN(n4715) );
  INV_X1 U5254 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U5255 ( .A1(n4743), .A2(n4711), .ZN(n4713) );
  NAND2_X1 U5256 ( .A1(n4872), .A2(n6534), .ZN(n4712) );
  NAND3_X1 U5257 ( .A1(n4713), .A2(n5337), .A3(n4712), .ZN(n4714) );
  AND2_X1 U5258 ( .A1(n4715), .A2(n4714), .ZN(n5515) );
  MUX2_X1 U5259 ( .A(n4729), .B(n5337), .S(EBX_REG_23__SCAN_IN), .Z(n4717) );
  OR2_X1 U5260 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4716)
         );
  NAND2_X1 U5261 ( .A1(n4717), .A2(n4716), .ZN(n5457) );
  MUX2_X1 U5262 ( .A(n4729), .B(n5337), .S(EBX_REG_25__SCAN_IN), .Z(n4719) );
  OR2_X1 U5263 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4718)
         );
  AND2_X1 U5264 ( .A1(n4719), .A2(n4718), .ZN(n5427) );
  OAI21_X1 U5265 ( .B1(n4750), .B2(n5754), .A(n4743), .ZN(n4721) );
  INV_X1 U5266 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5267 ( .A1(n4872), .A2(n4722), .ZN(n4720) );
  NAND2_X1 U5268 ( .A1(n4721), .A2(n4720), .ZN(n4724) );
  NAND2_X1 U5269 ( .A1(n4742), .A2(n4722), .ZN(n4723) );
  NAND2_X1 U5270 ( .A1(n4724), .A2(n4723), .ZN(n5446) );
  NAND2_X1 U5271 ( .A1(n5427), .A2(n5446), .ZN(n4725) );
  NAND2_X1 U5272 ( .A1(n4743), .A2(n5611), .ZN(n4726) );
  OAI211_X1 U5273 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5338), .A(n4726), .B(n5337), 
        .ZN(n4727) );
  OAI21_X1 U5274 ( .B1(n4728), .B2(EBX_REG_26__SCAN_IN), .A(n4727), .ZN(n5411)
         );
  MUX2_X1 U5275 ( .A(n4729), .B(n5337), .S(EBX_REG_27__SCAN_IN), .Z(n4731) );
  OR2_X1 U5276 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4730)
         );
  NAND2_X1 U5277 ( .A1(n4731), .A2(n4730), .ZN(n4732) );
  NAND2_X1 U5278 ( .A1(n5413), .A2(n4732), .ZN(n4733) );
  NAND2_X1 U5279 ( .A1(n3467), .A2(n4733), .ZN(n5506) );
  NAND2_X1 U5280 ( .A1(n4569), .A2(n4396), .ZN(n6576) );
  INV_X1 U5281 ( .A(n4734), .ZN(n4735) );
  NAND2_X1 U5282 ( .A1(n4735), .A2(n3763), .ZN(n4736) );
  AND2_X1 U5283 ( .A1(n6576), .A2(n4736), .ZN(n4737) );
  NAND2_X1 U5284 ( .A1(n6322), .A2(REIP_REG_27__SCAN_IN), .ZN(n5327) );
  OAI21_X1 U5285 ( .B1(n5506), .B2(n6339), .A(n5327), .ZN(n4739) );
  AOI211_X1 U5286 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5739), .A(n5738), .B(n4739), .ZN(n4740) );
  OAI21_X1 U5287 ( .B1(n5334), .B2(n6334), .A(n4740), .ZN(U2991) );
  NAND2_X1 U5288 ( .A1(n4741), .A2(n6327), .ZN(n4757) );
  INV_X1 U5289 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U5290 ( .A1(n4742), .A2(n5505), .ZN(n4746) );
  NAND2_X1 U5291 ( .A1(n4743), .A2(n5732), .ZN(n4744) );
  OAI211_X1 U5292 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5338), .A(n4744), .B(n5337), 
        .ZN(n4745) );
  AND2_X1 U5293 ( .A1(n4746), .A2(n4745), .ZN(n5392) );
  NOR2_X2 U5294 ( .A1(n3467), .A2(n5392), .ZN(n5393) );
  INV_X1 U5295 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5504) );
  AND2_X1 U5296 ( .A1(n4872), .A2(n5504), .ZN(n4748) );
  INV_X1 U5297 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5722) );
  AOI21_X1 U5298 ( .B1(n4747), .B2(n5722), .A(n4748), .ZN(n4749) );
  MUX2_X1 U5299 ( .A(n4748), .B(n4749), .S(n5337), .Z(n5388) );
  NAND2_X1 U5300 ( .A1(n5393), .A2(n5388), .ZN(n5387) );
  AOI22_X1 U5301 ( .A1(n5387), .A2(n4750), .B1(n5393), .B2(n4749), .ZN(n4751)
         );
  OAI22_X1 U5302 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n5338), .ZN(n5336) );
  AOI21_X1 U5303 ( .B1(n5817), .B2(n4752), .A(n5739), .ZN(n5721) );
  OAI21_X1 U5304 ( .B1(n5807), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5721), 
        .ZN(n5711) );
  NOR2_X1 U5305 ( .A1(n5731), .A2(n4752), .ZN(n5723) );
  AND3_X1 U5306 ( .A1(n5723), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5712), 
        .ZN(n4753) );
  AOI211_X1 U5307 ( .C1(n5711), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4754), .B(n4753), .ZN(n4755) );
  NAND2_X1 U5308 ( .A1(n4757), .A2(n3556), .ZN(U2988) );
  NAND3_X1 U5309 ( .A1(n3735), .A2(n6572), .A3(n5368), .ZN(n4766) );
  INV_X1 U5310 ( .A(n4766), .ZN(n4760) );
  INV_X1 U5311 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6629) );
  INV_X1 U5312 ( .A(n4758), .ZN(n5361) );
  INV_X1 U5313 ( .A(n5229), .ZN(n4759) );
  OAI211_X1 U5314 ( .C1(n4760), .C2(n6629), .A(n4778), .B(n4759), .ZN(U2788)
         );
  NAND2_X1 U5315 ( .A1(n3735), .A2(n5368), .ZN(n4761) );
  NAND2_X1 U5316 ( .A1(n4758), .A2(n4761), .ZN(n4762) );
  AND2_X1 U5317 ( .A1(n3483), .A2(n4762), .ZN(n5372) );
  AND2_X1 U5318 ( .A1(n5372), .A2(n6572), .ZN(n4765) );
  INV_X1 U5319 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n4764) );
  NAND3_X1 U5320 ( .A1(n6580), .A2(STATE2_REG_0__SCAN_IN), .A3(n6797), .ZN(
        n4763) );
  OAI21_X1 U5321 ( .B1(n4765), .B2(n4764), .A(n4763), .ZN(U2790) );
  NOR2_X1 U5322 ( .A1(n5229), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4768) );
  NAND3_X1 U5323 ( .A1(n6226), .A2(n6229), .A3(n5042), .ZN(n4767) );
  OAI21_X1 U5324 ( .B1(n6226), .B2(n4768), .A(n4767), .ZN(U3474) );
  INV_X1 U5325 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4786) );
  AOI21_X1 U5326 ( .B1(n6576), .B2(n6550), .A(n6221), .ZN(n4769) );
  NAND2_X1 U5327 ( .A1(n6049), .A2(n5370), .ZN(n4983) );
  AND2_X2 U5328 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5019), .ZN(n6228) );
  NOR2_X4 U5329 ( .A1(n6228), .A2(n6049), .ZN(n6061) );
  AOI22_X1 U5330 ( .A1(n6228), .A2(UWORD_REG_6__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4770) );
  OAI21_X1 U5331 ( .B1(n4786), .B2(n4983), .A(n4770), .ZN(U2901) );
  AOI22_X1 U5332 ( .A1(n6228), .A2(UWORD_REG_8__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4771) );
  OAI21_X1 U5333 ( .B1(n4790), .B2(n4983), .A(n4771), .ZN(U2899) );
  AOI22_X1 U5334 ( .A1(n6228), .A2(UWORD_REG_7__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4772) );
  OAI21_X1 U5335 ( .B1(n4784), .B2(n4983), .A(n4772), .ZN(U2900) );
  INV_X1 U5336 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4774) );
  AOI22_X1 U5337 ( .A1(n6228), .A2(UWORD_REG_5__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4773) );
  OAI21_X1 U5338 ( .B1(n4774), .B2(n4983), .A(n4773), .ZN(U2902) );
  AOI22_X1 U5339 ( .A1(n6228), .A2(UWORD_REG_9__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4775) );
  OAI21_X1 U5340 ( .B1(n4797), .B2(n4983), .A(n4775), .ZN(U2898) );
  INV_X1 U5341 ( .A(n6576), .ZN(n4776) );
  OR2_X1 U5342 ( .A1(n4779), .A2(n3725), .ZN(n4926) );
  INV_X1 U5343 ( .A(DATAI_7_), .ZN(n5141) );
  OR2_X1 U5344 ( .A1(n4926), .A2(n5141), .ZN(n4783) );
  NAND2_X1 U5345 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4847), .ZN(n4780) );
  OAI211_X1 U5346 ( .C1(n4800), .C2(n4781), .A(n4783), .B(n4780), .ZN(U2946)
         );
  NAND2_X1 U5347 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4847), .ZN(n4782) );
  OAI211_X1 U5348 ( .C1(n4800), .C2(n4784), .A(n4783), .B(n4782), .ZN(U2931)
         );
  NAND2_X1 U5349 ( .A1(n4815), .A2(DATAI_6_), .ZN(n4814) );
  NAND2_X1 U5350 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4847), .ZN(n4785) );
  OAI211_X1 U5351 ( .C1(n4800), .C2(n4786), .A(n4814), .B(n4785), .ZN(U2930)
         );
  NAND2_X1 U5352 ( .A1(n4815), .A2(DATAI_5_), .ZN(n4829) );
  NAND2_X1 U5353 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4847), .ZN(n4787) );
  OAI211_X1 U5354 ( .C1(n4800), .C2(n4788), .A(n4829), .B(n4787), .ZN(U2944)
         );
  NAND2_X1 U5355 ( .A1(n4815), .A2(DATAI_8_), .ZN(n4811) );
  NAND2_X1 U5356 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n4847), .ZN(n4789) );
  OAI211_X1 U5357 ( .C1(n4800), .C2(n4790), .A(n4811), .B(n4789), .ZN(U2932)
         );
  NAND2_X1 U5358 ( .A1(n4815), .A2(DATAI_3_), .ZN(n4823) );
  NAND2_X1 U5359 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n4847), .ZN(n4791) );
  OAI211_X1 U5360 ( .C1(n4800), .C2(n4792), .A(n4823), .B(n4791), .ZN(U2927)
         );
  INV_X1 U5361 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U5362 ( .A1(n4815), .A2(DATAI_2_), .ZN(n4809) );
  NAND2_X1 U5363 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n4847), .ZN(n4793) );
  OAI211_X1 U5364 ( .C1(n4800), .C2(n4975), .A(n4809), .B(n4793), .ZN(U2926)
         );
  NAND2_X1 U5365 ( .A1(n4815), .A2(DATAI_11_), .ZN(n4802) );
  NAND2_X1 U5366 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n4847), .ZN(n4794) );
  OAI211_X1 U5367 ( .C1(n4800), .C2(n4795), .A(n4802), .B(n4794), .ZN(U2935)
         );
  NAND2_X1 U5368 ( .A1(n4815), .A2(DATAI_9_), .ZN(n4805) );
  NAND2_X1 U5369 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n4847), .ZN(n4796) );
  OAI211_X1 U5370 ( .C1(n4800), .C2(n4797), .A(n4805), .B(n4796), .ZN(U2933)
         );
  NAND2_X1 U5371 ( .A1(n4815), .A2(DATAI_14_), .ZN(n4818) );
  NAND2_X1 U5372 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n4847), .ZN(n4798) );
  OAI211_X1 U5373 ( .C1(n4800), .C2(n4799), .A(n4818), .B(n4798), .ZN(U2953)
         );
  AOI22_X1 U5374 ( .A1(n4848), .A2(EAX_REG_11__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n4801) );
  NAND2_X1 U5375 ( .A1(n4802), .A2(n4801), .ZN(U2950) );
  NAND2_X1 U5376 ( .A1(n4815), .A2(DATAI_4_), .ZN(n4833) );
  AOI22_X1 U5377 ( .A1(n4848), .A2(EAX_REG_20__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4803) );
  NAND2_X1 U5378 ( .A1(n4833), .A2(n4803), .ZN(U2928) );
  AOI22_X1 U5379 ( .A1(n4848), .A2(EAX_REG_9__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U5380 ( .A1(n4805), .A2(n4804), .ZN(U2948) );
  NAND2_X1 U5381 ( .A1(n4815), .A2(DATAI_10_), .ZN(n4825) );
  AOI22_X1 U5382 ( .A1(n4848), .A2(EAX_REG_26__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U5383 ( .A1(n4825), .A2(n4806), .ZN(U2934) );
  NAND2_X1 U5384 ( .A1(n4815), .A2(DATAI_12_), .ZN(n4820) );
  AOI22_X1 U5385 ( .A1(n4848), .A2(EAX_REG_12__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U5386 ( .A1(n4820), .A2(n4807), .ZN(U2951) );
  AOI22_X1 U5387 ( .A1(n4848), .A2(EAX_REG_2__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4808) );
  NAND2_X1 U5388 ( .A1(n4809), .A2(n4808), .ZN(U2941) );
  AOI22_X1 U5389 ( .A1(n4848), .A2(EAX_REG_8__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U5390 ( .A1(n4811), .A2(n4810), .ZN(U2947) );
  INV_X1 U5391 ( .A(DATAI_0_), .ZN(n4930) );
  OR2_X1 U5392 ( .A1(n4926), .A2(n4930), .ZN(n4827) );
  AOI22_X1 U5393 ( .A1(n4848), .A2(EAX_REG_0__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U5394 ( .A1(n4827), .A2(n4812), .ZN(U2939) );
  AOI22_X1 U5395 ( .A1(n4848), .A2(EAX_REG_6__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U5396 ( .A1(n4814), .A2(n4813), .ZN(U2945) );
  NAND2_X1 U5397 ( .A1(n4815), .A2(DATAI_13_), .ZN(n4831) );
  AOI22_X1 U5398 ( .A1(n4848), .A2(EAX_REG_29__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n4816) );
  NAND2_X1 U5399 ( .A1(n4831), .A2(n4816), .ZN(U2937) );
  AOI22_X1 U5400 ( .A1(n4848), .A2(EAX_REG_30__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n4817) );
  NAND2_X1 U5401 ( .A1(n4818), .A2(n4817), .ZN(U2938) );
  AOI22_X1 U5402 ( .A1(n4848), .A2(EAX_REG_28__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4819) );
  NAND2_X1 U5403 ( .A1(n4820), .A2(n4819), .ZN(U2936) );
  INV_X1 U5404 ( .A(DATAI_1_), .ZN(n4934) );
  OR2_X1 U5405 ( .A1(n4926), .A2(n4934), .ZN(n4835) );
  AOI22_X1 U5406 ( .A1(n4848), .A2(EAX_REG_1__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5407 ( .A1(n4835), .A2(n4821), .ZN(U2940) );
  AOI22_X1 U5408 ( .A1(n4848), .A2(EAX_REG_3__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U5409 ( .A1(n4823), .A2(n4822), .ZN(U2942) );
  AOI22_X1 U5410 ( .A1(n4848), .A2(EAX_REG_10__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U5411 ( .A1(n4825), .A2(n4824), .ZN(U2949) );
  AOI22_X1 U5412 ( .A1(n4848), .A2(EAX_REG_16__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U5413 ( .A1(n4827), .A2(n4826), .ZN(U2924) );
  AOI22_X1 U5414 ( .A1(n4848), .A2(EAX_REG_21__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U5415 ( .A1(n4829), .A2(n4828), .ZN(U2929) );
  AOI22_X1 U5416 ( .A1(n4848), .A2(EAX_REG_13__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5417 ( .A1(n4831), .A2(n4830), .ZN(U2952) );
  AOI22_X1 U5418 ( .A1(n4848), .A2(EAX_REG_4__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U5419 ( .A1(n4833), .A2(n4832), .ZN(U2943) );
  AOI22_X1 U5420 ( .A1(n4848), .A2(EAX_REG_17__SCAN_IN), .B1(n4847), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U5421 ( .A1(n4835), .A2(n4834), .ZN(U2925) );
  INV_X1 U5422 ( .A(n4836), .ZN(n4837) );
  NAND3_X1 U5423 ( .A1(n3722), .A2(n4837), .A3(n3730), .ZN(n4838) );
  INV_X1 U5424 ( .A(n4922), .ZN(n4839) );
  NAND2_X1 U5425 ( .A1(n4839), .A2(n4872), .ZN(n4840) );
  OR2_X1 U5426 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4843)
         );
  NAND2_X1 U5427 ( .A1(n4843), .A2(n4842), .ZN(n6340) );
  INV_X1 U5428 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4846) );
  XNOR2_X1 U5429 ( .A(n4845), .B(n4844), .ZN(n6170) );
  OAI222_X1 U5430 ( .A1(n6157), .A2(n6340), .B1(n4846), .B2(n6162), .C1(n5558), 
        .C2(n6170), .ZN(U2859) );
  INV_X1 U5431 ( .A(DATAI_15_), .ZN(n5971) );
  AOI22_X1 U5432 ( .A1(n4848), .A2(EAX_REG_15__SCAN_IN), .B1(n4847), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n4849) );
  OAI21_X1 U5433 ( .B1(n4926), .B2(n5971), .A(n4849), .ZN(U2954) );
  INV_X1 U5434 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U5435 ( .A1(n6322), .A2(REIP_REG_1__SCAN_IN), .ZN(n5061) );
  OAI221_X1 U5436 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6216), .C1(n4850), 
        .C2(n6209), .A(n5061), .ZN(n4859) );
  NAND2_X1 U5437 ( .A1(n4851), .A2(n4852), .ZN(n4854) );
  INV_X1 U5438 ( .A(n6165), .ZN(n4853) );
  XNOR2_X1 U5439 ( .A(n4854), .B(n4853), .ZN(n5071) );
  OR2_X1 U5440 ( .A1(n4856), .A2(n4855), .ZN(n4857) );
  NAND2_X1 U5441 ( .A1(n4936), .A2(n4857), .ZN(n5079) );
  OAI22_X1 U5442 ( .A1(n6535), .A2(n5071), .B1(n6188), .B2(n5079), .ZN(n4858)
         );
  OR2_X1 U5443 ( .A1(n4859), .A2(n4858), .ZN(U2985) );
  XNOR2_X1 U5444 ( .A(n4861), .B(n5055), .ZN(n4862) );
  XNOR2_X1 U5445 ( .A(n4860), .B(n4862), .ZN(n5060) );
  NAND2_X1 U5446 ( .A1(n4864), .A2(n4865), .ZN(n4866) );
  NAND2_X1 U5447 ( .A1(n4863), .A2(n4866), .ZN(n5050) );
  INV_X1 U5448 ( .A(n5050), .ZN(n4870) );
  AND2_X1 U5449 ( .A1(n6322), .A2(REIP_REG_3__SCAN_IN), .ZN(n5056) );
  INV_X1 U5450 ( .A(n5056), .ZN(n4868) );
  NAND2_X1 U5451 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4867)
         );
  OAI211_X1 U5452 ( .C1(n6216), .C2(n5037), .A(n4868), .B(n4867), .ZN(n4869)
         );
  AOI21_X1 U5453 ( .B1(n6211), .B2(n4870), .A(n4869), .ZN(n4871) );
  OAI21_X1 U5454 ( .B1(n5060), .B2(n6535), .A(n4871), .ZN(U2983) );
  OR2_X1 U5455 ( .A1(n5075), .A2(n4872), .ZN(n4873) );
  NAND2_X1 U5456 ( .A1(n4874), .A2(n4873), .ZN(n5065) );
  AOI22_X1 U5457 ( .A1(n6150), .A2(n5065), .B1(EBX_REG_1__SCAN_IN), .B2(n5531), 
        .ZN(n4875) );
  OAI21_X1 U5458 ( .B1(n5558), .B2(n5079), .A(n4875), .ZN(U2858) );
  INV_X1 U5459 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5715) );
  AOI22_X1 U5460 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n5066), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n5715), .ZN(n4876) );
  INV_X1 U5461 ( .A(n4876), .ZN(n5833) );
  OR2_X1 U5462 ( .A1(n6585), .A2(n6346), .ZN(n5834) );
  INV_X1 U5463 ( .A(n5834), .ZN(n4892) );
  NOR2_X1 U5464 ( .A1(n6590), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4891)
         );
  INV_X1 U5465 ( .A(n4879), .ZN(n4882) );
  AND3_X1 U5466 ( .A1(n3507), .A2(n5109), .A3(n4880), .ZN(n4881) );
  NAND2_X1 U5467 ( .A1(n4882), .A2(n4881), .ZN(n5831) );
  NAND2_X1 U5468 ( .A1(n3455), .A2(n5831), .ZN(n4890) );
  XNOR2_X1 U5469 ( .A(n4877), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4887)
         );
  INV_X1 U5470 ( .A(n6550), .ZN(n5322) );
  NAND2_X1 U5471 ( .A1(n5322), .A2(n3567), .ZN(n5829) );
  NAND2_X1 U5472 ( .A1(n5322), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4883) );
  MUX2_X1 U5473 ( .A(n5829), .B(n4883), .S(n3824), .Z(n4886) );
  INV_X1 U5474 ( .A(n4884), .ZN(n5364) );
  OR2_X1 U5475 ( .A1(n4894), .A2(n5364), .ZN(n5098) );
  NAND2_X1 U5476 ( .A1(n5098), .A2(n4887), .ZN(n4885) );
  OAI211_X1 U5477 ( .C1(n4607), .C2(n4887), .A(n4886), .B(n4885), .ZN(n4888)
         );
  INV_X1 U5478 ( .A(n4888), .ZN(n4889) );
  NAND2_X1 U5479 ( .A1(n4890), .A2(n4889), .ZN(n5087) );
  AOI222_X1 U5480 ( .A1(n5833), .A2(n4892), .B1(n4877), .B2(n4891), .C1(n5087), 
        .C2(n6580), .ZN(n4909) );
  NAND2_X1 U5481 ( .A1(n4758), .A2(n6221), .ZN(n4893) );
  OAI211_X1 U5482 ( .C1(n5322), .C2(n4569), .A(n4893), .B(n6619), .ZN(n4904)
         );
  NAND2_X1 U5483 ( .A1(n5365), .A2(n4894), .ZN(n4897) );
  INV_X1 U5484 ( .A(n5109), .ZN(n4895) );
  NAND3_X1 U5485 ( .A1(n4895), .A2(n5368), .A3(n6619), .ZN(n4896) );
  INV_X1 U5486 ( .A(n4924), .ZN(n4903) );
  AND2_X1 U5487 ( .A1(n4899), .A2(n4898), .ZN(n4900) );
  AND2_X1 U5488 ( .A1(n4901), .A2(n4900), .ZN(n4902) );
  NOR2_X1 U5489 ( .A1(n6797), .A2(n6585), .ZN(n6587) );
  NAND2_X1 U5490 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6587), .ZN(n6586) );
  INV_X1 U5491 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6536) );
  OAI22_X1 U5492 ( .A1(n6555), .A2(n6598), .B1(n6586), .B2(n6536), .ZN(n6547)
         );
  AOI21_X1 U5493 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6594), .A(n6547), .ZN(
        n6542) );
  INV_X1 U5494 ( .A(n4877), .ZN(n4907) );
  INV_X1 U5495 ( .A(n6590), .ZN(n4906) );
  AOI21_X1 U5496 ( .B1(n4907), .B2(n4906), .A(n6542), .ZN(n4908) );
  OAI22_X1 U5497 ( .A1(n4909), .A2(n6542), .B1(n4908), .B2(n3824), .ZN(U3459)
         );
  OR2_X1 U5498 ( .A1(n4912), .A2(n4911), .ZN(n4913) );
  NAND2_X1 U5499 ( .A1(n4910), .A2(n4913), .ZN(n6368) );
  NAND2_X1 U5500 ( .A1(n6156), .A2(n4914), .ZN(n4915) );
  AND2_X1 U5501 ( .A1(n4965), .A2(n4915), .ZN(n6365) );
  AOI22_X1 U5502 ( .A1(n6150), .A2(n6365), .B1(EBX_REG_5__SCAN_IN), .B2(n5531), 
        .ZN(n4916) );
  OAI21_X1 U5503 ( .B1(n6368), .B2(n5558), .A(n4916), .ZN(U2854) );
  INV_X1 U5504 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4920) );
  AOI21_X1 U5505 ( .B1(n3490), .B2(n5151), .A(n4918), .ZN(n4919) );
  OR2_X1 U5506 ( .A1(n4919), .A2(n6154), .ZN(n5041) );
  OAI222_X1 U5507 ( .A1(n5050), .A2(n5558), .B1(n4920), .B2(n6162), .C1(n5041), 
        .C2(n6157), .ZN(U2856) );
  NOR2_X1 U5508 ( .A1(n4922), .A2(n4921), .ZN(n4923) );
  OR2_X1 U5509 ( .A1(n4927), .A2(n3722), .ZN(n4928) );
  INV_X1 U5510 ( .A(n4928), .ZN(n4929) );
  INV_X1 U5511 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6051) );
  OAI222_X1 U5512 ( .A1(n6635), .A2(n6170), .B1(n5255), .B2(n4930), .C1(n5564), 
        .C2(n6051), .ZN(U2891) );
  INV_X1 U5513 ( .A(n4931), .ZN(n4932) );
  XNOR2_X1 U5514 ( .A(n4932), .B(n4863), .ZN(n6357) );
  INV_X1 U5515 ( .A(n6357), .ZN(n4933) );
  INV_X1 U5516 ( .A(DATAI_4_), .ZN(n5938) );
  INV_X1 U5517 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6059) );
  OAI222_X1 U5518 ( .A1(n6635), .A2(n4933), .B1(n5255), .B2(n5938), .C1(n5564), 
        .C2(n6059), .ZN(U2887) );
  INV_X1 U5519 ( .A(DATAI_3_), .ZN(n5839) );
  INV_X1 U5520 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6057) );
  OAI222_X1 U5521 ( .A1(n5050), .A2(n6635), .B1(n5255), .B2(n5839), .C1(n5564), 
        .C2(n6057), .ZN(U2888) );
  INV_X1 U5522 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6053) );
  OAI222_X1 U5523 ( .A1(n5079), .A2(n6635), .B1(n5255), .B2(n4934), .C1(n5564), 
        .C2(n6053), .ZN(U2890) );
  INV_X1 U5524 ( .A(DATAI_5_), .ZN(n5937) );
  OAI222_X1 U5525 ( .A1(n6368), .A2(n6635), .B1(n5255), .B2(n5937), .C1(n5564), 
        .C2(n4788), .ZN(U2886) );
  INV_X1 U5526 ( .A(n4936), .ZN(n4937) );
  OAI21_X1 U5527 ( .B1(n4935), .B2(n4937), .A(n4864), .ZN(n6146) );
  INV_X1 U5528 ( .A(DATAI_2_), .ZN(n5840) );
  INV_X1 U5529 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6055) );
  OAI222_X1 U5530 ( .A1(n6146), .A2(n6635), .B1(n5255), .B2(n5840), .C1(n5564), 
        .C2(n6055), .ZN(U2889) );
  OR2_X1 U5531 ( .A1(n4938), .A2(n5126), .ZN(n4985) );
  INV_X1 U5532 ( .A(n4985), .ZN(n4940) );
  NAND2_X1 U5533 ( .A1(n4940), .A2(n4939), .ZN(n4950) );
  AND2_X1 U5534 ( .A1(n6808), .A2(n6817), .ZN(n6781) );
  AOI21_X1 U5535 ( .B1(n4950), .B2(n6211), .A(n6781), .ZN(n4946) );
  INV_X1 U5536 ( .A(n6713), .ZN(n6604) );
  AND2_X1 U5537 ( .A1(n3458), .A2(n6604), .ZN(n6690) );
  INV_X1 U5538 ( .A(n4942), .ZN(n6689) );
  NAND2_X1 U5539 ( .A1(n3455), .A2(n6689), .ZN(n6728) );
  INV_X1 U5540 ( .A(n6728), .ZN(n6715) );
  NOR2_X1 U5541 ( .A1(n4943), .A2(n5132), .ZN(n6994) );
  AOI21_X1 U5542 ( .B1(n6690), .B2(n6715), .A(n6994), .ZN(n4947) );
  INV_X1 U5543 ( .A(n4947), .ZN(n4945) );
  NAND2_X1 U5544 ( .A1(n6797), .A2(n6585), .ZN(n6591) );
  NAND3_X1 U5545 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4987) );
  NAND2_X1 U5546 ( .A1(n6768), .A2(n4987), .ZN(n4944) );
  OAI211_X1 U5547 ( .C1(n4946), .C2(n4945), .A(n6806), .B(n4944), .ZN(n6998)
         );
  INV_X1 U5548 ( .A(n6998), .ZN(n5280) );
  INV_X1 U5549 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U5550 ( .A1(DATAI_7_), .A2(n6680), .ZN(n7162) );
  OAI22_X1 U5551 ( .A1(n4947), .A2(n6768), .B1(n4987), .B2(n6797), .ZN(n6995)
         );
  INV_X1 U5552 ( .A(DATAI_23_), .ZN(n4948) );
  OR2_X1 U5553 ( .A1(n6188), .A2(n4948), .ZN(n7175) );
  NOR2_X2 U5554 ( .A1(n5274), .A2(n3722), .ZN(n7165) );
  NOR2_X2 U5555 ( .A1(n4950), .A2(n6799), .ZN(n6997) );
  INV_X1 U5556 ( .A(DATAI_31_), .ZN(n4951) );
  OR2_X1 U5557 ( .A1(n6188), .A2(n4951), .ZN(n7148) );
  INV_X1 U5558 ( .A(n7148), .ZN(n7170) );
  AOI22_X1 U5559 ( .A1(n7165), .A2(n6994), .B1(n6997), .B2(n7170), .ZN(n4952)
         );
  OAI21_X1 U5560 ( .B1(n7175), .B2(n7001), .A(n4952), .ZN(n4953) );
  AOI21_X1 U5561 ( .B1(n7167), .B2(n6995), .A(n4953), .ZN(n4954) );
  OAI21_X1 U5562 ( .B1(n5280), .B2(n4955), .A(n4954), .ZN(U3147) );
  INV_X1 U5563 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4960) );
  NAND2_X1 U5564 ( .A1(DATAI_0_), .A2(n6680), .ZN(n6811) );
  INV_X1 U5565 ( .A(DATAI_16_), .ZN(n5969) );
  OR2_X1 U5566 ( .A1(n6188), .A2(n5969), .ZN(n6792) );
  NOR2_X2 U5567 ( .A1(n5274), .A2(n3528), .ZN(n6827) );
  INV_X1 U5568 ( .A(DATAI_24_), .ZN(n4956) );
  OR2_X1 U5569 ( .A1(n6188), .A2(n4956), .ZN(n6764) );
  INV_X1 U5570 ( .A(n6764), .ZN(n6829) );
  AOI22_X1 U5571 ( .A1(n6827), .A2(n6994), .B1(n6997), .B2(n6829), .ZN(n4957)
         );
  OAI21_X1 U5572 ( .B1(n6792), .B2(n7001), .A(n4957), .ZN(n4958) );
  AOI21_X1 U5573 ( .B1(n6828), .B2(n6995), .A(n4958), .ZN(n4959) );
  OAI21_X1 U5574 ( .B1(n5280), .B2(n4960), .A(n4959), .ZN(U3140) );
  NAND2_X1 U5575 ( .A1(n4910), .A2(n4962), .ZN(n4963) );
  AND2_X1 U5576 ( .A1(n4961), .A2(n4963), .ZN(n6385) );
  INV_X1 U5577 ( .A(n6385), .ZN(n5018) );
  NAND2_X1 U5578 ( .A1(n4965), .A2(n4964), .ZN(n4966) );
  AND2_X1 U5579 ( .A1(n5138), .A2(n4966), .ZN(n6379) );
  AOI22_X1 U5580 ( .A1(n6150), .A2(n6379), .B1(EBX_REG_6__SCAN_IN), .B2(n5531), 
        .ZN(n4967) );
  OAI21_X1 U5581 ( .B1(n5018), .B2(n5558), .A(n4967), .ZN(U2853) );
  AOI22_X1 U5582 ( .A1(n6228), .A2(UWORD_REG_12__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4968) );
  OAI21_X1 U5583 ( .B1(n4334), .B2(n4983), .A(n4968), .ZN(U2895) );
  AOI22_X1 U5584 ( .A1(n6228), .A2(UWORD_REG_13__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4969) );
  OAI21_X1 U5585 ( .B1(n4360), .B2(n4983), .A(n4969), .ZN(U2894) );
  INV_X1 U5586 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4971) );
  AOI22_X1 U5587 ( .A1(n6228), .A2(UWORD_REG_14__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4970) );
  OAI21_X1 U5588 ( .B1(n4971), .B2(n4983), .A(n4970), .ZN(U2893) );
  INV_X1 U5589 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U5590 ( .A1(n6228), .A2(UWORD_REG_1__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4972) );
  OAI21_X1 U5591 ( .B1(n4973), .B2(n4983), .A(n4972), .ZN(U2906) );
  AOI22_X1 U5592 ( .A1(n6228), .A2(UWORD_REG_2__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4974) );
  OAI21_X1 U5593 ( .B1(n4975), .B2(n4983), .A(n4974), .ZN(U2905) );
  AOI22_X1 U5594 ( .A1(n6228), .A2(UWORD_REG_3__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4976) );
  OAI21_X1 U5595 ( .B1(n4792), .B2(n4983), .A(n4976), .ZN(U2904) );
  AOI22_X1 U5596 ( .A1(n6228), .A2(UWORD_REG_11__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4977) );
  OAI21_X1 U5597 ( .B1(n4795), .B2(n4983), .A(n4977), .ZN(U2896) );
  INV_X1 U5598 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4979) );
  AOI22_X1 U5599 ( .A1(n6228), .A2(UWORD_REG_4__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4978) );
  OAI21_X1 U5600 ( .B1(n4979), .B2(n4983), .A(n4978), .ZN(U2903) );
  INV_X1 U5601 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U5602 ( .A1(n6228), .A2(UWORD_REG_10__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4980) );
  OAI21_X1 U5603 ( .B1(n4981), .B2(n4983), .A(n4980), .ZN(U2897) );
  INV_X1 U5604 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4984) );
  AOI22_X1 U5605 ( .A1(n6228), .A2(UWORD_REG_0__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4982) );
  OAI21_X1 U5606 ( .B1(n4984), .B2(n4983), .A(n4982), .ZN(U2907) );
  NAND2_X1 U5607 ( .A1(n6728), .A2(n6808), .ZN(n6730) );
  INV_X1 U5608 ( .A(n7084), .ZN(n7038) );
  AOI211_X1 U5609 ( .C1(n6825), .C2(n6730), .A(n6997), .B(n7038), .ZN(n4986)
         );
  AOI21_X1 U5610 ( .B1(n6728), .B2(n6781), .A(n4986), .ZN(n4992) );
  NOR2_X1 U5611 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4987), .ZN(n5281)
         );
  INV_X1 U5612 ( .A(n5281), .ZN(n4990) );
  OR2_X1 U5613 ( .A1(n6727), .A2(n5132), .ZN(n6684) );
  INV_X1 U5614 ( .A(n6684), .ZN(n4988) );
  NOR2_X1 U5615 ( .A1(n4988), .A2(n6797), .ZN(n6681) );
  INV_X1 U5616 ( .A(n4993), .ZN(n4989) );
  NAND2_X1 U5617 ( .A1(n4989), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U5618 ( .A1(n6680), .A2(n6823), .ZN(n6755) );
  AOI211_X1 U5619 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4990), .A(n6681), .B(
        n6755), .ZN(n4991) );
  INV_X1 U5620 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U5621 ( .A1(DATAI_1_), .A2(n6680), .ZN(n6872) );
  NAND2_X1 U5622 ( .A1(n3458), .A2(n6808), .ZN(n6815) );
  NAND2_X1 U5623 ( .A1(n4993), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6751) );
  OAI22_X1 U5624 ( .A1(n6815), .A2(n6728), .B1(n6684), .B2(n6751), .ZN(n5284)
         );
  INV_X1 U5625 ( .A(DATAI_25_), .ZN(n4994) );
  OR2_X1 U5626 ( .A1(n6188), .A2(n4994), .ZN(n6860) );
  NOR2_X2 U5627 ( .A1(n5274), .A2(n3725), .ZN(n6873) );
  INV_X1 U5628 ( .A(DATAI_17_), .ZN(n5965) );
  OR2_X1 U5629 ( .A1(n6188), .A2(n5965), .ZN(n6869) );
  INV_X1 U5630 ( .A(n6869), .ZN(n6876) );
  AOI22_X1 U5631 ( .A1(n6873), .A2(n5281), .B1(n6997), .B2(n6876), .ZN(n4995)
         );
  OAI21_X1 U5632 ( .B1(n7084), .B2(n6860), .A(n4995), .ZN(n4996) );
  AOI21_X1 U5633 ( .B1(n6874), .B2(n5284), .A(n4996), .ZN(n4997) );
  OAI21_X1 U5634 ( .B1(n5287), .B2(n4998), .A(n4997), .ZN(U3133) );
  INV_X1 U5635 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U5636 ( .A1(DATAI_3_), .A2(n6680), .ZN(n6948) );
  INV_X1 U5637 ( .A(DATAI_27_), .ZN(n4999) );
  OR2_X1 U5638 ( .A1(n6188), .A2(n4999), .ZN(n6918) );
  NOR2_X2 U5639 ( .A1(n5274), .A2(n5000), .ZN(n6949) );
  INV_X1 U5640 ( .A(DATAI_19_), .ZN(n5959) );
  OR2_X1 U5641 ( .A1(n6188), .A2(n5959), .ZN(n6945) );
  INV_X1 U5642 ( .A(n6945), .ZN(n6952) );
  AOI22_X1 U5643 ( .A1(n6949), .A2(n5281), .B1(n6997), .B2(n6952), .ZN(n5001)
         );
  OAI21_X1 U5644 ( .B1(n7084), .B2(n6918), .A(n5001), .ZN(n5002) );
  AOI21_X1 U5645 ( .B1(n6950), .B2(n5284), .A(n5002), .ZN(n5003) );
  OAI21_X1 U5646 ( .B1(n5287), .B2(n5004), .A(n5003), .ZN(U3135) );
  INV_X1 U5647 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5008) );
  INV_X1 U5648 ( .A(n7175), .ZN(n7155) );
  AOI22_X1 U5649 ( .A1(n7165), .A2(n5281), .B1(n6997), .B2(n7155), .ZN(n5005)
         );
  OAI21_X1 U5650 ( .B1(n7084), .B2(n7148), .A(n5005), .ZN(n5006) );
  AOI21_X1 U5651 ( .B1(n7167), .B2(n5284), .A(n5006), .ZN(n5007) );
  OAI21_X1 U5652 ( .B1(n5287), .B2(n5008), .A(n5007), .ZN(U3139) );
  INV_X1 U5653 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U5654 ( .A1(DATAI_2_), .A2(n6680), .ZN(n6910) );
  INV_X1 U5655 ( .A(DATAI_26_), .ZN(n5944) );
  OR2_X1 U5656 ( .A1(n6188), .A2(n5944), .ZN(n6880) );
  INV_X1 U5657 ( .A(DATAI_18_), .ZN(n5956) );
  OR2_X1 U5658 ( .A1(n6188), .A2(n5956), .ZN(n6907) );
  INV_X1 U5659 ( .A(n6907), .ZN(n6914) );
  AOI22_X1 U5660 ( .A1(n6911), .A2(n5281), .B1(n6997), .B2(n6914), .ZN(n5010)
         );
  OAI21_X1 U5661 ( .B1(n7084), .B2(n6880), .A(n5010), .ZN(n5011) );
  AOI21_X1 U5662 ( .B1(n6912), .B2(n5284), .A(n5011), .ZN(n5012) );
  OAI21_X1 U5663 ( .B1(n5287), .B2(n5013), .A(n5012), .ZN(U3134) );
  INV_X1 U5664 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5017) );
  INV_X1 U5665 ( .A(n6792), .ZN(n6830) );
  AOI22_X1 U5666 ( .A1(n6827), .A2(n5281), .B1(n6997), .B2(n6830), .ZN(n5014)
         );
  OAI21_X1 U5667 ( .B1(n7084), .B2(n6764), .A(n5014), .ZN(n5015) );
  AOI21_X1 U5668 ( .B1(n6828), .B2(n5284), .A(n5015), .ZN(n5016) );
  OAI21_X1 U5669 ( .B1(n5287), .B2(n5017), .A(n5016), .ZN(U3132) );
  INV_X1 U5670 ( .A(DATAI_6_), .ZN(n5987) );
  OAI222_X1 U5671 ( .A1(n5018), .A2(n6635), .B1(n5255), .B2(n5987), .C1(n5564), 
        .C2(n3969), .ZN(U2885) );
  NAND3_X1 U5672 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6232), .ZN(n6596) );
  INV_X1 U5673 ( .A(n6596), .ZN(n5023) );
  NAND2_X1 U5674 ( .A1(n5020), .A2(n5019), .ZN(n6583) );
  INV_X1 U5675 ( .A(n6583), .ZN(n5021) );
  NOR2_X1 U5676 ( .A1(n5035), .A2(n6585), .ZN(n5024) );
  NAND2_X1 U5677 ( .A1(n5025), .A2(n6490), .ZN(n6369) );
  INV_X1 U5678 ( .A(n6369), .ZN(n5159) );
  INV_X1 U5679 ( .A(n6221), .ZN(n5026) );
  NAND2_X1 U5680 ( .A1(n5370), .A2(n5026), .ZN(n5027) );
  NOR2_X1 U5681 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n5039) );
  INV_X1 U5682 ( .A(n5039), .ZN(n5031) );
  AOI21_X1 U5683 ( .B1(n5338), .B2(n5027), .A(n5031), .ZN(n5028) );
  NAND2_X1 U5684 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5154) );
  INV_X1 U5685 ( .A(n5154), .ZN(n5030) );
  NAND2_X1 U5686 ( .A1(n5030), .A2(REIP_REG_3__SCAN_IN), .ZN(n6350) );
  INV_X1 U5687 ( .A(n6350), .ZN(n5228) );
  OAI21_X1 U5688 ( .B1(n6521), .B2(n5228), .A(n6402), .ZN(n6349) );
  AND2_X1 U5689 ( .A1(n6350), .A2(n5030), .ZN(n5034) );
  OR2_X1 U5690 ( .A1(n6221), .A2(n5031), .ZN(n6575) );
  NAND2_X1 U5691 ( .A1(n4396), .A2(n6575), .ZN(n5352) );
  INV_X1 U5692 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5502) );
  NAND3_X1 U5693 ( .A1(n5370), .A2(n5502), .A3(n5031), .ZN(n5032) );
  AND2_X1 U5694 ( .A1(n5352), .A2(n5032), .ZN(n5033) );
  NOR2_X2 U5695 ( .A1(n5043), .A2(n5033), .ZN(n6506) );
  AOI22_X1 U5696 ( .A1(n6434), .A2(n5034), .B1(n6506), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5047) );
  AND2_X2 U5697 ( .A1(n6402), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6524) );
  AND2_X1 U5698 ( .A1(n5035), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5036) );
  INV_X1 U5699 ( .A(n5037), .ZN(n5038) );
  AOI22_X1 U5700 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6524), .B1(n6528), 
        .B2(n5038), .ZN(n5046) );
  NOR2_X1 U5701 ( .A1(n5043), .A2(n5502), .ZN(n5350) );
  NOR2_X1 U5702 ( .A1(n5338), .A2(n5039), .ZN(n5040) );
  INV_X1 U5703 ( .A(n5041), .ZN(n5057) );
  NAND2_X1 U5704 ( .A1(n6526), .A2(n5057), .ZN(n5045) );
  NOR2_X1 U5705 ( .A1(n5043), .A2(n5042), .ZN(n6353) );
  NAND2_X1 U5706 ( .A1(n6353), .A2(n3458), .ZN(n5044) );
  NAND4_X1 U5707 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5048)
         );
  AOI21_X1 U5708 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6349), .A(n5048), .ZN(n5049)
         );
  OAI21_X1 U5709 ( .B1(n5159), .B2(n5050), .A(n5049), .ZN(U2824) );
  INV_X1 U5710 ( .A(n5176), .ZN(n5067) );
  OAI21_X1 U5711 ( .B1(n5051), .B2(n5054), .A(n5067), .ZN(n5052) );
  INV_X1 U5712 ( .A(n5052), .ZN(n6284) );
  OAI21_X1 U5713 ( .B1(n5053), .B2(n6288), .A(n6284), .ZN(n6269) );
  NAND2_X1 U5714 ( .A1(n6292), .A2(n5054), .ZN(n6268) );
  AOI22_X1 U5715 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n6269), .B1(n6276), 
        .B2(n5055), .ZN(n5059) );
  AOI21_X1 U5716 ( .B1(n6326), .B2(n5057), .A(n5056), .ZN(n5058) );
  OAI211_X1 U5717 ( .C1(n5060), .C2(n6334), .A(n5059), .B(n5058), .ZN(U3015)
         );
  INV_X1 U5718 ( .A(n5061), .ZN(n5064) );
  NOR3_X1 U5719 ( .A1(n5807), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5062), 
        .ZN(n5063) );
  AOI211_X1 U5720 ( .C1(n6326), .C2(n5065), .A(n5064), .B(n5063), .ZN(n5070)
         );
  OR2_X1 U5721 ( .A1(n6288), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6338)
         );
  AOI21_X1 U5722 ( .B1(n5067), .B2(n6338), .A(n5066), .ZN(n5068) );
  INV_X1 U5723 ( .A(n5068), .ZN(n5069) );
  OAI211_X1 U5724 ( .C1(n5071), .C2(n6334), .A(n5070), .B(n5069), .ZN(U3017)
         );
  NAND2_X1 U5725 ( .A1(n6506), .A2(EBX_REG_1__SCAN_IN), .ZN(n5073) );
  INV_X1 U5726 ( .A(n6402), .ZN(n5475) );
  AOI22_X1 U5727 ( .A1(n6524), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5475), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5072) );
  OAI211_X1 U5728 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6515), .A(n5073), 
        .B(n5072), .ZN(n5074) );
  AOI21_X1 U5729 ( .B1(n6526), .B2(n5075), .A(n5074), .ZN(n5078) );
  INV_X1 U5730 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5076) );
  AOI22_X1 U5731 ( .A1(n6434), .A2(n5076), .B1(n6353), .B2(n6689), .ZN(n5077)
         );
  OAI211_X1 U5732 ( .C1(n5159), .C2(n5079), .A(n5078), .B(n5077), .ZN(U2826)
         );
  NAND2_X1 U5733 ( .A1(n6521), .A2(n6402), .ZN(n5491) );
  INV_X1 U5734 ( .A(n6353), .ZN(n5081) );
  OAI21_X1 U5735 ( .B1(n6524), .B2(n6528), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5080) );
  OAI21_X1 U5736 ( .B1(n5081), .B2(n6713), .A(n5080), .ZN(n5082) );
  AOI21_X1 U5737 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5491), .A(n5082), .ZN(n5085)
         );
  INV_X1 U5738 ( .A(n6170), .ZN(n5083) );
  AOI22_X1 U5739 ( .A1(n6369), .A2(n5083), .B1(n6506), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5084) );
  OAI211_X1 U5740 ( .C1(n6510), .C2(n6340), .A(n5085), .B(n5084), .ZN(U2827)
         );
  AOI211_X1 U5741 ( .C1(n6585), .C2(n5101), .A(FLUSH_REG_SCAN_IN), .B(n4517), 
        .ZN(n5117) );
  NAND2_X1 U5742 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6536), .ZN(n5113) );
  INV_X1 U5743 ( .A(n5086), .ZN(n5112) );
  NAND2_X1 U5744 ( .A1(n5101), .A2(n5087), .ZN(n5089) );
  NAND2_X1 U5745 ( .A1(n6555), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5088) );
  INV_X1 U5746 ( .A(n6559), .ZN(n5104) );
  NAND2_X1 U5747 ( .A1(n3458), .A2(n5831), .ZN(n5100) );
  MUX2_X1 U5748 ( .A(n5090), .B(n6544), .S(n4877), .Z(n5091) );
  NOR2_X1 U5749 ( .A1(n5091), .A2(n5086), .ZN(n5097) );
  NAND2_X1 U5750 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5093) );
  INV_X1 U5751 ( .A(n5093), .ZN(n5092) );
  MUX2_X1 U5752 ( .A(n5093), .B(n5092), .S(n6544), .Z(n5095) );
  AOI21_X1 U5753 ( .B1(n4877), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3880), 
        .ZN(n5094) );
  NOR2_X1 U5754 ( .A1(n3459), .A2(n5094), .ZN(n6539) );
  OAI22_X1 U5755 ( .A1(n6550), .A2(n5095), .B1(n6539), .B2(n4607), .ZN(n5096)
         );
  AOI21_X1 U5756 ( .B1(n5098), .B2(n5097), .A(n5096), .ZN(n5099) );
  NAND2_X1 U5757 ( .A1(n5100), .A2(n5099), .ZN(n6538) );
  NAND2_X1 U5758 ( .A1(n5101), .A2(n6538), .ZN(n5103) );
  NAND2_X1 U5759 ( .A1(n6555), .A2(n6544), .ZN(n5102) );
  NAND2_X1 U5760 ( .A1(n5103), .A2(n5102), .ZN(n6560) );
  NAND3_X1 U5761 ( .A1(n5104), .A2(n6585), .A3(n6560), .ZN(n5111) );
  INV_X1 U5762 ( .A(n5105), .ZN(n5106) );
  NOR2_X1 U5763 ( .A1(n5107), .A2(n5106), .ZN(n5108) );
  XNOR2_X1 U5764 ( .A(n5108), .B(n4517), .ZN(n6352) );
  NOR2_X1 U5765 ( .A1(n5109), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U5766 ( .A1(n6352), .A2(n5110), .ZN(n6545) );
  OAI211_X1 U5767 ( .C1(n5113), .C2(n5112), .A(n5111), .B(n6545), .ZN(n5114)
         );
  OR2_X1 U5768 ( .A1(n5117), .A2(n5114), .ZN(n6569) );
  INV_X1 U5769 ( .A(n5115), .ZN(n5116) );
  OR2_X1 U5770 ( .A1(n5117), .A2(n5116), .ZN(n5118) );
  NAND2_X1 U5771 ( .A1(n6569), .A2(n5118), .ZN(n6588) );
  NAND2_X1 U5772 ( .A1(n6588), .A2(n6536), .ZN(n5120) );
  INV_X1 U5773 ( .A(n6586), .ZN(n5119) );
  NAND2_X1 U5774 ( .A1(n5120), .A2(n5119), .ZN(n5122) );
  NAND2_X1 U5775 ( .A1(n5122), .A2(n5121), .ZN(n6606) );
  NAND2_X1 U5776 ( .A1(n6606), .A2(n6808), .ZN(n6601) );
  NAND2_X1 U5777 ( .A1(n4939), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5123) );
  XNOR2_X1 U5778 ( .A(n4938), .B(n5123), .ZN(n5125) );
  INV_X1 U5779 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6734) );
  OAI21_X1 U5780 ( .B1(n6585), .B2(STATE2_REG_3__SCAN_IN), .A(n6606), .ZN(
        n6600) );
  INV_X1 U5781 ( .A(n3455), .ZN(n5124) );
  OAI222_X1 U5782 ( .A1(n6601), .A2(n5125), .B1(n6600), .B2(n5124), .C1(n6606), 
        .C2(n4482), .ZN(U3463) );
  NOR2_X1 U5783 ( .A1(n6718), .A2(n6817), .ZN(n6712) );
  INV_X1 U5784 ( .A(n6712), .ZN(n5129) );
  OAI21_X1 U5785 ( .B1(n4938), .B2(n6817), .A(n5127), .ZN(n5128) );
  NAND2_X1 U5786 ( .A1(n5129), .A2(n5128), .ZN(n5130) );
  AND2_X1 U5787 ( .A1(n6654), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6649) );
  NOR2_X1 U5788 ( .A1(n5130), .A2(n6649), .ZN(n5131) );
  OAI222_X1 U5789 ( .A1(n6606), .A2(n5132), .B1(n6600), .B2(n6785), .C1(n6601), 
        .C2(n5131), .ZN(U3462) );
  XNOR2_X1 U5790 ( .A(n4939), .B(STATEBS16_REG_SCAN_IN), .ZN(n5133) );
  AND2_X1 U5791 ( .A1(n4961), .A2(n5135), .ZN(n5136) );
  NOR2_X1 U5792 ( .A1(n5134), .A2(n5136), .ZN(n6397) );
  INV_X1 U5793 ( .A(n6397), .ZN(n5142) );
  AND2_X1 U5794 ( .A1(n5138), .A2(n5137), .ZN(n5139) );
  NOR2_X1 U5795 ( .A1(n5163), .A2(n5139), .ZN(n6391) );
  AOI22_X1 U5796 ( .A1(n6150), .A2(n6391), .B1(EBX_REG_7__SCAN_IN), .B2(n5531), 
        .ZN(n5140) );
  OAI21_X1 U5797 ( .B1(n5142), .B2(n5558), .A(n5140), .ZN(U2852) );
  OAI222_X1 U5798 ( .A1(n5142), .A2(n6635), .B1(n5255), .B2(n5141), .C1(n5564), 
        .C2(n4781), .ZN(U2884) );
  OAI21_X1 U5799 ( .B1(n5144), .B2(n5146), .A(n5145), .ZN(n5184) );
  INV_X1 U5800 ( .A(n5147), .ZN(n5148) );
  AOI21_X1 U5801 ( .B1(n5149), .B2(n5165), .A(n5148), .ZN(n6414) );
  AOI22_X1 U5802 ( .A1(n6150), .A2(n6414), .B1(EBX_REG_9__SCAN_IN), .B2(n5531), 
        .ZN(n5150) );
  OAI21_X1 U5803 ( .B1(n5184), .B2(n5558), .A(n5150), .ZN(U2850) );
  XNOR2_X1 U5804 ( .A(n4917), .B(n5151), .ZN(n6283) );
  AOI22_X1 U5805 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6524), .B1(n5475), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n5152) );
  OAI21_X1 U5806 ( .B1(n6515), .B2(n6177), .A(n5152), .ZN(n5153) );
  AOI21_X1 U5807 ( .B1(n6353), .B2(n3455), .A(n5153), .ZN(n5156) );
  OAI211_X1 U5808 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n6434), .B(n5154), .ZN(n5155) );
  OAI211_X1 U5809 ( .C1(n6533), .C2(n6148), .A(n5156), .B(n5155), .ZN(n5157)
         );
  AOI21_X1 U5810 ( .B1(n6526), .B2(n6283), .A(n5157), .ZN(n5158) );
  OAI21_X1 U5811 ( .B1(n5159), .B2(n6146), .A(n5158), .ZN(U2825) );
  INV_X1 U5812 ( .A(n5134), .ZN(n5161) );
  AOI21_X1 U5813 ( .B1(n3438), .B2(n5161), .A(n5144), .ZN(n6410) );
  INV_X1 U5814 ( .A(n6410), .ZN(n5173) );
  OR2_X1 U5815 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  NAND2_X1 U5816 ( .A1(n5165), .A2(n5164), .ZN(n6405) );
  INV_X1 U5817 ( .A(n6405), .ZN(n5166) );
  AOI22_X1 U5818 ( .A1(n6150), .A2(n5166), .B1(EBX_REG_8__SCAN_IN), .B2(n5531), 
        .ZN(n5167) );
  OAI21_X1 U5819 ( .B1(n5173), .B2(n5558), .A(n5167), .ZN(U2851) );
  XNOR2_X1 U5820 ( .A(n5168), .B(n5169), .ZN(n5209) );
  NAND2_X1 U5821 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5170)
         );
  NAND2_X1 U5822 ( .A1(n6322), .A2(REIP_REG_8__SCAN_IN), .ZN(n5202) );
  OAI211_X1 U5823 ( .C1(n6216), .C2(n6408), .A(n5170), .B(n5202), .ZN(n5171)
         );
  AOI21_X1 U5824 ( .B1(n6410), .B2(n6211), .A(n5171), .ZN(n5172) );
  OAI21_X1 U5825 ( .B1(n5209), .B2(n6535), .A(n5172), .ZN(U2978) );
  INV_X1 U5826 ( .A(DATAI_9_), .ZN(n5983) );
  INV_X1 U5827 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6067) );
  OAI222_X1 U5828 ( .A1(n5184), .A2(n6635), .B1(n5255), .B2(n5983), .C1(n5564), 
        .C2(n6067), .ZN(U2882) );
  INV_X1 U5829 ( .A(DATAI_8_), .ZN(n5940) );
  INV_X1 U5830 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6065) );
  OAI222_X1 U5831 ( .A1(n5173), .A2(n6635), .B1(n5255), .B2(n5940), .C1(n5564), 
        .C2(n6065), .ZN(U2883) );
  XNOR2_X1 U5832 ( .A(n5175), .B(n5174), .ZN(n5187) );
  OAI22_X1 U5833 ( .A1(n6269), .A2(n5177), .B1(n5176), .B2(n5817), .ZN(n6304)
         );
  OAI21_X1 U5834 ( .B1(n5203), .B2(n5807), .A(n6304), .ZN(n5217) );
  NAND4_X1 U5835 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6277), .A4(n6276), .ZN(n6301) );
  NOR2_X1 U5836 ( .A1(n5178), .A2(n6301), .ZN(n5197) );
  AOI22_X1 U5837 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n5217), .B1(n5197), 
        .B2(n5179), .ZN(n5181) );
  AND2_X1 U5838 ( .A1(n6322), .A2(REIP_REG_9__SCAN_IN), .ZN(n5183) );
  AOI21_X1 U5839 ( .B1(n6326), .B2(n6414), .A(n5183), .ZN(n5180) );
  OAI211_X1 U5840 ( .C1(n5187), .C2(n6334), .A(n5181), .B(n5180), .ZN(U3009)
         );
  AND2_X1 U5841 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5182)
         );
  AOI211_X1 U5842 ( .C1(n6206), .C2(n6418), .A(n5183), .B(n5182), .ZN(n5186)
         );
  INV_X1 U5843 ( .A(n5184), .ZN(n6419) );
  NAND2_X1 U5844 ( .A1(n6419), .A2(n6211), .ZN(n5185) );
  OAI211_X1 U5845 ( .C1(n5187), .C2(n6535), .A(n5186), .B(n5185), .ZN(U2977)
         );
  AND2_X1 U5846 ( .A1(n5145), .A2(n5189), .ZN(n5190) );
  OR2_X1 U5847 ( .A1(n5188), .A2(n5190), .ZN(n6427) );
  NAND2_X1 U5848 ( .A1(n5147), .A2(n5191), .ZN(n5192) );
  NAND2_X1 U5849 ( .A1(n5212), .A2(n5192), .ZN(n6423) );
  INV_X1 U5850 ( .A(n6423), .ZN(n5193) );
  AOI22_X1 U5851 ( .A1(n6150), .A2(n5193), .B1(EBX_REG_10__SCAN_IN), .B2(n5531), .ZN(n5194) );
  OAI21_X1 U5852 ( .B1(n6427), .B2(n5558), .A(n5194), .ZN(U2849) );
  XNOR2_X1 U5853 ( .A(n5196), .B(n5195), .ZN(n5226) );
  INV_X1 U5854 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6433) );
  OAI22_X1 U5855 ( .A1(n6339), .A2(n6423), .B1(n6433), .B2(n6262), .ZN(n5200)
         );
  OAI211_X1 U5856 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5197), .B(n5218), .ZN(n5198) );
  INV_X1 U5857 ( .A(n5198), .ZN(n5199) );
  AOI211_X1 U5858 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n5217), .A(n5200), .B(n5199), .ZN(n5201) );
  OAI21_X1 U5859 ( .B1(n5226), .B2(n6334), .A(n5201), .ZN(U3008) );
  INV_X1 U5860 ( .A(n6304), .ZN(n5207) );
  OAI21_X1 U5861 ( .B1(n6339), .B2(n6405), .A(n5202), .ZN(n5206) );
  AOI211_X1 U5862 ( .C1(n5204), .C2(n4459), .A(n5203), .B(n6301), .ZN(n5205)
         );
  AOI211_X1 U5863 ( .C1(n5207), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5206), 
        .B(n5205), .ZN(n5208) );
  OAI21_X1 U5864 ( .B1(n6334), .B2(n5209), .A(n5208), .ZN(U3010) );
  INV_X1 U5865 ( .A(DATAI_10_), .ZN(n5845) );
  INV_X1 U5866 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6069) );
  OAI222_X1 U5867 ( .A1(n6427), .A2(n6635), .B1(n5255), .B2(n5845), .C1(n5564), 
        .C2(n6069), .ZN(U2881) );
  OAI21_X1 U5868 ( .B1(n5188), .B2(n5211), .A(n5210), .ZN(n5241) );
  AOI21_X1 U5869 ( .B1(n5213), .B2(n5212), .A(n5232), .ZN(n6439) );
  AOI22_X1 U5870 ( .A1(n6150), .A2(n6439), .B1(EBX_REG_11__SCAN_IN), .B2(n5531), .ZN(n5214) );
  OAI21_X1 U5871 ( .B1(n5241), .B2(n5558), .A(n5214), .ZN(U2848) );
  INV_X1 U5872 ( .A(DATAI_11_), .ZN(n5844) );
  INV_X1 U5873 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6071) );
  OAI222_X1 U5874 ( .A1(n5241), .A2(n6635), .B1(n5255), .B2(n5844), .C1(n5564), 
        .C2(n6071), .ZN(U2880) );
  XNOR2_X1 U5875 ( .A(n5704), .B(n5250), .ZN(n5215) );
  XNOR2_X1 U5876 ( .A(n5216), .B(n5215), .ZN(n5244) );
  AOI21_X1 U5877 ( .B1(n5218), .B2(n5817), .A(n5217), .ZN(n5806) );
  INV_X1 U5878 ( .A(n5806), .ZN(n5816) );
  NAND2_X1 U5879 ( .A1(n5219), .A2(n6276), .ZN(n6320) );
  INV_X1 U5880 ( .A(n6320), .ZN(n5808) );
  AOI22_X1 U5881 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5816), .B1(n5808), .B2(n5250), .ZN(n5221) );
  AND2_X1 U5882 ( .A1(n6322), .A2(REIP_REG_11__SCAN_IN), .ZN(n5240) );
  AOI21_X1 U5883 ( .B1(n6326), .B2(n6439), .A(n5240), .ZN(n5220) );
  OAI211_X1 U5884 ( .C1(n5244), .C2(n6334), .A(n5221), .B(n5220), .ZN(U3007)
         );
  INV_X1 U5885 ( .A(n6427), .ZN(n5224) );
  AOI22_X1 U5886 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6322), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5222) );
  OAI21_X1 U5887 ( .B1(n6426), .B2(n6216), .A(n5222), .ZN(n5223) );
  AOI21_X1 U5888 ( .B1(n5224), .B2(n6211), .A(n5223), .ZN(n5225) );
  OAI21_X1 U5889 ( .B1(n5226), .B2(n6535), .A(n5225), .ZN(U2976) );
  XOR2_X1 U5890 ( .A(n5227), .B(n5210), .Z(n5260) );
  NAND2_X1 U5891 ( .A1(n5228), .A2(REIP_REG_4__SCAN_IN), .ZN(n6363) );
  INV_X1 U5892 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6362) );
  NOR2_X1 U5893 ( .A1(n6363), .A2(n6362), .ZN(n6377) );
  NAND4_X1 U5894 ( .A1(n6377), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n6415) );
  INV_X1 U5895 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6416) );
  NOR2_X1 U5896 ( .A1(n6415), .A2(n6416), .ZN(n6432) );
  NAND2_X1 U5897 ( .A1(n6432), .A2(REIP_REG_10__SCAN_IN), .ZN(n6440) );
  INV_X1 U5898 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6442) );
  NOR2_X1 U5899 ( .A1(n6440), .A2(n6442), .ZN(n5311) );
  OAI21_X1 U5900 ( .B1(n6521), .B2(n5311), .A(n6402), .ZN(n6454) );
  NAND2_X1 U5901 ( .A1(n6402), .A2(n5229), .ZN(n6455) );
  OAI22_X1 U5902 ( .A1(n5230), .A2(n6457), .B1(n4677), .B2(n6533), .ZN(n5235)
         );
  NAND2_X1 U5903 ( .A1(n6434), .A2(n5311), .ZN(n6465) );
  OR2_X1 U5904 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  NAND2_X1 U5905 ( .A1(n5295), .A2(n5233), .ZN(n5289) );
  OAI22_X1 U5906 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6465), .B1(n6510), .B2(
        n5289), .ZN(n5234) );
  NOR3_X1 U5907 ( .A1(n6499), .A2(n5235), .A3(n5234), .ZN(n5236) );
  OAI21_X1 U5908 ( .B1(n5258), .B2(n6515), .A(n5236), .ZN(n5237) );
  AOI21_X1 U5909 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6454), .A(n5237), .ZN(n5238) );
  OAI21_X1 U5910 ( .B1(n5288), .B2(n6490), .A(n5238), .ZN(U2815) );
  AND2_X1 U5911 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5239)
         );
  AOI211_X1 U5912 ( .C1(n6206), .C2(n6445), .A(n5240), .B(n5239), .ZN(n5243)
         );
  INV_X1 U5913 ( .A(n5241), .ZN(n6446) );
  NAND2_X1 U5914 ( .A1(n6446), .A2(n6211), .ZN(n5242) );
  OAI211_X1 U5915 ( .C1(n5244), .C2(n6535), .A(n5243), .B(n5242), .ZN(U2975)
         );
  NOR2_X1 U5916 ( .A1(n5245), .A2(n3486), .ZN(n5246) );
  XNOR2_X1 U5917 ( .A(n5247), .B(n5246), .ZN(n5262) );
  INV_X1 U5918 ( .A(n5248), .ZN(n5249) );
  OAI21_X1 U5919 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5249), .A(n5806), 
        .ZN(n5253) );
  NOR3_X1 U5920 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5250), .A3(n6320), 
        .ZN(n5252) );
  NAND2_X1 U5921 ( .A1(n6322), .A2(REIP_REG_12__SCAN_IN), .ZN(n5256) );
  OAI21_X1 U5922 ( .B1(n6339), .B2(n5289), .A(n5256), .ZN(n5251) );
  AOI211_X1 U5923 ( .C1(n5253), .C2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5252), .B(n5251), .ZN(n5254) );
  OAI21_X1 U5924 ( .B1(n5262), .B2(n6334), .A(n5254), .ZN(U3006) );
  INV_X1 U5925 ( .A(DATAI_12_), .ZN(n5978) );
  INV_X1 U5926 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6073) );
  OAI222_X1 U5927 ( .A1(n6635), .A2(n5288), .B1(n5255), .B2(n5978), .C1(n5564), 
        .C2(n6073), .ZN(U2879) );
  NAND2_X1 U5928 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5257)
         );
  OAI211_X1 U5929 ( .C1(n6216), .C2(n5258), .A(n5257), .B(n5256), .ZN(n5259)
         );
  AOI21_X1 U5930 ( .B1(n5260), .B2(n6211), .A(n5259), .ZN(n5261) );
  OAI21_X1 U5931 ( .B1(n5262), .B2(n6535), .A(n5261), .ZN(U2974) );
  INV_X1 U5932 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U5933 ( .A1(DATAI_5_), .A2(n6680), .ZN(n7030) );
  INV_X1 U5934 ( .A(DATAI_29_), .ZN(n5263) );
  OR2_X1 U5935 ( .A1(n6188), .A2(n5263), .ZN(n6996) );
  NOR2_X2 U5936 ( .A1(n5274), .A2(n5562), .ZN(n7031) );
  INV_X1 U5937 ( .A(DATAI_21_), .ZN(n5943) );
  OR2_X1 U5938 ( .A1(n6188), .A2(n5943), .ZN(n7027) );
  INV_X1 U5939 ( .A(n7027), .ZN(n7034) );
  AOI22_X1 U5940 ( .A1(n7031), .A2(n5281), .B1(n6997), .B2(n7034), .ZN(n5264)
         );
  OAI21_X1 U5941 ( .B1(n7084), .B2(n6996), .A(n5264), .ZN(n5265) );
  AOI21_X1 U5942 ( .B1(n7032), .B2(n5284), .A(n5265), .ZN(n5266) );
  OAI21_X1 U5943 ( .B1(n5287), .B2(n5267), .A(n5266), .ZN(U3137) );
  INV_X1 U5944 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U5945 ( .A1(DATAI_4_), .A2(n6680), .ZN(n6986) );
  INV_X1 U5946 ( .A(DATAI_28_), .ZN(n5268) );
  OR2_X1 U5947 ( .A1(n6188), .A2(n5268), .ZN(n6980) );
  NOR2_X2 U5948 ( .A1(n5274), .A2(n3763), .ZN(n6987) );
  INV_X1 U5949 ( .A(DATAI_20_), .ZN(n5958) );
  OR2_X1 U5950 ( .A1(n6188), .A2(n5958), .ZN(n6983) );
  INV_X1 U5951 ( .A(n6983), .ZN(n6990) );
  AOI22_X1 U5952 ( .A1(n6987), .A2(n5281), .B1(n6997), .B2(n6990), .ZN(n5269)
         );
  OAI21_X1 U5953 ( .B1(n7084), .B2(n6980), .A(n5269), .ZN(n5270) );
  AOI21_X1 U5954 ( .B1(n6988), .B2(n5284), .A(n5270), .ZN(n5271) );
  OAI21_X1 U5955 ( .B1(n5287), .B2(n5272), .A(n5271), .ZN(U3136) );
  INV_X1 U5956 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U5957 ( .A1(DATAI_6_), .A2(n6680), .ZN(n7070) );
  INV_X1 U5958 ( .A(DATAI_22_), .ZN(n5273) );
  OR2_X1 U5959 ( .A1(n6188), .A2(n5273), .ZN(n7067) );
  NOR2_X2 U5960 ( .A1(n5274), .A2(n3847), .ZN(n7071) );
  INV_X1 U5961 ( .A(DATAI_30_), .ZN(n5275) );
  OR2_X1 U5962 ( .A1(n6188), .A2(n5275), .ZN(n7064) );
  INV_X1 U5963 ( .A(n7064), .ZN(n7073) );
  AOI22_X1 U5964 ( .A1(n7071), .A2(n6994), .B1(n6997), .B2(n7073), .ZN(n5276)
         );
  OAI21_X1 U5965 ( .B1(n7067), .B2(n7001), .A(n5276), .ZN(n5277) );
  AOI21_X1 U5966 ( .B1(n7072), .B2(n6995), .A(n5277), .ZN(n5278) );
  OAI21_X1 U5967 ( .B1(n5280), .B2(n5279), .A(n5278), .ZN(U3146) );
  INV_X1 U5968 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5286) );
  INV_X1 U5969 ( .A(n7067), .ZN(n7074) );
  AOI22_X1 U5970 ( .A1(n7071), .A2(n5281), .B1(n6997), .B2(n7074), .ZN(n5282)
         );
  OAI21_X1 U5971 ( .B1(n7084), .B2(n7064), .A(n5282), .ZN(n5283) );
  AOI21_X1 U5972 ( .B1(n7072), .B2(n5284), .A(n5283), .ZN(n5285) );
  OAI21_X1 U5973 ( .B1(n5287), .B2(n5286), .A(n5285), .ZN(U3138) );
  OAI222_X1 U5974 ( .A1(n5289), .A2(n6157), .B1(n6162), .B2(n4677), .C1(n5558), 
        .C2(n5288), .ZN(U2847) );
  NAND2_X1 U5975 ( .A1(n5290), .A2(n5291), .ZN(n5292) );
  AND2_X1 U5976 ( .A1(n5293), .A2(n5292), .ZN(n6459) );
  INV_X1 U5977 ( .A(n6459), .ZN(n5298) );
  AOI22_X1 U5978 ( .A1(n5306), .A2(DATAI_13_), .B1(n6837), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5294) );
  OAI21_X1 U5979 ( .B1(n5298), .B2(n6635), .A(n5294), .ZN(U2878) );
  INV_X1 U5980 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5297) );
  INV_X1 U5981 ( .A(n5822), .ZN(n5309) );
  AOI21_X1 U5982 ( .B1(n5296), .B2(n5295), .A(n5309), .ZN(n6453) );
  INV_X1 U5983 ( .A(n6453), .ZN(n6249) );
  OAI222_X1 U5984 ( .A1(n5298), .A2(n5558), .B1(n5297), .B2(n6162), .C1(n6157), 
        .C2(n6249), .ZN(U2846) );
  OAI21_X1 U5985 ( .B1(n5299), .B2(n5301), .A(n5300), .ZN(n6149) );
  AOI22_X1 U5986 ( .A1(n5306), .A2(DATAI_14_), .B1(n6837), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5302) );
  OAI21_X1 U5987 ( .B1(n6149), .B2(n6635), .A(n5302), .ZN(U2877) );
  INV_X1 U5988 ( .A(n5300), .ZN(n5305) );
  OAI21_X1 U5989 ( .B1(n5305), .B2(n4109), .A(n5304), .ZN(n5702) );
  AOI22_X1 U5990 ( .A1(n5306), .A2(DATAI_15_), .B1(n6837), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5307) );
  OAI21_X1 U5991 ( .B1(n5702), .B2(n6635), .A(n5307), .ZN(U2876) );
  AOI21_X1 U5992 ( .B1(n5309), .B2(n5821), .A(n5308), .ZN(n5310) );
  NOR2_X1 U5993 ( .A1(n5310), .A2(n5552), .ZN(n6306) );
  INV_X1 U5994 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5559) );
  OAI22_X1 U5995 ( .A1(n6533), .A2(n5559), .B1(n5698), .B2(n6515), .ZN(n5315)
         );
  INV_X1 U5996 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6474) );
  NAND4_X1 U5997 ( .A1(n5311), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_14__SCAN_IN), .ZN(n5344) );
  INV_X1 U5998 ( .A(n5344), .ZN(n5488) );
  OR2_X1 U5999 ( .A1(n6521), .A2(n5488), .ZN(n5312) );
  AND2_X1 U6000 ( .A1(n5312), .A2(n6402), .ZN(n6477) );
  AOI21_X1 U6001 ( .B1(n6524), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6499), 
        .ZN(n5313) );
  NOR2_X1 U6002 ( .A1(n6521), .A2(n5344), .ZN(n5486) );
  NAND2_X1 U6003 ( .A1(n5486), .A2(n6474), .ZN(n6478) );
  OAI211_X1 U6004 ( .C1(n6474), .C2(n6477), .A(n5313), .B(n6478), .ZN(n5314)
         );
  AOI211_X1 U6005 ( .C1(n6306), .C2(n6526), .A(n5315), .B(n5314), .ZN(n5316)
         );
  OAI21_X1 U6006 ( .B1(n5702), .B2(n6490), .A(n5316), .ZN(U2812) );
  INV_X1 U6007 ( .A(n5831), .ZN(n5317) );
  OR2_X1 U6008 ( .A1(n6713), .A2(n5317), .ZN(n5320) );
  NAND2_X1 U6009 ( .A1(n5318), .A2(n3566), .ZN(n5319) );
  NAND2_X1 U6010 ( .A1(n5320), .A2(n5319), .ZN(n6552) );
  OAI22_X1 U6011 ( .A1(n6585), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6590), .ZN(n5321) );
  AOI21_X1 U6012 ( .B1(n6552), .B2(n6580), .A(n5321), .ZN(n5324) );
  AOI21_X1 U6013 ( .B1(n5322), .B2(n6580), .A(n6542), .ZN(n5323) );
  OAI22_X1 U6014 ( .A1(n5324), .A2(n6542), .B1(n5323), .B2(n3566), .ZN(U3461)
         );
  NAND3_X1 U6015 ( .A1(n5342), .A2(n3722), .A3(n5564), .ZN(n5326) );
  AND2_X1 U6016 ( .A1(n5564), .A2(n3555), .ZN(n6834) );
  AOI22_X1 U6017 ( .A1(n6834), .A2(DATAI_31_), .B1(n6837), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6018 ( .A1(n5326), .A2(n5325), .ZN(U2860) );
  OAI21_X1 U6019 ( .B1(n6209), .B2(n5328), .A(n5327), .ZN(n5332) );
  OAI21_X2 U6020 ( .B1(n3461), .B2(n5330), .A(n5329), .ZN(n5575) );
  NOR2_X1 U6021 ( .A1(n5575), .A2(n6188), .ZN(n5331) );
  OAI21_X1 U6022 ( .B1(n5334), .B2(n6535), .A(n5333), .ZN(U2959) );
  INV_X1 U6023 ( .A(n5387), .ZN(n5335) );
  MUX2_X1 U6024 ( .A(n5337), .B(n5336), .S(n5335), .Z(n5341) );
  OAI22_X1 U6025 ( .A1(n5339), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5338), .ZN(n5340) );
  NAND2_X1 U6026 ( .A1(n5342), .A2(n6530), .ZN(n5360) );
  NAND2_X1 U6027 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .ZN(
        n5356) );
  INV_X1 U6028 ( .A(n5356), .ZN(n5349) );
  INV_X1 U6029 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6108) );
  INV_X1 U6030 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6517) );
  NAND3_X1 U6031 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n5487) );
  NAND3_X1 U6032 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n5343) );
  NOR3_X1 U6033 ( .A1(n5344), .A2(n5487), .A3(n5343), .ZN(n5473) );
  NAND2_X1 U6034 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5473), .ZN(n6520) );
  NOR2_X1 U6035 ( .A1(n6517), .A2(n6520), .ZN(n5460) );
  NAND2_X1 U6036 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5460), .ZN(n5433) );
  NOR2_X1 U6037 ( .A1(n6108), .A2(n5433), .ZN(n5436) );
  NAND3_X1 U6038 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        n5436), .ZN(n5354) );
  INV_X1 U6039 ( .A(n5354), .ZN(n5345) );
  NAND2_X1 U6040 ( .A1(n6402), .A2(n5345), .ZN(n5346) );
  NAND2_X1 U6041 ( .A1(n5491), .A2(n5346), .ZN(n5416) );
  INV_X1 U6042 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6116) );
  INV_X1 U6043 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6111) );
  OR2_X1 U6044 ( .A1(n6116), .A2(n6111), .ZN(n5347) );
  NAND2_X1 U6045 ( .A1(n5491), .A2(n5347), .ZN(n5348) );
  OAI21_X1 U6046 ( .B1(n5349), .B2(n6521), .A(n5383), .ZN(n5380) );
  INV_X1 U6047 ( .A(n5350), .ZN(n5353) );
  OAI22_X1 U6048 ( .A1(n5353), .A2(n5352), .B1(n5351), .B2(n6457), .ZN(n5358)
         );
  OR2_X1 U6049 ( .A1(n6521), .A2(n5354), .ZN(n5406) );
  INV_X1 U6050 ( .A(n5406), .ZN(n5355) );
  NAND3_X1 U6051 ( .A1(n5355), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n5386) );
  NOR3_X1 U6052 ( .A1(n5386), .A2(REIP_REG_31__SCAN_IN), .A3(n5356), .ZN(n5357) );
  AOI211_X1 U6053 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5380), .A(n5358), .B(n5357), .ZN(n5359) );
  OAI211_X1 U6054 ( .C1(n5710), .C2(n6510), .A(n5360), .B(n5359), .ZN(U2796)
         );
  NOR2_X1 U6055 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  OR2_X1 U6056 ( .A1(n5365), .A2(n5363), .ZN(n5367) );
  NAND2_X1 U6057 ( .A1(n5365), .A2(n5364), .ZN(n5366) );
  OAI211_X1 U6058 ( .C1(n4586), .C2(n5368), .A(n5367), .B(n5366), .ZN(n6564)
         );
  NAND2_X1 U6059 ( .A1(n4396), .A2(n6221), .ZN(n5369) );
  OAI211_X1 U6060 ( .C1(n5371), .C2(n5370), .A(n5369), .B(n6619), .ZN(n6230)
         );
  NAND2_X1 U6061 ( .A1(n5372), .A2(n6230), .ZN(n6567) );
  AND2_X1 U6062 ( .A1(n6567), .A2(n6572), .ZN(n6537) );
  MUX2_X1 U6063 ( .A(MORE_REG_SCAN_IN), .B(n6564), .S(n6537), .Z(U3471) );
  INV_X1 U6064 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6030) );
  OAI21_X1 U6065 ( .B1(n5386), .B2(n6030), .A(n6118), .ZN(n5379) );
  INV_X1 U6066 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5503) );
  INV_X1 U6067 ( .A(n5374), .ZN(n5375) );
  AOI22_X1 U6068 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6524), .B1(n6528), 
        .B2(n5375), .ZN(n5376) );
  OAI21_X1 U6069 ( .B1(n6533), .B2(n5503), .A(n5376), .ZN(n5378) );
  AOI21_X1 U6070 ( .B1(n5382), .B2(n5395), .A(n5381), .ZN(n5596) );
  INV_X1 U6071 ( .A(n5596), .ZN(n5569) );
  INV_X1 U6072 ( .A(n5383), .ZN(n5402) );
  AOI22_X1 U6073 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6524), .B1(n6528), 
        .B2(n5595), .ZN(n5385) );
  NAND2_X1 U6074 ( .A1(n6506), .A2(EBX_REG_29__SCAN_IN), .ZN(n5384) );
  OAI211_X1 U6075 ( .C1(n5386), .C2(REIP_REG_29__SCAN_IN), .A(n5385), .B(n5384), .ZN(n5390) );
  OAI21_X1 U6076 ( .B1(n5393), .B2(n5388), .A(n5387), .ZN(n5726) );
  NOR2_X1 U6077 ( .A1(n5726), .A2(n6510), .ZN(n5389) );
  AOI211_X1 U6078 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5402), .A(n5390), .B(n5389), .ZN(n5391) );
  OAI21_X1 U6079 ( .B1(n5569), .B2(n6490), .A(n5391), .ZN(U2798) );
  AND2_X1 U6080 ( .A1(n3467), .A2(n5392), .ZN(n5394) );
  OR2_X1 U6081 ( .A1(n5394), .A2(n5393), .ZN(n5736) );
  INV_X1 U6082 ( .A(n5395), .ZN(n5396) );
  NAND2_X1 U6083 ( .A1(n5608), .A2(n6530), .ZN(n5404) );
  NAND2_X1 U6084 ( .A1(n6116), .A2(REIP_REG_27__SCAN_IN), .ZN(n5400) );
  AOI22_X1 U6085 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6524), .B1(n6528), 
        .B2(n5607), .ZN(n5399) );
  NAND2_X1 U6086 ( .A1(n6506), .A2(EBX_REG_28__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6087 ( .C1(n5406), .C2(n5400), .A(n5399), .B(n5398), .ZN(n5401)
         );
  AOI21_X1 U6088 ( .B1(n5402), .B2(REIP_REG_28__SCAN_IN), .A(n5401), .ZN(n5403) );
  OAI211_X1 U6089 ( .C1(n6510), .C2(n5736), .A(n5404), .B(n5403), .ZN(U2799)
         );
  AOI22_X1 U6090 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6524), .B1(
        EBX_REG_27__SCAN_IN), .B2(n6506), .ZN(n5405) );
  OAI221_X1 U6091 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5406), .C1(n6111), .C2(
        n5416), .A(n5405), .ZN(n5408) );
  NOR2_X1 U6092 ( .A1(n5506), .A2(n6510), .ZN(n5407) );
  AOI211_X1 U6093 ( .C1(n6528), .C2(n5409), .A(n5408), .B(n5407), .ZN(n5410)
         );
  OAI21_X1 U6094 ( .B1(n5575), .B2(n6490), .A(n5410), .ZN(U2800) );
  OR2_X1 U6095 ( .A1(n5426), .A2(n5411), .ZN(n5412) );
  NAND2_X1 U6096 ( .A1(n5413), .A2(n5412), .ZN(n5747) );
  INV_X1 U6097 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U6098 ( .A1(n5618), .A2(n6530), .ZN(n5425) );
  INV_X1 U6099 ( .A(n5416), .ZN(n5423) );
  NAND2_X1 U6100 ( .A1(n5436), .A2(REIP_REG_25__SCAN_IN), .ZN(n5418) );
  INV_X1 U6101 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5417) );
  OAI21_X1 U6102 ( .B1(n6521), .B2(n5418), .A(n5417), .ZN(n5422) );
  OAI22_X1 U6103 ( .A1(n5419), .A2(n6457), .B1(n6515), .B2(n5616), .ZN(n5421)
         );
  INV_X1 U6104 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5508) );
  NOR2_X1 U6105 ( .A1(n6533), .A2(n5508), .ZN(n5420) );
  AOI211_X1 U6106 ( .C1(n5423), .C2(n5422), .A(n5421), .B(n5420), .ZN(n5424)
         );
  OAI211_X1 U6107 ( .C1(n6510), .C2(n5747), .A(n5425), .B(n5424), .ZN(U2801)
         );
  INV_X1 U6108 ( .A(n5426), .ZN(n5431) );
  INV_X1 U6109 ( .A(n5446), .ZN(n5429) );
  INV_X1 U6110 ( .A(n5427), .ZN(n5428) );
  OAI21_X1 U6111 ( .B1(n5459), .B2(n5429), .A(n5428), .ZN(n5430) );
  NAND2_X1 U6112 ( .A1(n5431), .A2(n5430), .ZN(n6324) );
  INV_X1 U6113 ( .A(n5624), .ZN(n5432) );
  NAND2_X1 U6114 ( .A1(n5432), .A2(n6530), .ZN(n5443) );
  INV_X1 U6115 ( .A(n5433), .ZN(n5447) );
  NAND2_X1 U6116 ( .A1(n6402), .A2(n5447), .ZN(n5434) );
  NAND2_X1 U6117 ( .A1(n5491), .A2(n5434), .ZN(n5461) );
  INV_X1 U6118 ( .A(n5461), .ZN(n5441) );
  INV_X1 U6119 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5435) );
  AOI22_X1 U6120 ( .A1(n5436), .A2(n5435), .B1(REIP_REG_25__SCAN_IN), .B2(
        n6108), .ZN(n5439) );
  AOI22_X1 U6121 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6524), .B1(
        EBX_REG_25__SCAN_IN), .B2(n6506), .ZN(n5438) );
  NAND2_X1 U6122 ( .A1(n6528), .A2(n5627), .ZN(n5437) );
  OAI211_X1 U6123 ( .C1(n6521), .C2(n5439), .A(n5438), .B(n5437), .ZN(n5440)
         );
  AOI21_X1 U6124 ( .B1(n5441), .B2(REIP_REG_25__SCAN_IN), .A(n5440), .ZN(n5442) );
  OAI211_X1 U6125 ( .C1(n6324), .C2(n6510), .A(n5443), .B(n5442), .ZN(U2802)
         );
  INV_X1 U6126 ( .A(n5444), .ZN(n5455) );
  NOR2_X1 U6127 ( .A1(n3471), .A2(n3558), .ZN(n6836) );
  INV_X1 U6128 ( .A(n6836), .ZN(n5511) );
  XNOR2_X1 U6129 ( .A(n5459), .B(n5446), .ZN(n5757) );
  NAND3_X1 U6130 ( .A1(n6434), .A2(n6108), .A3(n5447), .ZN(n5449) );
  NAND2_X1 U6131 ( .A1(n6506), .A2(EBX_REG_24__SCAN_IN), .ZN(n5448) );
  OAI211_X1 U6132 ( .C1(n6515), .C2(n5635), .A(n5449), .B(n5448), .ZN(n5452)
         );
  INV_X1 U6133 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5450) );
  OAI22_X1 U6134 ( .A1(n5450), .A2(n6457), .B1(n6108), .B2(n5461), .ZN(n5451)
         );
  AOI211_X1 U6135 ( .C1(n6526), .C2(n5757), .A(n5452), .B(n5451), .ZN(n5453)
         );
  OAI21_X1 U6136 ( .B1(n5511), .B2(n6490), .A(n5453), .ZN(U2803) );
  INV_X1 U6137 ( .A(n3468), .ZN(n5513) );
  INV_X1 U6138 ( .A(n5454), .ZN(n5456) );
  OAI21_X1 U6139 ( .B1(n5513), .B2(n5456), .A(n5455), .ZN(n5646) );
  NAND2_X1 U6140 ( .A1(n5518), .A2(n5457), .ZN(n5458) );
  NAND2_X1 U6141 ( .A1(n5459), .A2(n5458), .ZN(n5761) );
  AOI21_X1 U6142 ( .B1(n6434), .B2(n5460), .A(REIP_REG_23__SCAN_IN), .ZN(n5462) );
  OAI22_X1 U6143 ( .A1(n5462), .A2(n5461), .B1(n5641), .B2(n6457), .ZN(n5463)
         );
  AOI21_X1 U6144 ( .B1(n6528), .B2(n5643), .A(n5463), .ZN(n5465) );
  NAND2_X1 U6145 ( .A1(n6506), .A2(EBX_REG_23__SCAN_IN), .ZN(n5464) );
  OAI211_X1 U6146 ( .C1(n5761), .C2(n6510), .A(n5465), .B(n5464), .ZN(n5466)
         );
  INV_X1 U6147 ( .A(n5466), .ZN(n5467) );
  OAI21_X1 U6148 ( .B1(n5646), .B2(n6490), .A(n5467), .ZN(U2804) );
  OAI21_X1 U6149 ( .B1(n5468), .B2(n5470), .A(n5469), .ZN(n5585) );
  OR2_X1 U6150 ( .A1(n5527), .A2(n5471), .ZN(n5472) );
  NAND2_X1 U6151 ( .A1(n5516), .A2(n5472), .ZN(n5780) );
  INV_X1 U6152 ( .A(n5780), .ZN(n5479) );
  INV_X1 U6153 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6041) );
  NAND3_X1 U6154 ( .A1(n6434), .A2(n5473), .A3(n6041), .ZN(n6519) );
  INV_X1 U6155 ( .A(n5473), .ZN(n5474) );
  OAI21_X1 U6156 ( .B1(n5475), .B2(n5474), .A(n5491), .ZN(n6518) );
  OAI22_X1 U6157 ( .A1(n5521), .A2(n6533), .B1(n6041), .B2(n6518), .ZN(n5476)
         );
  AOI21_X1 U6158 ( .B1(n6524), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5476), 
        .ZN(n5477) );
  OAI211_X1 U6159 ( .C1(n6515), .C2(n5657), .A(n6519), .B(n5477), .ZN(n5478)
         );
  AOI21_X1 U6160 ( .B1(n5479), .B2(n6526), .A(n5478), .ZN(n5480) );
  OAI21_X1 U6161 ( .B1(n5585), .B2(n6490), .A(n5480), .ZN(U2806) );
  AOI21_X1 U6162 ( .B1(n5483), .B2(n5481), .A(n5482), .ZN(n5484) );
  INV_X1 U6163 ( .A(n5484), .ZN(n5677) );
  AOI21_X1 U6164 ( .B1(n5485), .B2(n5538), .A(n5525), .ZN(n6237) );
  INV_X1 U6165 ( .A(n5674), .ZN(n5494) );
  INV_X1 U6166 ( .A(n5486), .ZN(n6475) );
  NOR2_X1 U6167 ( .A1(n6475), .A2(n5487), .ZN(n5495) );
  INV_X1 U6168 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U6169 ( .A1(n5495), .A2(n6496), .ZN(n6500) );
  INV_X1 U6170 ( .A(n5487), .ZN(n5489) );
  NAND3_X1 U6171 ( .A1(n6402), .A2(n5489), .A3(n5488), .ZN(n5490) );
  NAND2_X1 U6172 ( .A1(n5491), .A2(n5490), .ZN(n6495) );
  NAND2_X1 U6173 ( .A1(n6500), .A2(n6495), .ZN(n5492) );
  AOI21_X1 U6174 ( .B1(n5492), .B2(REIP_REG_19__SCAN_IN), .A(n6499), .ZN(n5493) );
  OAI21_X1 U6175 ( .B1(n5494), .B2(n6515), .A(n5493), .ZN(n5500) );
  INV_X1 U6176 ( .A(n5495), .ZN(n5496) );
  NOR2_X1 U6177 ( .A1(n5496), .A2(n6496), .ZN(n6508) );
  INV_X1 U6178 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6100) );
  AOI22_X1 U6179 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6524), .B1(n6508), 
        .B2(n6100), .ZN(n5497) );
  OAI21_X1 U6180 ( .B1(n5498), .B2(n6533), .A(n5497), .ZN(n5499) );
  AOI211_X1 U6181 ( .C1(n6237), .C2(n6526), .A(n5500), .B(n5499), .ZN(n5501)
         );
  OAI21_X1 U6182 ( .B1(n5677), .B2(n6490), .A(n5501), .ZN(U2808) );
  OAI22_X1 U6183 ( .A1(n5710), .A2(n6157), .B1(n6162), .B2(n5502), .ZN(U2828)
         );
  OAI222_X1 U6184 ( .A1(n5373), .A2(n5558), .B1(n5503), .B2(n6162), .C1(n6157), 
        .C2(n5377), .ZN(U2829) );
  OAI222_X1 U6185 ( .A1(n5558), .A2(n5569), .B1(n5504), .B2(n6162), .C1(n5726), 
        .C2(n6157), .ZN(U2830) );
  INV_X1 U6186 ( .A(n5608), .ZN(n5572) );
  OAI222_X1 U6187 ( .A1(n5558), .A2(n5572), .B1(n5505), .B2(n6162), .C1(n5736), 
        .C2(n6157), .ZN(U2831) );
  INV_X1 U6188 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5507) );
  OAI222_X1 U6189 ( .A1(n5558), .A2(n5575), .B1(n5507), .B2(n6162), .C1(n5506), 
        .C2(n6157), .ZN(U2832) );
  INV_X1 U6190 ( .A(n5618), .ZN(n5578) );
  OAI222_X1 U6191 ( .A1(n6157), .A2(n5747), .B1(n5508), .B2(n6162), .C1(n5578), 
        .C2(n5558), .ZN(U2833) );
  INV_X1 U6192 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5509) );
  OAI222_X1 U6193 ( .A1(n5558), .A2(n5624), .B1(n5509), .B2(n6162), .C1(n6324), 
        .C2(n6157), .ZN(U2834) );
  AOI22_X1 U6194 ( .A1(n5757), .A2(n6150), .B1(EBX_REG_24__SCAN_IN), .B2(n5531), .ZN(n5510) );
  OAI21_X1 U6195 ( .B1(n5511), .B2(n5558), .A(n5510), .ZN(U2835) );
  INV_X1 U6196 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5512) );
  OAI222_X1 U6197 ( .A1(n5558), .A2(n5646), .B1(n5512), .B2(n6162), .C1(n5761), 
        .C2(n6157), .ZN(U2836) );
  AOI21_X1 U6198 ( .B1(n5514), .B2(n5469), .A(n5513), .ZN(n6646) );
  INV_X1 U6199 ( .A(n5558), .ZN(n6159) );
  NAND2_X1 U6200 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U6201 ( .A1(n5518), .A2(n5517), .ZN(n6525) );
  OAI22_X1 U6202 ( .A1(n6525), .A2(n6157), .B1(n6534), .B2(n6162), .ZN(n5519)
         );
  AOI21_X1 U6203 ( .B1(n6646), .B2(n6159), .A(n5519), .ZN(n5520) );
  INV_X1 U6204 ( .A(n5520), .ZN(U2837) );
  INV_X1 U6205 ( .A(n5585), .ZN(n5659) );
  OAI22_X1 U6206 ( .A1(n5780), .A2(n6157), .B1(n5521), .B2(n6162), .ZN(n5522)
         );
  AOI21_X1 U6207 ( .B1(n5659), .B2(n6159), .A(n5522), .ZN(n5523) );
  INV_X1 U6208 ( .A(n5523), .ZN(U2838) );
  NOR2_X1 U6209 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  OR2_X1 U6210 ( .A1(n5527), .A2(n5526), .ZN(n6511) );
  NOR2_X1 U6211 ( .A1(n5482), .A2(n5528), .ZN(n5529) );
  OR2_X1 U6212 ( .A1(n5468), .A2(n5529), .ZN(n6507) );
  OAI222_X1 U6213 ( .A1(n6157), .A2(n6511), .B1(n5530), .B2(n6162), .C1(n6507), 
        .C2(n5558), .ZN(U2839) );
  AOI22_X1 U6214 ( .A1(n6237), .A2(n6150), .B1(EBX_REG_19__SCAN_IN), .B2(n5531), .ZN(n5532) );
  OAI21_X1 U6215 ( .B1(n5677), .B2(n5558), .A(n5532), .ZN(U2840) );
  NAND2_X1 U6216 ( .A1(n5544), .A2(n5534), .ZN(n5535) );
  AND2_X1 U6217 ( .A1(n5481), .A2(n5535), .ZN(n6640) );
  NAND2_X1 U6218 ( .A1(n5547), .A2(n5536), .ZN(n5537) );
  NAND2_X1 U6219 ( .A1(n5538), .A2(n5537), .ZN(n6505) );
  OAI22_X1 U6220 ( .A1(n6505), .A2(n6157), .B1(n6497), .B2(n6162), .ZN(n5539)
         );
  AOI21_X1 U6221 ( .B1(n6640), .B2(n6159), .A(n5539), .ZN(n5540) );
  INV_X1 U6222 ( .A(n5540), .ZN(U2841) );
  OR2_X1 U6223 ( .A1(n5541), .A2(n5542), .ZN(n5543) );
  NAND2_X1 U6224 ( .A1(n5544), .A2(n5543), .ZN(n6636) );
  INV_X1 U6225 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5548) );
  OR2_X1 U6226 ( .A1(n5554), .A2(n5545), .ZN(n5546) );
  AND2_X1 U6227 ( .A1(n5547), .A2(n5546), .ZN(n6315) );
  INV_X1 U6228 ( .A(n6315), .ZN(n6489) );
  OAI222_X1 U6229 ( .A1(n6636), .A2(n5558), .B1(n5548), .B2(n6162), .C1(n6489), 
        .C2(n6157), .ZN(U2842) );
  AND2_X1 U6230 ( .A1(n5304), .A2(n5549), .ZN(n5550) );
  NOR2_X1 U6231 ( .A1(n5541), .A2(n5550), .ZN(n6631) );
  NOR2_X1 U6232 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  OR2_X1 U6233 ( .A1(n5554), .A2(n5553), .ZN(n6484) );
  OAI22_X1 U6234 ( .A1(n6157), .A2(n6484), .B1(n5555), .B2(n6162), .ZN(n5556)
         );
  AOI21_X1 U6235 ( .B1(n6631), .B2(n6159), .A(n5556), .ZN(n5557) );
  INV_X1 U6236 ( .A(n5557), .ZN(U2843) );
  INV_X1 U6237 ( .A(n6306), .ZN(n5560) );
  OAI222_X1 U6238 ( .A1(n5560), .A2(n6157), .B1(n5559), .B2(n6162), .C1(n5702), 
        .C2(n5558), .ZN(U2844) );
  AOI22_X1 U6239 ( .A1(n6834), .A2(DATAI_30_), .B1(n6837), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5566) );
  AND2_X1 U6240 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U6241 ( .A1(n6838), .A2(DATAI_14_), .ZN(n5565) );
  OAI211_X1 U6242 ( .C1(n5373), .C2(n6635), .A(n5566), .B(n5565), .ZN(U2861)
         );
  AOI22_X1 U6243 ( .A1(n6834), .A2(DATAI_29_), .B1(n6837), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U6244 ( .A1(n6838), .A2(DATAI_13_), .ZN(n5567) );
  OAI211_X1 U6245 ( .C1(n5569), .C2(n6635), .A(n5568), .B(n5567), .ZN(U2862)
         );
  AOI22_X1 U6246 ( .A1(n6834), .A2(DATAI_28_), .B1(n6837), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U6247 ( .A1(n6838), .A2(DATAI_12_), .ZN(n5570) );
  OAI211_X1 U6248 ( .C1(n5572), .C2(n6635), .A(n5571), .B(n5570), .ZN(U2863)
         );
  AOI22_X1 U6249 ( .A1(n6834), .A2(DATAI_27_), .B1(n6837), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U6250 ( .A1(n6838), .A2(DATAI_11_), .ZN(n5573) );
  OAI211_X1 U6251 ( .C1(n5575), .C2(n6635), .A(n5574), .B(n5573), .ZN(U2864)
         );
  AOI22_X1 U6252 ( .A1(n6834), .A2(DATAI_26_), .B1(n6837), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U6253 ( .A1(n6838), .A2(DATAI_10_), .ZN(n5576) );
  OAI211_X1 U6254 ( .C1(n5578), .C2(n6635), .A(n5577), .B(n5576), .ZN(U2865)
         );
  AOI22_X1 U6255 ( .A1(n6834), .A2(DATAI_25_), .B1(n6837), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U6256 ( .A1(n6838), .A2(DATAI_9_), .ZN(n5579) );
  OAI211_X1 U6257 ( .C1(n5624), .C2(n6635), .A(n5580), .B(n5579), .ZN(U2866)
         );
  AOI22_X1 U6258 ( .A1(n6834), .A2(DATAI_23_), .B1(n6837), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U6259 ( .A1(n6838), .A2(DATAI_7_), .ZN(n5581) );
  OAI211_X1 U6260 ( .C1(n5646), .C2(n6635), .A(n5582), .B(n5581), .ZN(U2868)
         );
  AOI22_X1 U6261 ( .A1(n6834), .A2(DATAI_21_), .B1(n6837), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U6262 ( .A1(n6838), .A2(DATAI_5_), .ZN(n5583) );
  OAI211_X1 U6263 ( .C1(n5585), .C2(n6635), .A(n5584), .B(n5583), .ZN(U2870)
         );
  AOI22_X1 U6264 ( .A1(n6834), .A2(DATAI_19_), .B1(n6837), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U6265 ( .A1(n6838), .A2(DATAI_3_), .ZN(n5586) );
  OAI211_X1 U6266 ( .C1(n5677), .C2(n6635), .A(n5587), .B(n5586), .ZN(U2872)
         );
  AND2_X1 U6267 ( .A1(n5590), .A2(n5589), .ZN(n5591) );
  XNOR2_X1 U6268 ( .A(n5592), .B(n5591), .ZN(n5730) );
  NAND2_X1 U6269 ( .A1(n6322), .A2(REIP_REG_29__SCAN_IN), .ZN(n5725) );
  OAI21_X1 U6270 ( .B1(n6209), .B2(n5593), .A(n5725), .ZN(n5594) );
  AOI21_X1 U6271 ( .B1(n6206), .B2(n5595), .A(n5594), .ZN(n5598) );
  NAND2_X1 U6272 ( .A1(n5596), .A2(n6211), .ZN(n5597) );
  OAI211_X1 U6273 ( .C1(n5730), .C2(n6535), .A(n5598), .B(n5597), .ZN(U2957)
         );
  INV_X1 U6274 ( .A(n5600), .ZN(n5601) );
  XNOR2_X1 U6275 ( .A(n5704), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5603)
         );
  NAND2_X1 U6276 ( .A1(n6322), .A2(REIP_REG_28__SCAN_IN), .ZN(n5735) );
  OAI21_X1 U6277 ( .B1(n6209), .B2(n5605), .A(n5735), .ZN(n5606) );
  AOI21_X1 U6278 ( .B1(n6206), .B2(n5607), .A(n5606), .ZN(n5610) );
  NAND2_X1 U6279 ( .A1(n5608), .A2(n6211), .ZN(n5609) );
  OAI211_X1 U6280 ( .C1(n5742), .C2(n6535), .A(n5610), .B(n5609), .ZN(U2958)
         );
  NOR2_X1 U6281 ( .A1(n4466), .A2(n5611), .ZN(n5614) );
  XNOR2_X1 U6282 ( .A(n5704), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5613)
         );
  OAI22_X1 U6283 ( .A1(n4562), .A2(n5614), .B1(n5613), .B2(n5612), .ZN(n5751)
         );
  NAND2_X1 U6284 ( .A1(n6322), .A2(REIP_REG_26__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U6285 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5615)
         );
  OAI211_X1 U6286 ( .C1(n6216), .C2(n5616), .A(n5746), .B(n5615), .ZN(n5617)
         );
  AOI21_X1 U6287 ( .B1(n5618), .B2(n6211), .A(n5617), .ZN(n5619) );
  OAI21_X1 U6288 ( .B1(n5751), .B2(n6535), .A(n5619), .ZN(U2960) );
  OAI21_X1 U6289 ( .B1(n5622), .B2(n5621), .A(n5620), .ZN(n6323) );
  OAI22_X1 U6290 ( .A1(n6209), .A2(n5623), .B1(n6262), .B2(n5435), .ZN(n5626)
         );
  NOR2_X1 U6291 ( .A1(n5624), .A2(n6188), .ZN(n5625) );
  AOI211_X1 U6292 ( .C1(n6206), .C2(n5627), .A(n5626), .B(n5625), .ZN(n5628)
         );
  OAI21_X1 U6293 ( .B1(n6323), .B2(n6535), .A(n5628), .ZN(U2961) );
  XNOR2_X1 U6294 ( .A(n5629), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5668)
         );
  NAND4_X1 U6295 ( .A1(n5662), .A2(n5772), .A3(n5629), .A4(n5794), .ZN(n5639)
         );
  XNOR2_X1 U6296 ( .A(n5629), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5654)
         );
  NOR2_X1 U6297 ( .A1(n5689), .A2(n5794), .ZN(n5653) );
  NOR2_X1 U6298 ( .A1(n5654), .A2(n5653), .ZN(n5631) );
  AOI21_X1 U6299 ( .B1(n5787), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5629), 
        .ZN(n5630) );
  AOI21_X1 U6300 ( .B1(n5662), .B2(n5631), .A(n5630), .ZN(n5648) );
  NAND4_X1 U6301 ( .A1(n5648), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n5689), .ZN(n5632) );
  OAI21_X1 U6302 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5639), .A(n5632), 
        .ZN(n5633) );
  XNOR2_X1 U6303 ( .A(n5633), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5759)
         );
  NOR2_X1 U6304 ( .A1(n6262), .A2(n6108), .ZN(n5756) );
  AOI21_X1 U6305 ( .B1(n6210), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5756), 
        .ZN(n5634) );
  OAI21_X1 U6306 ( .B1(n5635), .B2(n6216), .A(n5634), .ZN(n5636) );
  AOI21_X1 U6307 ( .B1(n6836), .B2(n6211), .A(n5636), .ZN(n5637) );
  OAI21_X1 U6308 ( .B1(n5759), .B2(n6535), .A(n5637), .ZN(U2962) );
  NAND2_X1 U6309 ( .A1(n5704), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5682) );
  NOR2_X1 U6310 ( .A1(n3469), .A2(n5682), .ZN(n5796) );
  NAND3_X1 U6311 ( .A1(n5796), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5752), .ZN(n5638) );
  NAND2_X1 U6312 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  XNOR2_X1 U6313 ( .A(n5640), .B(n5768), .ZN(n5760) );
  NAND2_X1 U6314 ( .A1(n5760), .A2(n6212), .ZN(n5645) );
  INV_X1 U6315 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6105) );
  NOR2_X1 U6316 ( .A1(n6262), .A2(n6105), .ZN(n5764) );
  NOR2_X1 U6317 ( .A1(n6209), .A2(n5641), .ZN(n5642) );
  AOI211_X1 U6318 ( .C1(n6206), .C2(n5643), .A(n5764), .B(n5642), .ZN(n5644)
         );
  OAI211_X1 U6319 ( .C1(n6188), .C2(n5646), .A(n5645), .B(n5644), .ZN(U2963)
         );
  XNOR2_X1 U6320 ( .A(n5704), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5647)
         );
  XNOR2_X1 U6321 ( .A(n5648), .B(n5647), .ZN(n5777) );
  NAND2_X1 U6322 ( .A1(n6322), .A2(REIP_REG_22__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U6323 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5649)
         );
  OAI211_X1 U6324 ( .C1(n6216), .C2(n5650), .A(n5773), .B(n5649), .ZN(n5651)
         );
  AOI21_X1 U6325 ( .B1(n6646), .B2(n6211), .A(n5651), .ZN(n5652) );
  OAI21_X1 U6326 ( .B1(n5777), .B2(n6535), .A(n5652), .ZN(U2964) );
  INV_X1 U6327 ( .A(n5662), .ZN(n5669) );
  OAI22_X1 U6328 ( .A1(n5669), .A2(n5653), .B1(n5629), .B2(n5787), .ZN(n5655)
         );
  XNOR2_X1 U6329 ( .A(n5655), .B(n5654), .ZN(n5785) );
  NAND2_X1 U6330 ( .A1(n6322), .A2(REIP_REG_21__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U6331 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5656)
         );
  OAI211_X1 U6332 ( .C1(n6216), .C2(n5657), .A(n5779), .B(n5656), .ZN(n5658)
         );
  AOI21_X1 U6333 ( .B1(n5659), .B2(n6211), .A(n5658), .ZN(n5660) );
  OAI21_X1 U6334 ( .B1(n5785), .B2(n6535), .A(n5660), .ZN(U2965) );
  NOR2_X1 U6335 ( .A1(n5629), .A2(n5661), .ZN(n5663) );
  MUX2_X1 U6336 ( .A(n5663), .B(n5629), .S(n5662), .Z(n5664) );
  XNOR2_X1 U6337 ( .A(n5664), .B(n5794), .ZN(n5786) );
  NAND2_X1 U6338 ( .A1(n5786), .A2(n6212), .ZN(n5667) );
  NOR2_X1 U6339 ( .A1(n6262), .A2(n6102), .ZN(n5790) );
  NOR2_X1 U6340 ( .A1(n6216), .A2(n6516), .ZN(n5665) );
  AOI211_X1 U6341 ( .C1(n6210), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5790), 
        .B(n5665), .ZN(n5666) );
  OAI211_X1 U6342 ( .C1(n6188), .C2(n6507), .A(n5667), .B(n5666), .ZN(U2966)
         );
  INV_X1 U6343 ( .A(n3452), .ZN(n5671) );
  INV_X1 U6344 ( .A(n5668), .ZN(n5670) );
  OAI21_X1 U6345 ( .B1(n5671), .B2(n5670), .A(n5669), .ZN(n6238) );
  NAND2_X1 U6346 ( .A1(n6238), .A2(n6212), .ZN(n5676) );
  OAI22_X1 U6347 ( .A1(n6209), .A2(n5672), .B1(n6262), .B2(n6100), .ZN(n5673)
         );
  AOI21_X1 U6348 ( .B1(n6206), .B2(n5674), .A(n5673), .ZN(n5675) );
  OAI211_X1 U6349 ( .C1(n6188), .C2(n5677), .A(n5676), .B(n5675), .ZN(U2967)
         );
  OAI21_X1 U6350 ( .B1(n5689), .B2(n5678), .A(n3469), .ZN(n5683) );
  NAND2_X1 U6351 ( .A1(n5629), .A2(n4474), .ZN(n5679) );
  NOR2_X1 U6352 ( .A1(n5683), .A2(n5679), .ZN(n5797) );
  INV_X1 U6353 ( .A(n5797), .ZN(n5681) );
  NAND3_X1 U6354 ( .A1(n5683), .A2(n5682), .A3(n5679), .ZN(n5680) );
  OAI211_X1 U6355 ( .C1(n5683), .C2(n5682), .A(n5681), .B(n5680), .ZN(n6316)
         );
  NAND2_X1 U6356 ( .A1(n6316), .A2(n6212), .ZN(n5688) );
  INV_X1 U6357 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5684) );
  OAI22_X1 U6358 ( .A1(n6209), .A2(n5685), .B1(n6262), .B2(n5684), .ZN(n5686)
         );
  AOI21_X1 U6359 ( .B1(n6206), .B2(n6488), .A(n5686), .ZN(n5687) );
  OAI211_X1 U6360 ( .C1(n6188), .C2(n6636), .A(n5688), .B(n5687), .ZN(U2969)
         );
  MUX2_X1 U6361 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n5678), .S(n5689), 
        .Z(n5690) );
  XNOR2_X1 U6362 ( .A(n5691), .B(n5690), .ZN(n5814) );
  AOI22_X1 U6363 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6322), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5692) );
  OAI21_X1 U6364 ( .B1(n6216), .B2(n5693), .A(n5692), .ZN(n5694) );
  AOI21_X1 U6365 ( .B1(n6631), .B2(n6211), .A(n5694), .ZN(n5695) );
  OAI21_X1 U6366 ( .B1(n5814), .B2(n6535), .A(n5695), .ZN(U2970) );
  XNOR2_X1 U6367 ( .A(n5704), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5697)
         );
  XNOR2_X1 U6368 ( .A(n5696), .B(n5697), .ZN(n6308) );
  NAND2_X1 U6369 ( .A1(n6308), .A2(n6212), .ZN(n5701) );
  AND2_X1 U6370 ( .A1(n6322), .A2(REIP_REG_15__SCAN_IN), .ZN(n6305) );
  NOR2_X1 U6371 ( .A1(n6216), .A2(n5698), .ZN(n5699) );
  AOI211_X1 U6372 ( .C1(n6210), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6305), 
        .B(n5699), .ZN(n5700) );
  OAI211_X1 U6373 ( .C1(n6188), .C2(n5702), .A(n5701), .B(n5700), .ZN(U2971)
         );
  XNOR2_X1 U6374 ( .A(n5704), .B(n5819), .ZN(n5705) );
  XNOR2_X1 U6375 ( .A(n5703), .B(n5705), .ZN(n5815) );
  INV_X1 U6376 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5706) );
  OAI22_X1 U6377 ( .A1(n6209), .A2(n4092), .B1(n6262), .B2(n5706), .ZN(n5708)
         );
  NOR2_X1 U6378 ( .A1(n6149), .A2(n6188), .ZN(n5707) );
  AOI211_X1 U6379 ( .C1(n6206), .C2(n6468), .A(n5708), .B(n5707), .ZN(n5709)
         );
  OAI21_X1 U6380 ( .B1(n5815), .B2(n6535), .A(n5709), .ZN(U2972) );
  INV_X1 U6381 ( .A(n5710), .ZN(n5718) );
  AOI21_X1 U6382 ( .B1(n5817), .B2(n5712), .A(n5711), .ZN(n5716) );
  NAND4_X1 U6383 ( .A1(n5723), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n5715), .ZN(n5713) );
  OAI211_X1 U6384 ( .C1(n5716), .C2(n5715), .A(n5714), .B(n5713), .ZN(n5717)
         );
  AOI21_X1 U6385 ( .B1(n6326), .B2(n5718), .A(n5717), .ZN(n5719) );
  OAI21_X1 U6386 ( .B1(n5720), .B2(n6334), .A(n5719), .ZN(U2987) );
  INV_X1 U6387 ( .A(n5721), .ZN(n5728) );
  NAND2_X1 U6388 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  OAI211_X1 U6389 ( .C1(n5726), .C2(n6339), .A(n5725), .B(n5724), .ZN(n5727)
         );
  AOI21_X1 U6390 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5728), .A(n5727), 
        .ZN(n5729) );
  OAI21_X1 U6391 ( .B1(n5730), .B2(n6334), .A(n5729), .ZN(U2989) );
  INV_X1 U6392 ( .A(n5731), .ZN(n5733) );
  NAND3_X1 U6393 ( .A1(n5733), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5732), .ZN(n5734) );
  OAI211_X1 U6394 ( .C1(n5736), .C2(n6339), .A(n5735), .B(n5734), .ZN(n5737)
         );
  INV_X1 U6395 ( .A(n5737), .ZN(n5741) );
  OAI21_X1 U6396 ( .B1(n5739), .B2(n5738), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n5740) );
  OAI211_X1 U6397 ( .C1(n5742), .C2(n6334), .A(n5741), .B(n5740), .ZN(U2990)
         );
  INV_X1 U6398 ( .A(n6332), .ZN(n5749) );
  INV_X1 U6399 ( .A(n5743), .ZN(n5744) );
  OAI211_X1 U6400 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6321), .B(n5744), .ZN(n5745) );
  OAI211_X1 U6401 ( .C1(n5747), .C2(n6339), .A(n5746), .B(n5745), .ZN(n5748)
         );
  AOI21_X1 U6402 ( .B1(n5749), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5748), 
        .ZN(n5750) );
  OAI21_X1 U6403 ( .B1(n5751), .B2(n6334), .A(n5750), .ZN(U2992) );
  NAND3_X1 U6404 ( .A1(n5770), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5752), .ZN(n5753) );
  AOI21_X1 U6405 ( .B1(n5754), .B2(n5753), .A(n6332), .ZN(n5755) );
  AOI211_X1 U6406 ( .C1(n6326), .C2(n5757), .A(n5756), .B(n5755), .ZN(n5758)
         );
  OAI21_X1 U6407 ( .B1(n5759), .B2(n6334), .A(n5758), .ZN(U2994) );
  NAND2_X1 U6408 ( .A1(n5760), .A2(n6327), .ZN(n5767) );
  INV_X1 U6409 ( .A(n5761), .ZN(n5765) );
  INV_X1 U6410 ( .A(n5770), .ZN(n6241) );
  NOR3_X1 U6411 ( .A1(n6241), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5762), 
        .ZN(n5763) );
  AOI211_X1 U6412 ( .C1(n5765), .C2(n6326), .A(n5764), .B(n5763), .ZN(n5766)
         );
  OAI211_X1 U6413 ( .C1(n5769), .C2(n5768), .A(n5767), .B(n5766), .ZN(U2995)
         );
  INV_X1 U6414 ( .A(n6236), .ZN(n5795) );
  OAI21_X1 U6415 ( .B1(n5787), .B2(n5807), .A(n5795), .ZN(n5783) );
  NAND2_X1 U6416 ( .A1(n5770), .A2(n5787), .ZN(n5778) );
  NOR3_X1 U6417 ( .A1(n5778), .A2(n5772), .A3(n5771), .ZN(n5775) );
  OAI21_X1 U6418 ( .B1(n6525), .B2(n6339), .A(n5773), .ZN(n5774) );
  AOI211_X1 U6419 ( .C1(n5783), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5775), .B(n5774), .ZN(n5776) );
  OAI21_X1 U6420 ( .B1(n5777), .B2(n6334), .A(n5776), .ZN(U2996) );
  NOR2_X1 U6421 ( .A1(n5778), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5782)
         );
  OAI21_X1 U6422 ( .B1(n5780), .B2(n6339), .A(n5779), .ZN(n5781) );
  AOI211_X1 U6423 ( .C1(n5783), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5782), .B(n5781), .ZN(n5784) );
  OAI21_X1 U6424 ( .B1(n5785), .B2(n6334), .A(n5784), .ZN(U2997) );
  NAND2_X1 U6425 ( .A1(n5786), .A2(n6327), .ZN(n5793) );
  INV_X1 U6426 ( .A(n6511), .ZN(n5791) );
  NOR3_X1 U6427 ( .A1(n6241), .A2(n5788), .A3(n5787), .ZN(n5789) );
  AOI211_X1 U6428 ( .C1(n6326), .C2(n5791), .A(n5790), .B(n5789), .ZN(n5792)
         );
  OAI211_X1 U6429 ( .C1(n5795), .C2(n5794), .A(n5793), .B(n5792), .ZN(U2998)
         );
  NOR2_X1 U6430 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  XNOR2_X1 U6431 ( .A(n5798), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6213)
         );
  NOR3_X1 U6432 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5799), .A3(n6320), 
        .ZN(n5804) );
  OAI21_X1 U6433 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5800), .A(n6313), 
        .ZN(n5801) );
  AOI22_X1 U6434 ( .A1(n6322), .A2(REIP_REG_18__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5801), .ZN(n5802) );
  OAI21_X1 U6435 ( .B1(n6505), .B2(n6339), .A(n5802), .ZN(n5803) );
  AOI211_X1 U6436 ( .C1(n6213), .C2(n6327), .A(n5804), .B(n5803), .ZN(n5805)
         );
  INV_X1 U6437 ( .A(n5805), .ZN(U3000) );
  OAI21_X1 U6438 ( .B1(n5807), .B2(n5809), .A(n5806), .ZN(n6307) );
  INV_X1 U6439 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6479) );
  OAI22_X1 U6440 ( .A1(n6339), .A2(n6484), .B1(n6479), .B2(n6262), .ZN(n5812)
         );
  NAND2_X1 U6441 ( .A1(n5809), .A2(n5808), .ZN(n6311) );
  AOI221_X1 U6442 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n5678), .C2(n5810), .A(n6311), 
        .ZN(n5811) );
  AOI211_X1 U6443 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n6307), .A(n5812), .B(n5811), .ZN(n5813) );
  OAI21_X1 U6444 ( .B1(n5814), .B2(n6334), .A(n5813), .ZN(U3002) );
  NOR2_X1 U6445 ( .A1(n5815), .A2(n6334), .ZN(n5826) );
  AOI21_X1 U6447 ( .B1(n5817), .B2(n5818), .A(n5816), .ZN(n6260) );
  OAI33_X1 U6448 ( .A1(1'b0), .A2(n6260), .A3(n5819), .B1(
        INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5818), .B3(n6320), .ZN(n5825)
         );
  XNOR2_X1 U6449 ( .A(n5822), .B(n5821), .ZN(n6464) );
  INV_X1 U6450 ( .A(n6464), .ZN(n5823) );
  OAI22_X1 U6451 ( .A1(n6339), .A2(n5823), .B1(n5706), .B2(n6262), .ZN(n5824)
         );
  OR3_X1 U6452 ( .A1(n5826), .A2(n5825), .A3(n5824), .ZN(U3004) );
  NOR2_X1 U6453 ( .A1(n5828), .A2(n5827), .ZN(n5832) );
  INV_X1 U6454 ( .A(n6580), .ZN(n6540) );
  OAI21_X1 U6455 ( .B1(n5832), .B2(n3751), .A(n5829), .ZN(n5830) );
  AOI21_X1 U6456 ( .B1(n6689), .B2(n5831), .A(n5830), .ZN(n6554) );
  OAI222_X1 U6457 ( .A1(n5834), .A2(n5833), .B1(n5832), .B2(n6590), .C1(n6540), 
        .C2(n6554), .ZN(n5835) );
  MUX2_X1 U6458 ( .A(n5835), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n6542), 
        .Z(U3460) );
  INV_X1 U6459 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6615) );
  AOI21_X1 U6460 ( .B1(n6615), .B2(STATE_REG_1__SCAN_IN), .A(n4566), .ZN(n5836) );
  NOR2_X1 U6461 ( .A1(n6630), .A2(n5836), .ZN(n6612) );
  INV_X1 U6462 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6137) );
  INV_X1 U6463 ( .A(BS16_N), .ZN(n5999) );
  NAND2_X1 U6464 ( .A1(n6615), .A2(n4566), .ZN(n6218) );
  AOI21_X1 U6465 ( .B1(n5999), .B2(n6218), .A(n6046), .ZN(n6609) );
  AOI21_X1 U6466 ( .B1(n6046), .B2(n6137), .A(n6609), .ZN(U3451) );
  AND2_X1 U6467 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6046), .ZN(U3180) );
  AND2_X1 U6468 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6046), .ZN(U3179) );
  AND2_X1 U6469 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6046), .ZN(U3178) );
  AND2_X1 U6470 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6046), .ZN(U3177) );
  AND2_X1 U6471 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6046), .ZN(U3176) );
  AND2_X1 U6472 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6046), .ZN(U3175) );
  AND2_X1 U6473 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6046), .ZN(U3174) );
  AND2_X1 U6474 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6046), .ZN(U3173) );
  AND2_X1 U6475 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6046), .ZN(U3172) );
  AND2_X1 U6476 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6046), .ZN(U3171) );
  AND2_X1 U6477 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6046), .ZN(U3170) );
  AND2_X1 U6478 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6046), .ZN(U3169) );
  AND2_X1 U6479 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6046), .ZN(U3168) );
  AND2_X1 U6480 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6046), .ZN(U3167) );
  AND2_X1 U6481 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6046), .ZN(U3166) );
  AND2_X1 U6482 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6046), .ZN(U3165) );
  AND2_X1 U6483 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6046), .ZN(U3164) );
  AND2_X1 U6484 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6046), .ZN(U3163) );
  AND2_X1 U6485 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6046), .ZN(U3162) );
  AND2_X1 U6486 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6046), .ZN(U3161) );
  AND2_X1 U6487 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6046), .ZN(U3159) );
  AND2_X1 U6488 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6046), .ZN(U3158) );
  AND2_X1 U6489 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6046), .ZN(U3157) );
  AND2_X1 U6490 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6046), .ZN(U3156) );
  AND2_X1 U6491 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6046), .ZN(U3155) );
  AND2_X1 U6492 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6046), .ZN(U3154) );
  AND2_X1 U6493 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6046), .ZN(U3153) );
  AND2_X1 U6494 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6046), .ZN(U3152) );
  AND2_X1 U6495 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6046), .ZN(U3151) );
  INV_X1 U6496 ( .A(n6606), .ZN(n6608) );
  AND2_X1 U6497 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6608), .ZN(U3019)
         );
  AND2_X1 U6498 ( .A1(n6061), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6499 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6006) );
  AOI21_X1 U6500 ( .B1(n5836), .B2(n6006), .A(n6630), .ZN(U2789) );
  INV_X1 U6501 ( .A(keyinput_117), .ZN(n5920) );
  INV_X1 U6502 ( .A(keyinput_116), .ZN(n5918) );
  INV_X1 U6503 ( .A(keyinput_115), .ZN(n5916) );
  INV_X1 U6504 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6122) );
  INV_X1 U6505 ( .A(keyinput_111), .ZN(n5909) );
  INV_X1 U6506 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6019) );
  INV_X1 U6507 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6613) );
  OAI22_X1 U6508 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_103), .B1(
        ADS_N_REG_SCAN_IN), .B2(keyinput_102), .ZN(n5837) );
  AOI221_X1 U6509 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_103), .C1(
        keyinput_102), .C2(ADS_N_REG_SCAN_IN), .A(n5837), .ZN(n5898) );
  INV_X1 U6510 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n5896) );
  XNOR2_X1 U6511 ( .A(HOLD), .B(keyinput_100), .ZN(n5894) );
  INV_X1 U6512 ( .A(keyinput_99), .ZN(n5892) );
  INV_X1 U6513 ( .A(keyinput_98), .ZN(n5890) );
  INV_X1 U6514 ( .A(keyinput_97), .ZN(n5888) );
  INV_X1 U6515 ( .A(NA_N), .ZN(n6621) );
  INV_X1 U6516 ( .A(keyinput_96), .ZN(n5886) );
  AOI22_X1 U6517 ( .A1(n5840), .A2(keyinput_93), .B1(n5839), .B2(keyinput_92), 
        .ZN(n5838) );
  OAI221_X1 U6518 ( .B1(n5840), .B2(keyinput_93), .C1(n5839), .C2(keyinput_92), 
        .A(n5838), .ZN(n5883) );
  OAI22_X1 U6519 ( .A1(n5938), .A2(keyinput_91), .B1(DATAI_5_), .B2(
        keyinput_90), .ZN(n5841) );
  AOI221_X1 U6520 ( .B1(n5938), .B2(keyinput_91), .C1(keyinput_90), .C2(
        DATAI_5_), .A(n5841), .ZN(n5880) );
  OAI22_X1 U6521 ( .A1(n5940), .A2(keyinput_87), .B1(keyinput_88), .B2(
        DATAI_7_), .ZN(n5842) );
  AOI221_X1 U6522 ( .B1(n5940), .B2(keyinput_87), .C1(DATAI_7_), .C2(
        keyinput_88), .A(n5842), .ZN(n5877) );
  AOI22_X1 U6523 ( .A1(n5845), .A2(keyinput_85), .B1(n5844), .B2(keyinput_84), 
        .ZN(n5843) );
  OAI221_X1 U6524 ( .B1(n5845), .B2(keyinput_85), .C1(n5844), .C2(keyinput_84), 
        .A(n5843), .ZN(n5875) );
  INV_X1 U6525 ( .A(keyinput_83), .ZN(n5872) );
  INV_X1 U6526 ( .A(DATAI_14_), .ZN(n5972) );
  INV_X1 U6527 ( .A(DATAI_13_), .ZN(n5976) );
  OAI22_X1 U6528 ( .A1(n5976), .A2(keyinput_82), .B1(DATAI_15_), .B2(
        keyinput_80), .ZN(n5846) );
  AOI221_X1 U6529 ( .B1(n5976), .B2(keyinput_82), .C1(keyinput_80), .C2(
        DATAI_15_), .A(n5846), .ZN(n5869) );
  INV_X1 U6530 ( .A(keyinput_79), .ZN(n5867) );
  INV_X1 U6531 ( .A(keyinput_78), .ZN(n5865) );
  AOI22_X1 U6532 ( .A1(n5943), .A2(keyinput_74), .B1(n4956), .B2(keyinput_71), 
        .ZN(n5847) );
  OAI221_X1 U6533 ( .B1(n5943), .B2(keyinput_74), .C1(n4956), .C2(keyinput_71), 
        .A(n5847), .ZN(n5863) );
  OAI22_X1 U6534 ( .A1(DATAI_26_), .A2(keyinput_69), .B1(keyinput_70), .B2(
        DATAI_25_), .ZN(n5848) );
  AOI221_X1 U6535 ( .B1(DATAI_26_), .B2(keyinput_69), .C1(DATAI_25_), .C2(
        keyinput_70), .A(n5848), .ZN(n5858) );
  OAI22_X1 U6536 ( .A1(DATAI_27_), .A2(keyinput_68), .B1(keyinput_73), .B2(
        DATAI_22_), .ZN(n5849) );
  AOI221_X1 U6537 ( .B1(DATAI_27_), .B2(keyinput_68), .C1(DATAI_22_), .C2(
        keyinput_73), .A(n5849), .ZN(n5857) );
  INV_X1 U6538 ( .A(keyinput_67), .ZN(n5854) );
  INV_X1 U6539 ( .A(keyinput_64), .ZN(n5852) );
  OAI22_X1 U6540 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_29_), .B2(
        keyinput_66), .ZN(n5850) );
  AOI221_X1 U6541 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(keyinput_66), .C2(
        DATAI_29_), .A(n5850), .ZN(n5851) );
  OAI221_X1 U6542 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(n4951), .C2(n5852), 
        .A(n5851), .ZN(n5853) );
  OAI221_X1 U6543 ( .B1(DATAI_28_), .B2(keyinput_67), .C1(n5268), .C2(n5854), 
        .A(n5853), .ZN(n5856) );
  XNOR2_X1 U6544 ( .A(DATAI_23_), .B(keyinput_72), .ZN(n5855) );
  NAND4_X1 U6545 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n5862)
         );
  OAI22_X1 U6546 ( .A1(n5956), .A2(keyinput_77), .B1(DATAI_19_), .B2(
        keyinput_76), .ZN(n5859) );
  AOI221_X1 U6547 ( .B1(n5956), .B2(keyinput_77), .C1(keyinput_76), .C2(
        DATAI_19_), .A(n5859), .ZN(n5861) );
  XOR2_X1 U6548 ( .A(n5958), .B(keyinput_75), .Z(n5860) );
  OAI211_X1 U6549 ( .C1(n5863), .C2(n5862), .A(n5861), .B(n5860), .ZN(n5864)
         );
  OAI221_X1 U6550 ( .B1(DATAI_17_), .B2(keyinput_78), .C1(n5965), .C2(n5865), 
        .A(n5864), .ZN(n5866) );
  OAI221_X1 U6551 ( .B1(DATAI_16_), .B2(n5867), .C1(n5969), .C2(keyinput_79), 
        .A(n5866), .ZN(n5868) );
  OAI211_X1 U6552 ( .C1(n5972), .C2(keyinput_81), .A(n5869), .B(n5868), .ZN(
        n5870) );
  AOI21_X1 U6553 ( .B1(n5972), .B2(keyinput_81), .A(n5870), .ZN(n5871) );
  AOI221_X1 U6554 ( .B1(DATAI_12_), .B2(keyinput_83), .C1(n5978), .C2(n5872), 
        .A(n5871), .ZN(n5874) );
  NAND2_X1 U6555 ( .A1(DATAI_9_), .A2(keyinput_86), .ZN(n5873) );
  OAI221_X1 U6556 ( .B1(n5875), .B2(n5874), .C1(DATAI_9_), .C2(keyinput_86), 
        .A(n5873), .ZN(n5876) );
  AOI22_X1 U6557 ( .A1(keyinput_89), .A2(n5987), .B1(n5877), .B2(n5876), .ZN(
        n5878) );
  OAI21_X1 U6558 ( .B1(n5987), .B2(keyinput_89), .A(n5878), .ZN(n5879) );
  AOI22_X1 U6559 ( .A1(n5880), .A2(n5879), .B1(DATAI_1_), .B2(keyinput_94), 
        .ZN(n5881) );
  OAI21_X1 U6560 ( .B1(DATAI_1_), .B2(keyinput_94), .A(n5881), .ZN(n5882) );
  OAI22_X1 U6561 ( .A1(n5883), .A2(n5882), .B1(keyinput_95), .B2(DATAI_0_), 
        .ZN(n5884) );
  AOI21_X1 U6562 ( .B1(keyinput_95), .B2(DATAI_0_), .A(n5884), .ZN(n5885) );
  AOI221_X1 U6563 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5886), .C1(n6629), .C2(
        keyinput_96), .A(n5885), .ZN(n5887) );
  AOI221_X1 U6564 ( .B1(NA_N), .B2(n5888), .C1(n6621), .C2(keyinput_97), .A(
        n5887), .ZN(n5889) );
  AOI221_X1 U6565 ( .B1(BS16_N), .B2(n5890), .C1(n5999), .C2(keyinput_98), .A(
        n5889), .ZN(n5891) );
  AOI221_X1 U6566 ( .B1(READY_N), .B2(keyinput_99), .C1(n6619), .C2(n5892), 
        .A(n5891), .ZN(n5893) );
  OAI22_X1 U6567 ( .A1(n5894), .A2(n5893), .B1(n5896), .B2(keyinput_101), .ZN(
        n5895) );
  AOI21_X1 U6568 ( .B1(n5896), .B2(keyinput_101), .A(n5895), .ZN(n5897) );
  AOI22_X1 U6569 ( .A1(n5898), .A2(n5897), .B1(keyinput_106), .B2(n6613), .ZN(
        n5899) );
  OAI21_X1 U6570 ( .B1(keyinput_106), .B2(n6613), .A(n5899), .ZN(n5907) );
  INV_X1 U6571 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6010) );
  INV_X1 U6572 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6628) );
  AOI22_X1 U6573 ( .A1(n6010), .A2(keyinput_105), .B1(n6628), .B2(keyinput_104), .ZN(n5900) );
  OAI221_X1 U6574 ( .B1(n6010), .B2(keyinput_105), .C1(n6628), .C2(
        keyinput_104), .A(n5900), .ZN(n5906) );
  INV_X1 U6575 ( .A(MORE_REG_SCAN_IN), .ZN(n5902) );
  OAI22_X1 U6576 ( .A1(n5902), .A2(keyinput_108), .B1(keyinput_107), .B2(
        STATEBS16_REG_SCAN_IN), .ZN(n5901) );
  AOI221_X1 U6577 ( .B1(n5902), .B2(keyinput_108), .C1(STATEBS16_REG_SCAN_IN), 
        .C2(keyinput_107), .A(n5901), .ZN(n5905) );
  OAI22_X1 U6578 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_109), .B1(keyinput_110), .B2(W_R_N_REG_SCAN_IN), .ZN(n5903) );
  AOI221_X1 U6579 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_109), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput_110), .A(n5903), .ZN(n5904) );
  OAI211_X1 U6580 ( .C1(n5907), .C2(n5906), .A(n5905), .B(n5904), .ZN(n5908)
         );
  OAI221_X1 U6581 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(n5909), .C1(n6019), 
        .C2(keyinput_111), .A(n5908), .ZN(n5914) );
  INV_X1 U6582 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n5911) );
  OAI22_X1 U6583 ( .A1(n5911), .A2(keyinput_113), .B1(keyinput_112), .B2(
        BYTEENABLE_REG_1__SCAN_IN), .ZN(n5910) );
  AOI221_X1 U6584 ( .B1(n5911), .B2(keyinput_113), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_112), .A(n5910), .ZN(n5913)
         );
  NOR2_X1 U6585 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_114), .ZN(n5912) );
  AOI221_X1 U6586 ( .B1(n5914), .B2(n5913), .C1(keyinput_114), .C2(
        BYTEENABLE_REG_3__SCAN_IN), .A(n5912), .ZN(n5915) );
  AOI221_X1 U6587 ( .B1(REIP_REG_31__SCAN_IN), .B2(n5916), .C1(n6122), .C2(
        keyinput_115), .A(n5915), .ZN(n5917) );
  AOI221_X1 U6588 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5918), .C1(n6118), .C2(
        keyinput_116), .A(n5917), .ZN(n5919) );
  AOI221_X1 U6589 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5920), .C1(n6030), .C2(
        keyinput_117), .A(n5919), .ZN(n5927) );
  AOI22_X1 U6590 ( .A1(n6111), .A2(keyinput_119), .B1(n6116), .B2(keyinput_118), .ZN(n5921) );
  OAI221_X1 U6591 ( .B1(n6111), .B2(keyinput_119), .C1(n6116), .C2(
        keyinput_118), .A(n5921), .ZN(n5926) );
  OAI22_X1 U6592 ( .A1(n6105), .A2(keyinput_123), .B1(keyinput_120), .B2(
        REIP_REG_26__SCAN_IN), .ZN(n5922) );
  AOI221_X1 U6593 ( .B1(n6105), .B2(keyinput_123), .C1(REIP_REG_26__SCAN_IN), 
        .C2(keyinput_120), .A(n5922), .ZN(n5925) );
  OAI22_X1 U6594 ( .A1(n6108), .A2(keyinput_122), .B1(REIP_REG_25__SCAN_IN), 
        .B2(keyinput_121), .ZN(n5923) );
  AOI221_X1 U6595 ( .B1(n6108), .B2(keyinput_122), .C1(keyinput_121), .C2(
        REIP_REG_25__SCAN_IN), .A(n5923), .ZN(n5924) );
  OAI211_X1 U6596 ( .C1(n5927), .C2(n5926), .A(n5925), .B(n5924), .ZN(n5929)
         );
  XOR2_X1 U6597 ( .A(n6517), .B(keyinput_124), .Z(n5928) );
  OAI22_X1 U6598 ( .A1(n5929), .A2(n5928), .B1(keyinput_125), .B2(
        REIP_REG_21__SCAN_IN), .ZN(n5930) );
  AOI21_X1 U6599 ( .B1(keyinput_125), .B2(REIP_REG_21__SCAN_IN), .A(n5930), 
        .ZN(n6045) );
  INV_X1 U6600 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6102) );
  AOI22_X1 U6601 ( .A1(n6100), .A2(keyinput_127), .B1(n6102), .B2(keyinput_126), .ZN(n5931) );
  OAI221_X1 U6602 ( .B1(n6100), .B2(keyinput_127), .C1(n6102), .C2(
        keyinput_126), .A(n5931), .ZN(n6044) );
  OAI22_X1 U6603 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_54), .B1(
        REIP_REG_27__SCAN_IN), .B2(keyinput_55), .ZN(n5932) );
  AOI221_X1 U6604 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_54), .C1(
        keyinput_55), .C2(REIP_REG_27__SCAN_IN), .A(n5932), .ZN(n6036) );
  INV_X1 U6605 ( .A(keyinput_53), .ZN(n6029) );
  INV_X1 U6606 ( .A(keyinput_52), .ZN(n6027) );
  INV_X1 U6607 ( .A(keyinput_51), .ZN(n6025) );
  INV_X1 U6608 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6141) );
  OAI22_X1 U6609 ( .A1(n6141), .A2(keyinput_48), .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .ZN(n5933) );
  AOI221_X1 U6610 ( .B1(n6141), .B2(keyinput_48), .C1(keyinput_49), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n5933), .ZN(n6022) );
  INV_X1 U6611 ( .A(keyinput_47), .ZN(n6020) );
  OAI22_X1 U6612 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_37), .B1(
        CODEFETCH_REG_SCAN_IN), .B2(keyinput_39), .ZN(n5934) );
  AOI221_X1 U6613 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_37), .C1(
        keyinput_39), .C2(CODEFETCH_REG_SCAN_IN), .A(n5934), .ZN(n6008) );
  XOR2_X1 U6614 ( .A(HOLD), .B(keyinput_36), .Z(n6004) );
  INV_X1 U6615 ( .A(keyinput_35), .ZN(n6002) );
  INV_X1 U6616 ( .A(keyinput_34), .ZN(n6000) );
  INV_X1 U6617 ( .A(keyinput_33), .ZN(n5997) );
  INV_X1 U6618 ( .A(keyinput_32), .ZN(n5995) );
  AOI22_X1 U6619 ( .A1(DATAI_1_), .A2(keyinput_30), .B1(DATAI_3_), .B2(
        keyinput_28), .ZN(n5935) );
  OAI221_X1 U6620 ( .B1(DATAI_1_), .B2(keyinput_30), .C1(DATAI_3_), .C2(
        keyinput_28), .A(n5935), .ZN(n5992) );
  AOI22_X1 U6621 ( .A1(n5938), .A2(keyinput_27), .B1(n5937), .B2(keyinput_26), 
        .ZN(n5936) );
  OAI221_X1 U6622 ( .B1(n5938), .B2(keyinput_27), .C1(n5937), .C2(keyinput_26), 
        .A(n5936), .ZN(n5990) );
  AOI22_X1 U6623 ( .A1(DATAI_7_), .A2(keyinput_24), .B1(n5940), .B2(
        keyinput_23), .ZN(n5939) );
  OAI221_X1 U6624 ( .B1(DATAI_7_), .B2(keyinput_24), .C1(n5940), .C2(
        keyinput_23), .A(n5939), .ZN(n5985) );
  AOI22_X1 U6625 ( .A1(DATAI_10_), .A2(keyinput_21), .B1(DATAI_11_), .B2(
        keyinput_20), .ZN(n5941) );
  OAI221_X1 U6626 ( .B1(DATAI_10_), .B2(keyinput_21), .C1(DATAI_11_), .C2(
        keyinput_20), .A(n5941), .ZN(n5981) );
  INV_X1 U6627 ( .A(keyinput_19), .ZN(n5979) );
  INV_X1 U6628 ( .A(keyinput_15), .ZN(n5968) );
  INV_X1 U6629 ( .A(keyinput_14), .ZN(n5966) );
  XOR2_X1 U6630 ( .A(DATAI_23_), .B(keyinput_8), .Z(n5950) );
  AOI22_X1 U6631 ( .A1(n5944), .A2(keyinput_5), .B1(keyinput_10), .B2(n5943), 
        .ZN(n5942) );
  OAI221_X1 U6632 ( .B1(n5944), .B2(keyinput_5), .C1(n5943), .C2(keyinput_10), 
        .A(n5942), .ZN(n5949) );
  AOI22_X1 U6633 ( .A1(DATAI_22_), .A2(keyinput_9), .B1(DATAI_25_), .B2(
        keyinput_6), .ZN(n5945) );
  OAI221_X1 U6634 ( .B1(DATAI_22_), .B2(keyinput_9), .C1(DATAI_25_), .C2(
        keyinput_6), .A(n5945), .ZN(n5948) );
  AOI22_X1 U6635 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(DATAI_27_), .B2(
        keyinput_4), .ZN(n5946) );
  OAI221_X1 U6636 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(DATAI_27_), .C2(
        keyinput_4), .A(n5946), .ZN(n5947) );
  NOR4_X1 U6637 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(n5963)
         );
  INV_X1 U6638 ( .A(keyinput_3), .ZN(n5955) );
  INV_X1 U6639 ( .A(keyinput_0), .ZN(n5953) );
  OAI22_X1 U6640 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(keyinput_2), .B2(
        DATAI_29_), .ZN(n5951) );
  AOI221_X1 U6641 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_29_), .C2(
        keyinput_2), .A(n5951), .ZN(n5952) );
  OAI221_X1 U6642 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(n4951), .C2(n5953), 
        .A(n5952), .ZN(n5954) );
  OAI221_X1 U6643 ( .B1(DATAI_28_), .B2(n5955), .C1(n5268), .C2(keyinput_3), 
        .A(n5954), .ZN(n5962) );
  XNOR2_X1 U6644 ( .A(n5956), .B(keyinput_13), .ZN(n5961) );
  AOI22_X1 U6645 ( .A1(n5959), .A2(keyinput_12), .B1(n5958), .B2(keyinput_11), 
        .ZN(n5957) );
  OAI221_X1 U6646 ( .B1(n5959), .B2(keyinput_12), .C1(n5958), .C2(keyinput_11), 
        .A(n5957), .ZN(n5960) );
  AOI211_X1 U6647 ( .C1(n5963), .C2(n5962), .A(n5961), .B(n5960), .ZN(n5964)
         );
  AOI221_X1 U6648 ( .B1(DATAI_17_), .B2(n5966), .C1(n5965), .C2(keyinput_14), 
        .A(n5964), .ZN(n5967) );
  AOI221_X1 U6649 ( .B1(DATAI_16_), .B2(keyinput_15), .C1(n5969), .C2(n5968), 
        .A(n5967), .ZN(n5975) );
  OAI22_X1 U6650 ( .A1(n5972), .A2(keyinput_17), .B1(n5971), .B2(keyinput_16), 
        .ZN(n5970) );
  AOI221_X1 U6651 ( .B1(n5972), .B2(keyinput_17), .C1(keyinput_16), .C2(n5971), 
        .A(n5970), .ZN(n5973) );
  OAI21_X1 U6652 ( .B1(keyinput_18), .B2(n5976), .A(n5973), .ZN(n5974) );
  AOI211_X1 U6653 ( .C1(keyinput_18), .C2(n5976), .A(n5975), .B(n5974), .ZN(
        n5977) );
  AOI221_X1 U6654 ( .B1(DATAI_12_), .B2(n5979), .C1(n5978), .C2(keyinput_19), 
        .A(n5977), .ZN(n5980) );
  OAI22_X1 U6655 ( .A1(keyinput_22), .A2(n5983), .B1(n5981), .B2(n5980), .ZN(
        n5982) );
  AOI21_X1 U6656 ( .B1(keyinput_22), .B2(n5983), .A(n5982), .ZN(n5984) );
  OAI22_X1 U6657 ( .A1(keyinput_25), .A2(n5987), .B1(n5985), .B2(n5984), .ZN(
        n5986) );
  AOI21_X1 U6658 ( .B1(keyinput_25), .B2(n5987), .A(n5986), .ZN(n5989) );
  NAND2_X1 U6659 ( .A1(keyinput_29), .A2(DATAI_2_), .ZN(n5988) );
  OAI221_X1 U6660 ( .B1(n5990), .B2(n5989), .C1(keyinput_29), .C2(DATAI_2_), 
        .A(n5988), .ZN(n5991) );
  OAI22_X1 U6661 ( .A1(n5992), .A2(n5991), .B1(keyinput_31), .B2(DATAI_0_), 
        .ZN(n5993) );
  AOI21_X1 U6662 ( .B1(keyinput_31), .B2(DATAI_0_), .A(n5993), .ZN(n5994) );
  AOI221_X1 U6663 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_32), .C1(n6629), 
        .C2(n5995), .A(n5994), .ZN(n5996) );
  AOI221_X1 U6664 ( .B1(NA_N), .B2(n5997), .C1(n6621), .C2(keyinput_33), .A(
        n5996), .ZN(n5998) );
  AOI221_X1 U6665 ( .B1(BS16_N), .B2(n6000), .C1(n5999), .C2(keyinput_34), .A(
        n5998), .ZN(n6001) );
  AOI221_X1 U6666 ( .B1(READY_N), .B2(n6002), .C1(n6619), .C2(keyinput_35), 
        .A(n6001), .ZN(n6003) );
  OAI22_X1 U6667 ( .A1(n6004), .A2(n6003), .B1(n6006), .B2(keyinput_38), .ZN(
        n6005) );
  AOI21_X1 U6668 ( .B1(n6006), .B2(keyinput_38), .A(n6005), .ZN(n6007) );
  AOI22_X1 U6669 ( .A1(n6008), .A2(n6007), .B1(keyinput_41), .B2(n6010), .ZN(
        n6009) );
  OAI21_X1 U6670 ( .B1(keyinput_41), .B2(n6010), .A(n6009), .ZN(n6017) );
  AOI22_X1 U6671 ( .A1(keyinput_42), .A2(REQUESTPENDING_REG_SCAN_IN), .B1(
        n6628), .B2(keyinput_40), .ZN(n6011) );
  OAI221_X1 U6672 ( .B1(keyinput_42), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(
        n6628), .C2(keyinput_40), .A(n6011), .ZN(n6016) );
  INV_X1 U6673 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6219) );
  OAI22_X1 U6674 ( .A1(n6219), .A2(keyinput_46), .B1(MORE_REG_SCAN_IN), .B2(
        keyinput_44), .ZN(n6012) );
  AOI221_X1 U6675 ( .B1(n6219), .B2(keyinput_46), .C1(keyinput_44), .C2(
        MORE_REG_SCAN_IN), .A(n6012), .ZN(n6015) );
  OAI22_X1 U6676 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_43), .B1(
        FLUSH_REG_SCAN_IN), .B2(keyinput_45), .ZN(n6013) );
  AOI221_X1 U6677 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_43), .C1(
        keyinput_45), .C2(FLUSH_REG_SCAN_IN), .A(n6013), .ZN(n6014) );
  OAI211_X1 U6678 ( .C1(n6017), .C2(n6016), .A(n6015), .B(n6014), .ZN(n6018)
         );
  OAI221_X1 U6679 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(n6020), .C1(n6019), 
        .C2(keyinput_47), .A(n6018), .ZN(n6021) );
  AOI22_X1 U6680 ( .A1(n6022), .A2(n6021), .B1(keyinput_50), .B2(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U6681 ( .B1(keyinput_50), .B2(BYTEENABLE_REG_3__SCAN_IN), .A(n6023), 
        .ZN(n6024) );
  OAI221_X1 U6682 ( .B1(REIP_REG_31__SCAN_IN), .B2(n6025), .C1(n6122), .C2(
        keyinput_51), .A(n6024), .ZN(n6026) );
  OAI221_X1 U6683 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6027), .C1(n6118), .C2(
        keyinput_52), .A(n6026), .ZN(n6028) );
  OAI221_X1 U6684 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_53), .C1(n6030), 
        .C2(n6029), .A(n6028), .ZN(n6035) );
  AOI22_X1 U6685 ( .A1(n6105), .A2(keyinput_59), .B1(n6108), .B2(keyinput_58), 
        .ZN(n6031) );
  OAI221_X1 U6686 ( .B1(n6105), .B2(keyinput_59), .C1(n6108), .C2(keyinput_58), 
        .A(n6031), .ZN(n6034) );
  AOI22_X1 U6687 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_60), .B1(n5417), 
        .B2(keyinput_56), .ZN(n6032) );
  OAI221_X1 U6688 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_60), .C1(n5417), 
        .C2(keyinput_56), .A(n6032), .ZN(n6033) );
  AOI211_X1 U6689 ( .C1(n6036), .C2(n6035), .A(n6034), .B(n6033), .ZN(n6038)
         );
  XOR2_X1 U6690 ( .A(keyinput_57), .B(REIP_REG_25__SCAN_IN), .Z(n6037) );
  AOI22_X1 U6691 ( .A1(n6038), .A2(n6037), .B1(keyinput_61), .B2(n6041), .ZN(
        n6042) );
  AOI22_X1 U6692 ( .A1(n6100), .A2(keyinput_63), .B1(n6102), .B2(keyinput_62), 
        .ZN(n6039) );
  OAI221_X1 U6693 ( .B1(n6100), .B2(keyinput_63), .C1(n6102), .C2(keyinput_62), 
        .A(n6039), .ZN(n6040) );
  AOI221_X1 U6694 ( .B1(keyinput_61), .B2(n6042), .C1(n6041), .C2(n6042), .A(
        n6040), .ZN(n6043) );
  OAI21_X1 U6695 ( .B1(n6045), .B2(n6044), .A(n6043), .ZN(n6048) );
  NAND2_X1 U6696 ( .A1(n6046), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6047) );
  XOR2_X1 U6697 ( .A(n6048), .B(n6047), .Z(U3160) );
  AOI22_X1 U6698 ( .A1(n6228), .A2(LWORD_REG_0__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6050) );
  OAI21_X1 U6699 ( .B1(n6051), .B2(n6078), .A(n6050), .ZN(U2923) );
  AOI22_X1 U6700 ( .A1(n6228), .A2(LWORD_REG_1__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6052) );
  OAI21_X1 U6701 ( .B1(n6053), .B2(n6078), .A(n6052), .ZN(U2922) );
  AOI22_X1 U6702 ( .A1(n6228), .A2(LWORD_REG_2__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U6703 ( .B1(n6055), .B2(n6078), .A(n6054), .ZN(U2921) );
  AOI22_X1 U6704 ( .A1(n6228), .A2(LWORD_REG_3__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6056) );
  OAI21_X1 U6705 ( .B1(n6057), .B2(n6078), .A(n6056), .ZN(U2920) );
  AOI22_X1 U6706 ( .A1(n6228), .A2(LWORD_REG_4__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6058) );
  OAI21_X1 U6707 ( .B1(n6059), .B2(n6078), .A(n6058), .ZN(U2919) );
  AOI22_X1 U6708 ( .A1(n6228), .A2(LWORD_REG_5__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6060) );
  OAI21_X1 U6709 ( .B1(n4788), .B2(n6078), .A(n6060), .ZN(U2918) );
  AOI22_X1 U6710 ( .A1(n6228), .A2(LWORD_REG_6__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6062) );
  OAI21_X1 U6711 ( .B1(n3969), .B2(n6078), .A(n6062), .ZN(U2917) );
  AOI22_X1 U6712 ( .A1(n6228), .A2(LWORD_REG_7__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6063) );
  OAI21_X1 U6713 ( .B1(n4781), .B2(n6078), .A(n6063), .ZN(U2916) );
  AOI22_X1 U6714 ( .A1(n6228), .A2(LWORD_REG_8__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6064) );
  OAI21_X1 U6715 ( .B1(n6065), .B2(n6078), .A(n6064), .ZN(U2915) );
  AOI22_X1 U6716 ( .A1(n6228), .A2(LWORD_REG_9__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6066) );
  OAI21_X1 U6717 ( .B1(n6067), .B2(n6078), .A(n6066), .ZN(U2914) );
  AOI22_X1 U6718 ( .A1(n6228), .A2(LWORD_REG_10__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6068) );
  OAI21_X1 U6719 ( .B1(n6069), .B2(n6078), .A(n6068), .ZN(U2913) );
  AOI22_X1 U6720 ( .A1(n6228), .A2(LWORD_REG_11__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6070) );
  OAI21_X1 U6721 ( .B1(n6071), .B2(n6078), .A(n6070), .ZN(U2912) );
  AOI22_X1 U6722 ( .A1(n6228), .A2(LWORD_REG_12__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6072) );
  OAI21_X1 U6723 ( .B1(n6073), .B2(n6078), .A(n6072), .ZN(U2911) );
  INV_X1 U6724 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6075) );
  AOI22_X1 U6725 ( .A1(n6228), .A2(LWORD_REG_13__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6074) );
  OAI21_X1 U6726 ( .B1(n6075), .B2(n6078), .A(n6074), .ZN(U2910) );
  AOI22_X1 U6727 ( .A1(n6228), .A2(LWORD_REG_14__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6076) );
  OAI21_X1 U6728 ( .B1(n4799), .B2(n6078), .A(n6076), .ZN(U2909) );
  INV_X1 U6729 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6079) );
  AOI22_X1 U6730 ( .A1(n6228), .A2(LWORD_REG_15__SCAN_IN), .B1(n6061), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6077) );
  OAI21_X1 U6731 ( .B1(n6079), .B2(n6078), .A(n6077), .ZN(U2908) );
  INV_X2 U6732 ( .A(n6630), .ZN(n6627) );
  NOR2_X2 U6733 ( .A1(n6615), .A2(n6627), .ZN(n6119) );
  NAND2_X1 U6734 ( .A1(n6615), .A2(n6630), .ZN(n6121) );
  INV_X1 U6735 ( .A(n6121), .ZN(n6113) );
  AOI22_X1 U6736 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6627), .ZN(n6080) );
  OAI21_X1 U6737 ( .B1(n5076), .B2(n6115), .A(n6080), .ZN(U3184) );
  INV_X1 U6738 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6083) );
  AOI22_X1 U6739 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6627), .ZN(n6081) );
  OAI21_X1 U6740 ( .B1(n6083), .B2(n6121), .A(n6081), .ZN(U3185) );
  AOI22_X1 U6741 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6627), .ZN(n6082) );
  OAI21_X1 U6742 ( .B1(n6083), .B2(n6115), .A(n6082), .ZN(U3186) );
  AOI22_X1 U6743 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6627), .ZN(n6084) );
  OAI21_X1 U6744 ( .B1(n6362), .B2(n6121), .A(n6084), .ZN(U3187) );
  INV_X1 U6745 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6388) );
  AOI22_X1 U6746 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6627), .ZN(n6085) );
  OAI21_X1 U6747 ( .B1(n6388), .B2(n6121), .A(n6085), .ZN(U3188) );
  INV_X1 U6748 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6396) );
  AOI22_X1 U6749 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6627), .ZN(n6086) );
  OAI21_X1 U6750 ( .B1(n6396), .B2(n6121), .A(n6086), .ZN(U3189) );
  AOI22_X1 U6751 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6627), .ZN(n6087) );
  OAI21_X1 U6752 ( .B1(n6396), .B2(n6115), .A(n6087), .ZN(U3190) );
  AOI22_X1 U6753 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6627), .ZN(n6088) );
  OAI21_X1 U6754 ( .B1(n6416), .B2(n6121), .A(n6088), .ZN(U3191) );
  AOI22_X1 U6755 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6627), .ZN(n6089) );
  OAI21_X1 U6756 ( .B1(n6416), .B2(n6115), .A(n6089), .ZN(U3192) );
  AOI22_X1 U6757 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6627), .ZN(n6090) );
  OAI21_X1 U6758 ( .B1(n6433), .B2(n6115), .A(n6090), .ZN(U3193) );
  INV_X1 U6759 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6451) );
  AOI22_X1 U6760 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6627), .ZN(n6091) );
  OAI21_X1 U6761 ( .B1(n6451), .B2(n6121), .A(n6091), .ZN(U3194) );
  INV_X1 U6762 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6450) );
  AOI22_X1 U6763 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6627), .ZN(n6092) );
  OAI21_X1 U6764 ( .B1(n6450), .B2(n6121), .A(n6092), .ZN(U3195) );
  AOI22_X1 U6765 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6627), .ZN(n6093) );
  OAI21_X1 U6766 ( .B1(n5706), .B2(n6121), .A(n6093), .ZN(U3196) );
  AOI22_X1 U6767 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6627), .ZN(n6094) );
  OAI21_X1 U6768 ( .B1(n5706), .B2(n6115), .A(n6094), .ZN(U3197) );
  AOI22_X1 U6769 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6627), .ZN(n6095) );
  OAI21_X1 U6770 ( .B1(n6479), .B2(n6121), .A(n6095), .ZN(U3198) );
  AOI22_X1 U6771 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6627), .ZN(n6096) );
  OAI21_X1 U6772 ( .B1(n6479), .B2(n6115), .A(n6096), .ZN(U3199) );
  AOI22_X1 U6773 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6627), .ZN(n6097) );
  OAI21_X1 U6774 ( .B1(n6496), .B2(n6121), .A(n6097), .ZN(U3200) );
  AOI22_X1 U6775 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6627), .ZN(n6098) );
  OAI21_X1 U6776 ( .B1(n6100), .B2(n6121), .A(n6098), .ZN(U3201) );
  AOI22_X1 U6777 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6627), .ZN(n6099) );
  OAI21_X1 U6778 ( .B1(n6100), .B2(n6115), .A(n6099), .ZN(U3202) );
  AOI22_X1 U6779 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6627), .ZN(n6101) );
  OAI21_X1 U6780 ( .B1(n6102), .B2(n6115), .A(n6101), .ZN(U3203) );
  AOI22_X1 U6781 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6627), .ZN(n6103) );
  OAI21_X1 U6782 ( .B1(n6517), .B2(n6121), .A(n6103), .ZN(U3204) );
  AOI22_X1 U6783 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6627), .ZN(n6104) );
  OAI21_X1 U6784 ( .B1(n6105), .B2(n6121), .A(n6104), .ZN(U3205) );
  AOI22_X1 U6785 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6627), .ZN(n6106) );
  OAI21_X1 U6786 ( .B1(n6108), .B2(n6121), .A(n6106), .ZN(U3206) );
  AOI22_X1 U6787 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6627), .ZN(n6107) );
  OAI21_X1 U6788 ( .B1(n6108), .B2(n6115), .A(n6107), .ZN(U3207) );
  AOI22_X1 U6789 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6627), .ZN(n6109) );
  OAI21_X1 U6790 ( .B1(n5417), .B2(n6121), .A(n6109), .ZN(U3208) );
  AOI22_X1 U6791 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6627), .ZN(n6110) );
  OAI21_X1 U6792 ( .B1(n6111), .B2(n6121), .A(n6110), .ZN(U3209) );
  AOI22_X1 U6793 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6627), .ZN(n6112) );
  OAI21_X1 U6794 ( .B1(n6116), .B2(n6121), .A(n6112), .ZN(U3210) );
  AOI22_X1 U6795 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6113), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6627), .ZN(n6114) );
  OAI21_X1 U6796 ( .B1(n6116), .B2(n6115), .A(n6114), .ZN(U3211) );
  AOI22_X1 U6797 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6627), .ZN(n6117) );
  OAI21_X1 U6798 ( .B1(n6118), .B2(n6121), .A(n6117), .ZN(U3212) );
  AOI22_X1 U6799 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6119), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6627), .ZN(n6120) );
  OAI21_X1 U6800 ( .B1(n6122), .B2(n6121), .A(n6120), .ZN(U3213) );
  MUX2_X1 U6801 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6627), .Z(U3445) );
  NOR4_X1 U6802 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6132) );
  NOR4_X1 U6803 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6131) );
  INV_X1 U6804 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6611) );
  NOR4_X1 U6805 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U6806 ( .B1(n6137), .B2(n6611), .A(n6123), .ZN(n6129) );
  NOR4_X1 U6807 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6127) );
  NOR4_X1 U6808 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6126) );
  NOR4_X1 U6809 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6125) );
  NOR4_X1 U6810 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6124) );
  NAND4_X1 U6811 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n6128)
         );
  NOR4_X1 U6812 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_31__SCAN_IN), .A3(n6129), .A4(n6128), .ZN(n6130) );
  NAND3_X1 U6813 ( .A1(n6132), .A2(n6131), .A3(n6130), .ZN(n6140) );
  INV_X1 U6814 ( .A(n6140), .ZN(n6144) );
  INV_X1 U6815 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6133) );
  NOR2_X1 U6816 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6140), .ZN(n6142) );
  NAND2_X1 U6817 ( .A1(n6142), .A2(n6611), .ZN(n6138) );
  NOR2_X1 U6818 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6140), .ZN(n6134) );
  NAND3_X1 U6819 ( .A1(n6134), .A2(n6137), .A3(n6611), .ZN(n6139) );
  OAI211_X1 U6820 ( .C1(n6144), .C2(n6133), .A(n6138), .B(n6139), .ZN(U2795)
         );
  MUX2_X1 U6821 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6627), .Z(U3446) );
  NAND2_X1 U6822 ( .A1(n6134), .A2(n5076), .ZN(n6143) );
  NOR2_X1 U6823 ( .A1(n6140), .A2(n5076), .ZN(n6135) );
  AOI22_X1 U6824 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6140), .B1(
        REIP_REG_0__SCAN_IN), .B2(n6135), .ZN(n6136) );
  OAI221_X1 U6825 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6138), .C1(n6137), 
        .C2(n6143), .A(n6136), .ZN(U3468) );
  MUX2_X1 U6826 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6627), .Z(U3447) );
  OAI221_X1 U6827 ( .B1(n6142), .B2(n6141), .C1(n6142), .C2(n6140), .A(n6139), 
        .ZN(U2794) );
  MUX2_X1 U6828 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6627), .Z(U3448) );
  OAI21_X1 U6829 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(n6144), .A(n6143), .ZN(
        n6145) );
  INV_X1 U6830 ( .A(n6145), .ZN(U3469) );
  INV_X1 U6831 ( .A(n6146), .ZN(n6174) );
  AOI22_X1 U6832 ( .A1(n6174), .A2(n6159), .B1(n6150), .B2(n6283), .ZN(n6147)
         );
  OAI21_X1 U6833 ( .B1(n6162), .B2(n6148), .A(n6147), .ZN(U2857) );
  INV_X1 U6834 ( .A(n6149), .ZN(n6469) );
  AOI22_X1 U6835 ( .A1(n6469), .A2(n6159), .B1(n6150), .B2(n6464), .ZN(n6151)
         );
  OAI21_X1 U6836 ( .B1(n6162), .B2(n6152), .A(n6151), .ZN(U2845) );
  OR2_X1 U6837 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U6838 ( .A1(n6156), .A2(n6155), .ZN(n6355) );
  NOR2_X1 U6839 ( .A1(n6157), .A2(n6355), .ZN(n6158) );
  AOI21_X1 U6840 ( .B1(n6357), .B2(n6159), .A(n6158), .ZN(n6160) );
  OAI21_X1 U6841 ( .B1(n6162), .B2(n6161), .A(n6160), .ZN(U2855) );
  NOR2_X1 U6842 ( .A1(n6163), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6164)
         );
  OR2_X1 U6843 ( .A1(n6165), .A2(n6164), .ZN(n6333) );
  INV_X1 U6844 ( .A(n6333), .ZN(n6168) );
  NAND2_X1 U6845 ( .A1(n6166), .A2(n6209), .ZN(n6167) );
  AOI22_X1 U6846 ( .A1(n6212), .A2(n6168), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6167), .ZN(n6169) );
  NAND2_X1 U6847 ( .A1(n6322), .A2(REIP_REG_0__SCAN_IN), .ZN(n6337) );
  OAI211_X1 U6848 ( .C1(n6170), .C2(n6188), .A(n6169), .B(n6337), .ZN(U2986)
         );
  AOI22_X1 U6849 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6210), .B1(n6322), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6176) );
  XNOR2_X1 U6850 ( .A(n6172), .B(n6291), .ZN(n6173) );
  XNOR2_X1 U6851 ( .A(n6171), .B(n6173), .ZN(n6286) );
  AOI22_X1 U6852 ( .A1(n6211), .A2(n6174), .B1(n6286), .B2(n6212), .ZN(n6175)
         );
  OAI211_X1 U6853 ( .C1(n6216), .C2(n6177), .A(n6176), .B(n6175), .ZN(U2984)
         );
  AOI22_X1 U6854 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n6210), .B1(n6322), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U6855 ( .A1(n6178), .A2(n6179), .ZN(n6180) );
  AND2_X1 U6856 ( .A1(n6181), .A2(n6180), .ZN(n6264) );
  AOI22_X1 U6857 ( .A1(n6264), .A2(n6212), .B1(n6211), .B2(n6357), .ZN(n6182)
         );
  OAI211_X1 U6858 ( .C1(n6216), .C2(n6360), .A(n6183), .B(n6182), .ZN(U2982)
         );
  AOI22_X1 U6859 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6210), .B1(n6322), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n6191) );
  OR2_X1 U6860 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  AND2_X1 U6861 ( .A1(n6187), .A2(n6186), .ZN(n6278) );
  NOR2_X1 U6862 ( .A1(n6368), .A2(n6188), .ZN(n6189) );
  AOI21_X1 U6863 ( .B1(n6278), .B2(n6212), .A(n6189), .ZN(n6190) );
  OAI211_X1 U6864 ( .C1(n6216), .C2(n6376), .A(n6191), .B(n6190), .ZN(U2981)
         );
  AOI22_X1 U6865 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6210), .B1(n6322), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6196) );
  XNOR2_X1 U6866 ( .A(n6193), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6194)
         );
  XNOR2_X1 U6867 ( .A(n6192), .B(n6194), .ZN(n6272) );
  AOI22_X1 U6868 ( .A1(n6272), .A2(n6212), .B1(n6211), .B2(n6385), .ZN(n6195)
         );
  OAI211_X1 U6869 ( .C1(n6216), .C2(n6387), .A(n6196), .B(n6195), .ZN(U2980)
         );
  INV_X1 U6870 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6393) );
  INV_X1 U6871 ( .A(n6198), .ZN(n6199) );
  XNOR2_X1 U6872 ( .A(n6197), .B(n6199), .ZN(n6297) );
  INV_X1 U6873 ( .A(n6400), .ZN(n6200) );
  AOI222_X1 U6874 ( .A1(n6297), .A2(n6212), .B1(n6211), .B2(n6397), .C1(n6200), 
        .C2(n6206), .ZN(n6202) );
  AND2_X1 U6875 ( .A1(n6322), .A2(REIP_REG_7__SCAN_IN), .ZN(n6298) );
  INV_X1 U6876 ( .A(n6298), .ZN(n6201) );
  OAI211_X1 U6877 ( .C1(n6209), .C2(n6393), .A(n6202), .B(n6201), .ZN(U2979)
         );
  OAI21_X1 U6878 ( .B1(n6205), .B2(n6204), .A(n6203), .ZN(n6245) );
  INV_X1 U6879 ( .A(n6462), .ZN(n6207) );
  AOI222_X1 U6880 ( .A1(n6245), .A2(n6212), .B1(n6207), .B2(n6206), .C1(n6211), 
        .C2(n6459), .ZN(n6208) );
  NAND2_X1 U6881 ( .A1(n6322), .A2(REIP_REG_13__SCAN_IN), .ZN(n6248) );
  OAI211_X1 U6882 ( .C1(n6209), .C2(n4072), .A(n6208), .B(n6248), .ZN(U2973)
         );
  AOI22_X1 U6883 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6210), .B1(n6322), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n6215) );
  AOI22_X1 U6884 ( .A1(n6213), .A2(n6212), .B1(n6211), .B2(n6640), .ZN(n6214)
         );
  OAI211_X1 U6885 ( .C1(n6216), .C2(n6502), .A(n6215), .B(n6214), .ZN(U2968)
         );
  NOR2_X1 U6886 ( .A1(n6630), .A2(D_C_N_REG_SCAN_IN), .ZN(n6217) );
  AOI22_X1 U6887 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6630), .B1(n6218), .B2(
        n6217), .ZN(U2791) );
  AOI22_X1 U6888 ( .A1(n6630), .A2(READREQUEST_REG_SCAN_IN), .B1(n6219), .B2(
        n6627), .ZN(U3470) );
  AND2_X1 U6889 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6614) );
  NOR2_X1 U6890 ( .A1(n4566), .A2(n6613), .ZN(n6622) );
  AOI21_X1 U6891 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n6622), .ZN(n6222)
         );
  NOR2_X1 U6892 ( .A1(n6220), .A2(n6619), .ZN(n6616) );
  INV_X1 U6893 ( .A(n6616), .ZN(n6623) );
  OAI211_X1 U6894 ( .C1(n6614), .C2(n6222), .A(n6221), .B(n6623), .ZN(U3182)
         );
  NOR2_X1 U6895 ( .A1(READY_N), .A2(n6594), .ZN(n6223) );
  OAI21_X1 U6896 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6223), .A(n6586), .ZN(
        n6225) );
  OAI21_X1 U6897 ( .B1(n6232), .B2(n6225), .A(n6224), .ZN(U3150) );
  AOI211_X1 U6898 ( .C1(n6228), .C2(n6619), .A(n6227), .B(n6226), .ZN(n6235)
         );
  OAI21_X1 U6899 ( .B1(n6229), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U6900 ( .B1(n6231), .B2(n6230), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6234) );
  NOR2_X1 U6901 ( .A1(n6235), .A2(n6232), .ZN(n6233) );
  AOI22_X1 U6902 ( .A1(n6613), .A2(n6235), .B1(n6234), .B2(n6233), .ZN(U3472)
         );
  AOI22_X1 U6903 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6236), .B1(n6322), .B2(REIP_REG_19__SCAN_IN), .ZN(n6240) );
  AOI22_X1 U6904 ( .A1(n6238), .A2(n6327), .B1(n6326), .B2(n6237), .ZN(n6239)
         );
  OAI211_X1 U6905 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6241), .A(n6240), .B(n6239), .ZN(U2999) );
  NAND3_X1 U6906 ( .A1(n6259), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6246) );
  INV_X1 U6907 ( .A(n6246), .ZN(n6257) );
  NAND2_X1 U6908 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6242), .ZN(n6243)
         );
  OAI22_X1 U6909 ( .A1(n6288), .A2(n6244), .B1(n6247), .B2(n6243), .ZN(n6256)
         );
  INV_X1 U6910 ( .A(n6245), .ZN(n6254) );
  NOR2_X1 U6911 ( .A1(n6247), .A2(n6246), .ZN(n6251) );
  OAI21_X1 U6912 ( .B1(n6339), .B2(n6249), .A(n6248), .ZN(n6250) );
  AOI21_X1 U6913 ( .B1(n6252), .B2(n6251), .A(n6250), .ZN(n6253) );
  OAI21_X1 U6914 ( .B1(n6254), .B2(n6334), .A(n6253), .ZN(n6255) );
  AOI21_X1 U6915 ( .B1(n6257), .B2(n6256), .A(n6255), .ZN(n6258) );
  OAI21_X1 U6916 ( .B1(n6260), .B2(n6259), .A(n6258), .ZN(U3005) );
  INV_X1 U6917 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6261) );
  OAI22_X1 U6918 ( .A1(n6339), .A2(n6355), .B1(n6262), .B2(n6261), .ZN(n6263)
         );
  INV_X1 U6919 ( .A(n6263), .ZN(n6267) );
  AOI22_X1 U6920 ( .A1(n6269), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6327), 
        .B2(n6264), .ZN(n6266) );
  INV_X1 U6921 ( .A(n6277), .ZN(n6271) );
  OAI211_X1 U6922 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6276), .B(n6271), .ZN(n6265) );
  NAND3_X1 U6923 ( .A1(n6267), .A2(n6266), .A3(n6265), .ZN(U3014) );
  NAND3_X1 U6924 ( .A1(n6277), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6276), 
        .ZN(n6275) );
  INV_X1 U6925 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6274) );
  AOI21_X1 U6926 ( .B1(n6288), .B2(n6268), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6270) );
  AOI211_X1 U6927 ( .C1(n6271), .C2(n6276), .A(n6270), .B(n6269), .ZN(n6282)
         );
  AOI222_X1 U6928 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6322), .B1(n6326), .B2(
        n6379), .C1(n6327), .C2(n6272), .ZN(n6273) );
  OAI221_X1 U6929 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6275), .C1(n6274), .C2(n6282), .A(n6273), .ZN(U3012) );
  AOI21_X1 U6930 ( .B1(n6277), .B2(n6276), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6281) );
  AOI22_X1 U6931 ( .A1(n6278), .A2(n6327), .B1(n6326), .B2(n6365), .ZN(n6280)
         );
  NAND2_X1 U6932 ( .A1(n6322), .A2(REIP_REG_5__SCAN_IN), .ZN(n6279) );
  OAI211_X1 U6933 ( .C1(n6282), .C2(n6281), .A(n6280), .B(n6279), .ZN(U3013)
         );
  AOI22_X1 U6934 ( .A1(n6326), .A2(n6283), .B1(n6322), .B2(REIP_REG_2__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U6935 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6285) );
  OAI21_X1 U6936 ( .B1(n6285), .B2(n6288), .A(n6284), .ZN(n6287) );
  AOI22_X1 U6937 ( .A1(n6287), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6327), 
        .B2(n6286), .ZN(n6295) );
  INV_X1 U6938 ( .A(n6288), .ZN(n6290) );
  NAND2_X1 U6939 ( .A1(n6290), .A2(n6289), .ZN(n6294) );
  NAND3_X1 U6940 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6292), .A3(n6291), 
        .ZN(n6293) );
  NAND4_X1 U6941 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(U3016)
         );
  NAND2_X1 U6942 ( .A1(n6297), .A2(n6327), .ZN(n6300) );
  AOI21_X1 U6943 ( .B1(n6326), .B2(n6391), .A(n6298), .ZN(n6299) );
  OAI211_X1 U6944 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6301), .A(n6300), 
        .B(n6299), .ZN(n6302) );
  INV_X1 U6945 ( .A(n6302), .ZN(n6303) );
  OAI21_X1 U6946 ( .B1(n4459), .B2(n6304), .A(n6303), .ZN(U3011) );
  AOI21_X1 U6947 ( .B1(n6326), .B2(n6306), .A(n6305), .ZN(n6310) );
  AOI22_X1 U6948 ( .A1(n6308), .A2(n6327), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6307), .ZN(n6309) );
  OAI211_X1 U6949 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6311), .A(n6310), .B(n6309), .ZN(U3003) );
  NAND2_X1 U6950 ( .A1(n6312), .A2(n4474), .ZN(n6319) );
  INV_X1 U6951 ( .A(n6313), .ZN(n6314) );
  AOI22_X1 U6952 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6314), .B1(n6322), .B2(REIP_REG_17__SCAN_IN), .ZN(n6318) );
  AOI22_X1 U6953 ( .A1(n6316), .A2(n6327), .B1(n6326), .B2(n6315), .ZN(n6317)
         );
  OAI211_X1 U6954 ( .C1(n6320), .C2(n6319), .A(n6318), .B(n6317), .ZN(U3001)
         );
  AOI22_X1 U6955 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6322), .B1(n6321), .B2(
        n6331), .ZN(n6330) );
  INV_X1 U6956 ( .A(n6323), .ZN(n6328) );
  INV_X1 U6957 ( .A(n6324), .ZN(n6325) );
  AOI22_X1 U6958 ( .A1(n6328), .A2(n6327), .B1(n6326), .B2(n6325), .ZN(n6329)
         );
  OAI211_X1 U6959 ( .C1(n6332), .C2(n6331), .A(n6330), .B(n6329), .ZN(U2993)
         );
  OR2_X1 U6960 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  NAND2_X1 U6961 ( .A1(n6336), .A2(n6335), .ZN(n6342) );
  OAI211_X1 U6962 ( .C1(n6340), .C2(n6339), .A(n6338), .B(n6337), .ZN(n6341)
         );
  NOR2_X1 U6963 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  OAI221_X1 U6964 ( .B1(n6346), .B2(n6345), .C1(n6346), .C2(n6344), .A(n6343), 
        .ZN(U3018) );
  AOI22_X1 U6965 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n6524), .B1(
        EBX_REG_4__SCAN_IN), .B2(n6506), .ZN(n6347) );
  INV_X1 U6966 ( .A(n6347), .ZN(n6348) );
  AOI211_X1 U6967 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6349), .A(n6499), .B(n6348), 
        .ZN(n6359) );
  NOR3_X1 U6968 ( .A1(n6521), .A2(REIP_REG_4__SCAN_IN), .A3(n6350), .ZN(n6351)
         );
  AOI21_X1 U6969 ( .B1(n6353), .B2(n6352), .A(n6351), .ZN(n6354) );
  OAI21_X1 U6970 ( .B1(n6510), .B2(n6355), .A(n6354), .ZN(n6356) );
  AOI21_X1 U6971 ( .B1(n6357), .B2(n6369), .A(n6356), .ZN(n6358) );
  OAI211_X1 U6972 ( .C1(n6360), .C2(n6515), .A(n6359), .B(n6358), .ZN(U2823)
         );
  OR2_X1 U6973 ( .A1(n6521), .A2(n6377), .ZN(n6361) );
  AND2_X1 U6974 ( .A1(n6361), .A2(n6402), .ZN(n6389) );
  OAI21_X1 U6975 ( .B1(n6521), .B2(n6363), .A(n6362), .ZN(n6364) );
  INV_X1 U6976 ( .A(n6364), .ZN(n6373) );
  AOI22_X1 U6977 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6506), .B1(n6526), .B2(n6365), 
        .ZN(n6366) );
  NAND2_X1 U6978 ( .A1(n6455), .A2(n6366), .ZN(n6367) );
  AOI21_X1 U6979 ( .B1(n6524), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6367), 
        .ZN(n6372) );
  INV_X1 U6980 ( .A(n6368), .ZN(n6370) );
  NAND2_X1 U6981 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  OAI211_X1 U6982 ( .C1(n6389), .C2(n6373), .A(n6372), .B(n6371), .ZN(n6374)
         );
  INV_X1 U6983 ( .A(n6374), .ZN(n6375) );
  OAI21_X1 U6984 ( .B1(n6376), .B2(n6515), .A(n6375), .ZN(U2822) );
  AOI22_X1 U6985 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6524), .B1(
        EBX_REG_6__SCAN_IN), .B2(n6506), .ZN(n6383) );
  INV_X1 U6986 ( .A(n6377), .ZN(n6378) );
  OR2_X1 U6987 ( .A1(n6521), .A2(n6378), .ZN(n6390) );
  NAND2_X1 U6988 ( .A1(n6526), .A2(n6379), .ZN(n6380) );
  OAI211_X1 U6989 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6390), .A(n6380), .B(n6455), 
        .ZN(n6381) );
  INV_X1 U6990 ( .A(n6381), .ZN(n6382) );
  OAI211_X1 U6991 ( .C1(n6388), .C2(n6389), .A(n6383), .B(n6382), .ZN(n6384)
         );
  AOI21_X1 U6992 ( .B1(n6530), .B2(n6385), .A(n6384), .ZN(n6386) );
  OAI21_X1 U6993 ( .B1(n6387), .B2(n6515), .A(n6386), .ZN(U2821) );
  NOR2_X1 U6994 ( .A1(n6388), .A2(n6390), .ZN(n6404) );
  OAI21_X1 U6995 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6390), .A(n6389), .ZN(n6395)
         );
  AOI22_X1 U6996 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6506), .B1(n6526), .B2(n6391), 
        .ZN(n6392) );
  OAI211_X1 U6997 ( .C1(n6457), .C2(n6393), .A(n6392), .B(n6455), .ZN(n6394)
         );
  AOI221_X1 U6998 ( .B1(n6404), .B2(n6396), .C1(n6395), .C2(
        REIP_REG_7__SCAN_IN), .A(n6394), .ZN(n6399) );
  NAND2_X1 U6999 ( .A1(n6397), .A2(n6530), .ZN(n6398) );
  OAI211_X1 U7000 ( .C1(n6515), .C2(n6400), .A(n6399), .B(n6398), .ZN(U2820)
         );
  INV_X1 U7001 ( .A(n6415), .ZN(n6401) );
  OR2_X1 U7002 ( .A1(n6521), .A2(n6401), .ZN(n6403) );
  AND2_X1 U7003 ( .A1(n6403), .A2(n6402), .ZN(n6429) );
  AOI21_X1 U7004 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6404), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6413) );
  OAI22_X1 U7005 ( .A1(n6406), .A2(n6533), .B1(n6510), .B2(n6405), .ZN(n6407)
         );
  AOI211_X1 U7006 ( .C1(n6524), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6499), 
        .B(n6407), .ZN(n6412) );
  INV_X1 U7007 ( .A(n6408), .ZN(n6409) );
  AOI22_X1 U7008 ( .A1(n6410), .A2(n6530), .B1(n6528), .B2(n6409), .ZN(n6411)
         );
  OAI211_X1 U7009 ( .C1(n6429), .C2(n6413), .A(n6412), .B(n6411), .ZN(U2819)
         );
  AOI22_X1 U7010 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6524), .B1(n6526), 
        .B2(n6414), .ZN(n6422) );
  NOR3_X1 U7011 ( .A1(n6521), .A2(REIP_REG_9__SCAN_IN), .A3(n6415), .ZN(n6431)
         );
  NOR2_X1 U7012 ( .A1(n6429), .A2(n6416), .ZN(n6417) );
  AOI211_X1 U7013 ( .C1(n6506), .C2(EBX_REG_9__SCAN_IN), .A(n6431), .B(n6417), 
        .ZN(n6421) );
  AOI22_X1 U7014 ( .A1(n6419), .A2(n6530), .B1(n6528), .B2(n6418), .ZN(n6420)
         );
  NAND4_X1 U7015 ( .A1(n6422), .A2(n6421), .A3(n6420), .A4(n6455), .ZN(U2818)
         );
  OAI22_X1 U7016 ( .A1(n6424), .A2(n6533), .B1(n6510), .B2(n6423), .ZN(n6425)
         );
  AOI211_X1 U7017 ( .C1(n6524), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6499), 
        .B(n6425), .ZN(n6438) );
  OAI22_X1 U7018 ( .A1(n6427), .A2(n6490), .B1(n6426), .B2(n6515), .ZN(n6428)
         );
  INV_X1 U7019 ( .A(n6428), .ZN(n6437) );
  INV_X1 U7020 ( .A(n6429), .ZN(n6430) );
  OAI21_X1 U7021 ( .B1(n6431), .B2(n6430), .A(REIP_REG_10__SCAN_IN), .ZN(n6436) );
  NAND3_X1 U7022 ( .A1(n6434), .A2(n6433), .A3(n6432), .ZN(n6435) );
  NAND4_X1 U7023 ( .A1(n6438), .A2(n6437), .A3(n6436), .A4(n6435), .ZN(U2817)
         );
  AOI22_X1 U7024 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6524), .B1(n6526), 
        .B2(n6439), .ZN(n6449) );
  INV_X1 U7025 ( .A(n6454), .ZN(n6443) );
  OR3_X1 U7026 ( .A1(n6521), .A2(REIP_REG_11__SCAN_IN), .A3(n6440), .ZN(n6441)
         );
  OAI21_X1 U7027 ( .B1(n6443), .B2(n6442), .A(n6441), .ZN(n6444) );
  AOI21_X1 U7028 ( .B1(EBX_REG_11__SCAN_IN), .B2(n6506), .A(n6444), .ZN(n6448)
         );
  AOI22_X1 U7029 ( .A1(n6446), .A2(n6530), .B1(n6528), .B2(n6445), .ZN(n6447)
         );
  NAND4_X1 U7030 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6455), .ZN(U2816)
         );
  AOI21_X1 U7031 ( .B1(n6451), .B2(n6450), .A(n6465), .ZN(n6452) );
  NAND2_X1 U7032 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n6466) );
  AOI22_X1 U7033 ( .A1(n6526), .A2(n6453), .B1(n6452), .B2(n6466), .ZN(n6461)
         );
  AOI22_X1 U7034 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6506), .B1(
        REIP_REG_13__SCAN_IN), .B2(n6454), .ZN(n6456) );
  OAI211_X1 U7035 ( .C1(n6457), .C2(n4072), .A(n6456), .B(n6455), .ZN(n6458)
         );
  AOI21_X1 U7036 ( .B1(n6459), .B2(n6530), .A(n6458), .ZN(n6460) );
  OAI211_X1 U7037 ( .C1(n6462), .C2(n6515), .A(n6461), .B(n6460), .ZN(U2814)
         );
  INV_X1 U7038 ( .A(n6477), .ZN(n6463) );
  AOI22_X1 U7039 ( .A1(n6526), .A2(n6464), .B1(REIP_REG_14__SCAN_IN), .B2(
        n6463), .ZN(n6473) );
  AOI22_X1 U7040 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n6524), .B1(
        EBX_REG_14__SCAN_IN), .B2(n6506), .ZN(n6472) );
  NOR3_X1 U7041 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6466), .A3(n6465), .ZN(n6467) );
  NOR2_X1 U7042 ( .A1(n6467), .A2(n6499), .ZN(n6471) );
  AOI22_X1 U7043 ( .A1(n6469), .A2(n6530), .B1(n6468), .B2(n6528), .ZN(n6470)
         );
  NAND4_X1 U7044 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(U2813)
         );
  NOR2_X1 U7045 ( .A1(n6475), .A2(n6474), .ZN(n6485) );
  AOI22_X1 U7046 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6506), .B1(n6485), .B2(n6479), .ZN(n6476) );
  OAI221_X1 U7047 ( .B1(n6479), .B2(n6478), .C1(n6479), .C2(n6477), .A(n6476), 
        .ZN(n6480) );
  AOI211_X1 U7048 ( .C1(n6524), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6499), 
        .B(n6480), .ZN(n6483) );
  AOI22_X1 U7049 ( .A1(n6631), .A2(n6530), .B1(n6528), .B2(n6481), .ZN(n6482)
         );
  OAI211_X1 U7050 ( .C1(n6510), .C2(n6484), .A(n6483), .B(n6482), .ZN(U2811)
         );
  AOI21_X1 U7051 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6485), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6494) );
  AOI22_X1 U7052 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6524), .B1(
        EBX_REG_17__SCAN_IN), .B2(n6506), .ZN(n6486) );
  INV_X1 U7053 ( .A(n6486), .ZN(n6487) );
  AOI211_X1 U7054 ( .C1(n6528), .C2(n6488), .A(n6499), .B(n6487), .ZN(n6493)
         );
  OAI22_X1 U7055 ( .A1(n6636), .A2(n6490), .B1(n6510), .B2(n6489), .ZN(n6491)
         );
  INV_X1 U7056 ( .A(n6491), .ZN(n6492) );
  OAI211_X1 U7057 ( .C1(n6494), .C2(n6495), .A(n6493), .B(n6492), .ZN(U2810)
         );
  OAI22_X1 U7058 ( .A1(n6497), .A2(n6533), .B1(n6496), .B2(n6495), .ZN(n6498)
         );
  AOI211_X1 U7059 ( .C1(n6524), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6499), 
        .B(n6498), .ZN(n6501) );
  OAI211_X1 U7060 ( .C1(n6502), .C2(n6515), .A(n6501), .B(n6500), .ZN(n6503)
         );
  AOI21_X1 U7061 ( .B1(n6640), .B2(n6530), .A(n6503), .ZN(n6504) );
  OAI21_X1 U7062 ( .B1(n6505), .B2(n6510), .A(n6504), .ZN(U2809) );
  AOI22_X1 U7063 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6524), .B1(
        EBX_REG_20__SCAN_IN), .B2(n6506), .ZN(n6514) );
  INV_X1 U7064 ( .A(n6507), .ZN(n6643) );
  AOI21_X1 U7065 ( .B1(REIP_REG_19__SCAN_IN), .B2(n6508), .A(
        REIP_REG_20__SCAN_IN), .ZN(n6509) );
  OAI22_X1 U7066 ( .A1(n6511), .A2(n6510), .B1(n6518), .B2(n6509), .ZN(n6512)
         );
  AOI21_X1 U7067 ( .B1(n6643), .B2(n6530), .A(n6512), .ZN(n6513) );
  OAI211_X1 U7068 ( .C1(n6516), .C2(n6515), .A(n6514), .B(n6513), .ZN(U2807)
         );
  AOI21_X1 U7069 ( .B1(n6519), .B2(n6518), .A(n6517), .ZN(n6523) );
  NOR3_X1 U7070 ( .A1(n6521), .A2(REIP_REG_22__SCAN_IN), .A3(n6520), .ZN(n6522) );
  AOI211_X1 U7071 ( .C1(n6524), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n6523), 
        .B(n6522), .ZN(n6532) );
  INV_X1 U7072 ( .A(n6525), .ZN(n6527) );
  AOI222_X1 U7073 ( .A1(n6646), .A2(n6530), .B1(n6529), .B2(n6528), .C1(n6527), 
        .C2(n6526), .ZN(n6531) );
  OAI211_X1 U7074 ( .C1(n6534), .C2(n6533), .A(n6532), .B(n6531), .ZN(U2805)
         );
  OAI21_X1 U7075 ( .B1(n6537), .B2(n6536), .A(n6535), .ZN(U2793) );
  INV_X1 U7076 ( .A(n6538), .ZN(n6541) );
  OAI22_X1 U7077 ( .A1(n6541), .A2(n6540), .B1(n6539), .B2(n6590), .ZN(n6543)
         );
  INV_X1 U7078 ( .A(n6542), .ZN(n6549) );
  MUX2_X1 U7079 ( .A(n6544), .B(n6543), .S(n6549), .Z(U3456) );
  INV_X1 U7080 ( .A(n6545), .ZN(n6546) );
  NAND3_X1 U7081 ( .A1(n6547), .A2(n6734), .A3(n6546), .ZN(n6548) );
  OAI21_X1 U7082 ( .B1(n6549), .B2(n4517), .A(n6548), .ZN(U3455) );
  OAI21_X1 U7083 ( .B1(n6550), .B2(n3566), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .ZN(n6551) );
  NOR2_X1 U7084 ( .A1(n6552), .A2(n6551), .ZN(n6553) );
  INV_X1 U7085 ( .A(n6553), .ZN(n6557) );
  OAI22_X1 U7086 ( .A1(n6555), .A2(n6554), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6553), .ZN(n6556) );
  OAI21_X1 U7087 ( .B1(n6557), .B2(n6793), .A(n6556), .ZN(n6558) );
  AOI222_X1 U7088 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6559), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6558), .C1(n6559), .C2(n6558), 
        .ZN(n6561) );
  AOI222_X1 U7089 ( .A1(n6561), .A2(n6560), .B1(n6561), .B2(n5132), .C1(n6560), 
        .C2(n5132), .ZN(n6562) );
  OR2_X1 U7090 ( .A1(n6562), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6571)
         );
  NOR2_X1 U7091 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6566) );
  NOR2_X1 U7092 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  OAI21_X1 U7093 ( .B1(n6567), .B2(n6566), .A(n6565), .ZN(n6568) );
  NOR2_X1 U7094 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  NAND2_X1 U7095 ( .A1(n6599), .A2(n6572), .ZN(n6574) );
  NAND2_X1 U7096 ( .A1(READY_N), .A2(n6228), .ZN(n6573) );
  NAND2_X1 U7097 ( .A1(n6574), .A2(n6573), .ZN(n6578) );
  OR2_X1 U7098 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  OAI221_X1 U7099 ( .B1(n6579), .B2(READY_N), .C1(n6579), .C2(n6797), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6592) );
  NAND3_X1 U7100 ( .A1(n6580), .A2(STATE2_REG_0__SCAN_IN), .A3(n6619), .ZN(
        n6581) );
  NAND3_X1 U7101 ( .A1(n6581), .A2(n6598), .A3(n6589), .ZN(n6582) );
  OAI21_X1 U7102 ( .B1(n6587), .B2(n6589), .A(n6582), .ZN(n6584) );
  OAI211_X1 U7103 ( .C1(n6585), .C2(n6592), .A(n6584), .B(n6583), .ZN(U3149)
         );
  OAI221_X1 U7104 ( .B1(n6734), .B2(STATE2_REG_0__SCAN_IN), .C1(n6734), .C2(
        n6589), .A(n6586), .ZN(U3453) );
  NAND2_X1 U7105 ( .A1(n6588), .A2(n6587), .ZN(n6607) );
  OAI21_X1 U7106 ( .B1(n6591), .B2(n6590), .A(n6589), .ZN(n6593) );
  OAI221_X1 U7107 ( .B1(n6607), .B2(n6594), .C1(n6593), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6592), .ZN(n6595) );
  INV_X1 U7108 ( .A(n6595), .ZN(n6597) );
  OAI211_X1 U7109 ( .C1(n6599), .C2(n6598), .A(n6597), .B(n6596), .ZN(U3148)
         );
  INV_X1 U7110 ( .A(n6600), .ZN(n6603) );
  INV_X1 U7111 ( .A(n6601), .ZN(n6602) );
  AOI22_X1 U7112 ( .A1(n6604), .A2(n6603), .B1(n6602), .B2(n6799), .ZN(n6605)
         );
  OAI221_X1 U7113 ( .B1(n6608), .B2(n6607), .C1(n6606), .C2(n6794), .A(n6605), 
        .ZN(U3465) );
  INV_X1 U7114 ( .A(n6609), .ZN(n6610) );
  OAI21_X1 U7115 ( .B1(n6612), .B2(n6817), .A(n6610), .ZN(U2792) );
  OAI21_X1 U7116 ( .B1(n6612), .B2(n6611), .A(n6610), .ZN(U3452) );
  AOI211_X1 U7117 ( .C1(STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n6614), .B(n6613), 
        .ZN(n6618) );
  AOI221_X1 U7118 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6621), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6625) );
  AOI21_X1 U7119 ( .B1(n6616), .B2(n6615), .A(n6625), .ZN(n6617) );
  OAI21_X1 U7120 ( .B1(n6630), .B2(n6618), .A(n6617), .ZN(U3181) );
  AOI221_X1 U7121 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6619), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6620) );
  AOI221_X1 U7122 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6620), .C2(HOLD), .A(n4566), .ZN(n6626) );
  AOI21_X1 U7123 ( .B1(n6622), .B2(n6621), .A(STATE_REG_2__SCAN_IN), .ZN(n6624) );
  OAI22_X1 U7124 ( .A1(n6626), .A2(n6625), .B1(n6624), .B2(n6623), .ZN(U3183)
         );
  AOI22_X1 U7125 ( .A1(n6630), .A2(n6629), .B1(n6628), .B2(n6627), .ZN(U3473)
         );
  INV_X1 U7126 ( .A(n6635), .ZN(n6835) );
  AOI22_X1 U7127 ( .A1(n6631), .A2(n6835), .B1(n6834), .B2(DATAI_16_), .ZN(
        n6633) );
  AOI22_X1 U7128 ( .A1(n6838), .A2(DATAI_0_), .B1(n6837), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7129 ( .A1(n6633), .A2(n6632), .ZN(U2875) );
  INV_X1 U7130 ( .A(n6834), .ZN(n6634) );
  OAI22_X1 U7131 ( .A1(n6636), .A2(n6635), .B1(n6634), .B2(n5965), .ZN(n6637)
         );
  INV_X1 U7132 ( .A(n6637), .ZN(n6639) );
  AOI22_X1 U7133 ( .A1(n6838), .A2(DATAI_1_), .B1(n6837), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U7134 ( .A1(n6639), .A2(n6638), .ZN(U2874) );
  AOI22_X1 U7135 ( .A1(n6640), .A2(n6835), .B1(n6834), .B2(DATAI_18_), .ZN(
        n6642) );
  AOI22_X1 U7136 ( .A1(n6838), .A2(DATAI_2_), .B1(n6837), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7137 ( .A1(n6642), .A2(n6641), .ZN(U2873) );
  AOI22_X1 U7138 ( .A1(n6643), .A2(n6835), .B1(n6834), .B2(DATAI_20_), .ZN(
        n6645) );
  AOI22_X1 U7139 ( .A1(n6838), .A2(DATAI_4_), .B1(n6837), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U7140 ( .A1(n6645), .A2(n6644), .ZN(U2871) );
  AOI22_X1 U7141 ( .A1(n6646), .A2(n6835), .B1(n6834), .B2(DATAI_22_), .ZN(
        n6648) );
  AOI22_X1 U7142 ( .A1(n6838), .A2(DATAI_6_), .B1(n6837), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U7143 ( .A1(n6648), .A2(n6647), .ZN(U2869) );
  NAND3_X1 U7144 ( .A1(n6793), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6659) );
  NOR2_X1 U7145 ( .A1(n6649), .A2(n6768), .ZN(n6651) );
  INV_X1 U7146 ( .A(n6651), .ZN(n6650) );
  AND2_X1 U7147 ( .A1(n4942), .A2(n3455), .ZN(n6737) );
  NOR2_X1 U7148 ( .A1(n6794), .A2(n6659), .ZN(n7079) );
  AOI21_X1 U7149 ( .B1(n6690), .B2(n6737), .A(n7079), .ZN(n6652) );
  OAI22_X1 U7150 ( .A1(n6797), .A2(n6659), .B1(n6650), .B2(n6652), .ZN(n7080)
         );
  INV_X1 U7151 ( .A(n7080), .ZN(n6657) );
  AOI22_X1 U7152 ( .A1(n6827), .A2(n7079), .B1(n7038), .B2(n6830), .ZN(n6656)
         );
  AOI22_X1 U7153 ( .A1(n6652), .A2(n6651), .B1(n6768), .B2(n6659), .ZN(n6653)
         );
  NAND2_X1 U7154 ( .A1(n6806), .A2(n6653), .ZN(n7081) );
  AOI22_X1 U7155 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n7081), .B1(n6829), 
        .B2(n7078), .ZN(n6655) );
  OAI211_X1 U7156 ( .C1(n6657), .C2(n6811), .A(n6656), .B(n6655), .ZN(U3124)
         );
  NAND2_X1 U7157 ( .A1(n4938), .A2(n4939), .ZN(n6748) );
  INV_X1 U7158 ( .A(n6748), .ZN(n6658) );
  NAND2_X1 U7159 ( .A1(n6658), .A2(n5127), .ZN(n6668) );
  INV_X1 U7160 ( .A(n6737), .ZN(n6752) );
  AND2_X1 U7161 ( .A1(n6750), .A2(n6727), .ZN(n6661) );
  INV_X1 U7162 ( .A(n6661), .ZN(n6700) );
  OAI22_X1 U7163 ( .A1(n6752), .A2(n6815), .B1(n6751), .B2(n6700), .ZN(n7086)
         );
  INV_X1 U7164 ( .A(n6659), .ZN(n6660) );
  NAND2_X1 U7165 ( .A1(n6794), .A2(n6660), .ZN(n6662) );
  INV_X1 U7166 ( .A(n6662), .ZN(n7085) );
  AOI22_X1 U7167 ( .A1(n6828), .A2(n7086), .B1(n6827), .B2(n7085), .ZN(n6667)
         );
  NOR2_X1 U7168 ( .A1(n6661), .A2(n6797), .ZN(n6705) );
  AOI211_X1 U7169 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6662), .A(n6705), .B(
        n6755), .ZN(n6665) );
  INV_X1 U7170 ( .A(n6825), .ZN(n6663) );
  NOR2_X1 U7171 ( .A1(n6737), .A2(n6768), .ZN(n6757) );
  OAI211_X1 U7172 ( .C1(n6663), .C2(n6757), .A(n7090), .B(n7046), .ZN(n6664)
         );
  NAND2_X1 U7173 ( .A1(n6752), .A2(n6781), .ZN(n6759) );
  NAND3_X1 U7174 ( .A1(n6665), .A2(n6664), .A3(n6759), .ZN(n7087) );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n7087), .B1(n6830), 
        .B2(n7078), .ZN(n6666) );
  OAI211_X1 U7176 ( .C1(n6764), .C2(n7046), .A(n6667), .B(n6666), .ZN(U3116)
         );
  NAND3_X1 U7177 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4482), .ZN(n6676) );
  NOR2_X1 U7178 ( .A1(n6794), .A2(n6676), .ZN(n7092) );
  AOI22_X1 U7179 ( .A1(n6827), .A2(n7092), .B1(n6829), .B2(n7043), .ZN(n6675)
         );
  INV_X1 U7180 ( .A(n6676), .ZN(n6671) );
  OAI21_X1 U7181 ( .B1(n6668), .B2(n6817), .A(n6808), .ZN(n6673) );
  INV_X1 U7182 ( .A(n6673), .ZN(n6669) );
  OR2_X1 U7183 ( .A1(n3455), .A2(n4942), .ZN(n6776) );
  INV_X1 U7184 ( .A(n6776), .ZN(n6784) );
  AOI21_X1 U7185 ( .B1(n6690), .B2(n6784), .A(n7092), .ZN(n6672) );
  NAND2_X1 U7186 ( .A1(n6669), .A2(n6672), .ZN(n6670) );
  OAI211_X1 U7187 ( .C1(n6808), .C2(n6671), .A(n6670), .B(n6806), .ZN(n7094)
         );
  OAI22_X1 U7188 ( .A1(n6673), .A2(n6672), .B1(n6676), .B2(n6797), .ZN(n7093)
         );
  AOI22_X1 U7189 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n7094), .B1(n6828), 
        .B2(n7093), .ZN(n6674) );
  OAI211_X1 U7190 ( .C1(n6792), .C2(n7046), .A(n6675), .B(n6674), .ZN(U3108)
         );
  NOR2_X1 U7191 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6676), .ZN(n7097)
         );
  NAND2_X1 U7192 ( .A1(n5127), .A2(n6778), .ZN(n6692) );
  NOR2_X2 U7193 ( .A1(n6692), .A2(n6780), .ZN(n7105) );
  AOI22_X1 U7194 ( .A1(n6827), .A2(n7097), .B1(n6829), .B2(n7105), .ZN(n6688)
         );
  NAND2_X1 U7195 ( .A1(n7102), .A2(n6808), .ZN(n6679) );
  INV_X1 U7196 ( .A(n6781), .ZN(n6678) );
  OAI21_X1 U7197 ( .B1(n7105), .B2(n6679), .A(n6678), .ZN(n6683) );
  NAND2_X1 U7198 ( .A1(n6784), .A2(n3458), .ZN(n6685) );
  NAND2_X1 U7199 ( .A1(n6680), .A2(n6751), .ZN(n6787) );
  AOI211_X1 U7200 ( .C1(n6683), .C2(n6685), .A(n6681), .B(n6787), .ZN(n6682)
         );
  OAI21_X1 U7201 ( .B1(n7097), .B2(n6734), .A(n6682), .ZN(n7099) );
  INV_X1 U7202 ( .A(n6683), .ZN(n6686) );
  OAI22_X1 U7203 ( .A1(n6686), .A2(n6685), .B1(n6684), .B2(n6823), .ZN(n7098)
         );
  AOI22_X1 U7204 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n7099), .B1(n6828), 
        .B2(n7098), .ZN(n6687) );
  OAI211_X1 U7205 ( .C1(n7102), .C2(n6792), .A(n6688), .B(n6687), .ZN(U3100)
         );
  NAND3_X1 U7206 ( .A1(n4482), .A2(n6793), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6701) );
  OAI21_X1 U7207 ( .B1(n6692), .B2(n6817), .A(n6808), .ZN(n6696) );
  OR2_X1 U7208 ( .A1(n3455), .A2(n6689), .ZN(n6824) );
  INV_X1 U7209 ( .A(n6824), .ZN(n6795) );
  NOR2_X1 U7210 ( .A1(n6794), .A2(n6701), .ZN(n7104) );
  AOI21_X1 U7211 ( .B1(n6690), .B2(n6795), .A(n7104), .ZN(n6693) );
  OAI22_X1 U7212 ( .A1(n6797), .A2(n6701), .B1(n6696), .B2(n6693), .ZN(n6691)
         );
  AOI22_X1 U7213 ( .A1(n6827), .A2(n7104), .B1(n6829), .B2(n7103), .ZN(n6698)
         );
  INV_X1 U7214 ( .A(n6693), .ZN(n6695) );
  NAND2_X1 U7215 ( .A1(n6768), .A2(n6701), .ZN(n6694) );
  OAI211_X1 U7216 ( .C1(n6696), .C2(n6695), .A(n6806), .B(n6694), .ZN(n7106)
         );
  AOI22_X1 U7217 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n7106), .B1(n6830), 
        .B2(n7105), .ZN(n6697) );
  OAI211_X1 U7218 ( .C1(n7109), .C2(n6811), .A(n6698), .B(n6697), .ZN(U3092)
         );
  INV_X1 U7219 ( .A(n6718), .ZN(n6699) );
  NAND2_X1 U7220 ( .A1(n6699), .A2(n6799), .ZN(n6711) );
  OAI22_X1 U7221 ( .A1(n6815), .A2(n6824), .B1(n6823), .B2(n6700), .ZN(n7111)
         );
  INV_X1 U7222 ( .A(n6701), .ZN(n6702) );
  NAND2_X1 U7223 ( .A1(n6794), .A2(n6702), .ZN(n6706) );
  INV_X1 U7224 ( .A(n6706), .ZN(n7110) );
  AOI22_X1 U7225 ( .A1(n6828), .A2(n7111), .B1(n6827), .B2(n7110), .ZN(n6710)
         );
  NOR2_X1 U7226 ( .A1(n6825), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6704) );
  NAND2_X1 U7227 ( .A1(n6824), .A2(n6808), .ZN(n6814) );
  AOI211_X1 U7228 ( .C1(n6825), .C2(n6814), .A(n7116), .B(n7103), .ZN(n6703)
         );
  NOR2_X1 U7229 ( .A1(n6704), .A2(n6703), .ZN(n6708) );
  AOI211_X1 U7230 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6706), .A(n6705), .B(
        n6787), .ZN(n6707) );
  NAND2_X1 U7231 ( .A1(n6708), .A2(n6707), .ZN(n7112) );
  AOI22_X1 U7232 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n7112), .B1(n6830), 
        .B2(n7103), .ZN(n6709) );
  OAI211_X1 U7233 ( .C1(n6764), .C2(n6711), .A(n6710), .B(n6709), .ZN(U3084)
         );
  NAND2_X1 U7234 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6753), .ZN(n6729) );
  NOR2_X1 U7235 ( .A1(n6712), .A2(n6768), .ZN(n6720) );
  INV_X1 U7236 ( .A(n6720), .ZN(n6716) );
  NOR2_X1 U7237 ( .A1(n3458), .A2(n6713), .ZN(n6796) );
  INV_X1 U7238 ( .A(n6714), .ZN(n7117) );
  AOI21_X1 U7239 ( .B1(n6796), .B2(n6715), .A(n7117), .ZN(n6719) );
  OAI22_X1 U7240 ( .A1(n6797), .A2(n6729), .B1(n6716), .B2(n6719), .ZN(n6717)
         );
  AOI22_X1 U7241 ( .A1(n6827), .A2(n7117), .B1(n6829), .B2(n7118), .ZN(n6723)
         );
  AOI22_X1 U7242 ( .A1(n6720), .A2(n6719), .B1(n6768), .B2(n6729), .ZN(n6721)
         );
  NAND2_X1 U7243 ( .A1(n6806), .A2(n6721), .ZN(n7119) );
  AOI22_X1 U7244 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n7119), .B1(n6830), 
        .B2(n7116), .ZN(n6722) );
  OAI211_X1 U7245 ( .C1(n7122), .C2(n6811), .A(n6723), .B(n6722), .ZN(U3076)
         );
  INV_X1 U7246 ( .A(n6724), .ZN(n6726) );
  NOR2_X2 U7247 ( .A1(n6738), .A2(n6780), .ZN(n7131) );
  INV_X1 U7248 ( .A(n7131), .ZN(n6859) );
  INV_X1 U7249 ( .A(n6727), .ZN(n6749) );
  NAND2_X1 U7250 ( .A1(n6749), .A2(n5132), .ZN(n6775) );
  OAI22_X1 U7251 ( .A1(n6825), .A2(n6728), .B1(n6751), .B2(n6775), .ZN(n7124)
         );
  NOR2_X1 U7252 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6729), .ZN(n7123)
         );
  AOI22_X1 U7253 ( .A1(n6828), .A2(n7124), .B1(n6827), .B2(n7123), .ZN(n6736)
         );
  OAI21_X1 U7254 ( .B1(n7118), .B2(n7131), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6732) );
  NAND2_X1 U7255 ( .A1(n6815), .A2(n6730), .ZN(n6731) );
  AOI21_X1 U7256 ( .B1(n6732), .B2(n6731), .A(n6755), .ZN(n6733) );
  NAND2_X1 U7257 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6775), .ZN(n6788) );
  OAI211_X1 U7258 ( .C1(n7123), .C2(n6734), .A(n6733), .B(n6788), .ZN(n7125)
         );
  AOI22_X1 U7259 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n7125), .B1(n6830), 
        .B2(n7118), .ZN(n6735) );
  OAI211_X1 U7260 ( .C1(n6764), .C2(n6859), .A(n6736), .B(n6735), .ZN(U3068)
         );
  NAND2_X1 U7261 ( .A1(n6793), .A2(n6753), .ZN(n6741) );
  NOR2_X1 U7262 ( .A1(n6794), .A2(n6741), .ZN(n7130) );
  AOI21_X1 U7263 ( .B1(n6796), .B2(n6737), .A(n7130), .ZN(n6743) );
  INV_X1 U7264 ( .A(n6738), .ZN(n6745) );
  AOI21_X1 U7265 ( .B1(n6745), .B2(STATEBS16_REG_SCAN_IN), .A(n6768), .ZN(
        n6742) );
  INV_X1 U7266 ( .A(n6742), .ZN(n6739) );
  OAI22_X1 U7267 ( .A1(n6797), .A2(n6741), .B1(n6743), .B2(n6739), .ZN(n6740)
         );
  AOI22_X1 U7268 ( .A1(n6827), .A2(n7130), .B1(n6830), .B2(n7131), .ZN(n6747)
         );
  AOI22_X1 U7269 ( .A1(n6743), .A2(n6742), .B1(n6768), .B2(n6741), .ZN(n6744)
         );
  NAND2_X1 U7270 ( .A1(n6806), .A2(n6744), .ZN(n7132) );
  NAND2_X1 U7271 ( .A1(n6745), .A2(n6780), .ZN(n7141) );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n7132), .B1(n6829), 
        .B2(n7129), .ZN(n6746) );
  OAI211_X1 U7273 ( .C1(n7135), .C2(n6811), .A(n6747), .B(n6746), .ZN(U3060)
         );
  NOR2_X1 U7274 ( .A1(n6750), .A2(n6749), .ZN(n6754) );
  INV_X1 U7275 ( .A(n6754), .ZN(n6822) );
  OAI22_X1 U7276 ( .A1(n6825), .A2(n6752), .B1(n6751), .B2(n6822), .ZN(n7137)
         );
  NAND2_X1 U7277 ( .A1(n6753), .A2(n6813), .ZN(n6756) );
  INV_X1 U7278 ( .A(n6756), .ZN(n7136) );
  AOI22_X1 U7279 ( .A1(n6828), .A2(n7137), .B1(n6827), .B2(n7136), .ZN(n6763)
         );
  NOR2_X1 U7280 ( .A1(n6754), .A2(n6797), .ZN(n6821) );
  AOI211_X1 U7281 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6756), .A(n6821), .B(
        n6755), .ZN(n6761) );
  INV_X1 U7282 ( .A(n6815), .ZN(n6758) );
  OAI211_X1 U7283 ( .C1(n6758), .C2(n6757), .A(n7061), .B(n7141), .ZN(n6760)
         );
  NAND3_X1 U7284 ( .A1(n6761), .A2(n6760), .A3(n6759), .ZN(n7138) );
  AOI22_X1 U7285 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n7138), .B1(n6830), 
        .B2(n7129), .ZN(n6762) );
  OAI211_X1 U7286 ( .C1(n6764), .C2(n7061), .A(n6763), .B(n6762), .ZN(U3052)
         );
  NOR2_X1 U7287 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6812) );
  INV_X1 U7288 ( .A(n6812), .ZN(n6765) );
  NOR2_X1 U7289 ( .A1(n6766), .A2(n6765), .ZN(n7143) );
  INV_X1 U7290 ( .A(n7154), .ZN(n7022) );
  AOI22_X1 U7291 ( .A1(n6827), .A2(n7143), .B1(n7022), .B2(n6829), .ZN(n6774)
         );
  AOI21_X1 U7292 ( .B1(n6796), .B2(n6784), .A(n7143), .ZN(n6772) );
  AOI21_X1 U7293 ( .B1(n6767), .B2(STATEBS16_REG_SCAN_IN), .A(n6768), .ZN(
        n6770) );
  NAND2_X1 U7294 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6812), .ZN(n6777) );
  AOI22_X1 U7295 ( .A1(n6772), .A2(n6770), .B1(n6768), .B2(n6777), .ZN(n6769)
         );
  NAND2_X1 U7296 ( .A1(n6806), .A2(n6769), .ZN(n7145) );
  INV_X1 U7297 ( .A(n6770), .ZN(n6771) );
  OAI22_X1 U7298 ( .A1(n6772), .A2(n6771), .B1(n6797), .B2(n6777), .ZN(n7144)
         );
  AOI22_X1 U7299 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n7145), .B1(n6828), 
        .B2(n7144), .ZN(n6773) );
  OAI211_X1 U7300 ( .C1(n6792), .C2(n7061), .A(n6774), .B(n6773), .ZN(U3044)
         );
  OAI22_X1 U7301 ( .A1(n6825), .A2(n6776), .B1(n6823), .B2(n6775), .ZN(n7150)
         );
  NOR2_X1 U7302 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6777), .ZN(n7149)
         );
  AOI22_X1 U7303 ( .A1(n6828), .A2(n7150), .B1(n6827), .B2(n7149), .ZN(n6791)
         );
  INV_X1 U7304 ( .A(n5127), .ZN(n6779) );
  NAND2_X1 U7305 ( .A1(n6779), .A2(n6778), .ZN(n6800) );
  NOR2_X2 U7306 ( .A1(n6800), .A2(n6780), .ZN(n7156) );
  INV_X1 U7307 ( .A(n7156), .ZN(n6782) );
  AOI21_X1 U7308 ( .B1(n6782), .B2(n7154), .A(n6781), .ZN(n6783) );
  AOI21_X1 U7309 ( .B1(n6785), .B2(n6784), .A(n6783), .ZN(n6786) );
  NOR2_X1 U7310 ( .A1(n6786), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6789) );
  INV_X1 U7311 ( .A(n6787), .ZN(n6819) );
  AOI22_X1 U7312 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n7151), .B1(n6829), 
        .B2(n7156), .ZN(n6790) );
  OAI211_X1 U7313 ( .C1(n6792), .C2(n7154), .A(n6791), .B(n6790), .ZN(U3036)
         );
  NAND2_X1 U7314 ( .A1(n6793), .A2(n6812), .ZN(n6801) );
  OAI21_X1 U7315 ( .B1(n6800), .B2(n6817), .A(n6808), .ZN(n6802) );
  NOR2_X1 U7316 ( .A1(n6794), .A2(n6801), .ZN(n7157) );
  AOI21_X1 U7317 ( .B1(n6796), .B2(n6795), .A(n7157), .ZN(n6803) );
  OAI22_X1 U7318 ( .A1(n6797), .A2(n6801), .B1(n6802), .B2(n6803), .ZN(n6798)
         );
  AOI22_X1 U7319 ( .A1(n6827), .A2(n7157), .B1(n7158), .B2(n6829), .ZN(n6810)
         );
  INV_X1 U7320 ( .A(n6801), .ZN(n6807) );
  INV_X1 U7321 ( .A(n6802), .ZN(n6804) );
  NAND2_X1 U7322 ( .A1(n6804), .A2(n6803), .ZN(n6805) );
  OAI211_X1 U7323 ( .C1(n6808), .C2(n6807), .A(n6806), .B(n6805), .ZN(n7159)
         );
  AOI22_X1 U7324 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n7159), .B1(n6830), 
        .B2(n7156), .ZN(n6809) );
  OAI211_X1 U7325 ( .C1(n7163), .C2(n6811), .A(n6810), .B(n6809), .ZN(U3028)
         );
  NAND2_X1 U7326 ( .A1(n6813), .A2(n6812), .ZN(n6826) );
  NAND2_X1 U7327 ( .A1(n6815), .A2(n6814), .ZN(n6816) );
  OAI221_X1 U7328 ( .B1(n6817), .B2(n7001), .C1(n6817), .C2(n7174), .A(n6816), 
        .ZN(n6818) );
  NAND2_X1 U7329 ( .A1(n6819), .A2(n6818), .ZN(n6820) );
  AOI211_X2 U7330 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6826), .A(n6821), .B(
        n6820), .ZN(n7168) );
  INV_X1 U7331 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6833) );
  OAI22_X1 U7332 ( .A1(n6825), .A2(n6824), .B1(n6823), .B2(n6822), .ZN(n7166)
         );
  INV_X1 U7333 ( .A(n6826), .ZN(n7164) );
  AOI22_X1 U7334 ( .A1(n6828), .A2(n7166), .B1(n6827), .B2(n7164), .ZN(n6832)
         );
  AOI22_X1 U7335 ( .A1(n6830), .A2(n7158), .B1(n6829), .B2(n7169), .ZN(n6831)
         );
  OAI211_X1 U7336 ( .C1(n7168), .C2(n6833), .A(n6832), .B(n6831), .ZN(U3020)
         );
  AOI22_X1 U7337 ( .A1(n6836), .A2(n6835), .B1(n6834), .B2(DATAI_24_), .ZN(
        n6840) );
  AOI22_X1 U7338 ( .A1(n6838), .A2(DATAI_8_), .B1(n6837), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U7339 ( .A1(n6840), .A2(n6839), .ZN(U2867) );
  AOI22_X1 U7340 ( .A1(n6874), .A2(n6995), .B1(n6873), .B2(n6994), .ZN(n6842)
         );
  INV_X1 U7341 ( .A(n6860), .ZN(n6875) );
  AOI22_X1 U7342 ( .A1(n6998), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n6997), 
        .B2(n6875), .ZN(n6841) );
  OAI211_X1 U7343 ( .C1(n6869), .C2(n7001), .A(n6842), .B(n6841), .ZN(U3141)
         );
  AOI22_X1 U7344 ( .A1(n6873), .A2(n7079), .B1(n6875), .B2(n7078), .ZN(n6844)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n7081), .B1(n6874), 
        .B2(n7080), .ZN(n6843) );
  OAI211_X1 U7346 ( .C1(n6869), .C2(n7084), .A(n6844), .B(n6843), .ZN(U3125)
         );
  AOI22_X1 U7347 ( .A1(n6874), .A2(n7086), .B1(n6873), .B2(n7085), .ZN(n6846)
         );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n7087), .B1(n6875), 
        .B2(n7091), .ZN(n6845) );
  OAI211_X1 U7349 ( .C1(n6869), .C2(n7090), .A(n6846), .B(n6845), .ZN(U3117)
         );
  AOI22_X1 U7350 ( .A1(n6873), .A2(n7092), .B1(n6876), .B2(n7091), .ZN(n6848)
         );
  AOI22_X1 U7351 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n7094), .B1(n6874), 
        .B2(n7093), .ZN(n6847) );
  OAI211_X1 U7352 ( .C1(n7102), .C2(n6860), .A(n6848), .B(n6847), .ZN(U3109)
         );
  AOI22_X1 U7353 ( .A1(n6873), .A2(n7097), .B1(n6875), .B2(n7105), .ZN(n6850)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n7099), .B1(n6874), 
        .B2(n7098), .ZN(n6849) );
  OAI211_X1 U7355 ( .C1(n7102), .C2(n6869), .A(n6850), .B(n6849), .ZN(U3101)
         );
  AOI22_X1 U7356 ( .A1(n6873), .A2(n7104), .B1(n6875), .B2(n7103), .ZN(n6852)
         );
  AOI22_X1 U7357 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n7106), .B1(n7105), 
        .B2(n6876), .ZN(n6851) );
  OAI211_X1 U7358 ( .C1(n7109), .C2(n6872), .A(n6852), .B(n6851), .ZN(U3093)
         );
  AOI22_X1 U7359 ( .A1(n6874), .A2(n7111), .B1(n6873), .B2(n7110), .ZN(n6854)
         );
  AOI22_X1 U7360 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n7112), .B1(n6875), 
        .B2(n7116), .ZN(n6853) );
  OAI211_X1 U7361 ( .C1(n6869), .C2(n7115), .A(n6854), .B(n6853), .ZN(U3085)
         );
  AOI22_X1 U7362 ( .A1(n6873), .A2(n7117), .B1(n6876), .B2(n7116), .ZN(n6856)
         );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n7119), .B1(n6875), 
        .B2(n7118), .ZN(n6855) );
  OAI211_X1 U7364 ( .C1(n7122), .C2(n6872), .A(n6856), .B(n6855), .ZN(U3077)
         );
  AOI22_X1 U7365 ( .A1(n6874), .A2(n7124), .B1(n6873), .B2(n7123), .ZN(n6858)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n7125), .B1(n6876), 
        .B2(n7118), .ZN(n6857) );
  OAI211_X1 U7367 ( .C1(n6860), .C2(n6859), .A(n6858), .B(n6857), .ZN(U3069)
         );
  AOI22_X1 U7368 ( .A1(n6873), .A2(n7130), .B1(n6875), .B2(n7129), .ZN(n6862)
         );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n7132), .B1(n6876), 
        .B2(n7131), .ZN(n6861) );
  OAI211_X1 U7370 ( .C1(n7135), .C2(n6872), .A(n6862), .B(n6861), .ZN(U3061)
         );
  AOI22_X1 U7371 ( .A1(n6874), .A2(n7137), .B1(n6873), .B2(n7136), .ZN(n6864)
         );
  AOI22_X1 U7372 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n7138), .B1(n6875), 
        .B2(n7142), .ZN(n6863) );
  OAI211_X1 U7373 ( .C1(n6869), .C2(n7141), .A(n6864), .B(n6863), .ZN(U3053)
         );
  AOI22_X1 U7374 ( .A1(n6873), .A2(n7143), .B1(n7022), .B2(n6875), .ZN(n6866)
         );
  AOI22_X1 U7375 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n7145), .B1(n6874), 
        .B2(n7144), .ZN(n6865) );
  OAI211_X1 U7376 ( .C1(n6869), .C2(n7061), .A(n6866), .B(n6865), .ZN(U3045)
         );
  AOI22_X1 U7377 ( .A1(n6874), .A2(n7150), .B1(n6873), .B2(n7149), .ZN(n6868)
         );
  AOI22_X1 U7378 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n7151), .B1(n7156), 
        .B2(n6875), .ZN(n6867) );
  OAI211_X1 U7379 ( .C1(n7154), .C2(n6869), .A(n6868), .B(n6867), .ZN(U3037)
         );
  AOI22_X1 U7380 ( .A1(n6873), .A2(n7157), .B1(n7158), .B2(n6875), .ZN(n6871)
         );
  AOI22_X1 U7381 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n7159), .B1(n7156), 
        .B2(n6876), .ZN(n6870) );
  OAI211_X1 U7382 ( .C1(n7163), .C2(n6872), .A(n6871), .B(n6870), .ZN(U3029)
         );
  AOI22_X1 U7383 ( .A1(n6874), .A2(n7166), .B1(n6873), .B2(n7164), .ZN(n6878)
         );
  AOI22_X1 U7384 ( .A1(n6876), .A2(n7158), .B1(n6875), .B2(n7169), .ZN(n6877)
         );
  OAI211_X1 U7385 ( .C1(n7168), .C2(n6879), .A(n6878), .B(n6877), .ZN(U3021)
         );
  AOI22_X1 U7386 ( .A1(n6912), .A2(n6995), .B1(n6911), .B2(n6994), .ZN(n6882)
         );
  AOI22_X1 U7387 ( .A1(n6998), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n6997), 
        .B2(n6913), .ZN(n6881) );
  OAI211_X1 U7388 ( .C1(n6907), .C2(n7001), .A(n6882), .B(n6881), .ZN(U3142)
         );
  AOI22_X1 U7389 ( .A1(n6911), .A2(n7079), .B1(n6913), .B2(n7078), .ZN(n6884)
         );
  AOI22_X1 U7390 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n7081), .B1(n6912), 
        .B2(n7080), .ZN(n6883) );
  OAI211_X1 U7391 ( .C1(n6907), .C2(n7084), .A(n6884), .B(n6883), .ZN(U3126)
         );
  AOI22_X1 U7392 ( .A1(n6912), .A2(n7086), .B1(n6911), .B2(n7085), .ZN(n6886)
         );
  AOI22_X1 U7393 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n7087), .B1(n6913), 
        .B2(n7091), .ZN(n6885) );
  OAI211_X1 U7394 ( .C1(n6907), .C2(n7090), .A(n6886), .B(n6885), .ZN(U3118)
         );
  AOI22_X1 U7395 ( .A1(n6911), .A2(n7092), .B1(n6913), .B2(n7043), .ZN(n6888)
         );
  AOI22_X1 U7396 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n7094), .B1(n6912), 
        .B2(n7093), .ZN(n6887) );
  OAI211_X1 U7397 ( .C1(n6907), .C2(n7046), .A(n6888), .B(n6887), .ZN(U3110)
         );
  AOI22_X1 U7398 ( .A1(n6911), .A2(n7097), .B1(n6913), .B2(n7105), .ZN(n6890)
         );
  AOI22_X1 U7399 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n7099), .B1(n6912), 
        .B2(n7098), .ZN(n6889) );
  OAI211_X1 U7400 ( .C1(n7102), .C2(n6907), .A(n6890), .B(n6889), .ZN(U3102)
         );
  AOI22_X1 U7401 ( .A1(n6911), .A2(n7104), .B1(n6913), .B2(n7103), .ZN(n6892)
         );
  AOI22_X1 U7402 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n7106), .B1(n7105), 
        .B2(n6914), .ZN(n6891) );
  OAI211_X1 U7403 ( .C1(n7109), .C2(n6910), .A(n6892), .B(n6891), .ZN(U3094)
         );
  AOI22_X1 U7404 ( .A1(n6912), .A2(n7111), .B1(n6911), .B2(n7110), .ZN(n6894)
         );
  AOI22_X1 U7405 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n7112), .B1(n6913), 
        .B2(n7116), .ZN(n6893) );
  OAI211_X1 U7406 ( .C1(n6907), .C2(n7115), .A(n6894), .B(n6893), .ZN(U3086)
         );
  AOI22_X1 U7407 ( .A1(n6911), .A2(n7117), .B1(n6913), .B2(n7118), .ZN(n6896)
         );
  AOI22_X1 U7408 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n7119), .B1(n6914), 
        .B2(n7116), .ZN(n6895) );
  OAI211_X1 U7409 ( .C1(n7122), .C2(n6910), .A(n6896), .B(n6895), .ZN(U3078)
         );
  AOI22_X1 U7410 ( .A1(n6912), .A2(n7124), .B1(n6911), .B2(n7123), .ZN(n6898)
         );
  AOI22_X1 U7411 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n7125), .B1(n6913), 
        .B2(n7131), .ZN(n6897) );
  OAI211_X1 U7412 ( .C1(n6907), .C2(n7128), .A(n6898), .B(n6897), .ZN(U3070)
         );
  AOI22_X1 U7413 ( .A1(n6911), .A2(n7130), .B1(n6914), .B2(n7131), .ZN(n6900)
         );
  AOI22_X1 U7414 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n7132), .B1(n6913), 
        .B2(n7129), .ZN(n6899) );
  OAI211_X1 U7415 ( .C1(n7135), .C2(n6910), .A(n6900), .B(n6899), .ZN(U3062)
         );
  AOI22_X1 U7416 ( .A1(n6912), .A2(n7137), .B1(n6911), .B2(n7136), .ZN(n6902)
         );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(n7138), .B1(n6913), 
        .B2(n7142), .ZN(n6901) );
  OAI211_X1 U7418 ( .C1(n6907), .C2(n7141), .A(n6902), .B(n6901), .ZN(U3054)
         );
  AOI22_X1 U7419 ( .A1(n6911), .A2(n7143), .B1(n7022), .B2(n6913), .ZN(n6904)
         );
  AOI22_X1 U7420 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n7145), .B1(n6912), 
        .B2(n7144), .ZN(n6903) );
  OAI211_X1 U7421 ( .C1(n6907), .C2(n7061), .A(n6904), .B(n6903), .ZN(U3046)
         );
  AOI22_X1 U7422 ( .A1(n6912), .A2(n7150), .B1(n6911), .B2(n7149), .ZN(n6906)
         );
  AOI22_X1 U7423 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n7151), .B1(n7156), 
        .B2(n6913), .ZN(n6905) );
  OAI211_X1 U7424 ( .C1(n7154), .C2(n6907), .A(n6906), .B(n6905), .ZN(U3038)
         );
  AOI22_X1 U7425 ( .A1(n6911), .A2(n7157), .B1(n7156), .B2(n6914), .ZN(n6909)
         );
  AOI22_X1 U7426 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n7159), .B1(n6913), 
        .B2(n7158), .ZN(n6908) );
  OAI211_X1 U7427 ( .C1(n7163), .C2(n6910), .A(n6909), .B(n6908), .ZN(U3030)
         );
  INV_X1 U7428 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U7429 ( .A1(n6912), .A2(n7166), .B1(n6911), .B2(n7164), .ZN(n6916)
         );
  AOI22_X1 U7430 ( .A1(n6914), .A2(n7158), .B1(n6913), .B2(n7169), .ZN(n6915)
         );
  OAI211_X1 U7431 ( .C1(n7168), .C2(n6917), .A(n6916), .B(n6915), .ZN(U3022)
         );
  AOI22_X1 U7432 ( .A1(n6950), .A2(n6995), .B1(n6949), .B2(n6994), .ZN(n6920)
         );
  INV_X1 U7433 ( .A(n6918), .ZN(n6951) );
  AOI22_X1 U7434 ( .A1(n6998), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n6997), 
        .B2(n6951), .ZN(n6919) );
  OAI211_X1 U7435 ( .C1(n6945), .C2(n7001), .A(n6920), .B(n6919), .ZN(U3143)
         );
  AOI22_X1 U7436 ( .A1(n6949), .A2(n7079), .B1(n6951), .B2(n7078), .ZN(n6922)
         );
  AOI22_X1 U7437 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n7081), .B1(n6950), 
        .B2(n7080), .ZN(n6921) );
  OAI211_X1 U7438 ( .C1(n6945), .C2(n7084), .A(n6922), .B(n6921), .ZN(U3127)
         );
  AOI22_X1 U7439 ( .A1(n6950), .A2(n7086), .B1(n6949), .B2(n7085), .ZN(n6924)
         );
  AOI22_X1 U7440 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n7087), .B1(n6951), 
        .B2(n7091), .ZN(n6923) );
  OAI211_X1 U7441 ( .C1(n6945), .C2(n7090), .A(n6924), .B(n6923), .ZN(U3119)
         );
  AOI22_X1 U7442 ( .A1(n6949), .A2(n7092), .B1(n6951), .B2(n7043), .ZN(n6926)
         );
  AOI22_X1 U7443 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n7094), .B1(n6950), 
        .B2(n7093), .ZN(n6925) );
  OAI211_X1 U7444 ( .C1(n6945), .C2(n7046), .A(n6926), .B(n6925), .ZN(U3111)
         );
  AOI22_X1 U7445 ( .A1(n6949), .A2(n7097), .B1(n6951), .B2(n7105), .ZN(n6928)
         );
  AOI22_X1 U7446 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n7099), .B1(n6950), 
        .B2(n7098), .ZN(n6927) );
  OAI211_X1 U7447 ( .C1(n7102), .C2(n6945), .A(n6928), .B(n6927), .ZN(U3103)
         );
  AOI22_X1 U7448 ( .A1(n6949), .A2(n7104), .B1(n6951), .B2(n7103), .ZN(n6930)
         );
  AOI22_X1 U7449 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n7106), .B1(n7105), 
        .B2(n6952), .ZN(n6929) );
  OAI211_X1 U7450 ( .C1(n7109), .C2(n6948), .A(n6930), .B(n6929), .ZN(U3095)
         );
  AOI22_X1 U7451 ( .A1(n6950), .A2(n7111), .B1(n6949), .B2(n7110), .ZN(n6932)
         );
  AOI22_X1 U7452 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n7112), .B1(n6951), 
        .B2(n7116), .ZN(n6931) );
  OAI211_X1 U7453 ( .C1(n6945), .C2(n7115), .A(n6932), .B(n6931), .ZN(U3087)
         );
  AOI22_X1 U7454 ( .A1(n6949), .A2(n7117), .B1(n6951), .B2(n7118), .ZN(n6934)
         );
  AOI22_X1 U7455 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n7119), .B1(n6952), 
        .B2(n7116), .ZN(n6933) );
  OAI211_X1 U7456 ( .C1(n7122), .C2(n6948), .A(n6934), .B(n6933), .ZN(U3079)
         );
  AOI22_X1 U7457 ( .A1(n6950), .A2(n7124), .B1(n6949), .B2(n7123), .ZN(n6936)
         );
  AOI22_X1 U7458 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n7125), .B1(n6951), 
        .B2(n7131), .ZN(n6935) );
  OAI211_X1 U7459 ( .C1(n6945), .C2(n7128), .A(n6936), .B(n6935), .ZN(U3071)
         );
  AOI22_X1 U7460 ( .A1(n6949), .A2(n7130), .B1(n6952), .B2(n7131), .ZN(n6938)
         );
  AOI22_X1 U7461 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n7132), .B1(n6951), 
        .B2(n7129), .ZN(n6937) );
  OAI211_X1 U7462 ( .C1(n7135), .C2(n6948), .A(n6938), .B(n6937), .ZN(U3063)
         );
  AOI22_X1 U7463 ( .A1(n6950), .A2(n7137), .B1(n6949), .B2(n7136), .ZN(n6940)
         );
  AOI22_X1 U7464 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(n7138), .B1(n6951), 
        .B2(n7142), .ZN(n6939) );
  OAI211_X1 U7465 ( .C1(n6945), .C2(n7141), .A(n6940), .B(n6939), .ZN(U3055)
         );
  AOI22_X1 U7466 ( .A1(n6949), .A2(n7143), .B1(n7022), .B2(n6951), .ZN(n6942)
         );
  AOI22_X1 U7467 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n7145), .B1(n6950), 
        .B2(n7144), .ZN(n6941) );
  OAI211_X1 U7468 ( .C1(n6945), .C2(n7061), .A(n6942), .B(n6941), .ZN(U3047)
         );
  AOI22_X1 U7469 ( .A1(n6950), .A2(n7150), .B1(n6949), .B2(n7149), .ZN(n6944)
         );
  AOI22_X1 U7470 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n7151), .B1(n7156), 
        .B2(n6951), .ZN(n6943) );
  OAI211_X1 U7471 ( .C1(n7154), .C2(n6945), .A(n6944), .B(n6943), .ZN(U3039)
         );
  AOI22_X1 U7472 ( .A1(n6949), .A2(n7157), .B1(n7158), .B2(n6951), .ZN(n6947)
         );
  AOI22_X1 U7473 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n7159), .B1(n7156), 
        .B2(n6952), .ZN(n6946) );
  OAI211_X1 U7474 ( .C1(n7163), .C2(n6948), .A(n6947), .B(n6946), .ZN(U3031)
         );
  AOI22_X1 U7475 ( .A1(n6950), .A2(n7166), .B1(n6949), .B2(n7164), .ZN(n6954)
         );
  AOI22_X1 U7476 ( .A1(n6952), .A2(n7158), .B1(n6951), .B2(n7169), .ZN(n6953)
         );
  OAI211_X1 U7477 ( .C1(n7168), .C2(n6955), .A(n6954), .B(n6953), .ZN(U3023)
         );
  AOI22_X1 U7478 ( .A1(n6988), .A2(n6995), .B1(n6987), .B2(n6994), .ZN(n6957)
         );
  INV_X1 U7479 ( .A(n6980), .ZN(n6989) );
  AOI22_X1 U7480 ( .A1(n6998), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n6997), 
        .B2(n6989), .ZN(n6956) );
  OAI211_X1 U7481 ( .C1(n6983), .C2(n7001), .A(n6957), .B(n6956), .ZN(U3144)
         );
  AOI22_X1 U7482 ( .A1(n6987), .A2(n7079), .B1(n7038), .B2(n6990), .ZN(n6959)
         );
  AOI22_X1 U7483 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n7081), .B1(n6988), 
        .B2(n7080), .ZN(n6958) );
  OAI211_X1 U7484 ( .C1(n6980), .C2(n7090), .A(n6959), .B(n6958), .ZN(U3128)
         );
  AOI22_X1 U7485 ( .A1(n6988), .A2(n7086), .B1(n6987), .B2(n7085), .ZN(n6961)
         );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n7087), .B1(n6989), 
        .B2(n7091), .ZN(n6960) );
  OAI211_X1 U7487 ( .C1(n6983), .C2(n7090), .A(n6961), .B(n6960), .ZN(U3120)
         );
  AOI22_X1 U7488 ( .A1(n6987), .A2(n7092), .B1(n6989), .B2(n7043), .ZN(n6963)
         );
  AOI22_X1 U7489 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n7094), .B1(n6988), 
        .B2(n7093), .ZN(n6962) );
  OAI211_X1 U7490 ( .C1(n6983), .C2(n7046), .A(n6963), .B(n6962), .ZN(U3112)
         );
  AOI22_X1 U7491 ( .A1(n6987), .A2(n7097), .B1(n6989), .B2(n7105), .ZN(n6965)
         );
  AOI22_X1 U7492 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n7099), .B1(n6988), 
        .B2(n7098), .ZN(n6964) );
  OAI211_X1 U7493 ( .C1(n7102), .C2(n6983), .A(n6965), .B(n6964), .ZN(U3104)
         );
  AOI22_X1 U7494 ( .A1(n6987), .A2(n7104), .B1(n6990), .B2(n7105), .ZN(n6967)
         );
  AOI22_X1 U7495 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n7106), .B1(n6989), 
        .B2(n7103), .ZN(n6966) );
  OAI211_X1 U7496 ( .C1(n7109), .C2(n6986), .A(n6967), .B(n6966), .ZN(U3096)
         );
  AOI22_X1 U7497 ( .A1(n6988), .A2(n7111), .B1(n6987), .B2(n7110), .ZN(n6969)
         );
  AOI22_X1 U7498 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n7112), .B1(n6989), 
        .B2(n7116), .ZN(n6968) );
  OAI211_X1 U7499 ( .C1(n6983), .C2(n7115), .A(n6969), .B(n6968), .ZN(U3088)
         );
  AOI22_X1 U7500 ( .A1(n6987), .A2(n7117), .B1(n6989), .B2(n7118), .ZN(n6971)
         );
  AOI22_X1 U7501 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n7119), .B1(n6990), 
        .B2(n7116), .ZN(n6970) );
  OAI211_X1 U7502 ( .C1(n7122), .C2(n6986), .A(n6971), .B(n6970), .ZN(U3080)
         );
  AOI22_X1 U7503 ( .A1(n6988), .A2(n7124), .B1(n6987), .B2(n7123), .ZN(n6973)
         );
  AOI22_X1 U7504 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n7125), .B1(n6989), 
        .B2(n7131), .ZN(n6972) );
  OAI211_X1 U7505 ( .C1(n6983), .C2(n7128), .A(n6973), .B(n6972), .ZN(U3072)
         );
  AOI22_X1 U7506 ( .A1(n6987), .A2(n7130), .B1(n6989), .B2(n7129), .ZN(n6975)
         );
  AOI22_X1 U7507 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n7132), .B1(n6990), 
        .B2(n7131), .ZN(n6974) );
  OAI211_X1 U7508 ( .C1(n7135), .C2(n6986), .A(n6975), .B(n6974), .ZN(U3064)
         );
  AOI22_X1 U7509 ( .A1(n6988), .A2(n7137), .B1(n6987), .B2(n7136), .ZN(n6977)
         );
  AOI22_X1 U7510 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n7138), .B1(n6990), 
        .B2(n7129), .ZN(n6976) );
  OAI211_X1 U7511 ( .C1(n6980), .C2(n7061), .A(n6977), .B(n6976), .ZN(U3056)
         );
  AOI22_X1 U7512 ( .A1(n6987), .A2(n7143), .B1(n7142), .B2(n6990), .ZN(n6979)
         );
  AOI22_X1 U7513 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n7145), .B1(n6988), 
        .B2(n7144), .ZN(n6978) );
  OAI211_X1 U7514 ( .C1(n7154), .C2(n6980), .A(n6979), .B(n6978), .ZN(U3048)
         );
  AOI22_X1 U7515 ( .A1(n6988), .A2(n7150), .B1(n6987), .B2(n7149), .ZN(n6982)
         );
  AOI22_X1 U7516 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n7151), .B1(n7156), 
        .B2(n6989), .ZN(n6981) );
  OAI211_X1 U7517 ( .C1(n7154), .C2(n6983), .A(n6982), .B(n6981), .ZN(U3040)
         );
  AOI22_X1 U7518 ( .A1(n6987), .A2(n7157), .B1(n7156), .B2(n6990), .ZN(n6985)
         );
  AOI22_X1 U7519 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n7159), .B1(n6989), 
        .B2(n7158), .ZN(n6984) );
  OAI211_X1 U7520 ( .C1(n7163), .C2(n6986), .A(n6985), .B(n6984), .ZN(U3032)
         );
  INV_X1 U7521 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6993) );
  AOI22_X1 U7522 ( .A1(n6988), .A2(n7166), .B1(n6987), .B2(n7164), .ZN(n6992)
         );
  AOI22_X1 U7523 ( .A1(n6990), .A2(n7158), .B1(n6989), .B2(n7169), .ZN(n6991)
         );
  OAI211_X1 U7524 ( .C1(n7168), .C2(n6993), .A(n6992), .B(n6991), .ZN(U3024)
         );
  AOI22_X1 U7525 ( .A1(n7032), .A2(n6995), .B1(n7031), .B2(n6994), .ZN(n7000)
         );
  INV_X1 U7526 ( .A(n6996), .ZN(n7033) );
  AOI22_X1 U7527 ( .A1(n6998), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n6997), 
        .B2(n7033), .ZN(n6999) );
  OAI211_X1 U7528 ( .C1(n7027), .C2(n7001), .A(n7000), .B(n6999), .ZN(U3145)
         );
  AOI22_X1 U7529 ( .A1(n7031), .A2(n7079), .B1(n7033), .B2(n7078), .ZN(n7003)
         );
  AOI22_X1 U7530 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n7081), .B1(n7032), 
        .B2(n7080), .ZN(n7002) );
  OAI211_X1 U7531 ( .C1(n7027), .C2(n7084), .A(n7003), .B(n7002), .ZN(U3129)
         );
  AOI22_X1 U7532 ( .A1(n7032), .A2(n7086), .B1(n7031), .B2(n7085), .ZN(n7005)
         );
  AOI22_X1 U7533 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n7087), .B1(n7033), 
        .B2(n7091), .ZN(n7004) );
  OAI211_X1 U7534 ( .C1(n7027), .C2(n7090), .A(n7005), .B(n7004), .ZN(U3121)
         );
  AOI22_X1 U7535 ( .A1(n7031), .A2(n7092), .B1(n7033), .B2(n7043), .ZN(n7007)
         );
  AOI22_X1 U7536 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n7094), .B1(n7032), 
        .B2(n7093), .ZN(n7006) );
  OAI211_X1 U7537 ( .C1(n7027), .C2(n7046), .A(n7007), .B(n7006), .ZN(U3113)
         );
  AOI22_X1 U7538 ( .A1(n7031), .A2(n7097), .B1(n7033), .B2(n7105), .ZN(n7009)
         );
  AOI22_X1 U7539 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n7099), .B1(n7032), 
        .B2(n7098), .ZN(n7008) );
  OAI211_X1 U7540 ( .C1(n7102), .C2(n7027), .A(n7009), .B(n7008), .ZN(U3105)
         );
  AOI22_X1 U7541 ( .A1(n7031), .A2(n7104), .B1(n7034), .B2(n7105), .ZN(n7011)
         );
  AOI22_X1 U7542 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n7106), .B1(n7033), 
        .B2(n7103), .ZN(n7010) );
  OAI211_X1 U7543 ( .C1(n7109), .C2(n7030), .A(n7011), .B(n7010), .ZN(U3097)
         );
  AOI22_X1 U7544 ( .A1(n7032), .A2(n7111), .B1(n7031), .B2(n7110), .ZN(n7013)
         );
  AOI22_X1 U7545 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n7112), .B1(n7033), 
        .B2(n7116), .ZN(n7012) );
  OAI211_X1 U7546 ( .C1(n7027), .C2(n7115), .A(n7013), .B(n7012), .ZN(U3089)
         );
  AOI22_X1 U7547 ( .A1(n7031), .A2(n7117), .B1(n7034), .B2(n7116), .ZN(n7015)
         );
  AOI22_X1 U7548 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n7119), .B1(n7033), 
        .B2(n7118), .ZN(n7014) );
  OAI211_X1 U7549 ( .C1(n7122), .C2(n7030), .A(n7015), .B(n7014), .ZN(U3081)
         );
  AOI22_X1 U7550 ( .A1(n7032), .A2(n7124), .B1(n7031), .B2(n7123), .ZN(n7017)
         );
  AOI22_X1 U7551 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n7125), .B1(n7033), 
        .B2(n7131), .ZN(n7016) );
  OAI211_X1 U7552 ( .C1(n7027), .C2(n7128), .A(n7017), .B(n7016), .ZN(U3073)
         );
  AOI22_X1 U7553 ( .A1(n7031), .A2(n7130), .B1(n7034), .B2(n7131), .ZN(n7019)
         );
  AOI22_X1 U7554 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n7132), .B1(n7033), 
        .B2(n7129), .ZN(n7018) );
  OAI211_X1 U7555 ( .C1(n7135), .C2(n7030), .A(n7019), .B(n7018), .ZN(U3065)
         );
  AOI22_X1 U7556 ( .A1(n7032), .A2(n7137), .B1(n7031), .B2(n7136), .ZN(n7021)
         );
  AOI22_X1 U7557 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n7138), .B1(n7033), 
        .B2(n7142), .ZN(n7020) );
  OAI211_X1 U7558 ( .C1(n7027), .C2(n7141), .A(n7021), .B(n7020), .ZN(U3057)
         );
  AOI22_X1 U7559 ( .A1(n7031), .A2(n7143), .B1(n7022), .B2(n7033), .ZN(n7024)
         );
  AOI22_X1 U7560 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n7145), .B1(n7032), 
        .B2(n7144), .ZN(n7023) );
  OAI211_X1 U7561 ( .C1(n7027), .C2(n7061), .A(n7024), .B(n7023), .ZN(U3049)
         );
  AOI22_X1 U7562 ( .A1(n7032), .A2(n7150), .B1(n7031), .B2(n7149), .ZN(n7026)
         );
  AOI22_X1 U7563 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n7151), .B1(n7156), 
        .B2(n7033), .ZN(n7025) );
  OAI211_X1 U7564 ( .C1(n7154), .C2(n7027), .A(n7026), .B(n7025), .ZN(U3041)
         );
  AOI22_X1 U7565 ( .A1(n7031), .A2(n7157), .B1(n7158), .B2(n7033), .ZN(n7029)
         );
  AOI22_X1 U7566 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n7159), .B1(n7156), 
        .B2(n7034), .ZN(n7028) );
  OAI211_X1 U7567 ( .C1(n7163), .C2(n7030), .A(n7029), .B(n7028), .ZN(U3033)
         );
  AOI22_X1 U7568 ( .A1(n7032), .A2(n7166), .B1(n7031), .B2(n7164), .ZN(n7036)
         );
  AOI22_X1 U7569 ( .A1(n7034), .A2(n7158), .B1(n7033), .B2(n7169), .ZN(n7035)
         );
  OAI211_X1 U7570 ( .C1(n7168), .C2(n7037), .A(n7036), .B(n7035), .ZN(U3025)
         );
  AOI22_X1 U7571 ( .A1(n7071), .A2(n7079), .B1(n7038), .B2(n7074), .ZN(n7040)
         );
  AOI22_X1 U7572 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n7081), .B1(n7072), 
        .B2(n7080), .ZN(n7039) );
  OAI211_X1 U7573 ( .C1(n7064), .C2(n7090), .A(n7040), .B(n7039), .ZN(U3130)
         );
  AOI22_X1 U7574 ( .A1(n7072), .A2(n7086), .B1(n7071), .B2(n7085), .ZN(n7042)
         );
  AOI22_X1 U7575 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n7087), .B1(n7073), 
        .B2(n7091), .ZN(n7041) );
  OAI211_X1 U7576 ( .C1(n7067), .C2(n7090), .A(n7042), .B(n7041), .ZN(U3122)
         );
  AOI22_X1 U7577 ( .A1(n7071), .A2(n7092), .B1(n7073), .B2(n7043), .ZN(n7045)
         );
  AOI22_X1 U7578 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n7094), .B1(n7072), 
        .B2(n7093), .ZN(n7044) );
  OAI211_X1 U7579 ( .C1(n7067), .C2(n7046), .A(n7045), .B(n7044), .ZN(U3114)
         );
  AOI22_X1 U7580 ( .A1(n7071), .A2(n7097), .B1(n7073), .B2(n7105), .ZN(n7048)
         );
  AOI22_X1 U7581 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n7099), .B1(n7072), 
        .B2(n7098), .ZN(n7047) );
  OAI211_X1 U7582 ( .C1(n7102), .C2(n7067), .A(n7048), .B(n7047), .ZN(U3106)
         );
  AOI22_X1 U7583 ( .A1(n7071), .A2(n7104), .B1(n7074), .B2(n7105), .ZN(n7050)
         );
  AOI22_X1 U7584 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n7106), .B1(n7073), 
        .B2(n7103), .ZN(n7049) );
  OAI211_X1 U7585 ( .C1(n7109), .C2(n7070), .A(n7050), .B(n7049), .ZN(U3098)
         );
  AOI22_X1 U7586 ( .A1(n7072), .A2(n7111), .B1(n7071), .B2(n7110), .ZN(n7052)
         );
  AOI22_X1 U7587 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n7112), .B1(n7073), 
        .B2(n7116), .ZN(n7051) );
  OAI211_X1 U7588 ( .C1(n7067), .C2(n7115), .A(n7052), .B(n7051), .ZN(U3090)
         );
  AOI22_X1 U7589 ( .A1(n7071), .A2(n7117), .B1(n7073), .B2(n7118), .ZN(n7054)
         );
  AOI22_X1 U7590 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n7119), .B1(n7074), 
        .B2(n7116), .ZN(n7053) );
  OAI211_X1 U7591 ( .C1(n7122), .C2(n7070), .A(n7054), .B(n7053), .ZN(U3082)
         );
  AOI22_X1 U7592 ( .A1(n7072), .A2(n7124), .B1(n7071), .B2(n7123), .ZN(n7056)
         );
  AOI22_X1 U7593 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n7125), .B1(n7073), 
        .B2(n7131), .ZN(n7055) );
  OAI211_X1 U7594 ( .C1(n7067), .C2(n7128), .A(n7056), .B(n7055), .ZN(U3074)
         );
  AOI22_X1 U7595 ( .A1(n7071), .A2(n7130), .B1(n7073), .B2(n7129), .ZN(n7058)
         );
  AOI22_X1 U7596 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n7132), .B1(n7074), 
        .B2(n7131), .ZN(n7057) );
  OAI211_X1 U7597 ( .C1(n7135), .C2(n7070), .A(n7058), .B(n7057), .ZN(U3066)
         );
  AOI22_X1 U7598 ( .A1(n7072), .A2(n7137), .B1(n7071), .B2(n7136), .ZN(n7060)
         );
  AOI22_X1 U7599 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(n7138), .B1(n7074), 
        .B2(n7129), .ZN(n7059) );
  OAI211_X1 U7600 ( .C1(n7064), .C2(n7061), .A(n7060), .B(n7059), .ZN(U3058)
         );
  AOI22_X1 U7601 ( .A1(n7071), .A2(n7143), .B1(n7142), .B2(n7074), .ZN(n7063)
         );
  AOI22_X1 U7602 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n7145), .B1(n7072), 
        .B2(n7144), .ZN(n7062) );
  OAI211_X1 U7603 ( .C1(n7154), .C2(n7064), .A(n7063), .B(n7062), .ZN(U3050)
         );
  AOI22_X1 U7604 ( .A1(n7072), .A2(n7150), .B1(n7071), .B2(n7149), .ZN(n7066)
         );
  AOI22_X1 U7605 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n7151), .B1(n7156), 
        .B2(n7073), .ZN(n7065) );
  OAI211_X1 U7606 ( .C1(n7154), .C2(n7067), .A(n7066), .B(n7065), .ZN(U3042)
         );
  AOI22_X1 U7607 ( .A1(n7071), .A2(n7157), .B1(n7158), .B2(n7073), .ZN(n7069)
         );
  AOI22_X1 U7608 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n7159), .B1(n7156), 
        .B2(n7074), .ZN(n7068) );
  OAI211_X1 U7609 ( .C1(n7163), .C2(n7070), .A(n7069), .B(n7068), .ZN(U3034)
         );
  INV_X1 U7610 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n7077) );
  AOI22_X1 U7611 ( .A1(n7072), .A2(n7166), .B1(n7071), .B2(n7164), .ZN(n7076)
         );
  AOI22_X1 U7612 ( .A1(n7074), .A2(n7158), .B1(n7073), .B2(n7169), .ZN(n7075)
         );
  OAI211_X1 U7613 ( .C1(n7168), .C2(n7077), .A(n7076), .B(n7075), .ZN(U3026)
         );
  AOI22_X1 U7614 ( .A1(n7165), .A2(n7079), .B1(n7170), .B2(n7078), .ZN(n7083)
         );
  AOI22_X1 U7615 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n7081), .B1(n7167), 
        .B2(n7080), .ZN(n7082) );
  OAI211_X1 U7616 ( .C1(n7175), .C2(n7084), .A(n7083), .B(n7082), .ZN(U3131)
         );
  AOI22_X1 U7617 ( .A1(n7167), .A2(n7086), .B1(n7165), .B2(n7085), .ZN(n7089)
         );
  AOI22_X1 U7618 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n7087), .B1(n7170), 
        .B2(n7091), .ZN(n7088) );
  OAI211_X1 U7619 ( .C1(n7175), .C2(n7090), .A(n7089), .B(n7088), .ZN(U3123)
         );
  AOI22_X1 U7620 ( .A1(n7165), .A2(n7092), .B1(n7155), .B2(n7091), .ZN(n7096)
         );
  AOI22_X1 U7621 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n7094), .B1(n7167), 
        .B2(n7093), .ZN(n7095) );
  OAI211_X1 U7622 ( .C1(n7102), .C2(n7148), .A(n7096), .B(n7095), .ZN(U3115)
         );
  AOI22_X1 U7623 ( .A1(n7165), .A2(n7097), .B1(n7170), .B2(n7105), .ZN(n7101)
         );
  AOI22_X1 U7624 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n7099), .B1(n7167), 
        .B2(n7098), .ZN(n7100) );
  OAI211_X1 U7625 ( .C1(n7102), .C2(n7175), .A(n7101), .B(n7100), .ZN(U3107)
         );
  AOI22_X1 U7626 ( .A1(n7165), .A2(n7104), .B1(n7170), .B2(n7103), .ZN(n7108)
         );
  AOI22_X1 U7627 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n7106), .B1(n7105), 
        .B2(n7155), .ZN(n7107) );
  OAI211_X1 U7628 ( .C1(n7109), .C2(n7162), .A(n7108), .B(n7107), .ZN(U3099)
         );
  AOI22_X1 U7629 ( .A1(n7167), .A2(n7111), .B1(n7165), .B2(n7110), .ZN(n7114)
         );
  AOI22_X1 U7630 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n7112), .B1(n7170), 
        .B2(n7116), .ZN(n7113) );
  OAI211_X1 U7631 ( .C1(n7175), .C2(n7115), .A(n7114), .B(n7113), .ZN(U3091)
         );
  AOI22_X1 U7632 ( .A1(n7165), .A2(n7117), .B1(n7155), .B2(n7116), .ZN(n7121)
         );
  AOI22_X1 U7633 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n7119), .B1(n7170), 
        .B2(n7118), .ZN(n7120) );
  OAI211_X1 U7634 ( .C1(n7122), .C2(n7162), .A(n7121), .B(n7120), .ZN(U3083)
         );
  AOI22_X1 U7635 ( .A1(n7167), .A2(n7124), .B1(n7165), .B2(n7123), .ZN(n7127)
         );
  AOI22_X1 U7636 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n7125), .B1(n7170), 
        .B2(n7131), .ZN(n7126) );
  OAI211_X1 U7637 ( .C1(n7175), .C2(n7128), .A(n7127), .B(n7126), .ZN(U3075)
         );
  AOI22_X1 U7638 ( .A1(n7165), .A2(n7130), .B1(n7170), .B2(n7129), .ZN(n7134)
         );
  AOI22_X1 U7639 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n7132), .B1(n7155), 
        .B2(n7131), .ZN(n7133) );
  OAI211_X1 U7640 ( .C1(n7135), .C2(n7162), .A(n7134), .B(n7133), .ZN(U3067)
         );
  AOI22_X1 U7641 ( .A1(n7167), .A2(n7137), .B1(n7165), .B2(n7136), .ZN(n7140)
         );
  AOI22_X1 U7642 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n7138), .B1(n7170), 
        .B2(n7142), .ZN(n7139) );
  OAI211_X1 U7643 ( .C1(n7175), .C2(n7141), .A(n7140), .B(n7139), .ZN(U3059)
         );
  AOI22_X1 U7644 ( .A1(n7165), .A2(n7143), .B1(n7142), .B2(n7155), .ZN(n7147)
         );
  AOI22_X1 U7645 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n7145), .B1(n7167), 
        .B2(n7144), .ZN(n7146) );
  OAI211_X1 U7646 ( .C1(n7154), .C2(n7148), .A(n7147), .B(n7146), .ZN(U3051)
         );
  AOI22_X1 U7647 ( .A1(n7167), .A2(n7150), .B1(n7165), .B2(n7149), .ZN(n7153)
         );
  AOI22_X1 U7648 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n7151), .B1(n7156), 
        .B2(n7170), .ZN(n7152) );
  OAI211_X1 U7649 ( .C1(n7154), .C2(n7175), .A(n7153), .B(n7152), .ZN(U3043)
         );
  AOI22_X1 U7650 ( .A1(n7165), .A2(n7157), .B1(n7156), .B2(n7155), .ZN(n7161)
         );
  AOI22_X1 U7651 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n7159), .B1(n7170), 
        .B2(n7158), .ZN(n7160) );
  OAI211_X1 U7652 ( .C1(n7163), .C2(n7162), .A(n7161), .B(n7160), .ZN(U3035)
         );
  AOI22_X1 U7653 ( .A1(n7167), .A2(n7166), .B1(n7165), .B2(n7164), .ZN(n7173)
         );
  INV_X1 U7654 ( .A(n7168), .ZN(n7171) );
  AOI22_X1 U7655 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n7171), .B1(n7170), 
        .B2(n7169), .ZN(n7172) );
  OAI211_X1 U7656 ( .C1(n7175), .C2(n7174), .A(n7173), .B(n7172), .ZN(U3027)
         );
  CLKBUF_X1 U3503 ( .A(n4878), .Z(n3455) );
  CLKBUF_X1 U3744 ( .A(n3711), .Z(n4201) );
endmodule

