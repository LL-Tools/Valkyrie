

module b17_C_SARLock_k_128_7 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9747, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9793, n9794, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308;

  INV_X1 U11192 ( .A(n15205), .ZN(n9769) );
  NAND2_X1 U11193 ( .A1(n10191), .A2(n10189), .ZN(n15446) );
  AND2_X1 U11194 ( .A1(n9901), .A2(n9953), .ZN(n15451) );
  INV_X1 U11195 ( .A(n15209), .ZN(n10515) );
  NAND2_X1 U11196 ( .A1(n13722), .A2(n13082), .ZN(n13747) );
  NOR2_X1 U11198 ( .A1(n11579), .A2(n11578), .ZN(n18336) );
  OR2_X1 U11199 ( .A1(n10017), .A2(n10904), .ZN(n11321) );
  AND2_X1 U11201 ( .A1(n11066), .A2(n11065), .ZN(n11112) );
  CLKBUF_X1 U11202 ( .A(n10656), .Z(n14360) );
  AND2_X1 U11203 ( .A1(n11059), .A2(n11067), .ZN(n11125) );
  CLKBUF_X2 U11204 ( .A(n15808), .Z(n15871) );
  BUF_X1 U11205 ( .A(n10454), .Z(n14349) );
  NAND2_X1 U11206 ( .A1(n11182), .A2(n11181), .ZN(n11180) );
  CLKBUF_X1 U11207 ( .A(n12853), .Z(n14296) );
  CLKBUF_X1 U11208 ( .A(n14308), .Z(n9815) );
  CLKBUF_X1 U11209 ( .A(n11044), .Z(n11058) );
  BUF_X1 U11211 ( .A(n19990), .Z(n9772) );
  INV_X1 U11212 ( .A(n10639), .ZN(n13166) );
  INV_X1 U11213 ( .A(n10810), .ZN(n13165) );
  AND2_X1 U11214 ( .A1(n10375), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10603) );
  AND2_X1 U11215 ( .A1(n13998), .A2(n10595), .ZN(n13175) );
  AND2_X1 U11216 ( .A1(n9761), .A2(n10371), .ZN(n13173) );
  AND2_X1 U11217 ( .A1(n9760), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10736) );
  CLKBUF_X2 U11219 ( .A(n10286), .Z(n13352) );
  INV_X1 U11220 ( .A(n10373), .ZN(n10588) );
  INV_X1 U11222 ( .A(n9822), .ZN(n15894) );
  BUF_X2 U11223 ( .A(n10594), .Z(n13356) );
  INV_X1 U11224 ( .A(n11602), .ZN(n17224) );
  NAND2_X1 U11225 ( .A1(n10399), .A2(n14058), .ZN(n10983) );
  NOR2_X1 U11226 ( .A1(n11398), .A2(n17011), .ZN(n15826) );
  NOR2_X2 U11227 ( .A1(n11398), .A2(n18778), .ZN(n15808) );
  NAND2_X2 U11230 ( .A1(n10401), .A2(n10400), .ZN(n10433) );
  CLKBUF_X1 U11231 ( .A(n10385), .Z(n13539) );
  NOR2_X1 U11232 ( .A1(n10402), .A2(n10984), .ZN(n10390) );
  NAND2_X1 U11234 ( .A1(n10392), .A2(n13564), .ZN(n10402) );
  NAND2_X1 U11235 ( .A1(n10310), .A2(n10309), .ZN(n10984) );
  AND2_X4 U11236 ( .A1(n14025), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10286) );
  INV_X1 U11237 ( .A(n9753), .ZN(n9754) );
  AND2_X1 U11238 ( .A1(n11708), .A2(n11709), .ZN(n11854) );
  AND2_X1 U11239 ( .A1(n11709), .A2(n13621), .ZN(n11862) );
  INV_X1 U11240 ( .A(n9758), .ZN(n9760) );
  INV_X2 U11241 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10574) );
  CLKBUF_X1 U11242 ( .A(n18523), .Z(n9747) );
  NOR2_X1 U11243 ( .A1(n18532), .A2(n18480), .ZN(n18523) );
  NAND2_X4 U11244 ( .A1(n18747), .A2(n11640), .ZN(n18771) );
  INV_X2 U11245 ( .A(n17459), .ZN(n18343) );
  NOR2_X2 U11246 ( .A1(n18181), .A2(n18192), .ZN(n18230) );
  INV_X4 U11247 ( .A(n16230), .ZN(n20236) );
  INV_X1 U11250 ( .A(n15205), .ZN(n9750) );
  INV_X1 U11251 ( .A(n9754), .ZN(n9756) );
  NAND2_X1 U11252 ( .A1(n12847), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12759) );
  INV_X1 U11253 ( .A(n10357), .ZN(n9758) );
  INV_X1 U11254 ( .A(n9758), .ZN(n9761) );
  INV_X1 U11255 ( .A(n10464), .ZN(n10511) );
  INV_X1 U11256 ( .A(n9754), .ZN(n9755) );
  AND2_X1 U11257 ( .A1(n9798), .A2(n11709), .ZN(n12001) );
  INV_X1 U11258 ( .A(n10454), .ZN(n10508) );
  INV_X1 U11260 ( .A(n9758), .ZN(n9759) );
  INV_X1 U11261 ( .A(n9754), .ZN(n9757) );
  AND2_X1 U11262 ( .A1(n10286), .A2(n10355), .ZN(n13172) );
  AND2_X1 U11263 ( .A1(n10374), .A2(n10371), .ZN(n10666) );
  AND2_X1 U11264 ( .A1(n15764), .A2(n10072), .ZN(n11065) );
  NAND2_X1 U11265 ( .A1(n10298), .A2(n10903), .ZN(n10385) );
  NOR2_X1 U11266 ( .A1(n14387), .A2(n11026), .ZN(n14364) );
  NOR2_X1 U11267 ( .A1(n15609), .A2(n11364), .ZN(n15597) );
  AND2_X1 U11268 ( .A1(n10646), .A2(n10645), .ZN(n11094) );
  INV_X1 U11269 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10371) );
  AND2_X1 U11270 ( .A1(n11066), .A2(n11067), .ZN(n11124) );
  AND3_X1 U11271 ( .A1(n10394), .A2(n10405), .A3(n10393), .ZN(n10980) );
  CLKBUF_X2 U11272 ( .A(n11455), .Z(n17269) );
  NAND2_X1 U11273 ( .A1(n11506), .A2(n18074), .ZN(n17759) );
  CLKBUF_X2 U11274 ( .A(n13467), .Z(n9818) );
  NAND2_X1 U11275 ( .A1(n19990), .A2(n14103), .ZN(n11186) );
  OAI21_X1 U11276 ( .B1(n15420), .B2(n15419), .A(n15372), .ZN(n15411) );
  INV_X1 U11278 ( .A(n14103), .ZN(n14058) );
  INV_X1 U11279 ( .A(n17812), .ZN(n17802) );
  OR2_X1 U11280 ( .A1(n14746), .A2(n14745), .ZN(n14748) );
  AND2_X1 U11282 ( .A1(n9940), .A2(n9939), .ZN(n9788) );
  NAND2_X1 U11283 ( .A1(n15415), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9794) );
  NAND2_X2 U11284 ( .A1(n10350), .A2(n10349), .ZN(n19990) );
  NOR2_X2 U11285 ( .A1(n18961), .A2(n16654), .ZN(n17955) );
  INV_X1 U11286 ( .A(n20039), .ZN(n20107) );
  AOI211_X1 U11287 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15486), .A(
        n14392), .B(n14391), .ZN(n14393) );
  INV_X1 U11288 ( .A(n17950), .ZN(n17965) );
  INV_X2 U11289 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16981) );
  AND2_X2 U11290 ( .A1(n10161), .A2(n13621), .ZN(n9751) );
  NAND3_X1 U11291 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n9802) );
  NAND2_X2 U11293 ( .A1(n11002), .A2(n10443), .ZN(n11005) );
  OAI21_X2 U11294 ( .B1(n12686), .B2(n12687), .A(n10121), .ZN(n12696) );
  NAND2_X2 U11295 ( .A1(n11890), .A2(n11889), .ZN(n11912) );
  NOR2_X2 U11297 ( .A1(n11203), .A2(n10914), .ZN(n11182) );
  OAI21_X2 U11298 ( .B1(n14929), .B2(n10006), .A(n10125), .ZN(n12782) );
  NAND2_X2 U11299 ( .A1(n14967), .A2(n12770), .ZN(n14929) );
  NOR2_X2 U11301 ( .A1(n17919), .A2(n11498), .ZN(n17903) );
  AND2_X1 U11302 ( .A1(n10271), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9753) );
  AND2_X1 U11303 ( .A1(n10271), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10357) );
  AND2_X1 U11304 ( .A1(n13992), .A2(n10574), .ZN(n9762) );
  AND2_X1 U11305 ( .A1(n13992), .A2(n10574), .ZN(n9763) );
  BUF_X1 U11306 ( .A(n17532), .Z(n9764) );
  NOR4_X1 U11307 ( .A1(n18307), .A2(n12991), .A3(n17343), .A4(n11631), .ZN(
        n17532) );
  NOR2_X4 U11308 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14016) );
  CLKBUF_X3 U11309 ( .A(n13188), .Z(n10589) );
  AND2_X4 U11310 ( .A1(n13998), .A2(n10272), .ZN(n13188) );
  OAI21_X2 U11311 ( .B1(n12695), .B2(n11824), .A(n12694), .ZN(n12697) );
  OAI21_X4 U11312 ( .B1(n14677), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11928), 
        .ZN(n12695) );
  AND4_X1 U11313 ( .A1(n10751), .A2(n10750), .A3(n10749), .A4(n10748), .ZN(
        n9765) );
  AND2_X1 U11314 ( .A1(n10589), .A2(n10371), .ZN(n9766) );
  AND2_X1 U11315 ( .A1(n10589), .A2(n10371), .ZN(n10665) );
  XNOR2_X2 U11316 ( .A(n13202), .B(n13228), .ZN(n15138) );
  AND2_X4 U11317 ( .A1(n13992), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9767) );
  XNOR2_X1 U11318 ( .A(n14878), .B(n9809), .ZN(n9808) );
  OR2_X1 U11319 ( .A1(n15114), .A2(n13327), .ZN(n10066) );
  NAND2_X1 U11321 ( .A1(n15735), .A2(n11163), .ZN(n11168) );
  NOR2_X1 U11322 ( .A1(n15104), .A2(n14345), .ZN(n14351) );
  NAND2_X1 U11323 ( .A1(n15102), .A2(n15101), .ZN(n15104) );
  NAND2_X1 U11324 ( .A1(n13794), .A2(n12705), .ZN(n12712) );
  AND2_X1 U11325 ( .A1(n14729), .A2(n14535), .ZN(n14718) );
  NOR2_X2 U11326 ( .A1(n14748), .A2(n14581), .ZN(n14580) );
  AND2_X1 U11329 ( .A1(n11064), .A2(n11067), .ZN(n11115) );
  AND2_X1 U11330 ( .A1(n11064), .A2(n11053), .ZN(n11116) );
  AND2_X1 U11331 ( .A1(n11068), .A2(n11067), .ZN(n19338) );
  AND2_X1 U11332 ( .A1(n11064), .A2(n11065), .ZN(n11126) );
  NAND2_X1 U11333 ( .A1(n13819), .A2(n11944), .ZN(n13654) );
  OAI21_X1 U11334 ( .B1(n10072), .B2(n13069), .A(n13053), .ZN(n15775) );
  NAND2_X2 U11335 ( .A1(n11042), .A2(n11041), .ZN(n11049) );
  NAND2_X1 U11336 ( .A1(n14093), .A2(n9772), .ZN(n13596) );
  NAND2_X1 U11337 ( .A1(n16541), .A2(n16534), .ZN(n17838) );
  NAND2_X1 U11338 ( .A1(n10409), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10454) );
  AND2_X1 U11339 ( .A1(n10983), .A2(n10582), .ZN(n11002) );
  NAND2_X1 U11341 ( .A1(n10980), .A2(n10432), .ZN(n10464) );
  NAND2_X2 U11342 ( .A1(n14291), .A2(n13467), .ZN(n14301) );
  INV_X2 U11343 ( .A(n11654), .ZN(n10076) );
  NAND3_X2 U11344 ( .A1(n10647), .A2(n10625), .A3(n10904), .ZN(n10655) );
  INV_X2 U11345 ( .A(n18961), .ZN(n15915) );
  INV_X1 U11346 ( .A(n11826), .ZN(n11819) );
  NOR2_X1 U11347 ( .A1(n11823), .A2(n9802), .ZN(n13733) );
  OR2_X2 U11348 ( .A1(n11715), .A2(n11714), .ZN(n20284) );
  INV_X1 U11349 ( .A(n10984), .ZN(n19355) );
  INV_X1 U11350 ( .A(n10400), .ZN(n10381) );
  INV_X1 U11352 ( .A(n9822), .ZN(n17297) );
  BUF_X2 U11353 ( .A(n11860), .Z(n12596) );
  CLKBUF_X2 U11355 ( .A(n15826), .Z(n17295) );
  CLKBUF_X2 U11356 ( .A(n11455), .Z(n17298) );
  CLKBUF_X2 U11357 ( .A(n15819), .Z(n15868) );
  INV_X2 U11359 ( .A(n18289), .ZN(n9768) );
  NAND2_X1 U11360 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18778) );
  NAND2_X1 U11362 ( .A1(n12791), .A2(n12788), .ZN(n14867) );
  OR2_X1 U11363 ( .A1(n11388), .A2(n16456), .ZN(n11389) );
  INV_X1 U11364 ( .A(n9808), .ZN(n16162) );
  AOI211_X1 U11365 ( .C1(n19302), .C2(n19025), .A(n15407), .B(n15406), .ZN(
        n15408) );
  AND2_X1 U11367 ( .A1(n10145), .A2(n10144), .ZN(n11348) );
  MUX2_X1 U11368 ( .A(n13042), .B(n13041), .S(n16134), .Z(n13043) );
  OR2_X1 U11370 ( .A1(n9794), .A2(n15572), .ZN(n15392) );
  NAND2_X1 U11371 ( .A1(n10146), .A2(n11333), .ZN(n10143) );
  XNOR2_X1 U11372 ( .A(n12618), .B(n12617), .ZN(n14439) );
  INV_X1 U11373 ( .A(n16093), .ZN(n14811) );
  OR2_X1 U11374 ( .A1(n14507), .A2(n14704), .ZN(n16016) );
  NOR2_X1 U11375 ( .A1(n16412), .A2(n16472), .ZN(n16411) );
  AOI21_X1 U11376 ( .B1(n15441), .B2(n15437), .A(n15439), .ZN(n15429) );
  CLKBUF_X1 U11377 ( .A(n14506), .Z(n14507) );
  AND2_X1 U11378 ( .A1(n14506), .A2(n10174), .ZN(n14466) );
  AND2_X1 U11379 ( .A1(n14716), .A2(n14715), .ZN(n16093) );
  OR2_X1 U11380 ( .A1(n15446), .A2(n15673), .ZN(n16412) );
  OR2_X1 U11381 ( .A1(n13327), .A2(n10058), .ZN(n10057) );
  AOI21_X1 U11382 ( .B1(n15644), .B2(n15368), .A(n15645), .ZN(n15441) );
  NAND2_X1 U11384 ( .A1(n10153), .A2(n10154), .ZN(n15680) );
  XNOR2_X1 U11385 ( .A(n11168), .B(n11166), .ZN(n15470) );
  NAND2_X1 U11386 ( .A1(n15104), .A2(n15103), .ZN(n16347) );
  XNOR2_X1 U11387 ( .A(n15104), .B(n14345), .ZN(n11028) );
  NAND2_X1 U11388 ( .A1(n10056), .A2(n14314), .ZN(n13276) );
  NAND2_X1 U11389 ( .A1(n15726), .A2(n15725), .ZN(n9899) );
  NOR2_X1 U11390 ( .A1(n11172), .A2(n15710), .ZN(n10190) );
  NAND2_X1 U11391 ( .A1(n14316), .A2(n14315), .ZN(n14314) );
  XNOR2_X1 U11392 ( .A(n11212), .B(n15727), .ZN(n15726) );
  NAND2_X1 U11393 ( .A1(n11211), .A2(n19153), .ZN(n11212) );
  NOR2_X1 U11394 ( .A1(n16532), .A2(n17838), .ZN(n15924) );
  CLKBUF_X1 U11395 ( .A(n11161), .Z(n15747) );
  XNOR2_X1 U11396 ( .A(n11165), .B(n11169), .ZN(n11166) );
  AND2_X1 U11397 ( .A1(n14326), .A2(n14327), .ZN(n15125) );
  OAI21_X1 U11398 ( .B1(n16109), .B2(n12914), .A(n16134), .ZN(n10007) );
  NAND2_X1 U11399 ( .A1(n15744), .A2(n15742), .ZN(n11161) );
  AND2_X1 U11400 ( .A1(n16110), .A2(n10126), .ZN(n10125) );
  CLKBUF_X1 U11401 ( .A(n11164), .Z(n11165) );
  MUX2_X1 U11402 ( .A(n14456), .B(n9817), .S(n14451), .Z(n14310) );
  NAND2_X1 U11403 ( .A1(n9900), .A2(n11150), .ZN(n11164) );
  NOR2_X1 U11404 ( .A1(n14268), .A2(n10130), .ZN(n10129) );
  OR2_X1 U11405 ( .A1(n14487), .A2(n14486), .ZN(n14999) );
  NAND2_X1 U11406 ( .A1(n11179), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15743) );
  NAND2_X1 U11407 ( .A1(n9943), .A2(n9941), .ZN(n15741) );
  OR2_X1 U11408 ( .A1(n13436), .A2(n14386), .ZN(n14415) );
  OR2_X1 U11409 ( .A1(n14959), .A2(n14958), .ZN(n10004) );
  AND2_X1 U11410 ( .A1(n14943), .A2(n12773), .ZN(n16118) );
  AND2_X1 U11411 ( .A1(n12767), .A2(n12766), .ZN(n14268) );
  AND2_X1 U11412 ( .A1(n12737), .A2(n12736), .ZN(n16151) );
  NAND2_X1 U11414 ( .A1(n15231), .A2(n13437), .ZN(n13436) );
  NAND2_X1 U11415 ( .A1(n12071), .A2(n12070), .ZN(n13987) );
  NAND2_X1 U11416 ( .A1(n14706), .A2(n14705), .ZN(n14708) );
  OR2_X1 U11417 ( .A1(n12722), .A2(n12120), .ZN(n12071) );
  INV_X1 U11418 ( .A(n13961), .ZN(n13088) );
  NOR2_X2 U11419 ( .A1(n15233), .A2(n15232), .ZN(n15231) );
  NAND2_X1 U11420 ( .A1(n11149), .A2(n11148), .ZN(n11158) );
  OR2_X1 U11421 ( .A1(n15240), .A2(n14317), .ZN(n15233) );
  OR2_X1 U11422 ( .A1(n15050), .A2(n15242), .ZN(n15240) );
  AND2_X1 U11423 ( .A1(n14244), .A2(n14254), .ZN(n15207) );
  NAND2_X1 U11424 ( .A1(n12062), .A2(n12061), .ZN(n12092) );
  NAND2_X1 U11425 ( .A1(n9934), .A2(n11088), .ZN(n11090) );
  NAND2_X1 U11426 ( .A1(n10152), .A2(n11132), .ZN(n11134) );
  NAND2_X1 U11427 ( .A1(n14718), .A2(n14717), .ZN(n14720) );
  OR2_X1 U11428 ( .A1(n11146), .A2(n11145), .ZN(n11149) );
  AND3_X1 U11429 ( .A1(n11071), .A2(n11069), .A3(n11070), .ZN(n9859) );
  NAND4_X1 U11430 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n11120), .ZN(
        n10152) );
  AND2_X1 U11431 ( .A1(n15263), .A2(n15264), .ZN(n15262) );
  AND4_X1 U11432 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11086) );
  XNOR2_X1 U11433 ( .A(n13830), .B(n10160), .ZN(n20252) );
  AND2_X1 U11434 ( .A1(n11118), .A2(n10150), .ZN(n10149) );
  NAND2_X1 U11435 ( .A1(n14580), .A2(n14564), .ZN(n14566) );
  NOR2_X1 U11436 ( .A1(n15274), .A2(n15275), .ZN(n15263) );
  AOI22_X1 U11437 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n15795), .B1(
        n11113), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U11438 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11121), .B1(
        n11112), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11076) );
  AND2_X1 U11439 ( .A1(n15672), .A2(n11024), .ZN(n16473) );
  AND2_X1 U11440 ( .A1(n11059), .A2(n11053), .ZN(n11111) );
  AND2_X1 U11441 ( .A1(n11066), .A2(n11053), .ZN(n11113) );
  AND2_X1 U11442 ( .A1(n13081), .A2(n13080), .ZN(n13082) );
  NOR2_X2 U11443 ( .A1(n14396), .A2(n20259), .ZN(n14397) );
  AND2_X1 U11444 ( .A1(n13079), .A2(n13081), .ZN(n13723) );
  AND2_X1 U11445 ( .A1(n13560), .A2(n13061), .ZN(n13667) );
  AND2_X1 U11446 ( .A1(n11066), .A2(n11063), .ZN(n11123) );
  AND2_X1 U11447 ( .A1(n14221), .A2(n14120), .ZN(n11066) );
  AND2_X1 U11448 ( .A1(n11064), .A2(n11063), .ZN(n11121) );
  OR2_X1 U11449 ( .A1(n13078), .A2(n13077), .ZN(n13081) );
  AND2_X1 U11450 ( .A1(n11068), .A2(n11053), .ZN(n19375) );
  NAND2_X1 U11451 ( .A1(n14221), .A2(n13726), .ZN(n11060) );
  AND2_X1 U11452 ( .A1(n11068), .A2(n11063), .ZN(n15795) );
  AND2_X1 U11453 ( .A1(n12010), .A2(n12009), .ZN(n13829) );
  XNOR2_X1 U11454 ( .A(n9999), .B(n11963), .ZN(n11964) );
  NAND2_X2 U11455 ( .A1(n14861), .A2(n14135), .ZN(n14866) );
  NOR2_X1 U11456 ( .A1(n20119), .A2(n20979), .ZN(n20140) );
  OR2_X1 U11457 ( .A1(n13739), .A2(n13740), .ZN(n13737) );
  NOR2_X1 U11459 ( .A1(n15764), .A2(n19301), .ZN(n11067) );
  NOR2_X1 U11460 ( .A1(n13445), .A2(n10048), .ZN(n14145) );
  NOR2_X1 U11461 ( .A1(n13075), .A2(n13074), .ZN(n13078) );
  AND2_X1 U11462 ( .A1(n13669), .A2(n13726), .ZN(n11068) );
  OAI21_X1 U11463 ( .B1(n13669), .B2(n13069), .A(n13063), .ZN(n13067) );
  CLKBUF_X1 U11464 ( .A(n13654), .Z(n20690) );
  AND2_X1 U11465 ( .A1(n14120), .A2(n13669), .ZN(n11064) );
  NAND2_X1 U11466 ( .A1(n13444), .A2(n13446), .ZN(n13445) );
  NAND2_X2 U11467 ( .A1(n11052), .A2(n11051), .ZN(n15764) );
  NAND2_X1 U11468 ( .A1(n17960), .A2(n17864), .ZN(n17954) );
  CLKBUF_X1 U11469 ( .A(n14677), .Z(n20550) );
  NOR2_X1 U11470 ( .A1(n16501), .A2(n10459), .ZN(n15728) );
  CLKBUF_X1 U11471 ( .A(n11048), .Z(n11052) );
  AND2_X1 U11472 ( .A1(n19301), .A2(n11058), .ZN(n11053) );
  NOR2_X1 U11473 ( .A1(n11505), .A2(n18193), .ZN(n11682) );
  NAND2_X1 U11474 ( .A1(n11943), .A2(n11941), .ZN(n11939) );
  NAND2_X1 U11475 ( .A1(n10753), .A2(n10752), .ZN(n13689) );
  NOR2_X1 U11476 ( .A1(n10072), .A2(n11058), .ZN(n11063) );
  NAND2_X2 U11477 ( .A1(n15615), .A2(n9979), .ZN(n15762) );
  INV_X2 U11478 ( .A(n17434), .ZN(n17487) );
  NAND2_X1 U11479 ( .A1(n10449), .A2(n10448), .ZN(n11034) );
  NOR2_X1 U11480 ( .A1(n9920), .A2(n13413), .ZN(n16781) );
  NOR2_X2 U11481 ( .A1(n10625), .A2(n19367), .ZN(n19344) );
  AND2_X1 U11482 ( .A1(n10999), .A2(n16503), .ZN(n11351) );
  NAND2_X1 U11483 ( .A1(n11917), .A2(n11916), .ZN(n11920) );
  NAND2_X1 U11485 ( .A1(n11932), .A2(n11931), .ZN(n11941) );
  XNOR2_X1 U11486 ( .A(n10462), .B(n10461), .ZN(n11039) );
  NAND2_X1 U11487 ( .A1(n11942), .A2(n11940), .ZN(n11938) );
  NOR2_X1 U11488 ( .A1(n10661), .A2(n9829), .ZN(n10036) );
  OAI21_X1 U11489 ( .B1(n18758), .B2(n11642), .A(n18757), .ZN(n18192) );
  NAND2_X1 U11490 ( .A1(n10453), .A2(n10452), .ZN(n10462) );
  INV_X1 U11491 ( .A(n13775), .ZN(n9770) );
  AOI221_X1 U11492 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16507), .C1(n19983), .C2(
        n16507), .A(n19738), .ZN(n19977) );
  OAI21_X2 U11493 ( .B1(n19996), .B2(n13483), .A(n13597), .ZN(n13484) );
  CLKBUF_X1 U11494 ( .A(n11918), .Z(n11919) );
  OAI21_X1 U11495 ( .B1(n13005), .B2(n13004), .A(n18955), .ZN(n18217) );
  AND3_X1 U11496 ( .A1(n10429), .A2(n10428), .A3(n10427), .ZN(n10431) );
  AND2_X1 U11497 ( .A1(n11846), .A2(n11845), .ZN(n11921) );
  OAI21_X1 U11498 ( .B1(n10454), .B2(n10459), .A(n10458), .ZN(n10461) );
  NAND2_X2 U11499 ( .A1(n17531), .A2(n18798), .ZN(n17594) );
  AND2_X1 U11500 ( .A1(n13545), .A2(n13546), .ZN(n10650) );
  AND2_X1 U11501 ( .A1(n12622), .A2(n14308), .ZN(n12950) );
  NAND2_X1 U11502 ( .A1(n11766), .A2(n11825), .ZN(n11830) );
  OR2_X1 U11503 ( .A1(n13612), .A2(n12825), .ZN(n9853) );
  INV_X1 U11505 ( .A(n12988), .ZN(n18315) );
  NAND2_X1 U11506 ( .A1(n10336), .A2(n10335), .ZN(n10181) );
  AND2_X1 U11507 ( .A1(n11823), .A2(n11827), .ZN(n11766) );
  INV_X1 U11508 ( .A(n10433), .ZN(n9950) );
  NAND2_X2 U11509 ( .A1(n9843), .A2(n9994), .ZN(n17459) );
  INV_X1 U11510 ( .A(n11823), .ZN(n12847) );
  OR2_X1 U11511 ( .A1(n11882), .A2(n11881), .ZN(n12763) );
  NAND2_X1 U11512 ( .A1(n20272), .A2(n20284), .ZN(n12850) );
  AND2_X1 U11513 ( .A1(n11441), .A2(n10204), .ZN(n11654) );
  NAND3_X1 U11514 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n9803) );
  INV_X1 U11515 ( .A(n20284), .ZN(n9771) );
  NAND2_X1 U11516 ( .A1(n10404), .A2(n11186), .ZN(n11015) );
  AND3_X1 U11517 ( .A1(n9856), .A2(n11612), .A3(n11611), .ZN(n9994) );
  NOR2_X1 U11519 ( .A1(n11186), .A2(n16509), .ZN(n10432) );
  INV_X1 U11521 ( .A(n11186), .ZN(n11349) );
  AND2_X2 U11522 ( .A1(n9968), .A2(n9966), .ZN(n9855) );
  INV_X2 U11524 ( .A(U212), .ZN(n16602) );
  BUF_X2 U11525 ( .A(n10903), .Z(n11190) );
  NAND3_X2 U11527 ( .A1(n11781), .A2(n11780), .A3(n11779), .ZN(n20278) );
  NAND2_X2 U11528 ( .A1(n10322), .A2(n10321), .ZN(n13564) );
  AND3_X1 U11529 ( .A1(n11778), .A2(n11777), .A3(n11776), .ZN(n11779) );
  MUX2_X1 U11530 ( .A(n10333), .B(n10332), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19351) );
  INV_X2 U11531 ( .A(U214), .ZN(n16606) );
  AND4_X1 U11532 ( .A1(n11735), .A2(n11739), .A3(n11737), .A4(n11732), .ZN(
        n9820) );
  INV_X2 U11534 ( .A(n10965), .ZN(n13171) );
  INV_X2 U11535 ( .A(n10811), .ZN(n13164) );
  AND3_X1 U11536 ( .A1(n11757), .A2(n11754), .A3(n11762), .ZN(n10122) );
  NAND4_X1 U11537 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10296) );
  AND4_X1 U11538 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n11781) );
  NAND2_X1 U11539 ( .A1(n10343), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10350) );
  INV_X2 U11540 ( .A(n18956), .ZN(n17527) );
  BUF_X4 U11541 ( .A(n11606), .Z(n9773) );
  INV_X2 U11542 ( .A(n18832), .ZN(n18895) );
  BUF_X2 U11543 ( .A(n15808), .Z(n17289) );
  INV_X2 U11545 ( .A(n16634), .ZN(U215) );
  NAND2_X2 U11546 ( .A1(n20009), .A2(n19884), .ZN(n19926) );
  AND2_X2 U11548 ( .A1(n11706), .A2(n11708), .ZN(n11946) );
  OR2_X2 U11549 ( .A1(n11694), .A2(n11692), .ZN(n11945) );
  NOR2_X1 U11551 ( .A1(n11400), .A2(n11401), .ZN(n11477) );
  OR2_X1 U11552 ( .A1(n11397), .A2(n11401), .ZN(n9850) );
  BUF_X4 U11553 ( .A(n11413), .Z(n9775) );
  OR2_X1 U11554 ( .A1(n11402), .A2(n11401), .ZN(n9849) );
  BUF_X2 U11555 ( .A(n11392), .Z(n17249) );
  INV_X2 U11556 ( .A(n18970), .ZN(n18972) );
  INV_X2 U11557 ( .A(n16643), .ZN(n16645) );
  AND2_X2 U11558 ( .A1(n10270), .A2(n10563), .ZN(n10594) );
  AND3_X1 U11559 ( .A1(n13684), .A2(n12011), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11699) );
  AND2_X1 U11560 ( .A1(n10119), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11704) );
  AND2_X2 U11564 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13992) );
  AND2_X1 U11565 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13998) );
  AND2_X1 U11566 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10270) );
  NOR2_X1 U11567 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14025) );
  NOR2_X1 U11568 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10271) );
  AOI21_X1 U11572 ( .B1(n15680), .B2(n9825), .A(n9951), .ZN(n15355) );
  OAI21_X1 U11573 ( .B1(n14929), .B2(n10006), .A(n10125), .ZN(n9776) );
  NAND2_X1 U11574 ( .A1(n9771), .A2(n9777), .ZN(n9778) );
  NAND2_X1 U11575 ( .A1(n9778), .A2(n11830), .ZN(n11787) );
  INV_X1 U11576 ( .A(n12825), .ZN(n9777) );
  NAND2_X1 U11578 ( .A1(n14868), .A2(n9781), .ZN(n9782) );
  NAND2_X1 U11579 ( .A1(n9780), .A2(n14869), .ZN(n9783) );
  NAND2_X1 U11580 ( .A1(n9782), .A2(n9783), .ZN(n9847) );
  INV_X1 U11581 ( .A(n14868), .ZN(n9780) );
  INV_X1 U11582 ( .A(n14869), .ZN(n9781) );
  INV_X2 U11583 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9784) );
  INV_X1 U11584 ( .A(n13847), .ZN(n9785) );
  XNOR2_X1 U11585 ( .A(n11923), .B(n11921), .ZN(n11982) );
  AND2_X1 U11586 ( .A1(n15427), .A2(n15369), .ZN(n9786) );
  AND2_X1 U11587 ( .A1(n15427), .A2(n15369), .ZN(n15420) );
  XNOR2_X1 U11588 ( .A(n9787), .B(n9789), .ZN(n15594) );
  AND2_X1 U11589 ( .A1(n15410), .A2(n15409), .ZN(n9787) );
  INV_X1 U11590 ( .A(n11925), .ZN(n11924) );
  NOR2_X2 U11591 ( .A1(n15502), .A2(n15517), .ZN(n15481) );
  AND2_X2 U11592 ( .A1(n11699), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11852) );
  AOI211_X1 U11593 ( .C1(n11896), .C2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n12594), .B(n12593), .ZN(n12598) );
  AOI211_X1 U11594 ( .C1(n11896), .C2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n12561), .B(n12560), .ZN(n12563) );
  AND2_X1 U11595 ( .A1(n9940), .A2(n9939), .ZN(n15314) );
  OAI21_X1 U11596 ( .B1(n9786), .B2(n15419), .A(n15372), .ZN(n9789) );
  INV_X1 U11597 ( .A(n20349), .ZN(n9790) );
  OR2_X1 U11598 ( .A1(n11912), .A2(n11911), .ZN(n9791) );
  AND2_X1 U11600 ( .A1(n10192), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9793) );
  AND2_X1 U11601 ( .A1(n9798), .A2(n11709), .ZN(n9814) );
  INV_X1 U11602 ( .A(n15451), .ZN(n9796) );
  INV_X1 U11603 ( .A(n9796), .ZN(n9797) );
  AND2_X1 U11604 ( .A1(n9784), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9798) );
  XNOR2_X1 U11605 ( .A(n14377), .B(n14376), .ZN(n15304) );
  AOI21_X1 U11606 ( .B1(n9797), .B2(n15447), .A(n15449), .ZN(n9800) );
  AOI21_X2 U11607 ( .B1(n15451), .B2(n15447), .A(n15449), .ZN(n15644) );
  AND2_X2 U11608 ( .A1(n11108), .A2(n14150), .ZN(n15744) );
  AND2_X1 U11609 ( .A1(n11819), .A2(n9802), .ZN(n9801) );
  NAND3_X1 U11611 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n11821) );
  AND2_X1 U11612 ( .A1(n15415), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9804) );
  NAND2_X1 U11613 ( .A1(n9898), .A2(n10427), .ZN(n10451) );
  NAND2_X1 U11614 ( .A1(n10388), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9898) );
  OAI22_X1 U11615 ( .A1(n15304), .A2(n15479), .B1(n14378), .B2(n14379), .ZN(
        n10182) );
  INV_X4 U11616 ( .A(n10903), .ZN(n10904) );
  AOI21_X1 U11618 ( .B1(n15441), .B2(n15437), .A(n15439), .ZN(n9806) );
  NAND2_X1 U11619 ( .A1(n9791), .A2(n11913), .ZN(n9807) );
  AOI21_X2 U11621 ( .B1(n15345), .B2(n15346), .A(n11309), .ZN(n15333) );
  NAND2_X1 U11623 ( .A1(n11929), .A2(n11913), .ZN(n11972) );
  OR2_X2 U11624 ( .A1(n9794), .A2(n15574), .ZN(n15405) );
  NAND2_X1 U11625 ( .A1(n15734), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15735) );
  INV_X1 U11626 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9809) );
  NOR2_X4 U11627 ( .A1(n15446), .A2(n11174), .ZN(n15435) );
  NAND2_X1 U11628 ( .A1(n20173), .A2(n20172), .ZN(n9810) );
  INV_X1 U11629 ( .A(n12785), .ZN(n9811) );
  NOR2_X1 U11630 ( .A1(n11767), .A2(n11823), .ZN(n9812) );
  INV_X1 U11631 ( .A(n12785), .ZN(n14884) );
  NOR2_X1 U11632 ( .A1(n11767), .A2(n11823), .ZN(n11788) );
  AND2_X2 U11634 ( .A1(n14163), .A2(n14171), .ZN(n14172) );
  NOR2_X2 U11635 ( .A1(n14162), .A2(n14161), .ZN(n14163) );
  OAI21_X1 U11636 ( .B1(n13828), .B2(n12120), .A(n11970), .ZN(n11971) );
  AND2_X4 U11637 ( .A1(n14016), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9813) );
  NAND2_X2 U11638 ( .A1(n12786), .A2(n14902), .ZN(n12785) );
  NAND2_X2 U11639 ( .A1(n14903), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12786) );
  NAND2_X1 U11640 ( .A1(n11886), .A2(n11885), .ZN(n11980) );
  NAND2_X1 U11641 ( .A1(n12853), .A2(n12850), .ZN(n14308) );
  NOR2_X2 U11643 ( .A1(n11831), .A2(n11803), .ZN(n12831) );
  NAND2_X2 U11644 ( .A1(n11787), .A2(n11786), .ZN(n11831) );
  AOI21_X1 U11645 ( .B1(n11933), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11934), .ZN(n11942) );
  AND2_X2 U11646 ( .A1(n14887), .A2(n12787), .ZN(n9842) );
  INV_X1 U11647 ( .A(n12850), .ZN(n9817) );
  BUF_X4 U11648 ( .A(n12850), .Z(n14291) );
  NOR2_X2 U11651 ( .A1(n14520), .A2(n12452), .ZN(n14522) );
  AND2_X1 U11652 ( .A1(n20272), .A2(n20261), .ZN(n13467) );
  NOR2_X1 U11653 ( .A1(n19250), .A2(n20002), .ZN(n19279) );
  AND3_X1 U11655 ( .A1(n10983), .A2(n14070), .A3(n10443), .ZN(n10408) );
  NAND2_X1 U11656 ( .A1(n9950), .A2(n9948), .ZN(n9947) );
  AND2_X1 U11657 ( .A1(n19990), .A2(n13600), .ZN(n9948) );
  NOR2_X1 U11658 ( .A1(n10903), .A2(n10392), .ZN(n10405) );
  NAND2_X1 U11659 ( .A1(n9788), .A2(n9938), .ZN(n10146) );
  AND2_X1 U11660 ( .A1(n10210), .A2(n9863), .ZN(n9938) );
  AOI21_X1 U11661 ( .B1(n14346), .B2(P2_EBX_REG_3__SCAN_IN), .A(n10457), .ZN(
        n10458) );
  NAND3_X1 U11662 ( .A1(n9930), .A2(n11036), .A3(n9929), .ZN(n11040) );
  NAND2_X1 U11663 ( .A1(n10450), .A2(n11035), .ZN(n9930) );
  NOR3_X1 U11664 ( .A1(n9879), .A2(n10041), .A3(n10040), .ZN(n10039) );
  INV_X1 U11665 ( .A(n13437), .ZN(n10040) );
  INV_X1 U11666 ( .A(n10896), .ZN(n10041) );
  OR2_X1 U11667 ( .A1(n11868), .A2(n11867), .ZN(n12690) );
  OR2_X1 U11668 ( .A1(n10675), .A2(n10676), .ZN(n9982) );
  NAND2_X1 U11669 ( .A1(n11325), .A2(n11321), .ZN(n11314) );
  INV_X1 U11670 ( .A(n11478), .ZN(n11591) );
  NAND2_X1 U11671 ( .A1(n14197), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11992) );
  NAND3_X1 U11672 ( .A1(n11823), .A2(n20261), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12661) );
  NAND2_X1 U11673 ( .A1(n11314), .A2(n11324), .ZN(n11330) );
  NOR2_X1 U11674 ( .A1(n11257), .A2(n11256), .ZN(n11255) );
  NAND2_X1 U11675 ( .A1(n10828), .A2(n13981), .ZN(n10051) );
  CLKBUF_X1 U11676 ( .A(n10508), .Z(n10509) );
  NOR2_X1 U11677 ( .A1(n10051), .A2(n10050), .ZN(n10049) );
  INV_X1 U11678 ( .A(n15649), .ZN(n10050) );
  NAND2_X1 U11679 ( .A1(n11249), .A2(n15683), .ZN(n9955) );
  AOI21_X1 U11680 ( .B1(n9819), .B2(n11220), .A(n9830), .ZN(n10154) );
  NAND2_X1 U11681 ( .A1(n15468), .A2(n9819), .ZN(n10153) );
  AND2_X1 U11682 ( .A1(n13966), .A2(n13959), .ZN(n10016) );
  AND4_X1 U11683 ( .A1(n10724), .A2(n10723), .A3(n10722), .A4(n10721), .ZN(
        n10751) );
  AND4_X1 U11684 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        n10748) );
  NOR2_X1 U11685 ( .A1(n11399), .A2(n11397), .ZN(n11413) );
  INV_X2 U11686 ( .A(n15858), .ZN(n15895) );
  XOR2_X1 U11687 ( .A(n11500), .B(n17465), .Z(n11501) );
  NOR2_X1 U11688 ( .A1(n17940), .A2(n11491), .ZN(n11494) );
  NOR2_X1 U11689 ( .A1(n18278), .A2(n11490), .ZN(n11491) );
  OR2_X1 U11690 ( .A1(n9992), .A2(n11629), .ZN(n11639) );
  NAND2_X1 U11691 ( .A1(n14487), .A2(n14468), .ZN(n14451) );
  NAND4_X1 U11693 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10297) );
  OAI21_X1 U11694 ( .B1(n10143), .B2(n9960), .A(n9957), .ZN(n9961) );
  INV_X1 U11695 ( .A(n14374), .ZN(n9960) );
  AND2_X1 U11696 ( .A1(n14333), .A2(n9958), .ZN(n9957) );
  NOR2_X1 U11697 ( .A1(n15323), .A2(n11337), .ZN(n14374) );
  AND2_X1 U11698 ( .A1(n9839), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10192) );
  AND2_X1 U11699 ( .A1(n10467), .A2(n10466), .ZN(n13749) );
  OR2_X1 U11700 ( .A1(n14349), .A2(n15750), .ZN(n10467) );
  NAND2_X1 U11701 ( .A1(n11040), .A2(n10460), .ZN(n10010) );
  NOR2_X1 U11702 ( .A1(n16742), .A2(n9920), .ZN(n16734) );
  NAND2_X1 U11703 ( .A1(n10084), .A2(n17622), .ZN(n17612) );
  INV_X1 U11704 ( .A(n11520), .ZN(n10084) );
  NAND2_X1 U11705 ( .A1(n10938), .A2(n10937), .ZN(n10939) );
  NAND2_X1 U11706 ( .A1(n13374), .A2(n19182), .ZN(n10938) );
  NAND2_X1 U11707 ( .A1(n17606), .A2(n10198), .ZN(n16542) );
  INV_X1 U11708 ( .A(n12640), .ZN(n12658) );
  AND2_X1 U11709 ( .A1(n11117), .A2(n11130), .ZN(n10150) );
  NAND2_X1 U11710 ( .A1(n11136), .A2(n11135), .ZN(n11151) );
  INV_X1 U11711 ( .A(n11134), .ZN(n11135) );
  NAND2_X1 U11712 ( .A1(n11114), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11061) );
  AND2_X1 U11713 ( .A1(n11055), .A2(n11072), .ZN(n9937) );
  AOI22_X1 U11714 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n15795), .B1(
        n11123), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11072) );
  OR2_X1 U11716 ( .A1(n12060), .A2(n12059), .ZN(n12733) );
  NAND2_X1 U11717 ( .A1(n11923), .A2(n11922), .ZN(n11925) );
  OR2_X1 U11718 ( .A1(n12008), .A2(n12007), .ZN(n12716) );
  OAI21_X1 U11719 ( .B1(n10510), .B2(n15094), .A(n10441), .ZN(n10442) );
  OAI22_X1 U11720 ( .A1(n10464), .A2(n10439), .B1(n10456), .B2(n21219), .ZN(
        n10440) );
  NAND2_X1 U11721 ( .A1(n10414), .A2(n10413), .ZN(n10417) );
  NAND2_X1 U11722 ( .A1(n10012), .A2(n10397), .ZN(n10418) );
  NAND2_X1 U11723 ( .A1(n11085), .A2(n11086), .ZN(n9934) );
  AND4_X1 U11724 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11085) );
  NAND2_X1 U11725 ( .A1(n11087), .A2(n10625), .ZN(n11088) );
  INV_X1 U11726 ( .A(n10980), .ZN(n10978) );
  INV_X1 U11727 ( .A(n9982), .ZN(n11087) );
  INV_X1 U11728 ( .A(n10111), .ZN(n10109) );
  AND2_X1 U11729 ( .A1(n17479), .A2(n11652), .ZN(n11651) );
  NAND2_X1 U11730 ( .A1(n11630), .A2(n18321), .ZN(n9993) );
  AND2_X1 U11731 ( .A1(n13733), .A2(n11819), .ZN(n13469) );
  NOR2_X1 U11732 ( .A1(n10180), .A2(n14496), .ZN(n10179) );
  INV_X1 U11733 ( .A(n13045), .ZN(n10180) );
  NOR2_X1 U11734 ( .A1(n14552), .A2(n10165), .ZN(n10164) );
  INV_X1 U11735 ( .A(n10166), .ZN(n10165) );
  NOR2_X1 U11736 ( .A1(n14563), .A2(n10167), .ZN(n10166) );
  INV_X1 U11737 ( .A(n14579), .ZN(n10167) );
  OR2_X1 U11738 ( .A1(n15030), .A2(n20885), .ZN(n12574) );
  INV_X1 U11739 ( .A(n14755), .ZN(n12254) );
  AND2_X1 U11740 ( .A1(n10170), .A2(n9888), .ZN(n10169) );
  OR2_X1 U11741 ( .A1(n10171), .A2(n9875), .ZN(n10170) );
  XNOR2_X1 U11742 ( .A(n12761), .B(n12096), .ZN(n12743) );
  NAND3_X1 U11743 ( .A1(n10003), .A2(n12772), .A3(n10002), .ZN(n14928) );
  NAND2_X1 U11744 ( .A1(n12092), .A2(n12093), .ZN(n12732) );
  AND2_X1 U11745 ( .A1(n9817), .A2(n9818), .ZN(n14295) );
  NOR2_X2 U11746 ( .A1(n20284), .A2(n20278), .ZN(n13732) );
  OAI21_X1 U11747 ( .B1(n9982), .B2(n11186), .A(n9981), .ZN(n10943) );
  NAND2_X1 U11748 ( .A1(n10902), .A2(n11186), .ZN(n9981) );
  NAND2_X1 U11749 ( .A1(n10924), .A2(n11328), .ZN(n11340) );
  NOR2_X1 U11750 ( .A1(n10027), .A2(n11262), .ZN(n10026) );
  INV_X1 U11751 ( .A(n11265), .ZN(n10027) );
  INV_X1 U11752 ( .A(n11263), .ZN(n10025) );
  AND2_X1 U11753 ( .A1(n19111), .A2(n10918), .ZN(n10030) );
  NAND2_X1 U11754 ( .A1(n11241), .A2(n11245), .ZN(n11263) );
  NAND2_X1 U11755 ( .A1(n11246), .A2(n11321), .ZN(n11241) );
  AND2_X1 U11756 ( .A1(n11225), .A2(n10917), .ZN(n11232) );
  NAND2_X1 U11757 ( .A1(n11194), .A2(n11195), .ZN(n11196) );
  NAND2_X1 U11758 ( .A1(n9763), .A2(n10371), .ZN(n10639) );
  NAND2_X1 U11759 ( .A1(n9897), .A2(n13600), .ZN(n10427) );
  INV_X1 U11760 ( .A(n11001), .ZN(n9897) );
  NAND2_X1 U11761 ( .A1(n13278), .A2(n13277), .ZN(n10055) );
  INV_X1 U11762 ( .A(n10661), .ZN(n10034) );
  XNOR2_X1 U11763 ( .A(n11133), .B(n11134), .ZN(n11154) );
  INV_X1 U11764 ( .A(n10910), .ZN(n11097) );
  INV_X1 U11765 ( .A(n15188), .ZN(n10014) );
  AND2_X1 U11766 ( .A1(n10045), .A2(n15707), .ZN(n10044) );
  NOR2_X1 U11767 ( .A1(n16478), .A2(n10046), .ZN(n10045) );
  INV_X1 U11768 ( .A(n13688), .ZN(n10046) );
  NOR2_X1 U11769 ( .A1(n10137), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10134) );
  NAND2_X1 U11770 ( .A1(n10138), .A2(n10137), .ZN(n10136) );
  AND2_X1 U11771 ( .A1(n9945), .A2(n9882), .ZN(n9944) );
  NAND2_X1 U11772 ( .A1(n10406), .A2(n10401), .ZN(n10132) );
  OAI21_X1 U11773 ( .B1(n10958), .B2(n9984), .A(n9983), .ZN(n10960) );
  NAND2_X1 U11774 ( .A1(n10577), .A2(n16509), .ZN(n9983) );
  OR2_X1 U11775 ( .A1(n10975), .A2(n16509), .ZN(n9984) );
  NOR2_X1 U11776 ( .A1(n15922), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11606) );
  OR2_X1 U11777 ( .A1(n11400), .A2(n17011), .ZN(n10200) );
  NAND2_X1 U11778 ( .A1(n18934), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11401) );
  NAND2_X1 U11779 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11534), .ZN(
        n11400) );
  OR2_X1 U11780 ( .A1(n17011), .A2(n11402), .ZN(n10220) );
  OR2_X1 U11781 ( .A1(n11446), .A2(n11445), .ZN(n11451) );
  NOR2_X1 U11782 ( .A1(n17885), .A2(n11504), .ZN(n11505) );
  NOR2_X1 U11783 ( .A1(n17624), .A2(n11519), .ZN(n11520) );
  OR2_X1 U11784 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  INV_X1 U11785 ( .A(n9867), .ZN(n10101) );
  OR2_X1 U11786 ( .A1(n17670), .A2(n10103), .ZN(n10098) );
  NAND2_X1 U11787 ( .A1(n10100), .A2(n10102), .ZN(n10099) );
  INV_X1 U11788 ( .A(n17700), .ZN(n10100) );
  NOR2_X1 U11789 ( .A1(n18321), .A2(n18343), .ZN(n11638) );
  XNOR2_X1 U11790 ( .A(n10076), .B(n11646), .ZN(n11490) );
  AOI21_X1 U11791 ( .B1(n18747), .B2(n9858), .A(n15919), .ZN(n16011) );
  NAND2_X1 U11793 ( .A1(n14196), .A2(n14195), .ZN(n14636) );
  AOI21_X1 U11794 ( .B1(n14678), .B2(n9818), .A(n12854), .ZN(n13798) );
  AND2_X1 U11795 ( .A1(n12858), .A2(n12857), .ZN(n13797) );
  INV_X1 U11796 ( .A(n10007), .ZN(n10006) );
  NAND2_X1 U11797 ( .A1(n16121), .A2(n9893), .ZN(n10126) );
  CLKBUF_X1 U11798 ( .A(n14591), .Z(n14592) );
  AND2_X1 U11799 ( .A1(n14850), .A2(n14851), .ZN(n14852) );
  AOI21_X1 U11800 ( .B1(n12046), .B2(n12247), .A(n12045), .ZN(n14139) );
  INV_X1 U11801 ( .A(n12044), .ZN(n12045) );
  INV_X1 U11802 ( .A(n12714), .ZN(n12046) );
  NAND2_X1 U11803 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12013) );
  NAND2_X1 U11804 ( .A1(n13789), .A2(n11987), .ZN(n13922) );
  NAND2_X1 U11805 ( .A1(n9818), .A2(n14303), .ZN(n14304) );
  NOR2_X1 U11806 ( .A1(n14494), .A2(n14485), .ZN(n14487) );
  NAND2_X1 U11807 ( .A1(n9906), .A2(n9905), .ZN(n14494) );
  INV_X1 U11808 ( .A(n14492), .ZN(n9905) );
  NOR2_X2 U11809 ( .A1(n14720), .A2(n12938), .ZN(n14706) );
  OR2_X1 U11810 ( .A1(n16068), .A2(n9907), .ZN(n15014) );
  NAND2_X1 U11811 ( .A1(n9909), .A2(n9908), .ZN(n9907) );
  INV_X1 U11812 ( .A(n15013), .ZN(n9908) );
  INV_X1 U11813 ( .A(n16069), .ZN(n9909) );
  NAND2_X1 U11814 ( .A1(n14640), .A2(n14639), .ZN(n16068) );
  AOI21_X1 U11815 ( .B1(n10129), .B2(n16145), .A(n9870), .ZN(n10127) );
  INV_X1 U11816 ( .A(n16144), .ZN(n10131) );
  NAND2_X1 U11817 ( .A1(n20171), .A2(n12721), .ZN(n16158) );
  NAND2_X1 U11818 ( .A1(n16158), .A2(n16157), .ZN(n16156) );
  INV_X1 U11819 ( .A(n20226), .ZN(n20205) );
  AOI21_X1 U11820 ( .B1(n12688), .B2(n12758), .A(n20241), .ZN(n10121) );
  CLKBUF_X1 U11821 ( .A(n12831), .Z(n12832) );
  AND2_X1 U11823 ( .A1(n13831), .A2(n20349), .ZN(n20785) );
  AND2_X1 U11824 ( .A1(n13831), .A2(n12686), .ZN(n20650) );
  INV_X1 U11825 ( .A(n20759), .ZN(n20823) );
  AND2_X1 U11826 ( .A1(n11330), .A2(n11327), .ZN(n13430) );
  OR2_X1 U11827 ( .A1(n16381), .A2(n19192), .ZN(n9975) );
  AND2_X1 U11828 ( .A1(n9975), .A2(n9974), .ZN(n16370) );
  INV_X1 U11829 ( .A(n16372), .ZN(n9974) );
  NOR2_X1 U11830 ( .A1(n16382), .A2(n16383), .ZN(n16381) );
  NOR2_X1 U11831 ( .A1(n10020), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10019) );
  INV_X1 U11832 ( .A(n10021), .ZN(n10020) );
  AND2_X1 U11833 ( .A1(n11255), .A2(n11272), .ZN(n11271) );
  NOR2_X1 U11834 ( .A1(n10022), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10021) );
  NAND2_X1 U11835 ( .A1(n11301), .A2(n11321), .ZN(n11282) );
  OR2_X1 U11836 ( .A1(n14349), .A2(n16491), .ZN(n10484) );
  AND2_X1 U11837 ( .A1(n10480), .A2(n10479), .ZN(n13906) );
  OR2_X1 U11838 ( .A1(n14349), .A2(n16481), .ZN(n10480) );
  NOR2_X1 U11839 ( .A1(n13084), .A2(n13810), .ZN(n13085) );
  AND2_X1 U11840 ( .A1(n13302), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13746) );
  NAND2_X1 U11841 ( .A1(n10064), .A2(n13348), .ZN(n10061) );
  NOR2_X1 U11842 ( .A1(n15116), .A2(n15115), .ZN(n15114) );
  OAI21_X1 U11843 ( .B1(n15138), .B2(n10068), .A(n10067), .ZN(n15129) );
  NAND2_X1 U11844 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  INV_X1 U11845 ( .A(n15140), .ZN(n10069) );
  NOR2_X1 U11846 ( .A1(n15138), .A2(n15140), .ZN(n15139) );
  INV_X1 U11847 ( .A(n13202), .ZN(n15145) );
  NAND2_X1 U11848 ( .A1(n10234), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10236) );
  NAND2_X1 U11849 ( .A1(n10264), .A2(n9836), .ZN(n10239) );
  NAND2_X1 U11850 ( .A1(n10496), .A2(n13450), .ZN(n14245) );
  INV_X1 U11851 ( .A(n13451), .ZN(n10496) );
  NOR2_X1 U11852 ( .A1(n10254), .A2(n16461), .ZN(n10255) );
  XNOR2_X1 U11853 ( .A(n9852), .B(n14362), .ZN(n16334) );
  NOR2_X2 U11854 ( .A1(n15297), .A2(n15299), .ZN(n15298) );
  NAND2_X1 U11855 ( .A1(n13430), .A2(n10137), .ZN(n14378) );
  NOR2_X1 U11856 ( .A1(n11336), .A2(n15327), .ZN(n15323) );
  NAND2_X1 U11857 ( .A1(n15333), .A2(n11368), .ZN(n9939) );
  OAI21_X1 U11858 ( .B1(n15333), .B2(n11368), .A(n15334), .ZN(n9940) );
  INV_X1 U11859 ( .A(n9952), .ZN(n9951) );
  AOI21_X1 U11860 ( .B1(n10203), .B2(n9954), .A(n10211), .ZN(n9952) );
  NAND2_X1 U11861 ( .A1(n10049), .A2(n10868), .ZN(n10048) );
  AND2_X1 U11862 ( .A1(n15704), .A2(n11361), .ZN(n16467) );
  AND2_X1 U11863 ( .A1(n11224), .A2(n15460), .ZN(n10156) );
  AND2_X1 U11864 ( .A1(n10190), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10189) );
  NAND2_X1 U11865 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  AND2_X1 U11866 ( .A1(n10468), .A2(n10463), .ZN(n10009) );
  INV_X1 U11867 ( .A(n13749), .ZN(n10468) );
  NAND2_X1 U11868 ( .A1(n11200), .A2(n10459), .ZN(n9945) );
  NOR2_X1 U11869 ( .A1(n11200), .A2(n10459), .ZN(n9946) );
  XNOR2_X1 U11870 ( .A(n15775), .B(n13060), .ZN(n13558) );
  AOI21_X1 U11871 ( .B1(n15764), .B2(n13059), .A(n13058), .ZN(n13557) );
  OR2_X1 U11872 ( .A1(n19944), .A2(n19971), .ZN(n19744) );
  NAND2_X1 U11873 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19738), .ZN(n19367) );
  INV_X1 U11874 ( .A(n19738), .ZN(n19784) );
  INV_X1 U11875 ( .A(n11638), .ZN(n12991) );
  NAND3_X1 U11876 ( .A1(n18315), .A2(n18336), .A3(n18326), .ZN(n11631) );
  NOR2_X1 U11877 ( .A1(n16713), .A2(n9920), .ZN(n16705) );
  NAND2_X1 U11878 ( .A1(n16670), .A2(n9886), .ZN(n9913) );
  NOR2_X1 U11879 ( .A1(n11435), .A2(n11434), .ZN(n11441) );
  NAND2_X1 U11880 ( .A1(n17638), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13419) );
  NOR2_X2 U11881 ( .A1(n17749), .A2(n17750), .ZN(n17724) );
  OR2_X1 U11882 ( .A1(n17468), .A2(n11499), .ZN(n11500) );
  NAND2_X1 U11883 ( .A1(n10095), .A2(n10094), .ZN(n17636) );
  NAND2_X1 U11884 ( .A1(n10105), .A2(n10096), .ZN(n10095) );
  OR2_X1 U11885 ( .A1(n17670), .A2(n10103), .ZN(n10094) );
  NOR2_X1 U11886 ( .A1(n17700), .A2(n10103), .ZN(n10096) );
  AOI21_X1 U11887 ( .B1(n11515), .B2(n17650), .A(n11512), .ZN(n11513) );
  NAND2_X1 U11888 ( .A1(n17670), .A2(n10104), .ZN(n10107) );
  AOI211_X1 U11889 ( .C1(n17759), .C2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11510), .B(n17758), .ZN(n17754) );
  NOR2_X1 U11890 ( .A1(n11507), .A2(n17873), .ZN(n17834) );
  INV_X1 U11891 ( .A(n17461), .ZN(n16534) );
  NOR2_X1 U11892 ( .A1(n17890), .A2(n10112), .ZN(n10111) );
  INV_X1 U11893 ( .A(n10114), .ZN(n10112) );
  NAND2_X1 U11894 ( .A1(n17904), .A2(n10115), .ZN(n10114) );
  OAI21_X1 U11895 ( .B1(n17930), .B2(n10087), .A(n10086), .ZN(n17919) );
  NAND2_X1 U11896 ( .A1(n10090), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10087) );
  NAND2_X1 U11897 ( .A1(n11495), .A2(n10090), .ZN(n10086) );
  OR2_X1 U11898 ( .A1(n17930), .A2(n18246), .ZN(n10089) );
  OR3_X2 U11899 ( .A1(n11642), .A2(n11635), .A3(n11639), .ZN(n18747) );
  XNOR2_X1 U11900 ( .A(n12621), .B(n12620), .ZN(n14215) );
  XNOR2_X1 U11901 ( .A(n12795), .B(n12794), .ZN(n14313) );
  INV_X1 U11902 ( .A(n16291), .ZN(n20243) );
  OR2_X1 U11903 ( .A1(n16336), .A2(n19209), .ZN(n10033) );
  NOR2_X1 U11904 ( .A1(n11028), .A2(n19209), .ZN(n10940) );
  INV_X1 U11905 ( .A(n19178), .ZN(n19213) );
  INV_X1 U11906 ( .A(n16334), .ZN(n19217) );
  AND2_X1 U11907 ( .A1(n9852), .A2(n10897), .ZN(n13374) );
  AND2_X1 U11908 ( .A1(n19249), .A2(n13390), .ZN(n19221) );
  AND2_X1 U11909 ( .A1(n13372), .A2(n16503), .ZN(n19249) );
  NOR2_X1 U11910 ( .A1(n10181), .A2(n10433), .ZN(n13370) );
  AND2_X1 U11911 ( .A1(n16462), .A2(n19960), .ZN(n19302) );
  NAND2_X1 U11912 ( .A1(n14390), .A2(n15297), .ZN(n14402) );
  OR2_X1 U11913 ( .A1(n15102), .A2(n14384), .ZN(n16358) );
  INV_X1 U11914 ( .A(n19963), .ZN(n19961) );
  INV_X1 U11915 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20000) );
  OR2_X1 U11916 ( .A1(n19953), .A2(n19961), .ZN(n19937) );
  NAND2_X1 U11917 ( .A1(n14093), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16508) );
  NAND2_X1 U11918 ( .A1(n13722), .A2(n13725), .ZN(n19944) );
  OR2_X1 U11919 ( .A1(n13724), .A2(n13723), .ZN(n13725) );
  INV_X1 U11920 ( .A(n16686), .ZN(n9924) );
  NAND2_X1 U11921 ( .A1(n16699), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n9923) );
  XNOR2_X1 U11922 ( .A(n16683), .B(n9926), .ZN(n9925) );
  INV_X1 U11923 ( .A(n16684), .ZN(n9926) );
  INV_X1 U11924 ( .A(n9918), .ZN(n16724) );
  OR2_X1 U11925 ( .A1(n16733), .A2(n9920), .ZN(n9918) );
  NOR2_X1 U11926 ( .A1(n16762), .A2(n9920), .ZN(n16756) );
  NAND2_X1 U11927 ( .A1(n17426), .A2(n9840), .ZN(n17418) );
  NOR2_X1 U11928 ( .A1(n11408), .A2(n11407), .ZN(n17465) );
  NAND2_X1 U11929 ( .A1(n17488), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17486) );
  NOR2_X1 U11930 ( .A1(n16012), .A2(n17561), .ZN(n17488) );
  INV_X1 U11931 ( .A(n17480), .ZN(n17484) );
  NAND2_X1 U11932 ( .A1(n17607), .A2(n17608), .ZN(n17606) );
  NOR2_X2 U11933 ( .A1(n17461), .A2(n17964), .ZN(n17874) );
  AND2_X1 U11934 ( .A1(n10083), .A2(n10078), .ZN(n13025) );
  NAND2_X1 U11935 ( .A1(n12985), .A2(n12986), .ZN(n10083) );
  NAND2_X1 U11936 ( .A1(n10082), .A2(n10079), .ZN(n10078) );
  XNOR2_X1 U11937 ( .A(n11522), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15987) );
  NAND2_X1 U11938 ( .A1(n16550), .A2(n16549), .ZN(n16554) );
  AOI21_X1 U11939 ( .B1(n16548), .B2(n16547), .A(n16546), .ZN(n16550) );
  NAND2_X1 U11940 ( .A1(n10202), .A2(n17601), .ZN(n16552) );
  NAND2_X1 U11941 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13195) );
  AND2_X1 U11942 ( .A1(n11128), .A2(n11119), .ZN(n10147) );
  AND2_X1 U11943 ( .A1(n11127), .A2(n11129), .ZN(n10148) );
  AOI22_X1 U11944 ( .A1(n11112), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n19338), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U11945 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11121), .B1(
        n11126), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U11946 ( .A1(n11122), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11123), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U11947 ( .A1(n11111), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n19338), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U11948 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11125), .B1(
        n11116), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U11949 ( .A1(n19375), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11124), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11081) );
  AND2_X1 U11950 ( .A1(n11821), .A2(n11826), .ZN(n11782) );
  AND2_X1 U11951 ( .A1(n10172), .A2(n12164), .ZN(n10171) );
  OR2_X1 U11952 ( .A1(n12033), .A2(n12032), .ZN(n12723) );
  OR3_X1 U11953 ( .A1(n12658), .A2(n12657), .A3(n12816), .ZN(n12659) );
  INV_X1 U11955 ( .A(n11694), .ZN(n11707) );
  AND2_X1 U11956 ( .A1(n13684), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U11957 ( .A1(n10568), .A2(n10573), .ZN(n10580) );
  AND2_X1 U11958 ( .A1(n10566), .A2(n10565), .ZN(n10576) );
  OR2_X1 U11959 ( .A1(n10970), .A2(n10947), .ZN(n10566) );
  INV_X1 U11960 ( .A(n11090), .ZN(n10151) );
  NOR2_X1 U11961 ( .A1(n11089), .A2(n10691), .ZN(n9902) );
  INV_X1 U11962 ( .A(n15689), .ZN(n10155) );
  INV_X1 U11963 ( .A(n11151), .ZN(n9900) );
  OAI22_X1 U11964 ( .A1(n10810), .A2(n10606), .B1(n10605), .B2(n10604), .ZN(
        n10607) );
  AND2_X1 U11965 ( .A1(n10991), .A2(n13564), .ZN(n10323) );
  NAND2_X1 U11966 ( .A1(n16981), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11399) );
  NOR2_X1 U11967 ( .A1(n11398), .A2(n11399), .ZN(n11436) );
  NAND2_X1 U11968 ( .A1(n18918), .A2(n11534), .ZN(n11397) );
  OR2_X1 U11969 ( .A1(n11842), .A2(n11841), .ZN(n11843) );
  INV_X1 U11970 ( .A(n14467), .ZN(n10178) );
  NOR2_X1 U11971 ( .A1(n10173), .A2(n14635), .ZN(n10172) );
  INV_X1 U11972 ( .A(n14238), .ZN(n10173) );
  AND2_X1 U11973 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n12085), .ZN(
        n12097) );
  NOR2_X1 U11974 ( .A1(n12066), .A2(n20073), .ZN(n12085) );
  AND2_X1 U11975 ( .A1(n11829), .A2(n11840), .ZN(n12952) );
  NAND2_X1 U11976 ( .A1(n12782), .A2(n14921), .ZN(n14911) );
  INV_X1 U11977 ( .A(n12756), .ZN(n10130) );
  NOR2_X1 U11978 ( .A1(n12093), .A2(n12063), .ZN(n10005) );
  INV_X1 U11979 ( .A(n14301), .ZN(n12875) );
  OAI21_X1 U11980 ( .B1(n12692), .B2(n20982), .A(n10001), .ZN(n12693) );
  AND2_X1 U11981 ( .A1(n12691), .A2(n9803), .ZN(n10001) );
  NAND2_X1 U11982 ( .A1(n11827), .A2(n11826), .ZN(n12825) );
  NOR2_X1 U11983 ( .A1(n11961), .A2(n11960), .ZN(n12706) );
  NOR2_X1 U11984 ( .A1(n12661), .A2(n12758), .ZN(n12663) );
  AND2_X1 U11985 ( .A1(n12633), .A2(n12664), .ZN(n12820) );
  NOR2_X1 U11986 ( .A1(n12622), .A2(n11828), .ZN(n11820) );
  AOI22_X1 U11987 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12001), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U11988 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U11990 ( .A1(n20549), .A2(n20885), .ZN(n12010) );
  INV_X1 U11991 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20693) );
  OAI21_X1 U11992 ( .B1(n20983), .B2(n16324), .A(n15967), .ZN(n20260) );
  NAND2_X1 U11993 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19976), .ZN(
        n10947) );
  OR2_X1 U11994 ( .A1(n10601), .A2(n10600), .ZN(n10910) );
  AND2_X1 U11995 ( .A1(n14329), .A2(n10029), .ZN(n10028) );
  INV_X1 U11996 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U11997 ( .A1(n11305), .A2(n11304), .ZN(n11303) );
  NAND2_X1 U11998 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9963) );
  NOR2_X1 U11999 ( .A1(n10024), .A2(n11259), .ZN(n10023) );
  INV_X1 U12000 ( .A(n10026), .ZN(n10024) );
  OR2_X1 U12001 ( .A1(n11180), .A2(n11209), .ZN(n11219) );
  NAND2_X1 U12002 ( .A1(n10695), .A2(n13916), .ZN(n10037) );
  OR2_X1 U12003 ( .A1(n10705), .A2(n10704), .ZN(n10915) );
  NAND2_X1 U12004 ( .A1(n10906), .A2(n10905), .ZN(n11184) );
  NAND2_X1 U12005 ( .A1(n10912), .A2(n10911), .ZN(n11203) );
  INV_X1 U12006 ( .A(n11184), .ZN(n10912) );
  INV_X1 U12007 ( .A(n11196), .ZN(n10911) );
  OR2_X1 U12008 ( .A1(n10588), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10811) );
  NAND2_X1 U12009 ( .A1(n10587), .A2(n10355), .ZN(n10810) );
  NAND2_X1 U12010 ( .A1(n13256), .A2(n13255), .ZN(n10056) );
  INV_X1 U12011 ( .A(n13253), .ZN(n13256) );
  INV_X1 U12012 ( .A(n15130), .ZN(n10070) );
  INV_X1 U12013 ( .A(n15065), .ZN(n10052) );
  OR2_X1 U12014 ( .A1(n19990), .A2(n14103), .ZN(n10404) );
  NAND2_X1 U12015 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9971) );
  NOR2_X1 U12016 ( .A1(n15347), .A2(n9965), .ZN(n9964) );
  NOR3_X1 U12017 ( .A1(n10260), .A2(n19021), .A3(n9963), .ZN(n10242) );
  NOR2_X1 U12018 ( .A1(n9967), .A2(n15463), .ZN(n9966) );
  INV_X1 U12019 ( .A(n9969), .ZN(n9967) );
  NOR2_X1 U12020 ( .A1(n15473), .A2(n9970), .ZN(n9969) );
  INV_X1 U12021 ( .A(n10251), .ZN(n9968) );
  NAND2_X1 U12022 ( .A1(n10418), .A2(n10417), .ZN(n11035) );
  INV_X1 U12023 ( .A(n10418), .ZN(n10416) );
  OR2_X1 U12024 ( .A1(n11094), .A2(n10904), .ZN(n10908) );
  NAND2_X1 U12025 ( .A1(n14374), .A2(n9959), .ZN(n9958) );
  INV_X1 U12026 ( .A(n15502), .ZN(n10193) );
  AND2_X1 U12027 ( .A1(n16377), .A2(n10137), .ZN(n11335) );
  NOR2_X1 U12028 ( .A1(n15081), .A2(n10054), .ZN(n10053) );
  INV_X1 U12029 ( .A(n15570), .ZN(n10054) );
  AND2_X1 U12030 ( .A1(n16437), .A2(n16439), .ZN(n11173) );
  NAND2_X1 U12031 ( .A1(n11179), .A2(n11169), .ZN(n10142) );
  NOR2_X1 U12032 ( .A1(n10718), .A2(n10717), .ZN(n11147) );
  NAND2_X1 U12033 ( .A1(n9935), .A2(n11074), .ZN(n11089) );
  NOR2_X1 U12034 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  INV_X1 U12035 ( .A(n11088), .ZN(n9932) );
  INV_X1 U12036 ( .A(n11074), .ZN(n9933) );
  NAND2_X1 U12037 ( .A1(n9950), .A2(n11349), .ZN(n9949) );
  OAI21_X1 U12038 ( .B1(n10655), .B2(n10439), .A(n10629), .ZN(n10651) );
  INV_X1 U12039 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10272) );
  INV_X1 U12040 ( .A(n11065), .ZN(n9903) );
  NAND3_X1 U12041 ( .A1(n19942), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19738), 
        .ZN(n14105) );
  AND2_X1 U12042 ( .A1(n19355), .A2(n13564), .ZN(n10394) );
  NAND2_X1 U12043 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18918), .ZN(
        n11398) );
  NAND2_X1 U12044 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11431) );
  NOR2_X1 U12045 ( .A1(n18778), .A2(n11400), .ZN(n11479) );
  NOR2_X1 U12046 ( .A1(n17011), .A2(n11397), .ZN(n11478) );
  INV_X1 U12047 ( .A(n17759), .ZN(n11515) );
  CLKBUF_X1 U12048 ( .A(n11682), .Z(n16536) );
  AND2_X1 U12049 ( .A1(n11508), .A2(n10092), .ZN(n10091) );
  INV_X1 U12050 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10092) );
  INV_X1 U12051 ( .A(n16653), .ZN(n12998) );
  NAND2_X1 U12052 ( .A1(n10110), .A2(n10108), .ZN(n11503) );
  NAND2_X1 U12053 ( .A1(n10109), .A2(n9851), .ZN(n10108) );
  NOR2_X1 U12054 ( .A1(n11664), .A2(n17906), .ZN(n11666) );
  NAND2_X1 U12055 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U12056 ( .A1(n11933), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9998) );
  OR2_X1 U12057 ( .A1(n13637), .A2(n14128), .ZN(n13735) );
  AOI22_X1 U12058 ( .A1(n14490), .A2(n14192), .B1(n12546), .B2(n12545), .ZN(
        n13045) );
  AOI21_X1 U12059 ( .B1(n14459), .B2(n14192), .A(n12613), .ZN(n12804) );
  INV_X1 U12060 ( .A(n12547), .ZN(n12549) );
  OR2_X1 U12061 ( .A1(n12549), .A2(n12548), .ZN(n12619) );
  NOR2_X1 U12062 ( .A1(n10177), .A2(n10175), .ZN(n10174) );
  INV_X1 U12063 ( .A(n14508), .ZN(n10175) );
  NAND2_X1 U12064 ( .A1(n10179), .A2(n10178), .ZN(n10177) );
  INV_X1 U12065 ( .A(n10179), .ZN(n10176) );
  NAND2_X1 U12066 ( .A1(n12501), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12526) );
  NOR2_X1 U12067 ( .A1(n12453), .A2(n12435), .ZN(n12454) );
  NAND2_X1 U12068 ( .A1(n12454), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12479) );
  NOR2_X1 U12069 ( .A1(n12440), .A2(n12439), .ZN(n12449) );
  NAND2_X1 U12070 ( .A1(n12449), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12453) );
  NOR2_X1 U12071 ( .A1(n12369), .A2(n14914), .ZN(n12370) );
  AND2_X1 U12072 ( .A1(n10164), .A2(n14726), .ZN(n10163) );
  AND2_X1 U12073 ( .A1(n12330), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12331) );
  NAND2_X1 U12074 ( .A1(n12331), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12369) );
  NOR2_X1 U12075 ( .A1(n12294), .A2(n16044), .ZN(n12330) );
  NAND2_X1 U12076 ( .A1(n14928), .A2(n14931), .ZN(n12777) );
  NOR2_X1 U12077 ( .A1(n12780), .A2(n14941), .ZN(n16110) );
  NAND2_X1 U12078 ( .A1(n12214), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12215) );
  NOR2_X1 U12079 ( .A1(n21015), .A2(n12215), .ZN(n12273) );
  NOR2_X1 U12080 ( .A1(n12210), .A2(n16061), .ZN(n12214) );
  AND2_X1 U12081 ( .A1(n12158), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12159) );
  NAND2_X1 U12082 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n12159), .ZN(
        n12210) );
  AOI21_X1 U12083 ( .B1(n12732), .B2(n12247), .A(n12089), .ZN(n14234) );
  INV_X1 U12084 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20073) );
  NOR2_X1 U12085 ( .A1(n12013), .A2(n12012), .ZN(n12039) );
  AND2_X1 U12086 ( .A1(n13783), .A2(n11987), .ZN(n10162) );
  AND2_X1 U12087 ( .A1(n16134), .A2(n14885), .ZN(n10008) );
  INV_X1 U12088 ( .A(n9906), .ZN(n14517) );
  NAND2_X1 U12089 ( .A1(n9818), .A2(n14721), .ZN(n12934) );
  OAI21_X1 U12090 ( .B1(n9776), .B2(n12784), .A(n16121), .ZN(n14902) );
  NAND2_X1 U12091 ( .A1(n14757), .A2(n9868), .ZN(n14746) );
  INV_X1 U12092 ( .A(n14595), .ZN(n9904) );
  NAND2_X1 U12093 ( .A1(n14757), .A2(n14756), .ZN(n14759) );
  AND2_X1 U12094 ( .A1(n12899), .A2(n12898), .ZN(n16069) );
  AND2_X1 U12096 ( .A1(n16121), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12769) );
  NAND2_X1 U12097 ( .A1(n12889), .A2(n12888), .ZN(n14241) );
  OAI21_X1 U12098 ( .B1(n16158), .B2(n10118), .A(n10117), .ZN(n12741) );
  AND2_X1 U12099 ( .A1(n20087), .A2(n20085), .ZN(n12869) );
  AND2_X1 U12100 ( .A1(n12963), .A2(n12960), .ZN(n14277) );
  AND2_X1 U12101 ( .A1(n12963), .A2(n12947), .ZN(n20226) );
  AND3_X1 U12102 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20885), .A3(n20260), 
        .ZN(n20312) );
  INV_X1 U12103 ( .A(n20822), .ZN(n20829) );
  AND2_X1 U12104 ( .A1(n20884), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15963) );
  NAND2_X1 U12105 ( .A1(n10944), .A2(n9980), .ZN(n10974) );
  INV_X1 U12106 ( .A(n10943), .ZN(n9980) );
  OR2_X1 U12107 ( .A1(n16349), .A2(n10206), .ZN(n9976) );
  AND2_X1 U12108 ( .A1(n11340), .A2(n11331), .ZN(n16350) );
  OR2_X1 U12109 ( .A1(n13429), .A2(n15309), .ZN(n9978) );
  NOR2_X1 U12110 ( .A1(n16370), .A2(n19192), .ZN(n16360) );
  NOR2_X1 U12111 ( .A1(n16361), .A2(n16360), .ZN(n16359) );
  AND2_X1 U12112 ( .A1(n11303), .A2(n15136), .ZN(n11323) );
  NOR2_X1 U12113 ( .A1(n19192), .A2(n10265), .ZN(n15044) );
  AND2_X1 U12114 ( .A1(n15058), .A2(n15362), .ZN(n10265) );
  NAND2_X1 U12115 ( .A1(n11282), .A2(n11299), .ZN(n11305) );
  CLKBUF_X1 U12116 ( .A(n10242), .Z(n10263) );
  NAND2_X1 U12117 ( .A1(n10921), .A2(n10214), .ZN(n11257) );
  INV_X1 U12118 ( .A(n11266), .ZN(n10921) );
  NAND2_X1 U12119 ( .A1(n10025), .A2(n10026), .ZN(n11261) );
  NAND2_X1 U12120 ( .A1(n11232), .A2(n19111), .ZN(n11238) );
  INV_X1 U12121 ( .A(n11214), .ZN(n10018) );
  INV_X1 U12122 ( .A(n11202), .ZN(n10914) );
  INV_X1 U12123 ( .A(n10969), .ZN(n10989) );
  NAND2_X1 U12124 ( .A1(n10515), .A2(n9833), .ZN(n15190) );
  NAND2_X1 U12125 ( .A1(n10515), .A2(n10514), .ZN(n15201) );
  NOR2_X1 U12126 ( .A1(n15211), .A2(n15197), .ZN(n15192) );
  INV_X1 U12127 ( .A(n14167), .ZN(n10073) );
  OR2_X1 U12128 ( .A1(n14349), .A2(n15727), .ZN(n10476) );
  OAI22_X1 U12129 ( .A1(n10451), .A2(n10435), .B1(n10455), .B2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U12130 ( .A1(n10431), .A2(n10430), .ZN(n11042) );
  NAND2_X1 U12131 ( .A1(n10508), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10430) );
  NOR2_X1 U12132 ( .A1(n13436), .A2(n9879), .ZN(n14413) );
  OR2_X1 U12133 ( .A1(n13349), .A2(n10059), .ZN(n10058) );
  INV_X1 U12134 ( .A(n15115), .ZN(n10059) );
  INV_X1 U12135 ( .A(n15110), .ZN(n10065) );
  NAND2_X1 U12136 ( .A1(n15109), .A2(n13307), .ZN(n15116) );
  XNOR2_X1 U12137 ( .A(n13276), .B(n10219), .ZN(n15122) );
  XNOR2_X1 U12138 ( .A(n13253), .B(n13255), .ZN(n14316) );
  AND2_X1 U12139 ( .A1(n15262), .A2(n9884), .ZN(n15067) );
  INV_X1 U12140 ( .A(n13445), .ZN(n10047) );
  NAND2_X1 U12141 ( .A1(n9892), .A2(n10695), .ZN(n10035) );
  AND2_X1 U12142 ( .A1(n13599), .A2(n19989), .ZN(n19250) );
  NAND2_X1 U12143 ( .A1(n10264), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10266) );
  AND2_X1 U12144 ( .A1(n10240), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10264) );
  NAND2_X1 U12145 ( .A1(n10246), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10260) );
  NOR2_X1 U12146 ( .A1(n15611), .A2(n15633), .ZN(n10187) );
  NAND2_X1 U12147 ( .A1(n10259), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10258) );
  NOR2_X1 U12148 ( .A1(n10247), .A2(n15452), .ZN(n10259) );
  CLKBUF_X1 U12149 ( .A(n10247), .Z(n10257) );
  AND2_X1 U12150 ( .A1(n13960), .A2(n13959), .ZN(n13967) );
  NOR2_X1 U12151 ( .A1(n10251), .A2(n15473), .ZN(n10256) );
  INV_X1 U12152 ( .A(n15743), .ZN(n15746) );
  NAND2_X1 U12153 ( .A1(n9962), .A2(n9828), .ZN(n10254) );
  INV_X1 U12154 ( .A(n10252), .ZN(n9962) );
  INV_X1 U12155 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14185) );
  AOI21_X1 U12156 ( .B1(n11343), .B2(n9959), .A(n11342), .ZN(n10144) );
  OR3_X1 U12157 ( .A1(n11345), .A2(n11169), .A3(n11374), .ZN(n14334) );
  NOR2_X2 U12158 ( .A1(n9841), .A2(n14383), .ZN(n15102) );
  INV_X1 U12159 ( .A(n14378), .ZN(n14376) );
  NAND2_X1 U12160 ( .A1(n15526), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15517) );
  OR2_X1 U12161 ( .A1(n11335), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15322) );
  NAND2_X1 U12162 ( .A1(n10218), .A2(n9887), .ZN(n15134) );
  INV_X1 U12163 ( .A(n15048), .ZN(n10011) );
  OR2_X1 U12164 ( .A1(n15056), .A2(n11169), .ZN(n11307) );
  NAND2_X1 U12165 ( .A1(n9987), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15547) );
  AND2_X1 U12166 ( .A1(n10218), .A2(n15077), .ZN(n15079) );
  NAND2_X1 U12167 ( .A1(n15262), .A2(n10053), .ZN(n15083) );
  AND2_X1 U12168 ( .A1(n10529), .A2(n10528), .ZN(n15155) );
  AND2_X1 U12169 ( .A1(n10515), .A2(n9877), .ZN(n15180) );
  INV_X1 U12170 ( .A(n15179), .ZN(n10013) );
  NAND2_X1 U12171 ( .A1(n15180), .A2(n15173), .ZN(n15175) );
  INV_X1 U12172 ( .A(n15285), .ZN(n10873) );
  AND2_X1 U12173 ( .A1(n11270), .A2(n15369), .ZN(n15428) );
  CLKBUF_X1 U12174 ( .A(n15435), .Z(n15436) );
  NAND2_X1 U12175 ( .A1(n15680), .A2(n11249), .ZN(n9901) );
  AND2_X1 U12176 ( .A1(n10016), .A2(n14083), .ZN(n10015) );
  AND2_X1 U12177 ( .A1(n13960), .A2(n10016), .ZN(n14084) );
  NAND2_X1 U12178 ( .A1(n13689), .A2(n10044), .ZN(n15706) );
  AND2_X1 U12179 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  INV_X1 U12180 ( .A(n15693), .ZN(n10043) );
  AND2_X1 U12181 ( .A1(n10136), .A2(n10140), .ZN(n10135) );
  AOI21_X1 U12182 ( .B1(n9944), .B2(n9946), .A(n9942), .ZN(n9941) );
  NOR2_X1 U12183 ( .A1(n11204), .A2(n15750), .ZN(n9942) );
  NAND2_X1 U12184 ( .A1(n10624), .A2(n10623), .ZN(n13545) );
  NAND2_X1 U12185 ( .A1(n13356), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10965) );
  NOR2_X1 U12186 ( .A1(n13775), .A2(n10661), .ZN(n13929) );
  OR2_X1 U12187 ( .A1(n10960), .A2(n10959), .ZN(n14093) );
  NAND2_X1 U12188 ( .A1(n13665), .A2(n13068), .ZN(n13724) );
  AND3_X1 U12189 ( .A1(n10401), .A2(n10381), .A3(n10903), .ZN(n10382) );
  AOI22_X1 U12190 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10342) );
  INV_X1 U12191 ( .A(n14040), .ZN(n14264) );
  AND2_X1 U12192 ( .A1(n19944), .A2(n19971), .ZN(n19512) );
  AND2_X1 U12193 ( .A1(n19944), .A2(n19212), .ZN(n19546) );
  AND2_X1 U12194 ( .A1(n19953), .A2(n19961), .ZN(n19599) );
  INV_X1 U12195 ( .A(n19730), .ZN(n19745) );
  NOR2_X2 U12196 ( .A1(n14104), .A2(n14105), .ZN(n19366) );
  NOR2_X1 U12197 ( .A1(n19944), .A2(n19212), .ZN(n19694) );
  NAND2_X1 U12198 ( .A1(n10980), .A2(n10989), .ZN(n14070) );
  NOR2_X1 U12199 ( .A1(n9764), .A2(n15916), .ZN(n18748) );
  NOR2_X1 U12200 ( .A1(n16705), .A2(n16706), .ZN(n16704) );
  OAI21_X1 U12201 ( .B1(n16733), .B2(n9920), .A(n9916), .ZN(n13421) );
  NAND2_X1 U12202 ( .A1(n9921), .A2(n16725), .ZN(n9916) );
  NOR2_X1 U12204 ( .A1(n13421), .A2(n17630), .ZN(n16672) );
  OAI21_X1 U12206 ( .B1(n16762), .B2(n9920), .A(n9919), .ZN(n16743) );
  NAND2_X1 U12207 ( .A1(n9921), .A2(n17685), .ZN(n9919) );
  NOR2_X1 U12209 ( .A1(n16743), .A2(n17669), .ZN(n16742) );
  NOR2_X1 U12210 ( .A1(n16781), .A2(n17713), .ZN(n16774) );
  NOR2_X1 U12211 ( .A1(n17595), .A2(n9990), .ZN(n9989) );
  NOR2_X1 U12212 ( .A1(n11451), .A2(n11450), .ZN(n11454) );
  NOR2_X1 U12213 ( .A1(n16014), .A2(n18343), .ZN(n16013) );
  NAND2_X1 U12214 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11484) );
  NAND3_X1 U12215 ( .A1(n11589), .A2(n11588), .A3(n11587), .ZN(n17492) );
  AOI211_X1 U12216 ( .C1(n17289), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n11586), .B(n11585), .ZN(n11587) );
  NAND2_X1 U12217 ( .A1(n16670), .A2(n11677), .ZN(n16673) );
  NAND2_X1 U12218 ( .A1(n13420), .A2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17598) );
  INV_X1 U12220 ( .A(n17683), .ZN(n9927) );
  INV_X1 U12221 ( .A(n13412), .ZN(n13415) );
  NAND2_X1 U12222 ( .A1(n10216), .A2(n17863), .ZN(n17822) );
  NOR2_X1 U12223 ( .A1(n11676), .A2(n17870), .ZN(n17827) );
  INV_X1 U12224 ( .A(n17922), .ZN(n9928) );
  INV_X1 U12226 ( .A(n17960), .ZN(n17921) );
  NAND2_X1 U12227 ( .A1(n12982), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10082) );
  AND2_X1 U12228 ( .A1(n12983), .A2(n10080), .ZN(n10079) );
  NOR2_X1 U12229 ( .A1(n12981), .A2(n10081), .ZN(n10080) );
  INV_X1 U12230 ( .A(n12987), .ZN(n10081) );
  NAND2_X1 U12231 ( .A1(n17873), .A2(n12984), .ZN(n12982) );
  NAND2_X1 U12232 ( .A1(n11521), .A2(n17838), .ZN(n12983) );
  NAND2_X1 U12233 ( .A1(n15925), .A2(n16518), .ZN(n11521) );
  NOR2_X1 U12234 ( .A1(n17974), .A2(n13017), .ZN(n16517) );
  NOR2_X1 U12235 ( .A1(n11520), .A2(n10085), .ZN(n15925) );
  NAND2_X1 U12236 ( .A1(n17622), .A2(n16551), .ZN(n10085) );
  NOR2_X1 U12237 ( .A1(n17647), .A2(n11683), .ZN(n17976) );
  OAI211_X1 U12238 ( .C1(n10104), .C2(n10099), .A(n10098), .B(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U12239 ( .A1(n17625), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17624) );
  OR2_X1 U12240 ( .A1(n18010), .A2(n18007), .ZN(n17647) );
  NOR2_X1 U12241 ( .A1(n17873), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17744) );
  AND2_X1 U12242 ( .A1(n17834), .A2(n9891), .ZN(n17791) );
  NAND2_X1 U12243 ( .A1(n18230), .A2(n12989), .ZN(n15928) );
  OAI21_X1 U12244 ( .B1(n11548), .B2(n11547), .A(n11546), .ZN(n18746) );
  NOR2_X1 U12245 ( .A1(n17908), .A2(n17907), .ZN(n17906) );
  NOR2_X1 U12246 ( .A1(n11661), .A2(n17931), .ZN(n17915) );
  XNOR2_X1 U12247 ( .A(n11490), .B(n18278), .ZN(n17941) );
  XNOR2_X1 U12248 ( .A(n11654), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17953) );
  NAND2_X1 U12249 ( .A1(n18934), .A2(n16981), .ZN(n17011) );
  NAND2_X1 U12250 ( .A1(n18964), .A2(n15883), .ZN(n18781) );
  NAND2_X1 U12251 ( .A1(n10077), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15922) );
  INV_X1 U12252 ( .A(n11402), .ZN(n10077) );
  INV_X1 U12253 ( .A(n17492), .ZN(n18307) );
  NOR2_X2 U12254 ( .A1(n11532), .A2(n11531), .ZN(n18961) );
  NOR2_X1 U12255 ( .A1(n11559), .A2(n11558), .ZN(n18321) );
  INV_X1 U12256 ( .A(n13000), .ZN(n18326) );
  NOR2_X1 U12257 ( .A1(n11569), .A2(n11568), .ZN(n18331) );
  CLKBUF_X1 U12258 ( .A(n13574), .Z(n14104) );
  INV_X1 U12260 ( .A(n20976), .ZN(n14196) );
  NAND2_X1 U12261 ( .A1(n14659), .A2(n14198), .ZN(n20101) );
  AND2_X1 U12262 ( .A1(n14215), .A2(n14214), .ZN(n20039) );
  AND2_X1 U12263 ( .A1(n14636), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20051) );
  AND2_X1 U12264 ( .A1(n20115), .A2(n11828), .ZN(n20112) );
  CLKBUF_X1 U12265 ( .A(n14767), .Z(n14753) );
  INV_X1 U12266 ( .A(n20112), .ZN(n14769) );
  INV_X1 U12267 ( .A(n14782), .ZN(n14838) );
  OR2_X1 U12268 ( .A1(n14847), .A2(n14135), .ZN(n14864) );
  AND2_X1 U12269 ( .A1(n13464), .A2(n15960), .ZN(n20119) );
  BUF_X1 U12270 ( .A(n20140), .Z(n20132) );
  INV_X1 U12271 ( .A(n16016), .ZN(n16085) );
  NAND2_X1 U12272 ( .A1(n14578), .A2(n14579), .ZN(n14562) );
  CLKBUF_X1 U12273 ( .A(n14608), .Z(n14609) );
  AOI21_X1 U12274 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n16128) );
  XOR2_X1 U12275 ( .A(n14858), .B(n14857), .Z(n16139) );
  XNOR2_X1 U12276 ( .A(n14457), .B(n14456), .ZN(n14984) );
  XNOR2_X1 U12277 ( .A(n12803), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14987) );
  NAND2_X1 U12278 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  NAND2_X1 U12279 ( .A1(n12800), .A2(n16134), .ZN(n12801) );
  AND2_X1 U12280 ( .A1(n12972), .A2(n16223), .ZN(n16200) );
  NAND2_X1 U12281 ( .A1(n16143), .A2(n12756), .ZN(n14270) );
  NAND2_X1 U12282 ( .A1(n16156), .A2(n12731), .ZN(n16153) );
  NAND2_X1 U12283 ( .A1(n10120), .A2(n12688), .ZN(n13802) );
  NAND2_X1 U12284 ( .A1(n9790), .A2(n12742), .ZN(n10120) );
  INV_X1 U12285 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20611) );
  INV_X1 U12286 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20652) );
  INV_X1 U12287 ( .A(n15038), .ZN(n15967) );
  NOR2_X1 U12288 ( .A1(n20701), .A2(n13646), .ZN(n15038) );
  CLKBUF_X1 U12289 ( .A(n13616), .Z(n13617) );
  OAI21_X1 U12290 ( .B1(n20449), .B2(n20433), .A(n20794), .ZN(n20452) );
  INV_X1 U12291 ( .A(n20480), .ZN(n20468) );
  NAND2_X1 U12292 ( .A1(n20522), .A2(n20685), .ZN(n20480) );
  OAI211_X1 U12293 ( .C1(n20574), .C2(n20701), .A(n20614), .B(n20558), .ZN(
        n20577) );
  INV_X1 U12294 ( .A(n20571), .ZN(n20576) );
  OR2_X1 U12295 ( .A1(n20656), .A2(n20580), .ZN(n20639) );
  INV_X1 U12296 ( .A(n20619), .ZN(n20646) );
  OR2_X1 U12297 ( .A1(n20656), .A2(n20606), .ZN(n20684) );
  NAND2_X1 U12298 ( .A1(n20312), .A2(n9802), .ZN(n20732) );
  OAI211_X1 U12299 ( .C1(n20811), .C2(n20795), .A(n20794), .B(n20793), .ZN(
        n20814) );
  INV_X1 U12300 ( .A(n20808), .ZN(n20813) );
  INV_X1 U12301 ( .A(n20706), .ZN(n20835) );
  INV_X1 U12302 ( .A(n20713), .ZN(n20841) );
  INV_X1 U12303 ( .A(n20727), .ZN(n20853) );
  INV_X1 U12304 ( .A(n20882), .ZN(n20862) );
  INV_X1 U12305 ( .A(n20732), .ZN(n20859) );
  NAND2_X1 U12306 ( .A1(n20823), .A2(n20650), .ZN(n20882) );
  INV_X1 U12307 ( .A(n20865), .ZN(n20878) );
  INV_X1 U12308 ( .A(n20745), .ZN(n20874) );
  INV_X1 U12309 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20701) );
  INV_X1 U12310 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20885) );
  AND2_X1 U12311 ( .A1(n9976), .A2(n9977), .ZN(n16342) );
  AND2_X1 U12312 ( .A1(n9978), .A2(n9977), .ZN(n16349) );
  INV_X1 U12313 ( .A(n9976), .ZN(n16348) );
  INV_X1 U12314 ( .A(n9978), .ZN(n13428) );
  INV_X1 U12315 ( .A(n9975), .ZN(n16371) );
  AND2_X1 U12316 ( .A1(n11285), .A2(n11284), .ZN(n15086) );
  NAND2_X1 U12317 ( .A1(n11271), .A2(n10021), .ZN(n11283) );
  NAND2_X1 U12318 ( .A1(n10066), .A2(n15110), .ZN(n14411) );
  AND2_X1 U12319 ( .A1(n9832), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U12320 ( .A1(n13747), .A2(n9832), .ZN(n13904) );
  INV_X1 U12321 ( .A(n15178), .ZN(n15212) );
  CLKBUF_X1 U12322 ( .A(n13726), .Z(n13727) );
  AND2_X1 U12323 ( .A1(n15145), .A2(n13203), .ZN(n10071) );
  AND2_X1 U12324 ( .A1(n19249), .A2(n13384), .ZN(n19223) );
  AND2_X1 U12325 ( .A1(n19249), .A2(n13540), .ZN(n19245) );
  INV_X1 U12326 ( .A(n19971), .ZN(n19212) );
  XNOR2_X1 U12328 ( .A(n10227), .B(n10226), .ZN(n14353) );
  NAND2_X1 U12329 ( .A1(n10225), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10227) );
  AND2_X1 U12330 ( .A1(n10187), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10186) );
  INV_X1 U12331 ( .A(n13726), .ZN(n14120) );
  INV_X1 U12332 ( .A(n19302), .ZN(n19289) );
  NAND2_X1 U12333 ( .A1(n18987), .A2(n11381), .ZN(n16462) );
  CLKBUF_X1 U12334 ( .A(n13669), .Z(n13670) );
  INV_X1 U12335 ( .A(n16456), .ZN(n19300) );
  INV_X1 U12336 ( .A(n16453), .ZN(n19294) );
  INV_X1 U12337 ( .A(n16462), .ZN(n19296) );
  AOI21_X1 U12338 ( .B1(n14364), .B2(n9986), .A(n9985), .ZN(n14366) );
  AND2_X1 U12339 ( .A1(n14363), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9986) );
  OAI21_X1 U12340 ( .B1(n16334), .B2(n16466), .A(n14365), .ZN(n9985) );
  NAND2_X1 U12341 ( .A1(n9961), .A2(n14337), .ZN(n14343) );
  OAI21_X1 U12342 ( .B1(n11028), .B2(n19317), .A(n10201), .ZN(n11029) );
  AOI21_X1 U12343 ( .B1(n15299), .B2(n15297), .A(n15298), .ZN(n15478) );
  NAND2_X1 U12344 ( .A1(n9956), .A2(n14374), .ZN(n15295) );
  NAND2_X1 U12345 ( .A1(n10143), .A2(n11334), .ZN(n9956) );
  NOR2_X1 U12346 ( .A1(n15547), .A2(n15535), .ZN(n15526) );
  OR3_X1 U12347 ( .A1(n15546), .A2(n11369), .A3(n11368), .ZN(n15525) );
  CLKBUF_X1 U12348 ( .A(n15355), .Z(n15356) );
  INV_X1 U12349 ( .A(n9987), .ZN(n15558) );
  AND2_X1 U12350 ( .A1(n16467), .A2(n11363), .ZN(n15632) );
  NAND2_X1 U12351 ( .A1(n10157), .A2(n10156), .ZN(n15688) );
  AND2_X1 U12352 ( .A1(n16490), .A2(n11359), .ZN(n15704) );
  NOR2_X1 U12353 ( .A1(n11358), .A2(n16479), .ZN(n15711) );
  NAND2_X1 U12354 ( .A1(n15728), .A2(n9988), .ZN(n16479) );
  INV_X1 U12355 ( .A(n11357), .ZN(n9988) );
  CLKBUF_X1 U12356 ( .A(n15471), .Z(n15472) );
  INV_X1 U12357 ( .A(n15728), .ZN(n15748) );
  NAND2_X1 U12358 ( .A1(n11351), .A2(n11007), .ZN(n19317) );
  NAND2_X1 U12359 ( .A1(n10010), .A2(n10463), .ZN(n13750) );
  OAI21_X1 U12360 ( .B1(n11201), .B2(n9946), .A(n9945), .ZN(n14152) );
  INV_X1 U12361 ( .A(n19319), .ZN(n16496) );
  INV_X1 U12362 ( .A(n16466), .ZN(n19326) );
  AND2_X1 U12363 ( .A1(n11351), .A2(n14041), .ZN(n19314) );
  AND2_X1 U12364 ( .A1(n11351), .A2(n19981), .ZN(n19319) );
  INV_X1 U12365 ( .A(n19314), .ZN(n9979) );
  INV_X1 U12366 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19968) );
  INV_X1 U12367 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19950) );
  NAND2_X1 U12368 ( .A1(n13560), .A2(n13559), .ZN(n19963) );
  NAND2_X1 U12369 ( .A1(n13665), .A2(n13668), .ZN(n19953) );
  OR2_X1 U12370 ( .A1(n13666), .A2(n13667), .ZN(n13668) );
  INV_X1 U12371 ( .A(n19419), .ZN(n19428) );
  OAI21_X1 U12372 ( .B1(n19460), .B2(n19459), .A(n19458), .ZN(n19477) );
  INV_X1 U12373 ( .A(n19517), .ZN(n19566) );
  OAI21_X1 U12374 ( .B1(n19639), .B2(n19654), .A(n19738), .ZN(n19657) );
  INV_X1 U12375 ( .A(n19793), .ZN(n19747) );
  OR3_X1 U12376 ( .A1(n19785), .A2(n19784), .A3(n19783), .ZN(n19810) );
  OAI21_X1 U12377 ( .B1(n19789), .B2(n19788), .A(n19787), .ZN(n19809) );
  INV_X1 U12378 ( .A(n19754), .ZN(n19816) );
  INV_X1 U12379 ( .A(n19676), .ZN(n19822) );
  INV_X1 U12380 ( .A(n19679), .ZN(n19829) );
  INV_X1 U12381 ( .A(n19766), .ZN(n19842) );
  OR3_X1 U12382 ( .A1(n14097), .A2(n14100), .A3(n14096), .ZN(n19849) );
  AND2_X1 U12383 ( .A1(n10968), .A2(n10967), .ZN(n19983) );
  NOR2_X1 U12384 ( .A1(n11635), .A2(n18315), .ZN(n16653) );
  AOI21_X1 U12385 ( .B1(n18748), .B2(n18747), .A(n17530), .ZN(n18976) );
  INV_X1 U12387 ( .A(n17001), .ZN(n17015) );
  INV_X1 U12388 ( .A(n17012), .ZN(n17025) );
  AND3_X1 U12389 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17094), .ZN(n17093) );
  INV_X1 U12390 ( .A(n15888), .ZN(n17337) );
  NOR2_X1 U12391 ( .A1(n17558), .A2(n9845), .ZN(n17348) );
  NOR3_X1 U12392 ( .A1(n17368), .A2(n17552), .A3(n17554), .ZN(n17354) );
  NOR2_X1 U12393 ( .A1(n17368), .A2(n17552), .ZN(n17362) );
  INV_X1 U12394 ( .A(n17372), .ZN(n17369) );
  NAND2_X1 U12395 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17369), .ZN(n17368) );
  NOR2_X1 U12396 ( .A1(n17378), .A2(n17459), .ZN(n17373) );
  NAND2_X1 U12397 ( .A1(n17373), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17372) );
  NOR3_X1 U12398 ( .A1(n17418), .A2(n17545), .A3(n17390), .ZN(n17379) );
  NOR3_X1 U12399 ( .A1(n17454), .A2(n17339), .A3(n17579), .ZN(n17426) );
  NAND2_X1 U12400 ( .A1(n17426), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n17425) );
  NOR2_X1 U12401 ( .A1(n17486), .A2(n9996), .ZN(n17455) );
  NAND2_X1 U12402 ( .A1(n9997), .A2(P3_EAX_REG_2__SCAN_IN), .ZN(n9996) );
  INV_X1 U12403 ( .A(n17460), .ZN(n9997) );
  NAND2_X1 U12404 ( .A1(n17455), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n17454) );
  NOR2_X1 U12405 ( .A1(n11419), .A2(n11418), .ZN(n17468) );
  NOR2_X1 U12406 ( .A1(n17527), .A2(n17509), .ZN(n17519) );
  CLKBUF_X1 U12407 ( .A(n17519), .Z(n17526) );
  CLKBUF_X1 U12408 ( .A(n17592), .Z(n17589) );
  BUF_X1 U12409 ( .A(n17584), .Z(n17591) );
  NOR2_X1 U12410 ( .A1(n18961), .A2(n17591), .ZN(n17592) );
  OAI21_X1 U12411 ( .B1(n16533), .B2(n17838), .A(n17612), .ZN(n17607) );
  NAND2_X1 U12412 ( .A1(n17724), .A2(n10215), .ZN(n17711) );
  NAND2_X1 U12414 ( .A1(n17810), .A2(n10217), .ZN(n17786) );
  INV_X1 U12415 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17865) );
  NOR2_X1 U12416 ( .A1(n17883), .A2(n17865), .ZN(n17861) );
  INV_X1 U12417 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17896) );
  NOR2_X1 U12418 ( .A1(n17922), .A2(n17924), .ZN(n17901) );
  INV_X1 U12419 ( .A(n18411), .ZN(n18692) );
  INV_X1 U12420 ( .A(n17934), .ZN(n17958) );
  NAND2_X1 U12421 ( .A1(n10107), .A2(n17838), .ZN(n17635) );
  NAND2_X1 U12422 ( .A1(n17670), .A2(n11514), .ZN(n17657) );
  NAND2_X1 U12423 ( .A1(n17701), .A2(n13012), .ZN(n17671) );
  NAND2_X1 U12424 ( .A1(n17834), .A2(n9881), .ZN(n17776) );
  NAND2_X1 U12425 ( .A1(n17834), .A2(n11508), .ZN(n17820) );
  INV_X1 U12426 ( .A(n17877), .ZN(n18205) );
  NOR2_X1 U12427 ( .A1(n16534), .A2(n15928), .ZN(n18204) );
  NAND2_X1 U12428 ( .A1(n10113), .A2(n10114), .ZN(n17891) );
  NAND2_X1 U12429 ( .A1(n17903), .A2(n9823), .ZN(n10113) );
  NAND2_X1 U12430 ( .A1(n17903), .A2(n17904), .ZN(n17902) );
  INV_X1 U12431 ( .A(n11495), .ZN(n10088) );
  INV_X1 U12432 ( .A(n10089), .ZN(n17929) );
  INV_X1 U12433 ( .A(n18217), .ZN(n18288) );
  INV_X1 U12434 ( .A(n18224), .ZN(n18294) );
  INV_X1 U12435 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18934) );
  INV_X1 U12436 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18918) );
  AND2_X1 U12437 ( .A1(n13403), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20259)
         );
  CLKBUF_X1 U12438 ( .A(n16638), .Z(n16634) );
  OAI21_X1 U12439 ( .B1(n14313), .B2(n20198), .A(n12796), .ZN(P1_U2968) );
  NAND2_X1 U12440 ( .A1(n12849), .A2(n20243), .ZN(n12980) );
  OAI211_X1 U12441 ( .C1(n9821), .C2(n9883), .A(n9827), .B(n10032), .ZN(
        P2_U2824) );
  NAND2_X1 U12442 ( .A1(n19217), .A2(n19182), .ZN(n10032) );
  NOR2_X1 U12443 ( .A1(n10940), .A2(n10939), .ZN(n10941) );
  AOI21_X1 U12444 ( .B1(n13374), .B2(n13389), .A(n13388), .ZN(n13392) );
  NOR2_X1 U12445 ( .A1(n11387), .A2(n11386), .ZN(n11390) );
  INV_X1 U12446 ( .A(n10184), .ZN(n10183) );
  OAI21_X1 U12447 ( .B1(n14402), .B2(n16456), .A(n10185), .ZN(n10184) );
  AOI21_X1 U12448 ( .B1(n9925), .B2(n16987), .A(n9922), .ZN(n16689) );
  NAND2_X1 U12449 ( .A1(n9924), .A2(n9923), .ZN(n9922) );
  AND2_X1 U12450 ( .A1(n17485), .A2(BUF2_REG_1__SCAN_IN), .ZN(n10075) );
  AOI21_X1 U12451 ( .B1(n13034), .B2(n17950), .A(n13033), .ZN(n13035) );
  NAND2_X1 U12452 ( .A1(n13025), .A2(n17874), .ZN(n13036) );
  NOR2_X1 U12453 ( .A1(n11689), .A2(n11688), .ZN(n11690) );
  AOI21_X1 U12454 ( .B1(n16554), .B2(n16553), .A(n16552), .ZN(n16555) );
  NOR2_X2 U12455 ( .A1(n18778), .A2(n11402), .ZN(n11392) );
  INV_X1 U12456 ( .A(n11477), .ZN(n11466) );
  AND2_X1 U12457 ( .A1(n10156), .A2(n10155), .ZN(n9819) );
  NAND2_X1 U12458 ( .A1(n9804), .A2(n9839), .ZN(n15305) );
  OR2_X1 U12459 ( .A1(n10267), .A2(n10268), .ZN(n9821) );
  NAND2_X1 U12460 ( .A1(n10047), .A2(n10049), .ZN(n14143) );
  OAI21_X1 U12461 ( .B1(n11165), .B2(n11169), .A(n16491), .ZN(n16438) );
  INV_X1 U12462 ( .A(n11479), .ZN(n11602) );
  NAND2_X1 U12463 ( .A1(n15435), .A2(n10187), .ZN(n15422) );
  INV_X2 U12464 ( .A(n20272), .ZN(n11824) );
  INV_X2 U12465 ( .A(n14179), .ZN(n19192) );
  XNOR2_X1 U12466 ( .A(n11980), .B(n11979), .ZN(n12686) );
  NAND2_X1 U12467 ( .A1(n9855), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10248) );
  NAND2_X1 U12468 ( .A1(n9968), .A2(n9969), .ZN(n10250) );
  AND2_X1 U12469 ( .A1(n14172), .A2(n10172), .ZN(n14620) );
  NAND2_X1 U12470 ( .A1(n15262), .A2(n9885), .ZN(n15050) );
  NAND2_X1 U12471 ( .A1(n15262), .A2(n15570), .ZN(n15080) );
  OR2_X1 U12472 ( .A1(n18778), .A2(n11397), .ZN(n9822) );
  INV_X1 U12473 ( .A(n10695), .ZN(n13914) );
  AND2_X1 U12474 ( .A1(n14578), .A2(n10164), .ZN(n14551) );
  OR2_X1 U12475 ( .A1(n17904), .A2(n10115), .ZN(n9823) );
  NAND2_X1 U12476 ( .A1(n15143), .A2(n13163), .ZN(n13202) );
  INV_X1 U12477 ( .A(n11334), .ZN(n9959) );
  INV_X1 U12478 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10563) );
  AND2_X1 U12479 ( .A1(n10203), .A2(n11249), .ZN(n9825) );
  AND2_X1 U12480 ( .A1(n10188), .A2(n16438), .ZN(n15457) );
  NAND2_X1 U12481 ( .A1(n10131), .A2(n12752), .ZN(n16143) );
  AND2_X1 U12482 ( .A1(n9918), .A2(n17642), .ZN(n9826) );
  AND2_X1 U12483 ( .A1(n16335), .A2(n10033), .ZN(n9827) );
  AND2_X1 U12484 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9828) );
  OR2_X1 U12485 ( .A1(n10037), .A2(n10038), .ZN(n9829) );
  OR2_X1 U12486 ( .A1(n10213), .A2(n11237), .ZN(n9830) );
  AND2_X1 U12487 ( .A1(n11654), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9831) );
  NAND2_X1 U12488 ( .A1(n13088), .A2(n13087), .ZN(n14081) );
  NAND2_X1 U12489 ( .A1(n10218), .A2(n9880), .ZN(n15047) );
  AND2_X1 U12490 ( .A1(n13746), .A2(n13085), .ZN(n9832) );
  NAND2_X1 U12491 ( .A1(n10873), .A2(n10872), .ZN(n15274) );
  AND2_X1 U12492 ( .A1(n10514), .A2(n10014), .ZN(n9833) );
  AND2_X1 U12493 ( .A1(n13087), .A2(n10073), .ZN(n9834) );
  AND2_X1 U12494 ( .A1(n9834), .A2(n14249), .ZN(n9835) );
  AND2_X1 U12495 ( .A1(n9964), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9836) );
  OR2_X1 U12496 ( .A1(n17838), .A2(n10101), .ZN(n9837) );
  AND2_X1 U12497 ( .A1(n9835), .A2(n14253), .ZN(n9838) );
  NAND2_X1 U12498 ( .A1(n13689), .A2(n13688), .ZN(n13690) );
  INV_X1 U12499 ( .A(n11277), .ZN(n10022) );
  OR2_X1 U12500 ( .A1(n10679), .A2(n10678), .ZN(n13928) );
  AND2_X1 U12501 ( .A1(n11177), .A2(n10193), .ZN(n9839) );
  AND2_X1 U12502 ( .A1(n9989), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n9840) );
  OR2_X1 U12503 ( .A1(n13433), .A2(n13434), .ZN(n9841) );
  CLKBUF_X3 U12504 ( .A(n10455), .Z(n14346) );
  INV_X1 U12505 ( .A(n11436), .ZN(n15858) );
  NAND2_X1 U12506 ( .A1(n17753), .A2(n17838), .ZN(n17670) );
  AND2_X1 U12507 ( .A1(n11605), .A2(n11604), .ZN(n9843) );
  OR2_X1 U12508 ( .A1(n10617), .A2(n10616), .ZN(n10031) );
  OR2_X1 U12509 ( .A1(n14495), .A2(n10176), .ZN(n9844) );
  OR2_X1 U12510 ( .A1(n17368), .A2(n9995), .ZN(n9845) );
  INV_X1 U12511 ( .A(n10072), .ZN(n19301) );
  NAND2_X1 U12512 ( .A1(n11043), .A2(n11049), .ZN(n10072) );
  NAND2_X1 U12513 ( .A1(n11271), .A2(n11277), .ZN(n9846) );
  NAND2_X1 U12514 ( .A1(n15435), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15432) );
  NAND2_X1 U12515 ( .A1(n10188), .A2(n10190), .ZN(n15458) );
  AND3_X1 U12516 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10253) );
  OR2_X1 U12517 ( .A1(n11263), .A2(n11262), .ZN(n9848) );
  NAND2_X1 U12518 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11501), .ZN(
        n9851) );
  NAND2_X1 U12519 ( .A1(n9811), .A2(n16089), .ZN(n16080) );
  NAND2_X1 U12520 ( .A1(n15231), .A2(n10039), .ZN(n9852) );
  AND2_X1 U12521 ( .A1(n11068), .A2(n11065), .ZN(n11079) );
  OR2_X1 U12522 ( .A1(n11209), .A2(n11217), .ZN(n9854) );
  AND2_X1 U12523 ( .A1(n10157), .A2(n11224), .ZN(n15459) );
  NAND2_X1 U12524 ( .A1(n9804), .A2(n11177), .ZN(n15313) );
  NAND2_X1 U12525 ( .A1(n11000), .A2(n9950), .ZN(n10436) );
  AOI21_X1 U12526 ( .B1(n10654), .B2(n10653), .A(n10652), .ZN(n10659) );
  AND4_X1 U12527 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n9856) );
  AND4_X1 U12528 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n9857) );
  OR2_X1 U12529 ( .A1(n15914), .A2(n18961), .ZN(n9858) );
  AND2_X1 U12530 ( .A1(n9793), .A2(n15415), .ZN(n15306) );
  INV_X1 U12531 ( .A(n10017), .ZN(n11215) );
  OR2_X1 U12532 ( .A1(n11180), .A2(n9854), .ZN(n10017) );
  NAND2_X1 U12533 ( .A1(n17670), .A2(n17700), .ZN(n17701) );
  NAND2_X1 U12534 ( .A1(n11243), .A2(n11242), .ZN(n16406) );
  NAND2_X1 U12535 ( .A1(n14578), .A2(n10166), .ZN(n10168) );
  INV_X1 U12536 ( .A(n9954), .ZN(n9953) );
  NAND2_X1 U12537 ( .A1(n11253), .A2(n9955), .ZN(n9954) );
  INV_X2 U12538 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16509) );
  NAND2_X1 U12539 ( .A1(n16350), .A2(n10137), .ZN(n14380) );
  NAND2_X1 U12540 ( .A1(n15306), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15297) );
  OR2_X1 U12541 ( .A1(n9854), .A2(n10018), .ZN(n9860) );
  INV_X1 U12542 ( .A(n15681), .ZN(n11243) );
  NOR2_X1 U12543 ( .A1(n15129), .A2(n13229), .ZN(n13253) );
  NAND2_X1 U12544 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10252) );
  INV_X1 U12545 ( .A(n10105), .ZN(n10104) );
  NAND2_X1 U12546 ( .A1(n11514), .A2(n18010), .ZN(n10105) );
  OR2_X1 U12547 ( .A1(n12995), .A2(n11634), .ZN(n9861) );
  NOR2_X1 U12548 ( .A1(n15122), .A2(n15121), .ZN(n15120) );
  AND2_X1 U12549 ( .A1(n10407), .A2(n10221), .ZN(n9862) );
  NAND2_X1 U12550 ( .A1(n14378), .A2(n15479), .ZN(n9863) );
  AND2_X1 U12551 ( .A1(n11014), .A2(n10386), .ZN(n10425) );
  AND2_X1 U12552 ( .A1(n9851), .A2(n9823), .ZN(n9864) );
  INV_X1 U12553 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17924) );
  INV_X1 U12554 ( .A(n11169), .ZN(n10137) );
  INV_X2 U12555 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10456) );
  INV_X1 U12556 ( .A(n10455), .ZN(n10510) );
  AND2_X1 U12557 ( .A1(n10242), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10240) );
  NOR2_X1 U12558 ( .A1(n10258), .A2(n10224), .ZN(n10246) );
  NOR2_X1 U12559 ( .A1(n14252), .A2(n15210), .ZN(n15143) );
  NAND2_X1 U12560 ( .A1(n14172), .A2(n14238), .ZN(n14237) );
  AND2_X1 U12561 ( .A1(n17426), .A2(n9989), .ZN(n9865) );
  NOR2_X1 U12562 ( .A1(n10248), .A2(n16422), .ZN(n10249) );
  OR2_X1 U12563 ( .A1(n13445), .A2(n16463), .ZN(n9866) );
  OR2_X1 U12564 ( .A1(n17838), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9867) );
  NOR2_X1 U12565 ( .A1(n10260), .A2(n10243), .ZN(n10244) );
  INV_X1 U12566 ( .A(n20278), .ZN(n12691) );
  NAND2_X1 U12567 ( .A1(n13724), .A2(n13723), .ZN(n13722) );
  AND2_X1 U12568 ( .A1(n14756), .A2(n9904), .ZN(n9868) );
  NOR2_X1 U12569 ( .A1(n13445), .A2(n10051), .ZN(n13980) );
  NAND2_X1 U12570 ( .A1(n20272), .A2(n9803), .ZN(n12758) );
  NOR2_X1 U12571 ( .A1(n15139), .A2(n10071), .ZN(n9869) );
  OAI211_X1 U12572 ( .C1(n10383), .C2(n10384), .A(n14058), .B(n10398), .ZN(
        n11014) );
  AND2_X1 U12573 ( .A1(n12768), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9870) );
  NOR2_X1 U12574 ( .A1(n15134), .A2(n15133), .ZN(n14326) );
  AND2_X1 U12575 ( .A1(n10217), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9871) );
  OR2_X1 U12576 ( .A1(n10690), .A2(n10689), .ZN(n11110) );
  INV_X1 U12577 ( .A(n11220), .ZN(n10158) );
  NOR2_X1 U12578 ( .A1(n16756), .A2(n17685), .ZN(n9872) );
  INV_X1 U12579 ( .A(n15154), .ZN(n15162) );
  NOR2_X1 U12580 ( .A1(n15175), .A2(n15163), .ZN(n15154) );
  AND2_X1 U12581 ( .A1(n10264), .A2(n9964), .ZN(n9873) );
  INV_X1 U12582 ( .A(n13928), .ZN(n10038) );
  OR2_X1 U12583 ( .A1(n14566), .A2(n14554), .ZN(n9874) );
  NAND2_X1 U12584 ( .A1(n14172), .A2(n10171), .ZN(n14619) );
  NOR2_X1 U12585 ( .A1(n9949), .A2(n10181), .ZN(n11022) );
  AND2_X1 U12586 ( .A1(n10172), .A2(n12180), .ZN(n9875) );
  NOR2_X1 U12587 ( .A1(n10004), .A2(n14954), .ZN(n9876) );
  AND2_X1 U12588 ( .A1(n9833), .A2(n10013), .ZN(n9877) );
  INV_X1 U12589 ( .A(n10139), .ZN(n10138) );
  OR2_X1 U12590 ( .A1(n10260), .A2(n9963), .ZN(n9878) );
  INV_X1 U12591 ( .A(n13859), .ZN(n20144) );
  OAI22_X1 U12592 ( .A1(n16509), .A2(n14363), .B1(n14353), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14179) );
  INV_X1 U12593 ( .A(n19192), .ZN(n9977) );
  INV_X1 U12594 ( .A(n9920), .ZN(n9921) );
  NAND2_X1 U12595 ( .A1(n20086), .A2(n12869), .ZN(n13990) );
  NAND2_X1 U12596 ( .A1(n13747), .A2(n13746), .ZN(n13741) );
  NOR2_X1 U12597 ( .A1(n10236), .A2(n15307), .ZN(n10231) );
  NOR2_X1 U12598 ( .A1(n14245), .A2(n14246), .ZN(n14244) );
  INV_X1 U12599 ( .A(n17838), .ZN(n17873) );
  NOR2_X1 U12600 ( .A1(n10239), .A2(n16373), .ZN(n10234) );
  NAND2_X1 U12601 ( .A1(n13960), .A2(n10015), .ZN(n13451) );
  NOR2_X1 U12602 ( .A1(n13775), .A2(n10035), .ZN(n13913) );
  AND2_X1 U12603 ( .A1(n13689), .A2(n10045), .ZN(n15705) );
  AND2_X1 U12604 ( .A1(n13088), .A2(n9835), .ZN(n14247) );
  AND2_X1 U12605 ( .A1(n13088), .A2(n9834), .ZN(n14166) );
  AND2_X1 U12606 ( .A1(n13689), .A2(n10042), .ZN(n13444) );
  AND2_X1 U12607 ( .A1(n17834), .A2(n10091), .ZN(n17796) );
  OR2_X1 U12608 ( .A1(n14386), .A2(n14414), .ZN(n9879) );
  AND2_X1 U12609 ( .A1(n15077), .A2(n15063), .ZN(n9880) );
  AND2_X1 U12610 ( .A1(n10091), .A2(n18146), .ZN(n9881) );
  AND3_X1 U12611 ( .A1(n10132), .A2(n9862), .A3(n11015), .ZN(n11000) );
  XOR2_X1 U12612 ( .A(n19184), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n9882) );
  OR2_X1 U12613 ( .A1(n19192), .A2(n19216), .ZN(n9883) );
  INV_X1 U12614 ( .A(n10392), .ZN(n13541) );
  XNOR2_X1 U12615 ( .A(n10650), .B(n10651), .ZN(n13714) );
  NAND2_X1 U12616 ( .A1(n13915), .A2(n10719), .ZN(n13555) );
  AND2_X1 U12617 ( .A1(n10053), .A2(n10052), .ZN(n9884) );
  NOR3_X1 U12618 ( .A1(n10236), .A2(n9972), .A3(n9971), .ZN(n10225) );
  NOR2_X1 U12619 ( .A1(n10236), .A2(n9971), .ZN(n10228) );
  AND2_X1 U12620 ( .A1(n9884), .A2(n15051), .ZN(n9885) );
  AND2_X1 U12621 ( .A1(n11677), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9886) );
  AND2_X1 U12622 ( .A1(n9880), .A2(n10011), .ZN(n9887) );
  INV_X1 U12623 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9970) );
  INV_X1 U12624 ( .A(n10064), .ZN(n10063) );
  OR2_X1 U12625 ( .A1(n14410), .A2(n10065), .ZN(n10064) );
  AND2_X1 U12626 ( .A1(n14624), .A2(n14851), .ZN(n9888) );
  AND2_X1 U12627 ( .A1(n13203), .A2(n10070), .ZN(n9889) );
  AND2_X1 U12628 ( .A1(n10113), .A2(n10111), .ZN(n9890) );
  AND2_X1 U12629 ( .A1(n9881), .A2(n18160), .ZN(n9891) );
  AND2_X1 U12630 ( .A1(n10034), .A2(n13928), .ZN(n9892) );
  INV_X1 U12631 ( .A(n15200), .ZN(n10514) );
  NOR2_X1 U12632 ( .A1(n17942), .A2(n17941), .ZN(n17940) );
  NAND2_X1 U12633 ( .A1(n17810), .A2(n9871), .ZN(n9915) );
  NAND2_X1 U12634 ( .A1(n12775), .A2(n12914), .ZN(n9893) );
  AND2_X1 U12635 ( .A1(n10089), .A2(n10088), .ZN(n9894) );
  INV_X1 U12636 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9965) );
  INV_X1 U12637 ( .A(n10103), .ZN(n10102) );
  NAND2_X1 U12638 ( .A1(n13012), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10103) );
  INV_X1 U12639 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9910) );
  INV_X1 U12640 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9972) );
  INV_X1 U12641 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9973) );
  INV_X1 U12642 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n9991) );
  INV_X1 U12643 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n9990) );
  OR2_X1 U12644 ( .A1(n16318), .A2(n13840), .ZN(n20258) );
  NAND3_X2 U12645 ( .A1(n18974), .A2(n18973), .A3(n20997), .ZN(n18289) );
  CLKBUF_X1 U12646 ( .A(n18213), .Z(n9895) );
  NOR3_X1 U12647 ( .A1(n17461), .A2(n15928), .A3(n18217), .ZN(n18213) );
  OAI21_X2 U12648 ( .B1(n16508), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14095), 
        .ZN(n19738) );
  NOR3_X2 U12649 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18658), .A3(
        n18528), .ZN(n18497) );
  NOR3_X2 U12650 ( .A1(n18658), .A2(n18603), .A3(n18578), .ZN(n18573) );
  OAI22_X2 U12651 ( .A1(n20290), .A2(n20300), .B1(n20289), .B2(n20298), .ZN(
        n20855) );
  OAI22_X2 U12652 ( .A1(n20301), .A2(n20300), .B1(n20299), .B2(n20298), .ZN(
        n20861) );
  AOI22_X2 U12653 ( .A1(DATAI_23_), .A2(n20311), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20310), .ZN(n20883) );
  AOI22_X2 U12654 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20310), .B1(DATAI_26_), 
        .B2(n20311), .ZN(n20846) );
  AOI22_X2 U12655 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20310), .B1(DATAI_27_), 
        .B2(n20311), .ZN(n20852) );
  AOI22_X2 U12656 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20310), .B1(DATAI_29_), 
        .B2(n20311), .ZN(n20866) );
  AOI22_X2 U12657 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20310), .B1(DATAI_20_), 
        .B2(n20311), .ZN(n20858) );
  AOI22_X2 U12658 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20310), .B1(DATAI_25_), 
        .B2(n20311), .ZN(n20840) );
  NOR3_X4 U12659 ( .A1(n19239), .A2(n10402), .A3(n14106), .ZN(n19222) );
  AOI22_X2 U12660 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19365), .ZN(n19839) );
  NOR2_X2 U12661 ( .A1(n14106), .A2(n14105), .ZN(n19365) );
  NOR2_X2 U12662 ( .A1(n18411), .A2(n18319), .ZN(n18710) );
  NOR2_X2 U12663 ( .A1(n18921), .A2(n18813), .ZN(n16987) );
  OAI22_X2 U12664 ( .A1(n21017), .A2(n20298), .B1(n20275), .B2(n20300), .ZN(
        n20837) );
  NOR4_X4 U12665 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n10456), .ZN(n19174) );
  AOI22_X2 U12666 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20310), .B1(DATAI_16_), 
        .B2(n20311), .ZN(n20834) );
  NAND2_X1 U12667 ( .A1(n10438), .A2(n9896), .ZN(n11041) );
  NAND2_X2 U12668 ( .A1(n9899), .A2(n11213), .ZN(n15468) );
  AND2_X2 U12669 ( .A1(n11164), .A2(n11152), .ZN(n11208) );
  NAND2_X1 U12670 ( .A1(n9902), .A2(n10151), .ZN(n11133) );
  NAND4_X1 U12671 ( .A1(n9859), .A2(n9936), .A3(n11057), .A4(n9937), .ZN(n9935) );
  NOR2_X2 U12672 ( .A1(n11060), .A2(n9903), .ZN(n11114) );
  NOR2_X2 U12674 ( .A1(n15014), .A2(n14628), .ZN(n14629) );
  NOR2_X2 U12675 ( .A1(n14241), .A2(n14242), .ZN(n14640) );
  NOR3_X2 U12676 ( .A1(n14566), .A2(n14728), .A3(n14554), .ZN(n14729) );
  INV_X1 U12677 ( .A(n9913), .ZN(n16519) );
  XNOR2_X2 U12678 ( .A(n9911), .B(n9910), .ZN(n9920) );
  INV_X1 U12679 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9912) );
  INV_X1 U12680 ( .A(n9915), .ZN(n17763) );
  NAND2_X1 U12681 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9914) );
  NOR2_X1 U12682 ( .A1(n16694), .A2(n9920), .ZN(n16683) );
  NAND3_X1 U12684 ( .A1(n9928), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17832) );
  XNOR2_X2 U12685 ( .A(n11040), .B(n11039), .ZN(n13726) );
  NAND3_X1 U12686 ( .A1(n11049), .A2(n11035), .A3(n11032), .ZN(n9929) );
  AND2_X4 U12687 ( .A1(n14016), .A2(n10574), .ZN(n10373) );
  AND2_X1 U12688 ( .A1(n11056), .A2(n11054), .ZN(n9936) );
  NAND3_X1 U12689 ( .A1(n9935), .A2(n9934), .A3(n9931), .ZN(n11109) );
  NAND2_X2 U12690 ( .A1(n11091), .A2(n11109), .ZN(n14117) );
  NAND2_X1 U12691 ( .A1(n11201), .A2(n9944), .ZN(n9943) );
  NAND2_X1 U12692 ( .A1(n11201), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14113) );
  OR2_X1 U12693 ( .A1(n11201), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14114) );
  NOR2_X2 U12694 ( .A1(n9947), .A2(n10181), .ZN(n10455) );
  NOR2_X2 U12695 ( .A1(n15585), .A2(n15572), .ZN(n9987) );
  NAND3_X1 U12696 ( .A1(n9861), .A2(n11633), .A3(n9993), .ZN(n9992) );
  NAND3_X1 U12697 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(P3_EAX_REG_28__SCAN_IN), 
        .A3(P3_EAX_REG_27__SCAN_IN), .ZN(n9995) );
  INV_X1 U12698 ( .A(n17354), .ZN(n17359) );
  NAND2_X1 U12699 ( .A1(n11835), .A2(n11918), .ZN(n11933) );
  NAND3_X1 U12700 ( .A1(n11829), .A2(n12847), .A3(n11840), .ZN(n12835) );
  OAI21_X1 U12701 ( .B1(n11972), .B2(n12695), .A(n9791), .ZN(n10000) );
  INV_X1 U12702 ( .A(n10000), .ZN(n11965) );
  NAND2_X2 U12703 ( .A1(n11965), .A2(n11964), .ZN(n10160) );
  INV_X1 U12704 ( .A(n14954), .ZN(n10002) );
  OAI21_X1 U12705 ( .B1(n12771), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n14943), .ZN(n14959) );
  INV_X1 U12706 ( .A(n10004), .ZN(n10003) );
  NAND2_X1 U12707 ( .A1(n12062), .A2(n10005), .ZN(n12761) );
  AND2_X2 U12708 ( .A1(n12761), .A2(n12760), .ZN(n12771) );
  NOR2_X1 U12709 ( .A1(n14884), .A2(n10008), .ZN(n13040) );
  NAND2_X1 U12710 ( .A1(n10009), .A2(n10010), .ZN(n13752) );
  NAND2_X1 U12711 ( .A1(n10451), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10012) );
  NOR2_X2 U12712 ( .A1(n11180), .A2(n9860), .ZN(n11225) );
  NAND2_X1 U12713 ( .A1(n11271), .A2(n10019), .ZN(n11301) );
  NAND2_X1 U12714 ( .A1(n10025), .A2(n10023), .ZN(n11266) );
  NAND2_X1 U12715 ( .A1(n11323), .A2(n14329), .ZN(n11315) );
  NAND2_X1 U12716 ( .A1(n11323), .A2(n10028), .ZN(n11325) );
  NAND2_X1 U12717 ( .A1(n11232), .A2(n10030), .ZN(n11246) );
  INV_X1 U12718 ( .A(n10031), .ZN(n11188) );
  NAND2_X1 U12719 ( .A1(n10031), .A2(n10619), .ZN(n10624) );
  NAND2_X1 U12720 ( .A1(n10036), .A2(n9770), .ZN(n13915) );
  NAND2_X1 U12721 ( .A1(n9770), .A2(n9892), .ZN(n13912) );
  INV_X1 U12722 ( .A(n10055), .ZN(n13306) );
  NAND2_X2 U12723 ( .A1(n10055), .A2(n13304), .ZN(n15109) );
  NAND3_X1 U12724 ( .A1(n10060), .A2(n10061), .A3(n10057), .ZN(n13367) );
  NAND3_X1 U12725 ( .A1(n15109), .A2(n15116), .A3(n13348), .ZN(n10060) );
  INV_X1 U12726 ( .A(n10062), .ZN(n14409) );
  NAND2_X1 U12727 ( .A1(n10066), .A2(n10063), .ZN(n10062) );
  NAND2_X1 U12728 ( .A1(n15145), .A2(n9889), .ZN(n10067) );
  NAND2_X1 U12729 ( .A1(n13088), .A2(n9838), .ZN(n14252) );
  AND2_X2 U12730 ( .A1(n13747), .A2(n10074), .ZN(n13963) );
  NAND2_X1 U12731 ( .A1(n10076), .A2(n17959), .ZN(n11652) );
  NAND2_X1 U12732 ( .A1(n11646), .A2(n10076), .ZN(n11492) );
  AOI21_X1 U12733 ( .B1(n17484), .B2(n10076), .A(n10075), .ZN(n17490) );
  INV_X1 U12734 ( .A(n17920), .ZN(n10090) );
  XNOR2_X1 U12735 ( .A(n11494), .B(n11493), .ZN(n17930) );
  NAND2_X1 U12736 ( .A1(n10093), .A2(n9837), .ZN(n10097) );
  NAND3_X1 U12737 ( .A1(n17670), .A2(n9867), .A3(n10104), .ZN(n10093) );
  NAND2_X1 U12738 ( .A1(n10106), .A2(n10097), .ZN(n17625) );
  INV_X1 U12739 ( .A(n10107), .ZN(n17656) );
  NAND2_X1 U12740 ( .A1(n17903), .A2(n9864), .ZN(n10110) );
  INV_X1 U12741 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10115) );
  INV_X1 U12742 ( .A(n10116), .ZN(n10117) );
  OAI21_X1 U12743 ( .B1(n16157), .B2(n10118), .A(n12738), .ZN(n10116) );
  INV_X1 U12744 ( .A(n12731), .ZN(n10118) );
  NAND2_X1 U12746 ( .A1(n16144), .A2(n10129), .ZN(n10128) );
  NAND2_X1 U12747 ( .A1(n10128), .A2(n10127), .ZN(n14974) );
  NAND2_X1 U12748 ( .A1(n11179), .A2(n10134), .ZN(n10133) );
  OAI211_X1 U12749 ( .C1(n11179), .C2(n10139), .A(n10133), .B(n10135), .ZN(
        n15740) );
  NAND2_X1 U12750 ( .A1(n10142), .A2(n19165), .ZN(n11205) );
  NAND2_X1 U12751 ( .A1(n15740), .A2(n15741), .ZN(n11207) );
  NAND2_X1 U12752 ( .A1(n19165), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10139) );
  NAND2_X1 U12753 ( .A1(n10141), .A2(n15755), .ZN(n10140) );
  INV_X1 U12754 ( .A(n19165), .ZN(n10141) );
  NAND3_X1 U12755 ( .A1(n10146), .A2(n11333), .A3(n11343), .ZN(n10145) );
  NAND2_X1 U12756 ( .A1(n15314), .A2(n10210), .ZN(n14375) );
  INV_X1 U12757 ( .A(n15468), .ZN(n10159) );
  NAND2_X2 U12758 ( .A1(n11966), .A2(n10160), .ZN(n13828) );
  INV_X1 U12759 ( .A(n13986), .ZN(n12091) );
  NAND2_X1 U12760 ( .A1(n13988), .A2(n13987), .ZN(n13986) );
  NAND2_X1 U12762 ( .A1(n15037), .A2(n10161), .ZN(n13623) );
  NOR2_X1 U12763 ( .A1(n13625), .A2(n10161), .ZN(n13626) );
  NAND3_X1 U12764 ( .A1(n10162), .A2(n11971), .A3(n13784), .ZN(n13789) );
  NAND2_X1 U12765 ( .A1(n13784), .A2(n13783), .ZN(n13782) );
  NAND2_X1 U12766 ( .A1(n11971), .A2(n11987), .ZN(n13787) );
  NAND2_X1 U12767 ( .A1(n14578), .A2(n10163), .ZN(n14532) );
  INV_X1 U12768 ( .A(n10168), .ZN(n14550) );
  AND2_X2 U12769 ( .A1(n14172), .A2(n10169), .ZN(n14607) );
  NAND2_X1 U12770 ( .A1(n14506), .A2(n14508), .ZN(n14495) );
  NOR2_X2 U12771 ( .A1(n14495), .A2(n14496), .ZN(n13044) );
  NAND2_X1 U12772 ( .A1(n10181), .A2(n10401), .ZN(n10337) );
  OAI21_X1 U12773 ( .B1(n14405), .B2(n19305), .A(n10183), .ZN(P2_U2986) );
  XNOR2_X1 U12774 ( .A(n10182), .B(n14381), .ZN(n14405) );
  AOI21_X1 U12775 ( .B1(n14404), .B2(n19302), .A(n14403), .ZN(n10185) );
  AND2_X2 U12776 ( .A1(n15435), .A2(n10186), .ZN(n15415) );
  NAND2_X1 U12777 ( .A1(n15471), .A2(n11173), .ZN(n10191) );
  CLKBUF_X1 U12778 ( .A(n10191), .Z(n10188) );
  NAND2_X1 U12779 ( .A1(n12797), .A2(n16121), .ZN(n12788) );
  NAND2_X1 U12780 ( .A1(n17754), .A2(n18089), .ZN(n17753) );
  INV_X1 U12781 ( .A(n10903), .ZN(n10626) );
  INV_X1 U12782 ( .A(n11049), .ZN(n11050) );
  NAND2_X1 U12783 ( .A1(n10303), .A2(n10371), .ZN(n10310) );
  NAND2_X1 U12784 ( .A1(n10308), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10309) );
  INV_X1 U12785 ( .A(n11015), .ZN(n19991) );
  INV_X1 U12786 ( .A(n11034), .ZN(n10450) );
  NAND2_X1 U12788 ( .A1(n10626), .A2(n10392), .ZN(n10334) );
  INV_X1 U12789 ( .A(n10392), .ZN(n10298) );
  INV_X1 U12790 ( .A(n10234), .ZN(n10237) );
  OR2_X1 U12791 ( .A1(n13031), .A2(n17878), .ZN(n10194) );
  AND2_X2 U12792 ( .A1(n14133), .A2(n14132), .ZN(n14861) );
  INV_X1 U12793 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10355) );
  AND2_X1 U12794 ( .A1(n13563), .A2(n16503), .ZN(n15205) );
  OR2_X1 U12795 ( .A1(n16336), .A2(n19317), .ZN(n10195) );
  AND2_X1 U12796 ( .A1(n10372), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10196) );
  OR2_X1 U12797 ( .A1(n10979), .A2(n19996), .ZN(n10197) );
  AND2_X1 U12798 ( .A1(n18754), .A2(n16534), .ZN(n10198) );
  NAND2_X1 U12799 ( .A1(n19249), .A2(n19368), .ZN(n15276) );
  INV_X1 U12800 ( .A(n15276), .ZN(n13389) );
  AND2_X1 U12801 ( .A1(n11031), .A2(n11030), .ZN(n10199) );
  AND2_X1 U12802 ( .A1(n11027), .A2(n11384), .ZN(n10201) );
  OR3_X1 U12803 ( .A1(n17612), .A2(n18200), .A3(n17608), .ZN(n10202) );
  NOR2_X1 U12804 ( .A1(n11286), .A2(n15378), .ZN(n10203) );
  AND4_X1 U12805 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n10204) );
  AND3_X1 U12806 ( .A1(n11486), .A2(n11485), .A3(n11484), .ZN(n10205) );
  NOR2_X1 U12807 ( .A1(n10228), .A2(n10232), .ZN(n10206) );
  NOR2_X1 U12808 ( .A1(n15262), .A2(n15265), .ZN(n10207) );
  OR2_X1 U12809 ( .A1(n11827), .A2(n20888), .ZN(n10208) );
  AND4_X1 U12810 ( .A1(n11483), .A2(n11482), .A3(n11481), .A4(n11480), .ZN(
        n10209) );
  INV_X1 U12811 ( .A(n11827), .ZN(n11828) );
  AND2_X1 U12812 ( .A1(n15315), .A2(n15322), .ZN(n10210) );
  OR2_X1 U12813 ( .A1(n11298), .A2(n15389), .ZN(n10211) );
  AND4_X1 U12814 ( .A1(n11280), .A2(n15428), .A3(n15410), .A4(n15400), .ZN(
        n10212) );
  NOR2_X1 U12815 ( .A1(n11234), .A2(n11233), .ZN(n10213) );
  INV_X1 U12816 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12794) );
  NAND2_X1 U12817 ( .A1(n20885), .A2(n20260), .ZN(n20432) );
  OR2_X1 U12818 ( .A1(n11190), .A2(n19051), .ZN(n10214) );
  AND2_X1 U12819 ( .A1(n12678), .A2(n14128), .ZN(n20186) );
  INV_X1 U12820 ( .A(n12120), .ZN(n12247) );
  INV_X1 U12821 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15473) );
  AND2_X1 U12822 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10215) );
  AND3_X1 U12823 ( .A1(n17861), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U12824 ( .A1(n17680), .A2(n17960), .ZN(n17678) );
  AND2_X1 U12825 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10217) );
  AND2_X1 U12826 ( .A1(n15154), .A2(n10530), .ZN(n10218) );
  AND2_X1 U12827 ( .A1(n13275), .A2(n13302), .ZN(n10219) );
  NAND2_X2 U12828 ( .A1(n10364), .A2(n10363), .ZN(n14103) );
  INV_X1 U12829 ( .A(n11392), .ZN(n16967) );
  XNOR2_X1 U12830 ( .A(n13067), .B(n13065), .ZN(n13666) );
  AND2_X1 U12831 ( .A1(n10984), .A2(n13564), .ZN(n10221) );
  AND4_X1 U12833 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n10223) );
  NAND2_X1 U12834 ( .A1(n12639), .A2(n12638), .ZN(n12648) );
  OAI21_X1 U12836 ( .B1(n12940), .B2(n12821), .A(n9853), .ZN(n11822) );
  INV_X1 U12837 ( .A(n15388), .ZN(n11281) );
  AOI22_X1 U12838 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U12839 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U12840 ( .A1(n11281), .A2(n10212), .ZN(n11286) );
  NAND2_X1 U12841 ( .A1(n10904), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10905) );
  INV_X1 U12842 ( .A(n10991), .ZN(n10992) );
  INV_X1 U12843 ( .A(n14534), .ZN(n12391) );
  NAND2_X1 U12844 ( .A1(n12037), .A2(n12036), .ZN(n12064) );
  OR2_X1 U12845 ( .A1(n11907), .A2(n11906), .ZN(n12689) );
  AOI21_X1 U12846 ( .B1(n11767), .B2(n11826), .A(n11828), .ZN(n11840) );
  INV_X1 U12847 ( .A(n11919), .ZN(n11932) );
  AOI22_X1 U12848 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11734) );
  INV_X1 U12849 ( .A(n10396), .ZN(n10397) );
  INV_X1 U12850 ( .A(n11158), .ZN(n11150) );
  OR2_X1 U12851 ( .A1(n14523), .A2(n14714), .ZN(n12452) );
  INV_X1 U12852 ( .A(n14621), .ZN(n12164) );
  INV_X1 U12853 ( .A(n12063), .ZN(n12061) );
  NAND2_X1 U12854 ( .A1(n12691), .A2(n20284), .ZN(n12622) );
  INV_X1 U12855 ( .A(n12661), .ZN(n12669) );
  INV_X1 U12856 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10918) );
  INV_X1 U12857 ( .A(n13254), .ZN(n13255) );
  NOR2_X1 U12858 ( .A1(n10626), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10586) );
  INV_X1 U12859 ( .A(n11330), .ZN(n10924) );
  NAND2_X1 U12860 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U12861 ( .A1(n12824), .A2(n20261), .ZN(n12940) );
  NAND2_X1 U12862 ( .A1(n12824), .A2(n13467), .ZN(n14125) );
  NAND2_X1 U12863 ( .A1(n16134), .A2(n16275), .ZN(n12770) );
  AND2_X1 U12864 ( .A1(n12879), .A2(n12878), .ZN(n16297) );
  NOR2_X1 U12865 ( .A1(n10580), .A2(n10569), .ZN(n10570) );
  NAND2_X2 U12866 ( .A1(n10284), .A2(n10283), .ZN(n10392) );
  NAND2_X1 U12867 ( .A1(n10586), .A2(n10625), .ZN(n10618) );
  INV_X1 U12868 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10224) );
  INV_X1 U12869 ( .A(n16438), .ZN(n11172) );
  AOI22_X1 U12870 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U12871 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U12872 ( .A1(n11443), .A2(n11442), .ZN(n11446) );
  INV_X1 U12873 ( .A(n11513), .ZN(n11514) );
  NOR2_X1 U12874 ( .A1(n17475), .A2(n11492), .ZN(n11496) );
  INV_X1 U12875 ( .A(n12503), .ZN(n12501) );
  OR2_X1 U12876 ( .A1(n12619), .A2(n12806), .ZN(n12621) );
  INV_X1 U12877 ( .A(n12479), .ZN(n12478) );
  AND2_X1 U12878 ( .A1(n12372), .A2(n12371), .ZN(n14726) );
  INV_X1 U12879 ( .A(n14620), .ZN(n14634) );
  AND2_X1 U12880 ( .A1(n16118), .A2(n12774), .ZN(n14931) );
  INV_X1 U12881 ( .A(n14177), .ZN(n12888) );
  INV_X1 U12882 ( .A(n14295), .ZN(n14306) );
  NAND2_X1 U12883 ( .A1(n11991), .A2(n11990), .ZN(n20427) );
  AOI21_X1 U12884 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19950), .A(
        n10570), .ZN(n10578) );
  INV_X1 U12885 ( .A(n15155), .ZN(n10530) );
  NOR2_X1 U12886 ( .A1(n14080), .A2(n14079), .ZN(n13087) );
  AND2_X1 U12887 ( .A1(n10471), .A2(n10470), .ZN(n13742) );
  INV_X1 U12888 ( .A(n13305), .ZN(n13304) );
  INV_X1 U12889 ( .A(n14334), .ZN(n14336) );
  XNOR2_X1 U12890 ( .A(n11340), .B(n11339), .ZN(n11341) );
  AND2_X1 U12891 ( .A1(n14011), .A2(n14010), .ZN(n14040) );
  INV_X1 U12892 ( .A(n11591), .ZN(n17267) );
  CLKBUF_X3 U12893 ( .A(n15819), .Z(n17252) );
  INV_X1 U12894 ( .A(n17638), .ZN(n17639) );
  AND2_X1 U12895 ( .A1(n17873), .A2(n21097), .ZN(n11510) );
  AND2_X1 U12896 ( .A1(n18189), .A2(n17836), .ZN(n11508) );
  NAND2_X2 U12897 ( .A1(n18763), .A2(n18781), .ZN(n18181) );
  AND2_X1 U12899 ( .A1(n12525), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U12900 ( .A1(n12273), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12277) );
  NAND2_X1 U12901 ( .A1(n12121), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12140) );
  AND2_X1 U12902 ( .A1(n12097), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12121) );
  AND2_X1 U12903 ( .A1(n14636), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14659) );
  AND2_X1 U12904 ( .A1(n13641), .A2(n13640), .ZN(n14131) );
  NAND2_X1 U12905 ( .A1(n12478), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12503) );
  OR2_X1 U12906 ( .A1(n12277), .A2(n12276), .ZN(n12294) );
  NOR2_X1 U12907 ( .A1(n16121), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16120) );
  INV_X1 U12908 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12012) );
  AOI21_X1 U12909 ( .B1(n12791), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12790), .ZN(n12792) );
  INV_X2 U12910 ( .A(n12771), .ZN(n16134) );
  INV_X1 U12912 ( .A(n20432), .ZN(n20324) );
  OR2_X1 U12913 ( .A1(n9752), .A2(n20251), .ZN(n20389) );
  INV_X1 U12914 ( .A(n20394), .ZN(n20828) );
  AND2_X1 U12915 ( .A1(n15192), .A2(n15191), .ZN(n15193) );
  NOR2_X1 U12916 ( .A1(n14336), .A2(n14335), .ZN(n14337) );
  AND2_X1 U12917 ( .A1(n11297), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15389) );
  OR3_X1 U12918 ( .A1(n11292), .A2(n11169), .A3(n15633), .ZN(n15437) );
  AND2_X1 U12919 ( .A1(n10500), .A2(n10499), .ZN(n14246) );
  AND2_X1 U12920 ( .A1(n11011), .A2(n11010), .ZN(n14041) );
  INV_X1 U12921 ( .A(n19599), .ZN(n19601) );
  OR2_X1 U12922 ( .A1(n19953), .A2(n19963), .ZN(n19730) );
  AND2_X1 U12923 ( .A1(n14013), .A2(n14012), .ZN(n14064) );
  NOR2_X1 U12924 ( .A1(n11637), .A2(n12998), .ZN(n15916) );
  INV_X1 U12925 ( .A(n18331), .ZN(n17343) );
  OAI21_X1 U12926 ( .B1(n17018), .B2(n17678), .A(n18411), .ZN(n17809) );
  NAND2_X1 U12927 ( .A1(n17959), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17951) );
  NAND2_X1 U12928 ( .A1(n11507), .A2(n17872), .ZN(n17837) );
  NOR2_X1 U12929 ( .A1(n17871), .A2(n18193), .ZN(n17870) );
  NOR2_X1 U12930 ( .A1(n18238), .A2(n17894), .ZN(n17893) );
  NOR2_X1 U12931 ( .A1(n17952), .A2(n9831), .ZN(n17942) );
  INV_X1 U12932 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20991) );
  INV_X2 U12933 ( .A(n9849), .ZN(n17296) );
  INV_X1 U12934 ( .A(n13646), .ZN(n14128) );
  NAND2_X1 U12935 ( .A1(n14435), .A2(n14437), .ZN(n20976) );
  INV_X1 U12936 ( .A(n20101), .ZN(n16021) );
  AND2_X1 U12937 ( .A1(n14659), .A2(n14206), .ZN(n20071) );
  NOR2_X1 U12938 ( .A1(n12140), .A2(n12139), .ZN(n12158) );
  NOR2_X2 U12939 ( .A1(n14215), .A2(n14213), .ZN(n20066) );
  AND2_X1 U12940 ( .A1(n14659), .A2(n14202), .ZN(n20099) );
  INV_X1 U12941 ( .A(n14861), .ZN(n14847) );
  NAND2_X1 U12942 ( .A1(n12370), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12440) );
  AOI21_X1 U12944 ( .B1(n14610), .B2(n14623), .A(n12255), .ZN(n14951) );
  NAND2_X1 U12945 ( .A1(n12039), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12066) );
  AND2_X1 U12946 ( .A1(n20190), .A2(n12682), .ZN(n20185) );
  AND2_X1 U12948 ( .A1(n16200), .A2(n15995), .ZN(n16195) );
  AND2_X1 U12949 ( .A1(n12963), .A2(n15940), .ZN(n15999) );
  NOR2_X1 U12950 ( .A1(n16250), .A2(n12903), .ZN(n16223) );
  INV_X1 U12951 ( .A(n20239), .ZN(n16263) );
  NAND2_X1 U12952 ( .A1(n16300), .A2(n14159), .ZN(n14176) );
  AND2_X1 U12953 ( .A1(n12963), .A2(n12942), .ZN(n20238) );
  INV_X1 U12954 ( .A(n20379), .ZN(n20351) );
  INV_X1 U12955 ( .A(n20342), .ZN(n20345) );
  OAI21_X1 U12956 ( .B1(n20357), .B2(n20355), .A(n20354), .ZN(n20382) );
  INV_X1 U12957 ( .A(n20389), .ZN(n20385) );
  INV_X1 U12958 ( .A(n20513), .ZN(n20509) );
  INV_X1 U12959 ( .A(n20541), .ZN(n20544) );
  INV_X1 U12960 ( .A(n20457), .ZN(n20522) );
  INV_X1 U12961 ( .A(n20599), .ZN(n20602) );
  INV_X1 U12962 ( .A(n20639), .ZN(n20645) );
  INV_X1 U12963 ( .A(n20684), .ZN(n20670) );
  INV_X1 U12964 ( .A(n20686), .ZN(n20747) );
  INV_X1 U12965 ( .A(n20548), .ZN(n20685) );
  INV_X1 U12966 ( .A(n20580), .ZN(n20753) );
  INV_X1 U12967 ( .A(n20694), .ZN(n20819) );
  INV_X1 U12968 ( .A(n20720), .ZN(n20847) );
  INV_X1 U12969 ( .A(n20739), .ZN(n20867) );
  INV_X1 U12970 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20884) );
  INV_X1 U12971 ( .A(n19167), .ZN(n19204) );
  INV_X1 U12972 ( .A(n10240), .ZN(n10262) );
  AND2_X1 U12973 ( .A1(n20003), .A2(n10933), .ZN(n19167) );
  AND2_X1 U12974 ( .A1(n13589), .A2(n19781), .ZN(n19172) );
  INV_X1 U12975 ( .A(n15143), .ZN(n15211) );
  INV_X1 U12976 ( .A(n19249), .ZN(n19239) );
  INV_X1 U12977 ( .A(n13484), .ZN(n13591) );
  AND2_X1 U12978 ( .A1(n16462), .A2(n19295), .ZN(n16453) );
  OAI21_X1 U12979 ( .B1(n15390), .B2(n15388), .A(n15375), .ZN(n15380) );
  INV_X1 U12980 ( .A(n15761), .ZN(n19316) );
  AND2_X1 U12981 ( .A1(n19512), .A2(n19940), .ZN(n19446) );
  INV_X1 U12982 ( .A(n19481), .ZN(n19463) );
  INV_X1 U12983 ( .A(n19509), .ZN(n19497) );
  OR3_X1 U12984 ( .A1(n19516), .A2(n19784), .A3(n19515), .ZN(n19534) );
  INV_X1 U12985 ( .A(n19557), .ZN(n19567) );
  INV_X1 U12986 ( .A(n19937), .ZN(n19545) );
  INV_X1 U12987 ( .A(n19625), .ZN(n19626) );
  AND2_X1 U12988 ( .A1(n19953), .A2(n19963), .ZN(n19940) );
  NOR2_X1 U12989 ( .A1(n19695), .A2(n19730), .ZN(n19773) );
  INV_X1 U12990 ( .A(n19813), .ZN(n19801) );
  INV_X1 U12991 ( .A(n19683), .ZN(n19835) );
  AND2_X1 U12992 ( .A1(n19694), .A2(n19545), .ZN(n19859) );
  NAND2_X1 U12993 ( .A1(n18307), .A2(n15915), .ZN(n11637) );
  OAI22_X1 U12994 ( .A1(n18753), .A2(n15928), .B1(n12999), .B2(n18750), .ZN(
        n18755) );
  INV_X1 U12995 ( .A(n17006), .ZN(n17023) );
  INV_X1 U12996 ( .A(n17013), .ZN(n16903) );
  NOR3_X1 U12997 ( .A1(n17459), .A2(n17418), .A3(n17535), .ZN(n17410) );
  NAND2_X1 U12998 ( .A1(n13032), .A2(n10194), .ZN(n13033) );
  NOR2_X1 U12999 ( .A1(n18921), .A2(n17954), .ZN(n17812) );
  INV_X1 U13000 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17883) );
  OAI211_X1 U13001 ( .C1(n13021), .C2(n18217), .A(n13020), .B(n13019), .ZN(
        n13022) );
  NOR2_X1 U13002 ( .A1(n17465), .A2(n11500), .ZN(n16541) );
  NOR2_X1 U13003 ( .A1(n18161), .A2(n18217), .ZN(n18190) );
  NOR2_X1 U13004 ( .A1(n9768), .A2(n18288), .ZN(n18254) );
  NAND2_X1 U13005 ( .A1(n13461), .A2(n14128), .ZN(n14437) );
  AOI21_X1 U13006 ( .B1(n14695), .B2(n20099), .A(n14447), .ZN(n14448) );
  INV_X1 U13007 ( .A(n20051), .ZN(n20093) );
  INV_X1 U13008 ( .A(n20099), .ZN(n20061) );
  INV_X1 U13009 ( .A(n20066), .ZN(n14648) );
  AND2_X2 U13010 ( .A1(n13736), .A2(n14132), .ZN(n20115) );
  INV_X1 U13011 ( .A(n20119), .ZN(n20142) );
  NOR2_X1 U13012 ( .A1(n14437), .A2(n13692), .ZN(n13859) );
  OAI21_X1 U13013 ( .B1(n14852), .B2(n14624), .A(n14623), .ZN(n14966) );
  OR2_X1 U13014 ( .A1(n20186), .A2(n12679), .ZN(n20190) );
  INV_X1 U13015 ( .A(n20185), .ZN(n20179) );
  INV_X1 U13016 ( .A(n20186), .ZN(n20198) );
  AOI21_X1 U13017 ( .B1(n12978), .B2(n20238), .A(n12977), .ZN(n12979) );
  INV_X1 U13018 ( .A(n20238), .ZN(n20230) );
  INV_X1 U13019 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U13020 ( .A1(n20385), .A2(n20685), .ZN(n20342) );
  NAND2_X1 U13021 ( .A1(n20385), .A2(n20753), .ZN(n20379) );
  NAND2_X1 U13022 ( .A1(n20385), .A2(n20785), .ZN(n20426) );
  NAND2_X1 U13023 ( .A1(n20385), .A2(n20650), .ZN(n20446) );
  NAND2_X1 U13024 ( .A1(n20522), .A2(n20753), .ZN(n20513) );
  NAND2_X1 U13025 ( .A1(n20522), .A2(n20785), .ZN(n20541) );
  OR2_X1 U13026 ( .A1(n20656), .A2(n20548), .ZN(n20599) );
  OR2_X1 U13027 ( .A1(n20656), .A2(n20651), .ZN(n20686) );
  NAND2_X1 U13028 ( .A1(n20823), .A2(n20685), .ZN(n20783) );
  NAND2_X1 U13029 ( .A1(n20823), .A2(n20753), .ZN(n20808) );
  NAND2_X1 U13030 ( .A1(n20823), .A2(n20785), .ZN(n20865) );
  OR2_X1 U13031 ( .A1(n14043), .A2(n10584), .ZN(n13483) );
  INV_X1 U13032 ( .A(n19172), .ZN(n19209) );
  NAND2_X1 U13033 ( .A1(n13544), .A2(n13543), .ZN(n19971) );
  AND2_X1 U13034 ( .A1(n15282), .A2(n15276), .ZN(n19243) );
  INV_X1 U13035 ( .A(n19245), .ZN(n14148) );
  INV_X1 U13036 ( .A(n19250), .ZN(n19282) );
  INV_X1 U13037 ( .A(n13523), .ZN(n13597) );
  INV_X1 U13038 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16461) );
  INV_X1 U13039 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19976) );
  INV_X1 U13040 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19958) );
  NAND2_X1 U13041 ( .A1(n19599), .A2(n19512), .ZN(n19400) );
  INV_X1 U13042 ( .A(n19446), .ZN(n19442) );
  NAND2_X1 U13043 ( .A1(n19546), .A2(n19940), .ZN(n19481) );
  NAND2_X1 U13044 ( .A1(n19512), .A2(n19745), .ZN(n19509) );
  NAND2_X1 U13045 ( .A1(n19546), .A2(n19745), .ZN(n19537) );
  NAND2_X1 U13046 ( .A1(n19546), .A2(n19545), .ZN(n19598) );
  NAND2_X1 U13047 ( .A1(n19694), .A2(n19599), .ZN(n19625) );
  NAND2_X1 U13048 ( .A1(n19694), .A2(n19940), .ZN(n19693) );
  INV_X1 U13049 ( .A(n19773), .ZN(n19753) );
  AND2_X1 U13050 ( .A1(n19740), .A2(n19739), .ZN(n19771) );
  NAND2_X1 U13051 ( .A1(n19746), .A2(n19745), .ZN(n19813) );
  INV_X1 U13052 ( .A(n19859), .ZN(n19852) );
  AND2_X1 U13053 ( .A1(n14066), .A2(n14065), .ZN(n16515) );
  NAND2_X1 U13054 ( .A1(n18955), .A2(n18755), .ZN(n16654) );
  NAND2_X1 U13055 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17025), .ZN(n17013) );
  INV_X1 U13056 ( .A(n16977), .ZN(n17022) );
  AND2_X1 U13057 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17087), .ZN(n17083) );
  AND2_X1 U13058 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17093), .ZN(n17087) );
  AND2_X1 U13059 ( .A1(n17340), .A2(n17459), .ZN(n17434) );
  NOR2_X1 U13060 ( .A1(n11476), .A2(n11475), .ZN(n17461) );
  NOR2_X1 U13061 ( .A1(n11429), .A2(n11428), .ZN(n17475) );
  NAND2_X1 U13062 ( .A1(n15987), .A2(n17874), .ZN(n11691) );
  NAND2_X1 U13063 ( .A1(n18074), .A2(n17856), .ZN(n17771) );
  INV_X1 U13064 ( .A(n17874), .ZN(n17853) );
  NAND2_X1 U13065 ( .A1(n17461), .A2(n17955), .ZN(n17878) );
  OAI21_X2 U13066 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20992), .A(n16654), 
        .ZN(n17960) );
  INV_X1 U13067 ( .A(n17955), .ZN(n17964) );
  INV_X1 U13068 ( .A(n9895), .ZN(n18200) );
  INV_X1 U13069 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18579) );
  INV_X1 U13070 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18313) );
  INV_X1 U13071 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18910) );
  NAND2_X1 U13072 ( .A1(n12980), .A2(n12979), .ZN(P1_U3007) );
  NAND2_X1 U13073 ( .A1(n10942), .A2(n10941), .ZN(P2_U2825) );
  NAND2_X1 U13074 ( .A1(n11691), .A2(n11690), .ZN(P3_U2800) );
  NAND2_X1 U13075 ( .A1(n10255), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10251) );
  INV_X1 U13076 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15463) );
  INV_X1 U13077 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16422) );
  NAND2_X1 U13078 ( .A1(n10249), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10247) );
  INV_X1 U13079 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15452) );
  INV_X1 U13080 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10243) );
  INV_X1 U13081 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19021) );
  INV_X1 U13082 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15347) );
  INV_X1 U13083 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16373) );
  INV_X1 U13084 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10545) );
  INV_X1 U13085 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15307) );
  XNOR2_X1 U13086 ( .A(n10225), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11385) );
  INV_X1 U13087 ( .A(n11385), .ZN(n10267) );
  INV_X1 U13088 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14363) );
  INV_X1 U13089 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U13090 ( .A1(n10228), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10229) );
  OR2_X1 U13091 ( .A1(n10225), .A2(n10229), .ZN(n10230) );
  INV_X1 U13092 ( .A(n10230), .ZN(n16343) );
  NOR2_X1 U13093 ( .A1(n10231), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10232) );
  AND2_X1 U13094 ( .A1(n10236), .A2(n15307), .ZN(n10233) );
  NOR2_X1 U13095 ( .A1(n10231), .A2(n10233), .ZN(n15309) );
  NAND2_X1 U13096 ( .A1(n10237), .A2(n10545), .ZN(n10235) );
  NAND2_X1 U13097 ( .A1(n10236), .A2(n10235), .ZN(n15318) );
  INV_X1 U13098 ( .A(n15318), .ZN(n16361) );
  AOI21_X1 U13099 ( .B1(n16373), .B2(n10239), .A(n10234), .ZN(n16372) );
  OR2_X1 U13100 ( .A1(n9873), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10238) );
  NAND2_X1 U13101 ( .A1(n10239), .A2(n10238), .ZN(n15337) );
  INV_X1 U13102 ( .A(n15337), .ZN(n16383) );
  NOR2_X1 U13103 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10240), .ZN(
        n10241) );
  NOR2_X1 U13104 ( .A1(n10264), .A2(n10241), .ZN(n15384) );
  AOI21_X1 U13105 ( .B1(n19021), .B2(n9878), .A(n10263), .ZN(n19020) );
  AND2_X1 U13106 ( .A1(n10260), .A2(n10243), .ZN(n10245) );
  OR2_X1 U13107 ( .A1(n10245), .A2(n10244), .ZN(n19050) );
  INV_X1 U13108 ( .A(n19050), .ZN(n19041) );
  AOI21_X1 U13109 ( .B1(n10258), .B2(n10224), .A(n10246), .ZN(n19065) );
  AOI21_X1 U13110 ( .B1(n10257), .B2(n15452), .A(n10259), .ZN(n19093) );
  AOI21_X1 U13111 ( .B1(n16422), .B2(n10248), .A(n10249), .ZN(n16415) );
  AOI21_X1 U13112 ( .B1(n15463), .B2(n10250), .A(n9855), .ZN(n19125) );
  AOI21_X1 U13113 ( .B1(n15473), .B2(n10251), .A(n10256), .ZN(n19141) );
  AOI21_X1 U13114 ( .B1(n16461), .B2(n10254), .A(n10255), .ZN(n19170) );
  AOI21_X1 U13115 ( .B1(n14185), .B2(n10252), .A(n10253), .ZN(n14182) );
  INV_X1 U13116 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13676) );
  INV_X1 U13117 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19309) );
  AOI22_X1 U13118 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13676), .B1(n19309), 
        .B2(n16509), .ZN(n19198) );
  INV_X1 U13119 ( .A(n19198), .ZN(n14260) );
  INV_X1 U13120 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21219) );
  OAI22_X1 U13121 ( .A1(n16509), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21219), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14259) );
  AND2_X1 U13122 ( .A1(n14260), .A2(n14259), .ZN(n14219) );
  OAI21_X1 U13123 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10252), .ZN(n14427) );
  NAND2_X1 U13124 ( .A1(n14219), .A2(n14427), .ZN(n14180) );
  NOR2_X1 U13125 ( .A1(n14182), .A2(n14180), .ZN(n19191) );
  OAI21_X1 U13126 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10253), .A(
        n10254), .ZN(n19293) );
  NAND2_X1 U13127 ( .A1(n19191), .A2(n19293), .ZN(n19168) );
  NOR2_X1 U13128 ( .A1(n19170), .A2(n19168), .ZN(n19156) );
  OAI21_X1 U13129 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10255), .A(
        n10251), .ZN(n19157) );
  NAND2_X1 U13130 ( .A1(n19156), .A2(n19157), .ZN(n19140) );
  NOR2_X1 U13131 ( .A1(n19141), .A2(n19140), .ZN(n19133) );
  OAI21_X1 U13132 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10256), .A(
        n10250), .ZN(n19134) );
  NAND2_X1 U13133 ( .A1(n19133), .A2(n19134), .ZN(n19123) );
  NOR2_X1 U13134 ( .A1(n19125), .A2(n19123), .ZN(n19113) );
  OAI21_X1 U13135 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9855), .A(
        n10248), .ZN(n19114) );
  NAND2_X1 U13136 ( .A1(n19113), .A2(n19114), .ZN(n13443) );
  NOR2_X1 U13137 ( .A1(n16415), .A2(n13443), .ZN(n19102) );
  OAI21_X1 U13138 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10249), .A(
        n10257), .ZN(n19103) );
  NAND2_X1 U13139 ( .A1(n19102), .A2(n19103), .ZN(n19085) );
  NOR2_X1 U13140 ( .A1(n19093), .A2(n19085), .ZN(n19084) );
  OAI21_X1 U13141 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10259), .A(
        n10258), .ZN(n19075) );
  NAND2_X1 U13142 ( .A1(n19084), .A2(n19075), .ZN(n19064) );
  NOR2_X1 U13143 ( .A1(n19065), .A2(n19064), .ZN(n19057) );
  OAI21_X1 U13144 ( .B1(n10246), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n10260), .ZN(n19058) );
  NAND2_X1 U13145 ( .A1(n19057), .A2(n19058), .ZN(n19040) );
  NOR2_X1 U13146 ( .A1(n19041), .A2(n19040), .ZN(n19039) );
  OR2_X1 U13147 ( .A1(n10244), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10261) );
  NAND2_X1 U13148 ( .A1(n9878), .A2(n10261), .ZN(n19032) );
  NAND2_X1 U13149 ( .A1(n19039), .A2(n19032), .ZN(n19018) );
  NOR2_X1 U13150 ( .A1(n19020), .A2(n19018), .ZN(n19014) );
  OAI21_X1 U13151 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10263), .A(
        n10262), .ZN(n19017) );
  NAND2_X1 U13152 ( .A1(n19014), .A2(n19017), .ZN(n15072) );
  NOR2_X1 U13153 ( .A1(n15384), .A2(n15072), .ZN(n15058) );
  OAI21_X1 U13154 ( .B1(n10264), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n10266), .ZN(n15362) );
  AOI21_X1 U13155 ( .B1(n15347), .B2(n10266), .A(n9873), .ZN(n15349) );
  NOR2_X1 U13156 ( .A1(n15044), .A2(n15349), .ZN(n15043) );
  NOR2_X1 U13157 ( .A1(n19192), .A2(n15043), .ZN(n16382) );
  NOR2_X1 U13158 ( .A1(n19192), .A2(n16359), .ZN(n13429) );
  NOR2_X1 U13159 ( .A1(n16343), .A2(n16342), .ZN(n16341) );
  NOR2_X1 U13160 ( .A1(n19192), .A2(n16341), .ZN(n10268) );
  INV_X1 U13161 ( .A(n19174), .ZN(n19216) );
  AOI21_X1 U13162 ( .B1(n10268), .B2(n10267), .A(n19216), .ZN(n10269) );
  NAND2_X1 U13163 ( .A1(n9821), .A2(n10269), .ZN(n10942) );
  AOI22_X1 U13164 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13165 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10275) );
  AND2_X4 U13166 ( .A1(n13992), .A2(n10574), .ZN(n10375) );
  AOI22_X1 U13167 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10274) );
  AND2_X4 U13168 ( .A1(n14016), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10587) );
  AND2_X4 U13169 ( .A1(n13992), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10374) );
  AOI22_X1 U13170 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10273) );
  NAND4_X1 U13171 ( .A1(n10276), .A2(n10275), .A3(n10274), .A4(n10273), .ZN(
        n10277) );
  NAND2_X1 U13172 ( .A1(n10277), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10284) );
  AOI22_X1 U13173 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13174 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13175 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10279) );
  NAND4_X1 U13176 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  NAND2_X1 U13177 ( .A1(n10282), .A2(n10355), .ZN(n10283) );
  AOI22_X1 U13178 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10285) );
  AND2_X1 U13179 ( .A1(n10285), .A2(n10355), .ZN(n10290) );
  AOI22_X1 U13180 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13181 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13182 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13183 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10291) );
  AND2_X1 U13184 ( .A1(n10291), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10295) );
  AOI22_X1 U13185 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13186 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13187 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10292) );
  AND2_X4 U13188 ( .A1(n10297), .A2(n10296), .ZN(n10903) );
  AOI22_X1 U13189 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13190 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13191 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13192 ( .A1(n9756), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10299) );
  NAND4_X1 U13193 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10303) );
  AOI22_X1 U13194 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13195 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13196 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13197 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10304) );
  NAND4_X1 U13198 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10308) );
  NAND2_X1 U13199 ( .A1(n10385), .A2(n10984), .ZN(n10991) );
  AOI22_X1 U13200 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13201 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13202 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13203 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10311) );
  NAND4_X1 U13204 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10315) );
  NAND2_X1 U13205 ( .A1(n10315), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10322) );
  AOI22_X1 U13206 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13207 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13208 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9767), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13209 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9759), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10316) );
  NAND4_X1 U13210 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10320) );
  NAND2_X1 U13211 ( .A1(n10320), .A2(n10355), .ZN(n10321) );
  NAND2_X1 U13212 ( .A1(n10385), .A2(n10334), .ZN(n10988) );
  NAND2_X1 U13213 ( .A1(n10988), .A2(n19355), .ZN(n10982) );
  NAND2_X1 U13214 ( .A1(n10323), .A2(n10982), .ZN(n11012) );
  AOI22_X1 U13215 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13216 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13217 ( .A1(n9756), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13218 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9767), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10324) );
  NAND4_X1 U13219 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(
        n10333) );
  AOI22_X1 U13220 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13221 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13222 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9762), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13223 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10328) );
  NAND4_X1 U13224 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10332) );
  NAND2_X1 U13225 ( .A1(n11012), .A2(n19351), .ZN(n10338) );
  INV_X1 U13226 ( .A(n10334), .ZN(n10336) );
  NOR2_X1 U13227 ( .A1(n10984), .A2(n13564), .ZN(n10335) );
  INV_X2 U13228 ( .A(n19351), .ZN(n10401) );
  NAND2_X1 U13229 ( .A1(n10338), .A2(n10337), .ZN(n10423) );
  AOI22_X1 U13230 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13231 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10340) );
  NAND4_X1 U13232 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  AOI22_X1 U13233 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13234 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13235 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13236 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U13237 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10348) );
  NAND2_X1 U13238 ( .A1(n10348), .A2(n10371), .ZN(n10349) );
  AOI22_X1 U13239 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13240 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13241 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13242 ( .A1(n9756), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10351) );
  NAND4_X1 U13243 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10356) );
  NAND2_X1 U13244 ( .A1(n10356), .A2(n10355), .ZN(n10364) );
  AOI22_X1 U13245 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13246 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13247 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13248 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10358) );
  NAND4_X1 U13249 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10362) );
  NAND2_X1 U13250 ( .A1(n10362), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10363) );
  NAND2_X1 U13251 ( .A1(n10423), .A2(n11349), .ZN(n10387) );
  NAND2_X1 U13252 ( .A1(n13541), .A2(n19355), .ZN(n10366) );
  NAND2_X1 U13253 ( .A1(n10392), .A2(n11190), .ZN(n10365) );
  NAND2_X1 U13254 ( .A1(n10366), .A2(n10365), .ZN(n10384) );
  NAND2_X1 U13255 ( .A1(n10385), .A2(n19351), .ZN(n10407) );
  AOI22_X1 U13256 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13257 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13258 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13259 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10367) );
  NAND2_X1 U13260 ( .A1(n9857), .A2(n10371), .ZN(n10380) );
  AOI22_X1 U13261 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10286), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13262 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13263 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13264 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10376) );
  NAND4_X1 U13265 ( .A1(n10196), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10379) );
  NAND2_X2 U13266 ( .A1(n10380), .A2(n10379), .ZN(n10400) );
  AND2_X1 U13267 ( .A1(n10400), .A2(n13564), .ZN(n10985) );
  NAND2_X1 U13268 ( .A1(n10407), .A2(n10985), .ZN(n10383) );
  NAND2_X1 U13269 ( .A1(n10382), .A2(n10390), .ZN(n10398) );
  NAND2_X1 U13270 ( .A1(n13539), .A2(n10625), .ZN(n10424) );
  NAND2_X1 U13271 ( .A1(n10424), .A2(n14058), .ZN(n10386) );
  NAND2_X1 U13272 ( .A1(n10387), .A2(n10425), .ZN(n10388) );
  AND3_X1 U13273 ( .A1(n10400), .A2(n19351), .A3(n10903), .ZN(n10389) );
  NAND2_X1 U13274 ( .A1(n10390), .A2(n10389), .ZN(n14057) );
  NOR2_X1 U13275 ( .A1(n10625), .A2(n10381), .ZN(n10391) );
  NAND2_X1 U13276 ( .A1(n14057), .A2(n10391), .ZN(n10395) );
  AND2_X1 U13277 ( .A1(n10400), .A2(n19351), .ZN(n10393) );
  NAND2_X1 U13278 ( .A1(n10395), .A2(n10978), .ZN(n11001) );
  AND2_X1 U13279 ( .A1(n14103), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13600) );
  OAI21_X1 U13280 ( .B1(n19958), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10456), 
        .ZN(n10396) );
  INV_X1 U13281 ( .A(n10398), .ZN(n10399) );
  NAND2_X1 U13282 ( .A1(n10625), .A2(n14103), .ZN(n10969) );
  INV_X1 U13283 ( .A(n10404), .ZN(n13369) );
  INV_X1 U13284 ( .A(n10402), .ZN(n10403) );
  NAND4_X1 U13285 ( .A1(n9950), .A2(n13369), .A3(n10904), .A4(n10403), .ZN(
        n10443) );
  NAND2_X1 U13286 ( .A1(n10405), .A2(n14058), .ZN(n10406) );
  NAND2_X1 U13287 ( .A1(n10408), .A2(n10436), .ZN(n10409) );
  NAND2_X1 U13288 ( .A1(n10508), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10414) );
  INV_X1 U13289 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13290 ( .A1(n10511), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10410) );
  OAI21_X1 U13291 ( .B1(n10510), .B2(n10411), .A(n10410), .ZN(n10412) );
  INV_X1 U13292 ( .A(n10412), .ZN(n10413) );
  INV_X1 U13293 ( .A(n10417), .ZN(n10415) );
  NAND2_X1 U13294 ( .A1(n10416), .A2(n10415), .ZN(n11036) );
  INV_X1 U13295 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10421) );
  NOR2_X1 U13296 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14067) );
  INV_X1 U13297 ( .A(n14067), .ZN(n10420) );
  NAND2_X1 U13298 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10419) );
  OAI211_X1 U13299 ( .C1(n10464), .C2(n10421), .A(n10420), .B(n10419), .ZN(
        n10422) );
  AOI21_X1 U13300 ( .B1(n10455), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10422), .ZN(
        n10429) );
  NAND2_X1 U13301 ( .A1(n10423), .A2(n10424), .ZN(n11021) );
  NAND2_X1 U13302 ( .A1(n11021), .A2(n10425), .ZN(n10426) );
  NAND2_X1 U13303 ( .A1(n10426), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10428) );
  INV_X1 U13304 ( .A(n10432), .ZN(n10434) );
  NOR2_X1 U13305 ( .A1(n10434), .A2(n10433), .ZN(n10435) );
  INV_X1 U13306 ( .A(n10436), .ZN(n10437) );
  AOI22_X1 U13307 ( .A1(n10437), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n14067), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10438) );
  INV_X1 U13308 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10439) );
  INV_X1 U13309 ( .A(n10440), .ZN(n10441) );
  AOI21_X2 U13310 ( .B1(n10508), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10442), .ZN(n10448) );
  INV_X1 U13311 ( .A(n10448), .ZN(n10446) );
  NAND2_X1 U13312 ( .A1(n10451), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10445) );
  NAND2_X1 U13313 ( .A1(n10980), .A2(n14103), .ZN(n10582) );
  AOI22_X1 U13314 ( .A1(n11005), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n14067), .ZN(n10444) );
  NAND2_X1 U13315 ( .A1(n10445), .A2(n10444), .ZN(n10447) );
  NAND2_X1 U13316 ( .A1(n10446), .A2(n10447), .ZN(n11032) );
  INV_X1 U13317 ( .A(n10447), .ZN(n10449) );
  NAND2_X1 U13318 ( .A1(n10451), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13319 ( .A1(n14067), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10452) );
  INV_X1 U13320 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10459) );
  INV_X1 U13321 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10663) );
  OAI22_X1 U13322 ( .A1(n10464), .A2(n10663), .B1(n10456), .B2(n14185), .ZN(
        n10457) );
  INV_X1 U13323 ( .A(n11039), .ZN(n10460) );
  OR2_X1 U13324 ( .A1(n10462), .A2(n10461), .ZN(n10463) );
  INV_X1 U13325 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15750) );
  INV_X1 U13326 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10694) );
  INV_X1 U13327 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19179) );
  OAI22_X1 U13328 ( .A1(n10556), .A2(n10694), .B1(n10456), .B2(n19179), .ZN(
        n10465) );
  AOI21_X1 U13329 ( .B1(n14346), .B2(P2_EBX_REG_4__SCAN_IN), .A(n10465), .ZN(
        n10466) );
  INV_X1 U13330 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15755) );
  OR2_X1 U13331 ( .A1(n14349), .A2(n15755), .ZN(n10471) );
  INV_X1 U13332 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15751) );
  OAI22_X1 U13333 ( .A1(n10556), .A2(n15751), .B1(n10456), .B2(n16461), .ZN(
        n10469) );
  AOI21_X1 U13334 ( .B1(n14346), .B2(P2_EBX_REG_5__SCAN_IN), .A(n10469), .ZN(
        n10470) );
  NOR2_X2 U13335 ( .A1(n13752), .A2(n13742), .ZN(n13808) );
  INV_X1 U13336 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15727) );
  INV_X1 U13337 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10473) );
  INV_X1 U13338 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10472) );
  OAI22_X1 U13339 ( .A1(n10556), .A2(n10473), .B1(n10456), .B2(n10472), .ZN(
        n10474) );
  AOI21_X1 U13340 ( .B1(n14346), .B2(P2_EBX_REG_6__SCAN_IN), .A(n10474), .ZN(
        n10475) );
  NAND2_X1 U13341 ( .A1(n10476), .A2(n10475), .ZN(n13807) );
  NAND2_X1 U13342 ( .A1(n13808), .A2(n13807), .ZN(n13905) );
  INV_X1 U13343 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16481) );
  INV_X1 U13344 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10477) );
  OAI22_X1 U13345 ( .A1(n10556), .A2(n10477), .B1(n10456), .B2(n15473), .ZN(
        n10478) );
  AOI21_X1 U13346 ( .B1(n14346), .B2(P2_EBX_REG_7__SCAN_IN), .A(n10478), .ZN(
        n10479) );
  NOR2_X2 U13347 ( .A1(n13905), .A2(n13906), .ZN(n13960) );
  INV_X1 U13348 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16491) );
  INV_X1 U13349 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10481) );
  OAI22_X1 U13350 ( .A1(n10556), .A2(n10481), .B1(n10456), .B2(n9970), .ZN(
        n10482) );
  AOI21_X1 U13351 ( .B1(n14346), .B2(P2_EBX_REG_8__SCAN_IN), .A(n10482), .ZN(
        n10483) );
  NAND2_X1 U13352 ( .A1(n10484), .A2(n10483), .ZN(n13959) );
  INV_X1 U13353 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15710) );
  OR2_X1 U13354 ( .A1(n14349), .A2(n15710), .ZN(n10487) );
  INV_X1 U13355 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15464) );
  OAI22_X1 U13356 ( .A1(n10556), .A2(n15464), .B1(n10456), .B2(n15463), .ZN(
        n10485) );
  AOI21_X1 U13357 ( .B1(n14346), .B2(P2_EBX_REG_9__SCAN_IN), .A(n10485), .ZN(
        n10486) );
  NAND2_X1 U13358 ( .A1(n10487), .A2(n10486), .ZN(n13966) );
  INV_X1 U13359 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15696) );
  OR2_X1 U13360 ( .A1(n14349), .A2(n15696), .ZN(n10492) );
  INV_X1 U13361 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10489) );
  INV_X1 U13362 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10488) );
  OAI22_X1 U13363 ( .A1(n10556), .A2(n10489), .B1(n10456), .B2(n10488), .ZN(
        n10490) );
  AOI21_X1 U13364 ( .B1(n14346), .B2(P2_EBX_REG_10__SCAN_IN), .A(n10490), .ZN(
        n10491) );
  NAND2_X1 U13365 ( .A1(n10492), .A2(n10491), .ZN(n14083) );
  INV_X1 U13366 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15673) );
  OR2_X1 U13367 ( .A1(n14349), .A2(n15673), .ZN(n10495) );
  INV_X1 U13368 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10808) );
  OAI22_X1 U13369 ( .A1(n10556), .A2(n10808), .B1(n10456), .B2(n16422), .ZN(
        n10493) );
  AOI21_X1 U13370 ( .B1(n14346), .B2(P2_EBX_REG_11__SCAN_IN), .A(n10493), .ZN(
        n10494) );
  NAND2_X1 U13371 ( .A1(n10495), .A2(n10494), .ZN(n13450) );
  INV_X1 U13372 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16472) );
  OR2_X1 U13373 ( .A1(n14349), .A2(n16472), .ZN(n10500) );
  INV_X1 U13374 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10827) );
  INV_X1 U13375 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10497) );
  OAI22_X1 U13376 ( .A1(n10556), .A2(n10827), .B1(n10456), .B2(n10497), .ZN(
        n10498) );
  AOI21_X1 U13377 ( .B1(n14346), .B2(P2_EBX_REG_12__SCAN_IN), .A(n10498), .ZN(
        n10499) );
  INV_X1 U13378 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15661) );
  OR2_X1 U13379 ( .A1(n14349), .A2(n15661), .ZN(n10503) );
  INV_X1 U13380 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10842) );
  OAI22_X1 U13381 ( .A1(n10556), .A2(n10842), .B1(n10456), .B2(n15452), .ZN(
        n10501) );
  AOI21_X1 U13382 ( .B1(n14346), .B2(P2_EBX_REG_13__SCAN_IN), .A(n10501), .ZN(
        n10502) );
  NAND2_X1 U13383 ( .A1(n10503), .A2(n10502), .ZN(n14254) );
  INV_X1 U13384 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15655) );
  OR2_X1 U13385 ( .A1(n14349), .A2(n15655), .ZN(n10507) );
  INV_X1 U13386 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10855) );
  INV_X1 U13387 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10504) );
  OAI22_X1 U13388 ( .A1(n10556), .A2(n10855), .B1(n10456), .B2(n10504), .ZN(
        n10505) );
  AOI21_X1 U13389 ( .B1(n14346), .B2(P2_EBX_REG_14__SCAN_IN), .A(n10505), .ZN(
        n10506) );
  NAND2_X1 U13390 ( .A1(n10507), .A2(n10506), .ZN(n15206) );
  NAND2_X1 U13391 ( .A1(n15207), .A2(n15206), .ZN(n15209) );
  INV_X1 U13392 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13393 ( .A1(n10511), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10512) );
  OAI21_X1 U13394 ( .B1(n10510), .B2(n10920), .A(n10512), .ZN(n10513) );
  AOI21_X1 U13395 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10513), .ZN(n15200) );
  INV_X1 U13396 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19051) );
  AOI22_X1 U13397 ( .A1(n10511), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10516) );
  OAI21_X1 U13398 ( .B1(n10510), .B2(n19051), .A(n10516), .ZN(n10517) );
  AOI21_X1 U13399 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10517), .ZN(n15188) );
  INV_X1 U13400 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13401 ( .A1(n10511), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10518) );
  OAI21_X1 U13402 ( .B1(n10510), .B2(n10922), .A(n10518), .ZN(n10519) );
  AOI21_X1 U13403 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10519), .ZN(n15179) );
  INV_X1 U13404 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15596) );
  OR2_X1 U13405 ( .A1(n14349), .A2(n15596), .ZN(n10522) );
  INV_X1 U13406 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19904) );
  INV_X1 U13407 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15414) );
  OAI22_X1 U13408 ( .A1(n10556), .A2(n19904), .B1(n10456), .B2(n15414), .ZN(
        n10520) );
  AOI21_X1 U13409 ( .B1(n14346), .B2(P2_EBX_REG_18__SCAN_IN), .A(n10520), .ZN(
        n10521) );
  NAND2_X1 U13410 ( .A1(n10522), .A2(n10521), .ZN(n15173) );
  INV_X1 U13411 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15574) );
  OR2_X1 U13412 ( .A1(n14349), .A2(n15574), .ZN(n10525) );
  INV_X1 U13413 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19906) );
  OAI22_X1 U13414 ( .A1(n10556), .A2(n19906), .B1(n10456), .B2(n19021), .ZN(
        n10523) );
  AOI21_X1 U13415 ( .B1(n14346), .B2(P2_EBX_REG_19__SCAN_IN), .A(n10523), .ZN(
        n10524) );
  AND2_X1 U13416 ( .A1(n10525), .A2(n10524), .ZN(n15163) );
  INV_X1 U13417 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15575) );
  OR2_X1 U13418 ( .A1(n14349), .A2(n15575), .ZN(n10529) );
  INV_X1 U13419 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19908) );
  INV_X1 U13420 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10526) );
  OAI22_X1 U13421 ( .A1(n10556), .A2(n19908), .B1(n10456), .B2(n10526), .ZN(
        n10527) );
  AOI21_X1 U13422 ( .B1(n14346), .B2(P2_EBX_REG_20__SCAN_IN), .A(n10527), .ZN(
        n10528) );
  INV_X1 U13423 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15564) );
  OR2_X1 U13424 ( .A1(n14349), .A2(n15564), .ZN(n10533) );
  INV_X1 U13425 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19910) );
  INV_X1 U13426 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15382) );
  OAI22_X1 U13427 ( .A1(n10556), .A2(n19910), .B1(n10456), .B2(n15382), .ZN(
        n10531) );
  AOI21_X1 U13428 ( .B1(n14346), .B2(P2_EBX_REG_21__SCAN_IN), .A(n10531), .ZN(
        n10532) );
  NAND2_X1 U13429 ( .A1(n10533), .A2(n10532), .ZN(n15077) );
  INV_X1 U13430 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11175) );
  OR2_X1 U13431 ( .A1(n14349), .A2(n11175), .ZN(n10536) );
  INV_X1 U13432 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15361) );
  OAI22_X1 U13433 ( .A1(n10556), .A2(n15361), .B1(n10456), .B2(n9965), .ZN(
        n10534) );
  AOI21_X1 U13434 ( .B1(n14346), .B2(P2_EBX_REG_22__SCAN_IN), .A(n10534), .ZN(
        n10535) );
  NAND2_X1 U13435 ( .A1(n10536), .A2(n10535), .ZN(n15063) );
  INV_X1 U13436 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11308) );
  OR2_X1 U13437 ( .A1(n14349), .A2(n11308), .ZN(n10539) );
  INV_X1 U13438 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19913) );
  OAI22_X1 U13439 ( .A1(n10556), .A2(n19913), .B1(n10456), .B2(n15347), .ZN(
        n10537) );
  AOI21_X1 U13440 ( .B1(n14346), .B2(P2_EBX_REG_23__SCAN_IN), .A(n10537), .ZN(
        n10538) );
  AND2_X1 U13441 ( .A1(n10539), .A2(n10538), .ZN(n15048) );
  INV_X1 U13442 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15136) );
  AOI22_X1 U13443 ( .A1(n10511), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10540) );
  OAI21_X1 U13444 ( .B1(n10510), .B2(n15136), .A(n10540), .ZN(n10541) );
  AOI21_X1 U13445 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10541), .ZN(n15133) );
  INV_X1 U13446 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15327) );
  OR2_X1 U13447 ( .A1(n14349), .A2(n15327), .ZN(n10544) );
  INV_X1 U13448 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19916) );
  OAI22_X1 U13449 ( .A1(n10556), .A2(n19916), .B1(n10456), .B2(n16373), .ZN(
        n10542) );
  AOI21_X1 U13450 ( .B1(n14346), .B2(P2_EBX_REG_25__SCAN_IN), .A(n10542), .ZN(
        n10543) );
  NAND2_X1 U13451 ( .A1(n10544), .A2(n10543), .ZN(n14327) );
  INV_X1 U13452 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15508) );
  OR2_X1 U13453 ( .A1(n14349), .A2(n15508), .ZN(n10548) );
  INV_X1 U13454 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19918) );
  OAI22_X1 U13455 ( .A1(n10556), .A2(n19918), .B1(n10456), .B2(n10545), .ZN(
        n10546) );
  AOI21_X1 U13456 ( .B1(n14346), .B2(P2_EBX_REG_26__SCAN_IN), .A(n10546), .ZN(
        n10547) );
  NAND2_X1 U13457 ( .A1(n10548), .A2(n10547), .ZN(n15124) );
  NAND2_X1 U13458 ( .A1(n15125), .A2(n15124), .ZN(n13433) );
  INV_X1 U13459 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15479) );
  OR2_X1 U13460 ( .A1(n14349), .A2(n15479), .ZN(n10551) );
  INV_X1 U13461 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19919) );
  OAI22_X1 U13462 ( .A1(n10556), .A2(n19919), .B1(n10456), .B2(n15307), .ZN(
        n10549) );
  AOI21_X1 U13463 ( .B1(n14346), .B2(P2_EBX_REG_27__SCAN_IN), .A(n10549), .ZN(
        n10550) );
  AND2_X1 U13464 ( .A1(n10551), .A2(n10550), .ZN(n13434) );
  INV_X1 U13465 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21140) );
  OR2_X1 U13466 ( .A1(n14349), .A2(n21140), .ZN(n10555) );
  INV_X1 U13467 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n10552) );
  OAI22_X1 U13468 ( .A1(n10556), .A2(n10552), .B1(n10456), .B2(n9973), .ZN(
        n10553) );
  AOI21_X1 U13469 ( .B1(n14346), .B2(P2_EBX_REG_28__SCAN_IN), .A(n10553), .ZN(
        n10554) );
  AND2_X1 U13470 ( .A1(n10555), .A2(n10554), .ZN(n14383) );
  INV_X1 U13471 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15299) );
  OR2_X1 U13472 ( .A1(n14349), .A2(n15299), .ZN(n10559) );
  INV_X1 U13473 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19921) );
  OAI22_X1 U13474 ( .A1(n10556), .A2(n19921), .B1(n10456), .B2(n9972), .ZN(
        n10557) );
  AOI21_X1 U13475 ( .B1(n14346), .B2(P2_EBX_REG_29__SCAN_IN), .A(n10557), .ZN(
        n10558) );
  NAND2_X1 U13476 ( .A1(n10559), .A2(n10558), .ZN(n15101) );
  INV_X1 U13477 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13478 ( .A1(n10511), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10560) );
  OAI21_X1 U13479 ( .B1(n10510), .B2(n10561), .A(n10560), .ZN(n10562) );
  AOI21_X1 U13480 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10562), .ZN(n14345) );
  NAND2_X1 U13481 ( .A1(n19968), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10565) );
  NAND2_X1 U13482 ( .A1(n10563), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U13483 ( .A1(n10565), .A2(n10564), .ZN(n10970) );
  NAND2_X1 U13484 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19958), .ZN(
        n10567) );
  NAND2_X1 U13485 ( .A1(n10576), .A2(n10567), .ZN(n10568) );
  NAND2_X1 U13486 ( .A1(n10574), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10573) );
  XNOR2_X1 U13487 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10579) );
  INV_X1 U13488 ( .A(n10579), .ZN(n10569) );
  INV_X1 U13489 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n10577) );
  INV_X1 U13490 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16008) );
  NOR2_X1 U13491 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16008), .ZN(
        n10571) );
  AOI221_X1 U13492 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10578), 
        .C1(n10577), .C2(n10578), .A(n10571), .ZN(n10975) );
  INV_X1 U13493 ( .A(n10947), .ZN(n10572) );
  XNOR2_X1 U13494 ( .A(n10970), .B(n10572), .ZN(n10948) );
  OAI21_X1 U13495 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n10574), .A(
        n10573), .ZN(n10575) );
  XNOR2_X1 U13496 ( .A(n10576), .B(n10575), .ZN(n10950) );
  NAND3_X1 U13497 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10578), .A3(
        n10577), .ZN(n10913) );
  XNOR2_X1 U13498 ( .A(n10580), .B(n10579), .ZN(n10901) );
  NAND2_X1 U13499 ( .A1(n10913), .A2(n10901), .ZN(n10945) );
  NOR2_X1 U13500 ( .A1(n10950), .A2(n10945), .ZN(n10961) );
  AND2_X1 U13501 ( .A1(n10948), .A2(n10961), .ZN(n10581) );
  OR2_X1 U13502 ( .A1(n10975), .A2(n10581), .ZN(n14043) );
  INV_X1 U13503 ( .A(n10582), .ZN(n10583) );
  NOR2_X1 U13504 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16509), .ZN(n14076) );
  AND2_X1 U13505 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n14076), .ZN(n16503) );
  NAND2_X1 U13506 ( .A1(n10583), .A2(n16503), .ZN(n10584) );
  NAND2_X1 U13507 ( .A1(READY12_REG_SCAN_IN), .A2(READY21_REG_SCAN_IN), .ZN(
        n20001) );
  NAND2_X1 U13508 ( .A1(n9772), .A2(n20001), .ZN(n10585) );
  NOR2_X1 U13509 ( .A1(n13483), .A2(n10585), .ZN(n13589) );
  INV_X1 U13510 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19781) );
  AOI22_X1 U13511 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13165), .B1(
        n13164), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10593) );
  AND2_X2 U13512 ( .A1(n10587), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10730) );
  INV_X1 U13513 ( .A(n10374), .ZN(n13993) );
  AOI22_X1 U13514 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13515 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10665), .B1(
        n13166), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10591) );
  AND2_X2 U13516 ( .A1(n10589), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10680) );
  AOI22_X1 U13517 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10680), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10590) );
  NAND4_X1 U13518 ( .A1(n10593), .A2(n10592), .A3(n10591), .A4(n10590), .ZN(
        n10601) );
  AND2_X2 U13519 ( .A1(n13352), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10725) );
  AOI22_X1 U13520 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13173), .B1(
        n10725), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13521 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n13171), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10597) );
  NAND2_X1 U13523 ( .A1(n13356), .A2(n10371), .ZN(n10741) );
  INV_X2 U13524 ( .A(n10741), .ZN(n13174) );
  AND2_X1 U13525 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13526 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n13175), .ZN(n10596) );
  NAND4_X1 U13527 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(
        n10600) );
  NAND2_X1 U13528 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10602) );
  INV_X1 U13529 ( .A(n13539), .ZN(n13373) );
  AND2_X2 U13530 ( .A1(n19990), .A2(n20000), .ZN(n10657) );
  NAND2_X1 U13531 ( .A1(n13373), .A2(n10657), .ZN(n10622) );
  OAI211_X1 U13532 ( .C1(n10618), .C2(n11097), .A(n10602), .B(n10622), .ZN(
        n10660) );
  AOI22_X1 U13533 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13166), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13534 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13535 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10609) );
  INV_X1 U13536 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10606) );
  INV_X1 U13537 ( .A(n10730), .ZN(n10605) );
  INV_X1 U13538 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10604) );
  INV_X1 U13539 ( .A(n10607), .ZN(n10608) );
  NAND4_X1 U13540 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10617) );
  AOI22_X1 U13541 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13542 ( .A1(n13171), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13543 ( .A1(n13172), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13175), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13544 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10725), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10612) );
  NAND4_X1 U13545 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10616) );
  INV_X1 U13546 ( .A(n10618), .ZN(n10619) );
  AND2_X1 U13547 ( .A1(n13564), .A2(n20000), .ZN(n10647) );
  INV_X1 U13548 ( .A(n10647), .ZN(n10620) );
  OAI21_X1 U13549 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20000), .A(
        n10620), .ZN(n10621) );
  AND2_X1 U13550 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  AOI21_X1 U13551 ( .B1(n9772), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10628) );
  INV_X1 U13552 ( .A(n13564), .ZN(n19368) );
  NAND2_X1 U13553 ( .A1(n19368), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10627) );
  OAI211_X1 U13554 ( .C1(n10655), .C2(n10421), .A(n10628), .B(n10627), .ZN(
        n13546) );
  NOR2_X1 U13555 ( .A1(n13564), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13556 ( .A1(n10656), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10629) );
  INV_X1 U13557 ( .A(n13714), .ZN(n10654) );
  INV_X1 U13558 ( .A(n10664), .ZN(n10632) );
  INV_X1 U13559 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10631) );
  INV_X1 U13560 ( .A(n13175), .ZN(n13997) );
  INV_X1 U13561 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13055) );
  INV_X1 U13562 ( .A(n13172), .ZN(n10732) );
  INV_X1 U13563 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10630) );
  OAI222_X1 U13564 ( .A1(n10632), .A2(n10631), .B1(n13997), .B2(n13055), .C1(
        n10732), .C2(n10630), .ZN(n10638) );
  AOI22_X1 U13565 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9766), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13566 ( .A1(n13171), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10725), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13567 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10666), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13568 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10633) );
  NAND4_X1 U13569 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n10637) );
  AOI211_X1 U13570 ( .C1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n10680), .A(
        n10638), .B(n10637), .ZN(n10646) );
  INV_X1 U13571 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10640) );
  INV_X1 U13572 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13204) );
  OAI22_X1 U13573 ( .A1(n10640), .A2(n10810), .B1(n10639), .B2(n13204), .ZN(
        n10644) );
  INV_X1 U13574 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10642) );
  INV_X1 U13575 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10641) );
  OAI22_X1 U13576 ( .A1(n10811), .A2(n10642), .B1(n10741), .B2(n10641), .ZN(
        n10643) );
  NOR2_X1 U13577 ( .A1(n10644), .A2(n10643), .ZN(n10645) );
  OR2_X1 U13578 ( .A1(n11094), .A2(n10618), .ZN(n10649) );
  AOI22_X1 U13579 ( .A1(n13539), .A2(n10647), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10648) );
  NAND2_X1 U13580 ( .A1(n10649), .A2(n10648), .ZN(n13715) );
  INV_X1 U13581 ( .A(n13715), .ZN(n10653) );
  NOR2_X1 U13582 ( .A1(n10650), .A2(n10651), .ZN(n10652) );
  XNOR2_X1 U13583 ( .A(n10660), .B(n10659), .ZN(n13774) );
  INV_X1 U13584 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U13585 ( .A1(n14360), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10658) );
  OAI21_X1 U13586 ( .B1(n10655), .B2(n19885), .A(n10658), .ZN(n13773) );
  NOR2_X1 U13587 ( .A1(n13774), .A2(n13773), .ZN(n13775) );
  NOR2_X1 U13588 ( .A1(n10659), .A2(n10660), .ZN(n10661) );
  AOI22_X1 U13589 ( .A1(n10657), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10662) );
  OAI21_X1 U13590 ( .B1(n10655), .B2(n10663), .A(n10662), .ZN(n10679) );
  AOI22_X1 U13591 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10730), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13592 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10665), .B1(
        n13166), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13593 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10680), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10667) );
  NAND4_X1 U13594 ( .A1(n10670), .A2(n10669), .A3(n10668), .A4(n10667), .ZN(
        n10676) );
  AOI22_X1 U13595 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13174), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13596 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13597 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13173), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13598 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13175), .ZN(n10671) );
  NAND4_X1 U13599 ( .A1(n10674), .A2(n10673), .A3(n10672), .A4(n10671), .ZN(
        n10675) );
  NAND2_X1 U13600 ( .A1(n14360), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10677) );
  OAI21_X1 U13601 ( .B1(n10618), .B2(n11087), .A(n10677), .ZN(n10678) );
  AOI22_X1 U13602 ( .A1(n14360), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13603 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13604 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13605 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13166), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13606 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10680), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10681) );
  NAND4_X1 U13607 ( .A1(n10684), .A2(n10683), .A3(n10682), .A4(n10681), .ZN(
        n10690) );
  AOI22_X1 U13608 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13174), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13609 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13610 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13173), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13611 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n13175), .ZN(n10685) );
  NAND4_X1 U13612 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10689) );
  INV_X1 U13613 ( .A(n11110), .ZN(n10691) );
  OR2_X1 U13614 ( .A1(n10618), .A2(n10691), .ZN(n10692) );
  OAI211_X1 U13615 ( .C1(n10655), .C2(n10694), .A(n10693), .B(n10692), .ZN(
        n10695) );
  AOI22_X1 U13616 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13165), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13617 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13618 ( .A1(n10666), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13166), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13619 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10696) );
  NAND4_X1 U13620 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n10705) );
  AOI22_X1 U13621 ( .A1(n13171), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13174), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13622 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13623 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13624 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13175), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10700) );
  NAND4_X1 U13625 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10704) );
  INV_X1 U13626 ( .A(n10915), .ZN(n11131) );
  OAI22_X1 U13627 ( .A1(n11131), .A2(n10618), .B1(n10655), .B2(n15751), .ZN(
        n10706) );
  INV_X1 U13628 ( .A(n10706), .ZN(n10708) );
  AOI22_X1 U13629 ( .A1(n14360), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10707) );
  NAND2_X1 U13630 ( .A1(n10708), .A2(n10707), .ZN(n13916) );
  AOI22_X1 U13631 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13632 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13633 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10666), .B1(
        n13166), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13634 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10680), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10709) );
  NAND4_X1 U13635 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10718) );
  AOI22_X1 U13636 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13174), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13637 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13638 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13172), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13639 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n13175), .ZN(n10713) );
  NAND4_X1 U13640 ( .A1(n10716), .A2(n10715), .A3(n10714), .A4(n10713), .ZN(
        n10717) );
  OR2_X1 U13641 ( .A1(n10618), .A2(n11147), .ZN(n10719) );
  AOI22_X1 U13642 ( .A1(n14360), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10720) );
  OAI21_X1 U13643 ( .B1(n10655), .B2(n10473), .A(n10720), .ZN(n13556) );
  NAND2_X1 U13644 ( .A1(n13555), .A2(n13556), .ZN(n10753) );
  NAND2_X1 U13645 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10724) );
  NAND2_X1 U13646 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10723) );
  NAND2_X1 U13647 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U13648 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10721) );
  INV_X1 U13649 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10729) );
  INV_X1 U13650 ( .A(n13173), .ZN(n10728) );
  INV_X1 U13651 ( .A(n10725), .ZN(n10727) );
  INV_X1 U13652 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10726) );
  OAI22_X1 U13653 ( .A1(n10729), .A2(n10728), .B1(n10727), .B2(n10726), .ZN(
        n10735) );
  INV_X1 U13654 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10733) );
  INV_X1 U13655 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10731) );
  OAI22_X1 U13656 ( .A1(n10605), .A2(n10733), .B1(n10732), .B2(n10731), .ZN(
        n10734) );
  NOR2_X1 U13657 ( .A1(n10735), .A2(n10734), .ZN(n10750) );
  INV_X1 U13658 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10739) );
  INV_X1 U13659 ( .A(n10736), .ZN(n10738) );
  INV_X1 U13660 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10737) );
  OAI22_X1 U13661 ( .A1(n10739), .A2(n10965), .B1(n10738), .B2(n10737), .ZN(
        n10743) );
  INV_X1 U13662 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10740) );
  INV_X1 U13663 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13086) );
  OAI22_X1 U13664 ( .A1(n10741), .A2(n10740), .B1(n13086), .B2(n13997), .ZN(
        n10742) );
  NOR2_X1 U13665 ( .A1(n10743), .A2(n10742), .ZN(n10749) );
  NAND2_X1 U13666 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10747) );
  NAND2_X1 U13667 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10746) );
  NAND2_X1 U13668 ( .A1(n10666), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10745) );
  NAND2_X1 U13669 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10744) );
  AND4_X2 U13670 ( .A1(n10751), .A2(n10750), .A3(n10749), .A4(n10748), .ZN(
        n11169) );
  OR2_X1 U13671 ( .A1(n10618), .A2(n11169), .ZN(n10752) );
  AOI22_X1 U13672 ( .A1(n14360), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10754) );
  OAI21_X1 U13673 ( .B1(n10655), .B2(n10477), .A(n10754), .ZN(n13688) );
  INV_X1 U13674 ( .A(n10655), .ZN(n14361) );
  AOI22_X1 U13675 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13166), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10761) );
  INV_X1 U13676 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10756) );
  INV_X1 U13677 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10755) );
  OAI22_X1 U13678 ( .A1(n10811), .A2(n10756), .B1(n10810), .B2(n10755), .ZN(
        n10757) );
  INV_X1 U13679 ( .A(n10757), .ZN(n10760) );
  AOI22_X1 U13680 ( .A1(n10666), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13681 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10758) );
  NAND4_X1 U13682 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n10767) );
  AOI22_X1 U13683 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13684 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13175), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13685 ( .A1(n13173), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13686 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10725), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10762) );
  NAND4_X1 U13687 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n10766) );
  OR2_X1 U13688 ( .A1(n10767), .A2(n10766), .ZN(n13962) );
  INV_X1 U13689 ( .A(n13962), .ZN(n10769) );
  AOI22_X1 U13690 ( .A1(n14360), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10768) );
  OAI21_X1 U13691 ( .B1(n10618), .B2(n10769), .A(n10768), .ZN(n10770) );
  AOI21_X1 U13692 ( .B1(n14361), .B2(P2_REIP_REG_8__SCAN_IN), .A(n10770), .ZN(
        n16478) );
  AOI22_X1 U13693 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13694 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13695 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13696 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10680), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U13697 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10780) );
  AOI22_X1 U13698 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13699 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13175), .ZN(n10777) );
  AOI22_X1 U13700 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13701 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13172), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10775) );
  NAND4_X1 U13702 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10779) );
  NOR2_X1 U13703 ( .A1(n10780), .A2(n10779), .ZN(n14080) );
  OAI22_X1 U13704 ( .A1(n14080), .A2(n10618), .B1(n10655), .B2(n15464), .ZN(
        n10781) );
  INV_X1 U13705 ( .A(n10781), .ZN(n10783) );
  AOI22_X1 U13706 ( .A1(n14360), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10657), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10782) );
  NAND2_X1 U13707 ( .A1(n10783), .A2(n10782), .ZN(n15707) );
  AOI22_X1 U13708 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13709 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10786) );
  AOI22_X1 U13710 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13711 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10680), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10784) );
  NAND4_X1 U13712 ( .A1(n10787), .A2(n10786), .A3(n10785), .A4(n10784), .ZN(
        n10793) );
  AOI22_X1 U13713 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13714 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13175), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13715 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13716 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13172), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10788) );
  NAND4_X1 U13717 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .ZN(
        n10792) );
  NOR2_X1 U13718 ( .A1(n10793), .A2(n10792), .ZN(n14079) );
  AOI22_X1 U13719 ( .A1(n14360), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10794) );
  OAI21_X1 U13720 ( .B1(n10618), .B2(n14079), .A(n10794), .ZN(n10795) );
  AOI21_X1 U13721 ( .B1(n14361), .B2(P2_REIP_REG_10__SCAN_IN), .A(n10795), 
        .ZN(n15693) );
  AOI22_X1 U13722 ( .A1(n14360), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13723 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13724 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U13725 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13726 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10680), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10796) );
  NAND4_X1 U13727 ( .A1(n10799), .A2(n10798), .A3(n10797), .A4(n10796), .ZN(
        n10805) );
  AOI22_X1 U13728 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13729 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n13175), .ZN(n10802) );
  AOI22_X1 U13730 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13731 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13172), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10800) );
  NAND4_X1 U13732 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10804) );
  NOR2_X1 U13733 ( .A1(n10805), .A2(n10804), .ZN(n14167) );
  OR2_X1 U13734 ( .A1(n10618), .A2(n14167), .ZN(n10806) );
  OAI211_X1 U13735 ( .C1(n10655), .C2(n10808), .A(n10807), .B(n10806), .ZN(
        n13446) );
  AOI22_X1 U13736 ( .A1(n14360), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10826) );
  INV_X1 U13737 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10812) );
  INV_X1 U13738 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10809) );
  OAI22_X1 U13739 ( .A1(n10812), .A2(n10811), .B1(n10810), .B2(n10809), .ZN(
        n10813) );
  INV_X1 U13740 ( .A(n10813), .ZN(n10817) );
  AOI22_X1 U13741 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13742 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13743 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10680), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10814) );
  NAND4_X1 U13744 ( .A1(n10817), .A2(n10816), .A3(n10815), .A4(n10814), .ZN(
        n10823) );
  AOI22_X1 U13745 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10725), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13746 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13747 ( .A1(n13171), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13748 ( .A1(n13173), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13175), .ZN(n10818) );
  NAND4_X1 U13749 ( .A1(n10821), .A2(n10820), .A3(n10819), .A4(n10818), .ZN(
        n10822) );
  OR2_X1 U13750 ( .A1(n10823), .A2(n10822), .ZN(n14249) );
  INV_X1 U13751 ( .A(n14249), .ZN(n10824) );
  OR2_X1 U13752 ( .A1(n10618), .A2(n10824), .ZN(n10825) );
  OAI211_X1 U13753 ( .C1(n10655), .C2(n10827), .A(n10826), .B(n10825), .ZN(
        n10828) );
  INV_X1 U13754 ( .A(n10828), .ZN(n16463) );
  AOI22_X1 U13755 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13756 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13757 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13758 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10829) );
  NAND4_X1 U13759 ( .A1(n10832), .A2(n10831), .A3(n10830), .A4(n10829), .ZN(
        n10838) );
  AOI22_X1 U13760 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13761 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13175), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13762 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13763 ( .A1(n13173), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10833) );
  NAND4_X1 U13764 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10837) );
  OR2_X1 U13765 ( .A1(n10838), .A2(n10837), .ZN(n14253) );
  INV_X1 U13766 ( .A(n14253), .ZN(n10839) );
  OR2_X1 U13767 ( .A1(n10618), .A2(n10839), .ZN(n10841) );
  AOI22_X1 U13768 ( .A1(n14360), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10840) );
  OAI211_X1 U13769 ( .C1(n10655), .C2(n10842), .A(n10841), .B(n10840), .ZN(
        n13981) );
  AOI22_X1 U13770 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10664), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13771 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13772 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13773 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10680), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10843) );
  NAND4_X1 U13774 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10852) );
  AOI22_X1 U13775 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13776 ( .A1(n13171), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U13777 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10725), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U13778 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n13175), .ZN(n10847) );
  NAND4_X1 U13779 ( .A1(n10850), .A2(n10849), .A3(n10848), .A4(n10847), .ZN(
        n10851) );
  NOR2_X1 U13780 ( .A1(n10852), .A2(n10851), .ZN(n15210) );
  OR2_X1 U13781 ( .A1(n10618), .A2(n15210), .ZN(n10854) );
  AOI22_X1 U13782 ( .A1(n14360), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10853) );
  OAI211_X1 U13783 ( .C1(n10655), .C2(n10855), .A(n10854), .B(n10853), .ZN(
        n15649) );
  INV_X1 U13784 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U13785 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13786 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13787 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13788 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10680), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10856) );
  NAND4_X1 U13789 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10865) );
  AOI22_X1 U13790 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13791 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13175), .ZN(n10862) );
  AOI22_X1 U13792 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13793 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13172), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10860) );
  NAND4_X1 U13794 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10864) );
  NOR2_X1 U13795 ( .A1(n10865), .A2(n10864), .ZN(n15197) );
  OR2_X1 U13796 ( .A1(n10618), .A2(n15197), .ZN(n10867) );
  AOI22_X1 U13797 ( .A1(n14360), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10866) );
  OAI211_X1 U13798 ( .C1(n10655), .C2(n19899), .A(n10867), .B(n10866), .ZN(
        n10868) );
  INV_X1 U13799 ( .A(n10868), .ZN(n14144) );
  INV_X1 U13800 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13801 ( .A1(n14360), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10869) );
  OAI21_X1 U13802 ( .B1(n10655), .B2(n10870), .A(n10869), .ZN(n15621) );
  NAND2_X1 U13803 ( .A1(n14145), .A2(n15621), .ZN(n15285) );
  INV_X1 U13804 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U13805 ( .A1(n14360), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10871) );
  OAI21_X1 U13806 ( .B1(n10655), .B2(n19902), .A(n10871), .ZN(n10872) );
  INV_X1 U13807 ( .A(n10872), .ZN(n15287) );
  NAND2_X1 U13808 ( .A1(n14361), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13809 ( .A1(n14360), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10874) );
  AND2_X1 U13810 ( .A1(n10875), .A2(n10874), .ZN(n15275) );
  AOI22_X1 U13811 ( .A1(n14360), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10876) );
  OAI21_X1 U13812 ( .B1(n10655), .B2(n19906), .A(n10876), .ZN(n15264) );
  AOI22_X1 U13813 ( .A1(n14360), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10877) );
  OAI21_X1 U13814 ( .B1(n10655), .B2(n19908), .A(n10877), .ZN(n15570) );
  NAND2_X1 U13815 ( .A1(n14361), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13816 ( .A1(n14360), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10878) );
  AND2_X1 U13817 ( .A1(n10879), .A2(n10878), .ZN(n15081) );
  NAND2_X1 U13818 ( .A1(n14361), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13819 ( .A1(n14360), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10880) );
  AND2_X1 U13820 ( .A1(n10881), .A2(n10880), .ZN(n15065) );
  AOI22_X1 U13821 ( .A1(n10656), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10882) );
  OAI21_X1 U13822 ( .B1(n10655), .B2(n19913), .A(n10882), .ZN(n15051) );
  NAND2_X1 U13823 ( .A1(n14361), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13824 ( .A1(n10656), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10883) );
  AND2_X1 U13825 ( .A1(n10884), .A2(n10883), .ZN(n15242) );
  NAND2_X1 U13826 ( .A1(n14361), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13827 ( .A1(n10656), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10885) );
  AND2_X1 U13828 ( .A1(n10886), .A2(n10885), .ZN(n14317) );
  NAND2_X1 U13829 ( .A1(n14361), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13830 ( .A1(n10656), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10887) );
  AND2_X1 U13831 ( .A1(n10888), .A2(n10887), .ZN(n15232) );
  AOI22_X1 U13832 ( .A1(n10656), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10889) );
  OAI21_X1 U13833 ( .B1(n10655), .B2(n19919), .A(n10889), .ZN(n13437) );
  NAND2_X1 U13834 ( .A1(n14361), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13835 ( .A1(n10656), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10890) );
  AND2_X1 U13836 ( .A1(n10891), .A2(n10890), .ZN(n14386) );
  NAND2_X1 U13837 ( .A1(n14361), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13838 ( .A1(n10656), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10892) );
  AND2_X1 U13839 ( .A1(n10893), .A2(n10892), .ZN(n14414) );
  NAND2_X1 U13840 ( .A1(n14361), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13841 ( .A1(n14360), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10657), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U13842 ( .A1(n10895), .A2(n10894), .ZN(n10896) );
  OR2_X1 U13843 ( .A1(n14413), .A2(n10896), .ZN(n10897) );
  OR2_X1 U13844 ( .A1(n14043), .A2(n11002), .ZN(n14052) );
  INV_X1 U13845 ( .A(n14052), .ZN(n10898) );
  NAND2_X1 U13846 ( .A1(n10898), .A2(n16503), .ZN(n20003) );
  INV_X1 U13847 ( .A(n20001), .ZN(n19996) );
  INV_X1 U13848 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19872) );
  NAND2_X1 U13849 ( .A1(n19872), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20007) );
  INV_X2 U13850 ( .A(n20007), .ZN(n20009) );
  NAND2_X2 U13851 ( .A1(n20009), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19923) );
  NOR2_X1 U13852 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19868) );
  INV_X1 U13853 ( .A(n19868), .ZN(n19878) );
  NAND3_X1 U13854 ( .A1(n19872), .A2(n19923), .A3(n19878), .ZN(n19875) );
  NOR2_X1 U13855 ( .A1(n19996), .A2(n19875), .ZN(n14048) );
  NAND2_X1 U13856 ( .A1(n14048), .A2(n19781), .ZN(n14069) );
  INV_X1 U13857 ( .A(n14069), .ZN(n10899) );
  NAND2_X1 U13858 ( .A1(n10989), .A2(n10899), .ZN(n10900) );
  OR2_X1 U13859 ( .A1(n20003), .A2(n10900), .ZN(n19203) );
  INV_X1 U13860 ( .A(n19203), .ZN(n19182) );
  INV_X1 U13861 ( .A(n10901), .ZN(n10902) );
  NAND2_X1 U13862 ( .A1(n10943), .A2(n10903), .ZN(n10906) );
  NOR2_X1 U13863 ( .A1(n10903), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11189) );
  INV_X1 U13864 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15094) );
  NAND2_X1 U13865 ( .A1(n11189), .A2(n15094), .ZN(n10907) );
  NAND2_X1 U13866 ( .A1(n10908), .A2(n10907), .ZN(n11194) );
  INV_X1 U13867 ( .A(n10950), .ZN(n10909) );
  MUX2_X1 U13868 ( .A(n10910), .B(n10909), .S(n11186), .Z(n10972) );
  MUX2_X1 U13869 ( .A(n10972), .B(n10411), .S(n10904), .Z(n11195) );
  INV_X1 U13870 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n21133) );
  MUX2_X1 U13871 ( .A(n10913), .B(n11110), .S(n11349), .Z(n10944) );
  MUX2_X1 U13872 ( .A(n21133), .B(n10944), .S(n10903), .Z(n11202) );
  INV_X1 U13873 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10916) );
  MUX2_X1 U13874 ( .A(n10916), .B(n10915), .S(n10903), .Z(n11181) );
  MUX2_X1 U13875 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11147), .S(n10903), .Z(
        n11209) );
  MUX2_X1 U13876 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n9765), .S(n11190), .Z(n11217) );
  NAND2_X1 U13877 ( .A1(n10904), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11214) );
  INV_X1 U13878 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10917) );
  INV_X1 U13879 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19111) );
  NAND2_X1 U13880 ( .A1(n10904), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11245) );
  INV_X1 U13881 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10919) );
  NOR2_X1 U13882 ( .A1(n10903), .A2(n10919), .ZN(n11262) );
  NAND2_X1 U13883 ( .A1(n10904), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11265) );
  NOR2_X1 U13884 ( .A1(n11190), .A2(n10920), .ZN(n11259) );
  NOR2_X1 U13885 ( .A1(n11190), .A2(n10922), .ZN(n11256) );
  NAND2_X1 U13886 ( .A1(n10904), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U13887 ( .A1(n10904), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11277) );
  NAND2_X1 U13888 ( .A1(n10904), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11299) );
  INV_X1 U13889 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10923) );
  NOR2_X1 U13890 ( .A1(n11190), .A2(n10923), .ZN(n11304) );
  INV_X1 U13891 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14329) );
  NAND2_X1 U13892 ( .A1(n10904), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U13893 ( .A1(n10904), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11328) );
  INV_X1 U13894 ( .A(n11340), .ZN(n10925) );
  NAND2_X1 U13895 ( .A1(n10904), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U13896 ( .A1(n10925), .A2(n11338), .ZN(n14338) );
  NAND2_X1 U13897 ( .A1(n10904), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10926) );
  XNOR2_X1 U13898 ( .A(n14338), .B(n10926), .ZN(n11344) );
  INV_X1 U13899 ( .A(n11344), .ZN(n11345) );
  INV_X1 U13900 ( .A(n13483), .ZN(n10928) );
  NAND2_X1 U13901 ( .A1(n20001), .A2(n19781), .ZN(n10927) );
  NAND2_X1 U13902 ( .A1(n10928), .A2(n10927), .ZN(n10929) );
  INV_X1 U13903 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16330) );
  OR3_X1 U13904 ( .A1(n10929), .A2(n10625), .A3(n16330), .ZN(n19201) );
  NOR2_X2 U13905 ( .A1(n13483), .A2(n9772), .ZN(n13523) );
  NAND2_X1 U13906 ( .A1(n13523), .A2(n14069), .ZN(n16329) );
  OR2_X1 U13907 ( .A1(n10929), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n10930) );
  NAND2_X1 U13908 ( .A1(n16329), .A2(n10930), .ZN(n19207) );
  NAND2_X1 U13909 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19207), .ZN(n10935) );
  NOR2_X1 U13910 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19941) );
  INV_X1 U13911 ( .A(n19941), .ZN(n15787) );
  NOR2_X1 U13912 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15787), .ZN(n14372) );
  AND2_X1 U13913 ( .A1(n14372), .A2(n16509), .ZN(n11352) );
  INV_X1 U13914 ( .A(n11352), .ZN(n19151) );
  INV_X1 U13915 ( .A(n19151), .ZN(n15730) );
  INV_X1 U13916 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19995) );
  NAND2_X1 U13917 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19995), .ZN(n14075) );
  INV_X1 U13918 ( .A(n14075), .ZN(n19510) );
  AND2_X1 U13919 ( .A1(n14076), .A2(n19510), .ZN(n16504) );
  INV_X1 U13920 ( .A(n16504), .ZN(n10931) );
  NAND2_X1 U13921 ( .A1(n19216), .A2(n10931), .ZN(n10932) );
  NOR2_X1 U13922 ( .A1(n15730), .A2(n10932), .ZN(n10933) );
  OR2_X1 U13923 ( .A1(n19167), .A2(n20000), .ZN(n19178) );
  AOI22_X1 U13924 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19167), .ZN(n10934) );
  OAI211_X1 U13925 ( .C1(n11345), .C2(n19201), .A(n10935), .B(n10934), .ZN(
        n10936) );
  INV_X1 U13926 ( .A(n10936), .ZN(n10937) );
  NAND2_X1 U13927 ( .A1(n10381), .A2(n14048), .ZN(n10998) );
  INV_X1 U13928 ( .A(n10945), .ZN(n10957) );
  NAND2_X1 U13929 ( .A1(n14058), .A2(n9772), .ZN(n10946) );
  MUX2_X1 U13930 ( .A(n11186), .B(n10946), .S(n10950), .Z(n10955) );
  OAI21_X1 U13931 ( .B1(n19976), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10947), .ZN(n11187) );
  INV_X1 U13932 ( .A(n11187), .ZN(n10962) );
  OAI21_X1 U13933 ( .B1(n9772), .B2(n10962), .A(n10948), .ZN(n10949) );
  OAI21_X1 U13934 ( .B1(n10950), .B2(n19990), .A(n10949), .ZN(n10951) );
  NAND2_X1 U13935 ( .A1(n10951), .A2(n14058), .ZN(n10953) );
  OAI21_X1 U13936 ( .B1(n11187), .B2(n10970), .A(n11349), .ZN(n10952) );
  NAND2_X1 U13937 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  NAND2_X1 U13938 ( .A1(n10955), .A2(n10954), .ZN(n10956) );
  AOI22_X1 U13939 ( .A1(n10974), .A2(n11186), .B1(n10957), .B2(n10956), .ZN(
        n10958) );
  AND2_X1 U13940 ( .A1(n10975), .A2(n13600), .ZN(n10959) );
  OAI211_X1 U13941 ( .C1(n14103), .C2(n10960), .A(n13596), .B(n10984), .ZN(
        n10997) );
  AOI21_X1 U13942 ( .B1(n10962), .B2(n10961), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n10963) );
  INV_X1 U13943 ( .A(n10963), .ZN(n10964) );
  OR2_X1 U13944 ( .A1(n14043), .A2(n10964), .ZN(n10968) );
  AOI21_X1 U13945 ( .B1(n13998), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15788) );
  NAND2_X1 U13946 ( .A1(n10965), .A2(n15788), .ZN(n10966) );
  INV_X1 U13947 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18988) );
  AOI21_X1 U13948 ( .B1(n10966), .B2(n18988), .A(n10456), .ZN(n19973) );
  INV_X1 U13949 ( .A(n19973), .ZN(n10967) );
  OR2_X1 U13950 ( .A1(n14057), .A2(n10625), .ZN(n10977) );
  OR2_X1 U13951 ( .A1(n14057), .A2(n10969), .ZN(n11178) );
  NOR2_X1 U13952 ( .A1(n10970), .A2(n11187), .ZN(n10971) );
  NOR2_X1 U13953 ( .A1(n10972), .A2(n10971), .ZN(n10973) );
  NOR2_X1 U13954 ( .A1(n10974), .A2(n10973), .ZN(n10976) );
  OR2_X1 U13955 ( .A1(n10976), .A2(n10975), .ZN(n19980) );
  OAI22_X1 U13956 ( .A1(n19983), .A2(n10977), .B1(n11178), .B2(n19980), .ZN(
        n11379) );
  MUX2_X1 U13957 ( .A(n10978), .B(n10400), .S(n10625), .Z(n10979) );
  NAND2_X1 U13958 ( .A1(n10980), .A2(n14048), .ZN(n10981) );
  OR2_X1 U13959 ( .A1(n14043), .A2(n10981), .ZN(n10994) );
  NAND2_X1 U13960 ( .A1(n10625), .A2(n10984), .ZN(n11009) );
  NAND2_X1 U13961 ( .A1(n11009), .A2(n14058), .ZN(n10986) );
  NAND2_X1 U13962 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  NAND2_X1 U13963 ( .A1(n10983), .A2(n10987), .ZN(n10990) );
  OAI21_X1 U13964 ( .B1(n10988), .B2(n19368), .A(n10989), .ZN(n11013) );
  NAND4_X1 U13965 ( .A1(n10982), .A2(n10990), .A3(n10433), .A4(n11013), .ZN(
        n11008) );
  NOR2_X1 U13966 ( .A1(n11008), .A2(n10992), .ZN(n10993) );
  AND2_X1 U13967 ( .A1(n10994), .A2(n10993), .ZN(n14007) );
  OAI21_X1 U13968 ( .B1(n14043), .B2(n10197), .A(n14007), .ZN(n10995) );
  NOR2_X1 U13969 ( .A1(n11379), .A2(n10995), .ZN(n10996) );
  OAI211_X1 U13970 ( .C1(n10998), .C2(n13596), .A(n10997), .B(n10996), .ZN(
        n10999) );
  NAND2_X1 U13971 ( .A1(n11000), .A2(n11001), .ZN(n13561) );
  INV_X1 U13972 ( .A(n11002), .ZN(n14042) );
  NAND2_X1 U13973 ( .A1(n14042), .A2(n9772), .ZN(n11003) );
  NAND2_X1 U13974 ( .A1(n13561), .A2(n11003), .ZN(n11004) );
  NAND2_X1 U13975 ( .A1(n11351), .A2(n11004), .ZN(n16466) );
  NAND2_X1 U13976 ( .A1(n13374), .A2(n19326), .ZN(n11031) );
  NAND2_X1 U13977 ( .A1(n11005), .A2(n10625), .ZN(n11006) );
  NAND2_X1 U13978 ( .A1(n11006), .A2(n10436), .ZN(n11007) );
  NAND2_X1 U13979 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15502) );
  AND2_X1 U13980 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15672) );
  NOR2_X1 U13981 ( .A1(n16481), .A2(n16491), .ZN(n16480) );
  INV_X1 U13982 ( .A(n16480), .ZN(n11358) );
  NOR2_X1 U13983 ( .A1(n15755), .A2(n15750), .ZN(n15749) );
  NAND2_X1 U13984 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15749), .ZN(
        n11357) );
  INV_X1 U13985 ( .A(n11008), .ZN(n11011) );
  NOR2_X1 U13986 ( .A1(n13539), .A2(n11009), .ZN(n11010) );
  INV_X1 U13987 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19330) );
  NAND2_X1 U13988 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19322) );
  NOR2_X1 U13989 ( .A1(n19330), .A2(n19322), .ZN(n19311) );
  NAND2_X1 U13990 ( .A1(n19330), .A2(n19322), .ZN(n11355) );
  NAND2_X1 U13991 ( .A1(n11012), .A2(n9772), .ZN(n14014) );
  NAND2_X1 U13992 ( .A1(n14014), .A2(n11013), .ZN(n11019) );
  NAND2_X1 U13993 ( .A1(n10433), .A2(n19355), .ZN(n11016) );
  AOI22_X1 U13994 ( .A1(n19991), .A2(n11016), .B1(n14103), .B2(n10381), .ZN(
        n11017) );
  NAND2_X1 U13995 ( .A1(n11014), .A2(n11017), .ZN(n11018) );
  AOI21_X1 U13996 ( .B1(n19351), .B2(n11019), .A(n11018), .ZN(n11020) );
  OAI21_X1 U13997 ( .B1(n11021), .B2(n10433), .A(n11020), .ZN(n14021) );
  OR2_X1 U13998 ( .A1(n14021), .A2(n11022), .ZN(n11023) );
  NAND2_X1 U13999 ( .A1(n11351), .A2(n11023), .ZN(n15615) );
  OAI211_X1 U14000 ( .C1(n19314), .C2(n19311), .A(n11355), .B(n15762), .ZN(
        n16501) );
  NAND2_X1 U14001 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15711), .ZN(
        n15697) );
  INV_X1 U14002 ( .A(n15697), .ZN(n11024) );
  NAND3_X1 U14003 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11362) );
  INV_X1 U14004 ( .A(n11362), .ZN(n11025) );
  NAND2_X1 U14005 ( .A1(n16473), .A2(n11025), .ZN(n15609) );
  NAND3_X1 U14006 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11364) );
  NAND2_X1 U14007 ( .A1(n15597), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15585) );
  NAND2_X1 U14008 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15572) );
  NAND2_X1 U14009 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15535) );
  NAND2_X1 U14010 ( .A1(n15481), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14387) );
  AND2_X1 U14011 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11372) );
  INV_X1 U14012 ( .A(n11372), .ZN(n11026) );
  INV_X1 U14013 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11374) );
  NAND2_X1 U14014 ( .A1(n14364), .A2(n11374), .ZN(n11027) );
  NAND2_X1 U14015 ( .A1(n15730), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11384) );
  INV_X1 U14016 ( .A(n11029), .ZN(n11030) );
  INV_X1 U14017 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11046) );
  NAND2_X1 U14018 ( .A1(n11032), .A2(n11034), .ZN(n11044) );
  INV_X1 U14019 ( .A(n11044), .ZN(n11033) );
  NAND2_X1 U14020 ( .A1(n11033), .A2(n11049), .ZN(n11048) );
  NAND2_X1 U14021 ( .A1(n11048), .A2(n11034), .ZN(n11038) );
  NAND2_X1 U14022 ( .A1(n11036), .A2(n11035), .ZN(n11037) );
  XNOR2_X2 U14023 ( .A(n11038), .B(n11037), .ZN(n13669) );
  INV_X1 U14024 ( .A(n13669), .ZN(n14221) );
  OR2_X1 U14025 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  INV_X1 U14026 ( .A(n11113), .ZN(n19737) );
  NAND2_X1 U14027 ( .A1(n11116), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11045) );
  OAI211_X1 U14028 ( .C1(n11046), .C2(n19737), .A(n11045), .B(n9772), .ZN(
        n11047) );
  INV_X1 U14029 ( .A(n11047), .ZN(n11057) );
  NAND2_X1 U14030 ( .A1(n11050), .A2(n11058), .ZN(n11051) );
  AOI22_X1 U14031 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11079), .B1(
        n11124), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11056) );
  INV_X1 U14032 ( .A(n11060), .ZN(n11059) );
  AOI22_X1 U14033 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11111), .B1(
        n19375), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14034 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11125), .B1(
        n11115), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11054) );
  NAND2_X1 U14036 ( .A1(n11122), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11062) );
  AND2_X1 U14037 ( .A1(n11062), .A2(n11061), .ZN(n11071) );
  NOR2_X1 U14038 ( .A1(n11188), .A2(n11094), .ZN(n11073) );
  NAND2_X1 U14039 ( .A1(n10625), .A2(n11073), .ZN(n11098) );
  NAND2_X1 U14040 ( .A1(n11098), .A2(n11097), .ZN(n11074) );
  AOI22_X1 U14041 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11079), .B1(
        n11114), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11080) );
  AND2_X1 U14042 ( .A1(n11080), .A2(n9772), .ZN(n11084) );
  AOI22_X1 U14043 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11115), .B1(
        n11126), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U14044 ( .A1(n11090), .A2(n11089), .ZN(n11091) );
  NOR2_X1 U14045 ( .A1(n10031), .A2(n13676), .ZN(n13675) );
  INV_X1 U14046 ( .A(n11094), .ZN(n11092) );
  NAND2_X1 U14047 ( .A1(n13675), .A2(n11092), .ZN(n11096) );
  NOR2_X1 U14048 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n10031), .ZN(
        n11093) );
  XOR2_X1 U14049 ( .A(n11094), .B(n11093), .Z(n13534) );
  NAND2_X1 U14050 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13534), .ZN(
        n11095) );
  NAND2_X1 U14051 ( .A1(n11096), .A2(n11095), .ZN(n11099) );
  XOR2_X1 U14052 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11099), .Z(
        n14432) );
  XNOR2_X1 U14053 ( .A(n11098), .B(n11097), .ZN(n14430) );
  NAND2_X1 U14054 ( .A1(n14432), .A2(n14430), .ZN(n11101) );
  NAND2_X1 U14055 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11099), .ZN(
        n11100) );
  NAND2_X1 U14056 ( .A1(n11101), .A2(n11100), .ZN(n11102) );
  XNOR2_X1 U14057 ( .A(n11102), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14118) );
  NAND2_X1 U14058 ( .A1(n11102), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11103) );
  OAI21_X2 U14059 ( .B1(n14117), .B2(n14118), .A(n11103), .ZN(n11104) );
  XNOR2_X1 U14060 ( .A(n11109), .B(n11110), .ZN(n11105) );
  NAND2_X1 U14061 ( .A1(n11104), .A2(n11105), .ZN(n14149) );
  NAND2_X1 U14062 ( .A1(n14149), .A2(n15750), .ZN(n11108) );
  INV_X1 U14063 ( .A(n11104), .ZN(n11107) );
  INV_X1 U14064 ( .A(n11105), .ZN(n11106) );
  NAND2_X1 U14065 ( .A1(n11107), .A2(n11106), .ZN(n14150) );
  AOI22_X1 U14066 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19338), .B1(
        n11111), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14067 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n11112), .B1(
        n11113), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14068 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n11114), .B1(
        n11115), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14069 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n11079), .B1(
        n11116), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14070 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n15795), .B1(
        n11121), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14071 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11122), .B1(
        n11123), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14072 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19375), .B1(
        n11124), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14073 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n11125), .B1(
        n11126), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U14074 ( .A1(n11131), .A2(n10625), .ZN(n11132) );
  NAND2_X1 U14075 ( .A1(n11154), .A2(n15755), .ZN(n15742) );
  INV_X1 U14076 ( .A(n11161), .ZN(n11153) );
  INV_X1 U14077 ( .A(n11133), .ZN(n11136) );
  AOI22_X1 U14078 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19338), .B1(
        n11112), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U14079 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11122), .B1(
        n11121), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14080 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11115), .B1(
        n11126), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11138) );
  AOI22_X1 U14081 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11079), .B1(
        n11116), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11137) );
  NAND4_X1 U14082 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n11146) );
  AOI22_X1 U14083 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11111), .B1(
        n11113), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14084 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11123), .B1(
        n15795), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14085 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19375), .B1(
        n11124), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14086 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11114), .B1(
        n11125), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11141) );
  NAND4_X1 U14087 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11145) );
  NAND2_X1 U14088 ( .A1(n11147), .A2(n10625), .ZN(n11148) );
  NAND2_X1 U14089 ( .A1(n11151), .A2(n11158), .ZN(n11152) );
  NAND2_X1 U14090 ( .A1(n11153), .A2(n11208), .ZN(n11157) );
  INV_X1 U14091 ( .A(n11154), .ZN(n11179) );
  NAND2_X1 U14092 ( .A1(n11208), .A2(n15743), .ZN(n11155) );
  NAND2_X1 U14093 ( .A1(n11155), .A2(n11161), .ZN(n11156) );
  NAND2_X1 U14094 ( .A1(n11157), .A2(n11156), .ZN(n11160) );
  NAND2_X1 U14095 ( .A1(n15746), .A2(n11158), .ZN(n11159) );
  NAND2_X1 U14096 ( .A1(n11160), .A2(n11159), .ZN(n15734) );
  NAND2_X1 U14097 ( .A1(n15747), .A2(n15743), .ZN(n11162) );
  NAND2_X1 U14098 ( .A1(n11162), .A2(n11208), .ZN(n11163) );
  NAND2_X1 U14099 ( .A1(n15470), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15471) );
  INV_X1 U14100 ( .A(n11166), .ZN(n11167) );
  NAND2_X1 U14101 ( .A1(n11168), .A2(n11167), .ZN(n16437) );
  INV_X1 U14102 ( .A(n11165), .ZN(n11171) );
  AND2_X1 U14103 ( .A1(n10137), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11170) );
  NAND2_X1 U14104 ( .A1(n11171), .A2(n11170), .ZN(n16439) );
  OR2_X1 U14105 ( .A1(n11362), .A2(n15673), .ZN(n11174) );
  INV_X1 U14106 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15611) );
  INV_X1 U14107 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15423) );
  OR2_X1 U14108 ( .A1(n11175), .A2(n15564), .ZN(n15342) );
  OR2_X1 U14109 ( .A1(n11308), .A2(n15342), .ZN(n11176) );
  NOR2_X1 U14110 ( .A1(n11176), .A2(n15572), .ZN(n15332) );
  AND2_X1 U14111 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15332), .ZN(
        n11177) );
  XNOR2_X1 U14112 ( .A(n15298), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11388) );
  INV_X1 U14113 ( .A(n11178), .ZN(n19981) );
  OR2_X1 U14114 ( .A1(n11388), .A2(n16496), .ZN(n11377) );
  OR2_X1 U14115 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  NAND2_X1 U14116 ( .A1(n11180), .A2(n11183), .ZN(n19165) );
  NAND2_X1 U14117 ( .A1(n11196), .A2(n11184), .ZN(n11185) );
  NAND2_X1 U14118 ( .A1(n11203), .A2(n11185), .ZN(n14184) );
  OAI21_X1 U14119 ( .B1(n14117), .B2(n10137), .A(n14184), .ZN(n11201) );
  MUX2_X1 U14120 ( .A(n11188), .B(n11187), .S(n11186), .Z(n11191) );
  AOI21_X1 U14121 ( .B1(n11191), .B2(n11190), .A(n11189), .ZN(n19199) );
  NAND2_X1 U14122 ( .A1(n19199), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13673) );
  AND3_X1 U14123 ( .A1(n10904), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11192) );
  OR2_X1 U14124 ( .A1(n11194), .A2(n11192), .ZN(n15089) );
  NOR2_X1 U14125 ( .A1(n13673), .A2(n15089), .ZN(n11193) );
  NAND2_X1 U14126 ( .A1(n13673), .A2(n15089), .ZN(n13532) );
  OAI21_X1 U14127 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11193), .A(
        n13532), .ZN(n14423) );
  OR2_X1 U14128 ( .A1(n11195), .A2(n11194), .ZN(n11197) );
  NAND2_X1 U14129 ( .A1(n11197), .A2(n11196), .ZN(n14222) );
  XNOR2_X1 U14130 ( .A(n14222), .B(n19330), .ZN(n14422) );
  OR2_X1 U14131 ( .A1(n14423), .A2(n14422), .ZN(n14425) );
  INV_X1 U14132 ( .A(n14222), .ZN(n11198) );
  NAND2_X1 U14133 ( .A1(n11198), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11199) );
  NAND2_X1 U14134 ( .A1(n14425), .A2(n11199), .ZN(n14115) );
  INV_X1 U14135 ( .A(n14115), .ZN(n11200) );
  XNOR2_X1 U14136 ( .A(n11203), .B(n11202), .ZN(n19184) );
  INV_X1 U14137 ( .A(n19184), .ZN(n11204) );
  NAND2_X1 U14138 ( .A1(n11205), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11206) );
  NAND2_X1 U14139 ( .A1(n11207), .A2(n11206), .ZN(n15725) );
  NAND2_X1 U14140 ( .A1(n11208), .A2(n11169), .ZN(n11211) );
  NAND2_X1 U14141 ( .A1(n11180), .A2(n11209), .ZN(n11210) );
  NAND2_X1 U14142 ( .A1(n11219), .A2(n11210), .ZN(n19153) );
  NAND2_X1 U14143 ( .A1(n11212), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11213) );
  NOR2_X1 U14144 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  OR2_X1 U14145 ( .A1(n11225), .A2(n11216), .ZN(n19131) );
  NOR2_X1 U14146 ( .A1(n19131), .A2(n11169), .ZN(n11221) );
  NAND2_X1 U14147 ( .A1(n11221), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16431) );
  INV_X1 U14148 ( .A(n11217), .ZN(n11218) );
  XNOR2_X1 U14149 ( .A(n11219), .B(n11218), .ZN(n19143) );
  NAND2_X1 U14150 ( .A1(n19143), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16432) );
  NAND2_X1 U14151 ( .A1(n16431), .A2(n16432), .ZN(n11220) );
  INV_X1 U14152 ( .A(n11221), .ZN(n11222) );
  NAND2_X1 U14153 ( .A1(n11222), .A2(n16491), .ZN(n16430) );
  INV_X1 U14154 ( .A(n19143), .ZN(n11223) );
  NAND2_X1 U14155 ( .A1(n11223), .A2(n16481), .ZN(n16434) );
  AND2_X1 U14156 ( .A1(n16430), .A2(n16434), .ZN(n11224) );
  INV_X1 U14157 ( .A(n11232), .ZN(n11228) );
  NAND2_X1 U14158 ( .A1(n10904), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11226) );
  MUX2_X1 U14159 ( .A(n11226), .B(n10904), .S(n11225), .Z(n11227) );
  NAND2_X1 U14160 ( .A1(n11228), .A2(n11227), .ZN(n19120) );
  OAI21_X1 U14161 ( .B1(n19120), .B2(n11169), .A(n15710), .ZN(n15460) );
  NOR2_X1 U14162 ( .A1(n11232), .A2(n19111), .ZN(n11229) );
  NAND2_X1 U14163 ( .A1(n10904), .A2(n11229), .ZN(n11230) );
  NAND2_X1 U14164 ( .A1(n11321), .A2(n11230), .ZN(n11231) );
  AOI21_X1 U14165 ( .B1(n11232), .B2(n19111), .A(n11231), .ZN(n19109) );
  AOI21_X1 U14166 ( .B1(n19109), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15689) );
  INV_X1 U14167 ( .A(n19109), .ZN(n11234) );
  OR2_X1 U14168 ( .A1(n11169), .A2(n15696), .ZN(n11233) );
  INV_X1 U14169 ( .A(n19120), .ZN(n11236) );
  NOR2_X1 U14170 ( .A1(n11169), .A2(n15710), .ZN(n11235) );
  NAND2_X1 U14171 ( .A1(n11236), .A2(n11235), .ZN(n15687) );
  INV_X1 U14172 ( .A(n15687), .ZN(n11237) );
  NAND2_X1 U14173 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n11238), .ZN(n11239) );
  NOR2_X1 U14174 ( .A1(n10903), .A2(n11239), .ZN(n11240) );
  NOR2_X1 U14175 ( .A1(n11241), .A2(n11240), .ZN(n13448) );
  NAND2_X1 U14176 ( .A1(n13448), .A2(n10137), .ZN(n11244) );
  NOR2_X1 U14177 ( .A1(n11244), .A2(n15673), .ZN(n15683) );
  INV_X1 U14178 ( .A(n15683), .ZN(n11242) );
  NAND2_X1 U14179 ( .A1(n11244), .A2(n15673), .ZN(n16407) );
  INV_X1 U14180 ( .A(n11245), .ZN(n11247) );
  NAND2_X1 U14181 ( .A1(n11247), .A2(n11246), .ZN(n11248) );
  AND2_X1 U14182 ( .A1(n11263), .A2(n11248), .ZN(n19098) );
  NAND2_X1 U14183 ( .A1(n19098), .A2(n10137), .ZN(n11251) );
  NAND2_X1 U14184 ( .A1(n11251), .A2(n16472), .ZN(n11250) );
  AND2_X1 U14185 ( .A1(n16407), .A2(n11250), .ZN(n11249) );
  INV_X1 U14186 ( .A(n11250), .ZN(n11252) );
  XNOR2_X1 U14187 ( .A(n11251), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16409) );
  OR2_X1 U14188 ( .A1(n11252), .A2(n16409), .ZN(n11253) );
  NAND2_X1 U14189 ( .A1(n10904), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11254) );
  XNOR2_X1 U14190 ( .A(n9846), .B(n11254), .ZN(n19006) );
  NAND2_X1 U14191 ( .A1(n19006), .A2(n10137), .ZN(n11296) );
  AND2_X1 U14192 ( .A1(n11296), .A2(n15575), .ZN(n15388) );
  INV_X1 U14193 ( .A(n11255), .ZN(n11274) );
  NAND2_X1 U14194 ( .A1(n11257), .A2(n11256), .ZN(n11258) );
  NAND2_X1 U14195 ( .A1(n11274), .A2(n11258), .ZN(n19043) );
  NOR2_X1 U14196 ( .A1(n19043), .A2(n11169), .ZN(n11291) );
  NOR2_X1 U14197 ( .A1(n11291), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15370) );
  INV_X1 U14198 ( .A(n11259), .ZN(n11260) );
  XNOR2_X1 U14199 ( .A(n11261), .B(n11260), .ZN(n19067) );
  AOI21_X1 U14200 ( .B1(n19067), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15439) );
  NAND2_X1 U14201 ( .A1(n11263), .A2(n11262), .ZN(n11264) );
  AND2_X1 U14202 ( .A1(n9848), .A2(n11264), .ZN(n19086) );
  AOI21_X1 U14203 ( .B1(n19086), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15449) );
  XNOR2_X1 U14204 ( .A(n9848), .B(n11265), .ZN(n19077) );
  AOI21_X1 U14205 ( .B1(n19077), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15646) );
  NOR4_X1 U14206 ( .A1(n15370), .A2(n15439), .A3(n15449), .A4(n15646), .ZN(
        n11280) );
  MUX2_X1 U14207 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n10214), .S(n11266), .Z(
        n11267) );
  NAND2_X1 U14208 ( .A1(n11267), .A2(n11321), .ZN(n19052) );
  OAI21_X1 U14209 ( .B1(n19052), .B2(n11169), .A(n15611), .ZN(n11270) );
  INV_X1 U14210 ( .A(n19052), .ZN(n11269) );
  NOR2_X1 U14211 ( .A1(n11169), .A2(n15611), .ZN(n11268) );
  NAND2_X1 U14212 ( .A1(n11269), .A2(n11268), .ZN(n15369) );
  INV_X1 U14213 ( .A(n11271), .ZN(n11278) );
  INV_X1 U14214 ( .A(n11272), .ZN(n11273) );
  NAND2_X1 U14215 ( .A1(n11274), .A2(n11273), .ZN(n11275) );
  NAND2_X1 U14216 ( .A1(n11278), .A2(n11275), .ZN(n19030) );
  OR2_X1 U14217 ( .A1(n19030), .A2(n11169), .ZN(n11276) );
  NAND2_X1 U14218 ( .A1(n11276), .A2(n15596), .ZN(n15410) );
  NAND2_X1 U14219 ( .A1(n11278), .A2(n10022), .ZN(n11279) );
  NAND2_X1 U14220 ( .A1(n9846), .A2(n11279), .ZN(n19022) );
  OAI21_X1 U14221 ( .B1(n19022), .B2(n11169), .A(n15574), .ZN(n15400) );
  INV_X1 U14222 ( .A(n11282), .ZN(n11285) );
  NAND3_X1 U14223 ( .A1(n11283), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n10904), 
        .ZN(n11284) );
  AOI21_X1 U14224 ( .B1(n15086), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15378) );
  NOR2_X1 U14225 ( .A1(n11169), .A2(n15564), .ZN(n11287) );
  NAND2_X1 U14226 ( .A1(n15086), .A2(n11287), .ZN(n15376) );
  INV_X1 U14227 ( .A(n19022), .ZN(n11289) );
  NOR2_X1 U14228 ( .A1(n11169), .A2(n15574), .ZN(n11288) );
  NAND2_X1 U14229 ( .A1(n11289), .A2(n11288), .ZN(n15399) );
  OR2_X1 U14230 ( .A1(n11169), .A2(n15596), .ZN(n11290) );
  OR2_X1 U14231 ( .A1(n19030), .A2(n11290), .ZN(n15409) );
  AND2_X1 U14232 ( .A1(n15399), .A2(n15409), .ZN(n15373) );
  NAND2_X1 U14233 ( .A1(n11291), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15372) );
  INV_X1 U14234 ( .A(n19067), .ZN(n11292) );
  INV_X1 U14235 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15633) );
  NOR2_X1 U14236 ( .A1(n11169), .A2(n15655), .ZN(n11293) );
  NAND2_X1 U14237 ( .A1(n19077), .A2(n11293), .ZN(n15367) );
  NOR2_X1 U14238 ( .A1(n11169), .A2(n15661), .ZN(n11294) );
  NAND2_X1 U14239 ( .A1(n19086), .A2(n11294), .ZN(n15447) );
  AND4_X1 U14240 ( .A1(n15372), .A2(n15437), .A3(n15367), .A4(n15447), .ZN(
        n11295) );
  NAND4_X1 U14241 ( .A1(n15376), .A2(n15373), .A3(n11295), .A4(n15369), .ZN(
        n11298) );
  INV_X1 U14242 ( .A(n11296), .ZN(n11297) );
  INV_X1 U14243 ( .A(n11299), .ZN(n11300) );
  NAND2_X1 U14244 ( .A1(n11301), .A2(n11300), .ZN(n11302) );
  AND2_X1 U14245 ( .A1(n11305), .A2(n11302), .ZN(n15057) );
  AOI21_X1 U14246 ( .B1(n15057), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15358) );
  NAND3_X1 U14247 ( .A1(n15057), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n10137), .ZN(n15357) );
  OAI21_X2 U14248 ( .B1(n15355), .B2(n15358), .A(n15357), .ZN(n15345) );
  INV_X1 U14249 ( .A(n11303), .ZN(n11310) );
  NAND2_X1 U14250 ( .A1(n11305), .A2(n11304), .ZN(n11306) );
  NAND2_X1 U14251 ( .A1(n11310), .A2(n11306), .ZN(n15056) );
  XNOR2_X1 U14252 ( .A(n11307), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15346) );
  NOR3_X1 U14253 ( .A1(n15056), .A2(n11169), .A3(n11308), .ZN(n11309) );
  NOR2_X1 U14254 ( .A1(n10903), .A2(n15136), .ZN(n11311) );
  MUX2_X1 U14255 ( .A(n15136), .B(n11311), .S(n11310), .Z(n11313) );
  INV_X1 U14256 ( .A(n11321), .ZN(n11312) );
  NOR2_X1 U14257 ( .A1(n11313), .A2(n11312), .ZN(n16387) );
  NAND2_X1 U14258 ( .A1(n16387), .A2(n10137), .ZN(n15334) );
  INV_X1 U14259 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11368) );
  INV_X1 U14260 ( .A(n11314), .ZN(n14340) );
  NAND3_X1 U14261 ( .A1(n10904), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n11315), 
        .ZN(n11316) );
  NAND2_X1 U14262 ( .A1(n14340), .A2(n11316), .ZN(n16365) );
  NOR3_X1 U14263 ( .A1(n16365), .A2(n11169), .A3(n15508), .ZN(n11337) );
  INV_X1 U14264 ( .A(n16365), .ZN(n11317) );
  AOI21_X1 U14265 ( .B1(n11317), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11318) );
  NOR2_X1 U14266 ( .A1(n11337), .A2(n11318), .ZN(n15315) );
  NOR2_X1 U14267 ( .A1(n11323), .A2(n14329), .ZN(n11319) );
  NAND2_X1 U14268 ( .A1(n10904), .A2(n11319), .ZN(n11320) );
  NAND2_X1 U14269 ( .A1(n11321), .A2(n11320), .ZN(n11322) );
  AOI21_X1 U14270 ( .B1(n11323), .B2(n14329), .A(n11322), .ZN(n16377) );
  INV_X1 U14271 ( .A(n11324), .ZN(n11326) );
  NAND2_X1 U14272 ( .A1(n11326), .A2(n11325), .ZN(n11327) );
  INV_X1 U14273 ( .A(n11328), .ZN(n11329) );
  NAND2_X1 U14274 ( .A1(n11330), .A2(n11329), .ZN(n11331) );
  AOI21_X1 U14275 ( .B1(n21140), .B2(n15479), .A(n14380), .ZN(n11332) );
  INV_X1 U14276 ( .A(n11332), .ZN(n11333) );
  NAND2_X1 U14277 ( .A1(n14380), .A2(n21140), .ZN(n11334) );
  INV_X1 U14278 ( .A(n11335), .ZN(n11336) );
  INV_X1 U14279 ( .A(n11338), .ZN(n11339) );
  INV_X1 U14280 ( .A(n11341), .ZN(n16337) );
  NAND3_X1 U14281 ( .A1(n16337), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10137), .ZN(n15293) );
  AND2_X1 U14282 ( .A1(n14374), .A2(n15293), .ZN(n11343) );
  OAI21_X1 U14283 ( .B1(n11341), .B2(n11169), .A(n15299), .ZN(n15294) );
  INV_X1 U14284 ( .A(n15294), .ZN(n11342) );
  AOI21_X1 U14285 ( .B1(n11344), .B2(n10137), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14332) );
  INV_X1 U14286 ( .A(n14332), .ZN(n11346) );
  NAND2_X1 U14287 ( .A1(n11346), .A2(n14334), .ZN(n11347) );
  XNOR2_X1 U14288 ( .A(n11348), .B(n11347), .ZN(n11380) );
  INV_X1 U14289 ( .A(n14057), .ZN(n11350) );
  AND2_X1 U14290 ( .A1(n11350), .A2(n11349), .ZN(n19982) );
  NAND2_X1 U14291 ( .A1(n11351), .A2(n19982), .ZN(n15761) );
  INV_X1 U14292 ( .A(n15615), .ZN(n11354) );
  INV_X1 U14293 ( .A(n11351), .ZN(n11353) );
  NAND2_X1 U14294 ( .A1(n11353), .A2(n19151), .ZN(n13672) );
  INV_X1 U14295 ( .A(n13672), .ZN(n15766) );
  AOI21_X1 U14296 ( .B1(n11354), .B2(n19322), .A(n15766), .ZN(n19331) );
  NAND2_X1 U14297 ( .A1(n11354), .A2(n19330), .ZN(n19323) );
  INV_X1 U14298 ( .A(n11355), .ZN(n19312) );
  NAND2_X1 U14299 ( .A1(n19314), .A2(n19312), .ZN(n11356) );
  NAND4_X1 U14300 ( .A1(n19331), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19323), .A4(n11356), .ZN(n16492) );
  INV_X1 U14301 ( .A(n15762), .ZN(n15616) );
  NAND2_X1 U14302 ( .A1(n15616), .A2(n19331), .ZN(n14154) );
  OAI21_X1 U14303 ( .B1(n16492), .B2(n11357), .A(n14154), .ZN(n16490) );
  NAND2_X1 U14304 ( .A1(n15762), .A2(n11358), .ZN(n11359) );
  NAND2_X1 U14305 ( .A1(n15672), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11360) );
  NAND2_X1 U14306 ( .A1(n15762), .A2(n11360), .ZN(n11361) );
  NAND2_X1 U14307 ( .A1(n15762), .A2(n11362), .ZN(n11363) );
  OAI21_X1 U14308 ( .B1(n11364), .B2(n15596), .A(n15762), .ZN(n11365) );
  NAND2_X1 U14309 ( .A1(n15632), .A2(n11365), .ZN(n15602) );
  AND2_X1 U14310 ( .A1(n15762), .A2(n15572), .ZN(n11366) );
  NOR2_X1 U14311 ( .A1(n15602), .A2(n11366), .ZN(n15565) );
  NAND2_X1 U14312 ( .A1(n15762), .A2(n15564), .ZN(n11367) );
  NAND2_X1 U14313 ( .A1(n15565), .A2(n11367), .ZN(n15546) );
  AND2_X1 U14314 ( .A1(n15762), .A2(n15535), .ZN(n11369) );
  NAND2_X1 U14315 ( .A1(n15565), .A2(n15616), .ZN(n11370) );
  NAND2_X1 U14316 ( .A1(n15525), .A2(n11370), .ZN(n15515) );
  NAND2_X1 U14317 ( .A1(n11370), .A2(n15502), .ZN(n11371) );
  NAND2_X1 U14318 ( .A1(n15515), .A2(n11371), .ZN(n15497) );
  AOI21_X1 U14319 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11372), .A(
        n15616), .ZN(n11373) );
  NOR2_X1 U14320 ( .A1(n15497), .A2(n11373), .ZN(n14358) );
  NOR2_X1 U14321 ( .A1(n14358), .A2(n11374), .ZN(n11375) );
  AOI21_X1 U14322 ( .B1(n11380), .B2(n19316), .A(n11375), .ZN(n11376) );
  NAND3_X1 U14323 ( .A1(n10199), .A2(n11377), .A3(n11376), .ZN(P2_U3016) );
  AND2_X1 U14324 ( .A1(n14103), .A2(n16503), .ZN(n11378) );
  NAND2_X1 U14325 ( .A1(n11379), .A2(n11378), .ZN(n18987) );
  OR2_X1 U14326 ( .A1(n18987), .A2(n10625), .ZN(n19305) );
  INV_X1 U14327 ( .A(n19305), .ZN(n19283) );
  NAND2_X1 U14328 ( .A1(n11380), .A2(n19283), .ZN(n11391) );
  NOR2_X2 U14329 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19942) );
  OR2_X1 U14330 ( .A1(n19942), .A2(n19941), .ZN(n19959) );
  NAND2_X1 U14331 ( .A1(n19959), .A2(n16509), .ZN(n11381) );
  AND2_X1 U14332 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19960) );
  NOR2_X1 U14333 ( .A1(n11028), .A2(n19289), .ZN(n11387) );
  NAND2_X1 U14334 ( .A1(n16509), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13069) );
  NAND2_X1 U14335 ( .A1(n19781), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U14336 ( .A1(n13069), .A2(n11382), .ZN(n19295) );
  NAND2_X1 U14337 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11383) );
  OAI211_X1 U14338 ( .C1(n19294), .C2(n11385), .A(n11384), .B(n11383), .ZN(
        n11386) );
  OR2_X1 U14339 ( .A1(n18987), .A2(n9772), .ZN(n16456) );
  NAND3_X1 U14340 ( .A1(n11391), .A2(n11390), .A3(n11389), .ZN(P2_U2984) );
  AOI22_X1 U14341 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11396) );
  INV_X2 U14342 ( .A(n10220), .ZN(n15891) );
  AOI22_X1 U14343 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14344 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11394) );
  INV_X2 U14345 ( .A(n11591), .ZN(n17294) );
  AOI22_X1 U14346 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11393) );
  NAND4_X1 U14347 ( .A1(n11396), .A2(n11395), .A3(n11394), .A4(n11393), .ZN(
        n11408) );
  AOI22_X1 U14348 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14349 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11405) );
  INV_X2 U14350 ( .A(n10200), .ZN(n17286) );
  NOR2_X2 U14351 ( .A1(n11398), .A2(n11401), .ZN(n15819) );
  AOI22_X1 U14352 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11404) );
  NOR2_X1 U14353 ( .A1(n11400), .A2(n11399), .ZN(n11455) );
  AOI22_X1 U14354 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11403) );
  NAND4_X1 U14355 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11407) );
  AOI22_X1 U14356 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14357 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14358 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14359 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11409) );
  NAND4_X1 U14360 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n11419) );
  AOI22_X1 U14361 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14362 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14363 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11415) );
  INV_X2 U14364 ( .A(n9850), .ZN(n17287) );
  AOI22_X1 U14365 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11414) );
  NAND4_X1 U14366 ( .A1(n11417), .A2(n11416), .A3(n11415), .A4(n11414), .ZN(
        n11418) );
  AOI22_X1 U14367 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14368 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14369 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14370 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11420) );
  NAND4_X1 U14371 ( .A1(n11423), .A2(n11422), .A3(n11421), .A4(n11420), .ZN(
        n11429) );
  INV_X2 U14372 ( .A(n9849), .ZN(n17276) );
  AOI22_X1 U14373 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14374 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14375 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17249), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14376 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U14377 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11428) );
  AOI22_X1 U14378 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11430) );
  OAI21_X1 U14379 ( .B1(n16967), .B2(n18313), .A(n11430), .ZN(n11435) );
  AOI22_X1 U14380 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14381 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11477), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11432) );
  NAND3_X1 U14382 ( .A1(n11433), .A2(n11432), .A3(n11431), .ZN(n11434) );
  AOI22_X1 U14383 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11436), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14384 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14385 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14386 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14387 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11443) );
  INV_X1 U14388 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21223) );
  AOI22_X1 U14389 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11444) );
  OAI21_X1 U14390 ( .B1(n11591), .B2(n21223), .A(n11444), .ZN(n11445) );
  INV_X2 U14391 ( .A(n11466), .ZN(n17275) );
  AOI22_X1 U14392 ( .A1(n17275), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14393 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14394 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11447) );
  NAND3_X1 U14395 ( .A1(n11449), .A2(n11448), .A3(n11447), .ZN(n11450) );
  INV_X2 U14396 ( .A(n11602), .ZN(n17259) );
  AOI22_X1 U14397 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14398 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11452) );
  NAND3_X1 U14399 ( .A1(n11454), .A2(n11453), .A3(n11452), .ZN(n11646) );
  AOI22_X1 U14400 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14401 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11464) );
  INV_X1 U14402 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21134) );
  AOI22_X1 U14403 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11456) );
  OAI21_X1 U14404 ( .B1(n11466), .B2(n21134), .A(n11456), .ZN(n11462) );
  AOI22_X1 U14405 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14406 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14407 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14408 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U14409 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11461) );
  AOI211_X1 U14410 ( .C1(n17269), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n11462), .B(n11461), .ZN(n11463) );
  NAND3_X1 U14411 ( .A1(n11465), .A2(n11464), .A3(n11463), .ZN(n11647) );
  NAND2_X1 U14412 ( .A1(n11496), .A2(n11647), .ZN(n11499) );
  INV_X2 U14413 ( .A(n15858), .ZN(n17288) );
  AOI22_X1 U14414 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17288), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11470) );
  INV_X2 U14415 ( .A(n11466), .ZN(n17250) );
  AOI22_X1 U14416 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11469) );
  INV_X2 U14417 ( .A(n10220), .ZN(n17270) );
  AOI22_X1 U14418 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14419 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11467) );
  NAND4_X1 U14420 ( .A1(n11470), .A2(n11469), .A3(n11468), .A4(n11467), .ZN(
        n11476) );
  AOI22_X1 U14421 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14422 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17269), .ZN(n11473) );
  AOI22_X1 U14423 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14424 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17249), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11471) );
  NAND4_X1 U14425 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11475) );
  INV_X1 U14426 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17622) );
  INV_X1 U14427 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16551) );
  NOR2_X1 U14428 ( .A1(n17622), .A2(n16551), .ZN(n16527) );
  NAND2_X1 U14429 ( .A1(n16527), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13017) );
  INV_X1 U14430 ( .A(n13017), .ZN(n11684) );
  INV_X1 U14431 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17996) );
  INV_X1 U14432 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18246) );
  AOI22_X1 U14433 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14434 ( .A1(n11478), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11477), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14435 ( .A1(n11479), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14436 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14437 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14438 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11485) );
  INV_X1 U14439 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n21158) );
  AOI22_X1 U14440 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11487) );
  OAI21_X1 U14441 ( .B1(n9822), .B2(n21158), .A(n11487), .ZN(n11488) );
  INV_X1 U14442 ( .A(n11488), .ZN(n11489) );
  NAND3_X1 U14443 ( .A1(n10209), .A2(n10205), .A3(n11489), .ZN(n17959) );
  NOR2_X1 U14444 ( .A1(n17951), .A2(n17953), .ZN(n17952) );
  INV_X1 U14445 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18923) );
  INV_X1 U14446 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18278) );
  XNOR2_X1 U14447 ( .A(n11492), .B(n17475), .ZN(n11493) );
  NOR2_X1 U14448 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  INV_X1 U14449 ( .A(n11647), .ZN(n17471) );
  XNOR2_X1 U14450 ( .A(n11496), .B(n17471), .ZN(n11497) );
  XNOR2_X1 U14451 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11497), .ZN(
        n17920) );
  AND2_X1 U14452 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11497), .ZN(
        n11498) );
  INV_X1 U14453 ( .A(n17468), .ZN(n11648) );
  XOR2_X1 U14454 ( .A(n11499), .B(n11648), .Z(n17904) );
  XNOR2_X1 U14455 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11501), .ZN(
        n17890) );
  OAI21_X1 U14456 ( .B1(n16541), .B2(n16534), .A(n17838), .ZN(n11502) );
  XNOR2_X1 U14457 ( .A(n11503), .B(n11502), .ZN(n17886) );
  INV_X1 U14458 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18222) );
  NOR2_X1 U14459 ( .A1(n17886), .A2(n18222), .ZN(n17885) );
  NOR2_X1 U14460 ( .A1(n11503), .A2(n11502), .ZN(n11504) );
  INV_X1 U14461 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18193) );
  NAND2_X1 U14462 ( .A1(n11505), .A2(n18193), .ZN(n11507) );
  INV_X2 U14463 ( .A(n11682), .ZN(n18170) );
  NAND2_X1 U14464 ( .A1(n18170), .A2(n11507), .ZN(n17877) );
  NAND2_X1 U14465 ( .A1(n18205), .A2(n17873), .ZN(n17872) );
  INV_X1 U14466 ( .A(n17837), .ZN(n11506) );
  INV_X1 U14467 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18160) );
  INV_X1 U14468 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18189) );
  INV_X1 U14469 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17836) );
  NOR2_X1 U14470 ( .A1(n18189), .A2(n17836), .ZN(n18174) );
  NAND2_X1 U14471 ( .A1(n18174), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18159) );
  INV_X1 U14472 ( .A(n18159), .ZN(n18141) );
  NAND3_X1 U14473 ( .A1(n18141), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17777) );
  OR2_X1 U14474 ( .A1(n18160), .A2(n17777), .ZN(n18126) );
  INV_X1 U14475 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18115) );
  NOR2_X1 U14476 ( .A1(n18126), .A2(n18115), .ZN(n18074) );
  INV_X1 U14477 ( .A(n18074), .ZN(n16538) );
  INV_X1 U14478 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21097) );
  INV_X1 U14479 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18146) );
  NOR2_X1 U14480 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11509) );
  AOI21_X1 U14481 ( .B1(n17791), .B2(n11509), .A(n17873), .ZN(n17758) );
  INV_X1 U14482 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18089) );
  NOR2_X1 U14483 ( .A1(n21097), .A2(n18089), .ZN(n17743) );
  NAND2_X1 U14484 ( .A1(n17743), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18043) );
  INV_X1 U14485 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17707) );
  NAND2_X1 U14486 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17704) );
  NOR2_X1 U14487 ( .A1(n17707), .A2(n17704), .ZN(n13013) );
  NAND2_X1 U14488 ( .A1(n13013), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11516) );
  NOR2_X1 U14489 ( .A1(n18043), .A2(n11516), .ZN(n18018) );
  AND2_X1 U14490 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18018), .ZN(
        n17650) );
  INV_X1 U14491 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18070) );
  NAND2_X1 U14492 ( .A1(n17744), .A2(n18070), .ZN(n11511) );
  NOR2_X1 U14493 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11511), .ZN(
        n17702) );
  NAND2_X1 U14494 ( .A1(n17702), .A2(n17707), .ZN(n17687) );
  NOR3_X1 U14495 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17687), .ZN(n11512) );
  NAND2_X1 U14496 ( .A1(n17743), .A2(n11515), .ZN(n17700) );
  INV_X1 U14497 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17737) );
  NOR2_X1 U14498 ( .A1(n17737), .A2(n11516), .ZN(n13012) );
  INV_X1 U14499 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18023) );
  NOR2_X1 U14500 ( .A1(n17636), .A2(n17838), .ZN(n11518) );
  INV_X1 U14501 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17985) );
  NOR2_X1 U14502 ( .A1(n17996), .A2(n17985), .ZN(n17972) );
  INV_X1 U14503 ( .A(n17972), .ZN(n11683) );
  AND2_X1 U14504 ( .A1(n17873), .A2(n11683), .ZN(n11517) );
  NAND2_X1 U14505 ( .A1(n11520), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16532) );
  NAND2_X1 U14506 ( .A1(n11684), .A2(n15924), .ZN(n12984) );
  INV_X1 U14507 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16518) );
  NAND2_X1 U14508 ( .A1(n12982), .A2(n12983), .ZN(n11522) );
  AOI22_X1 U14509 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14510 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11525) );
  BUF_X1 U14511 ( .A(n15826), .Z(n15869) );
  AOI22_X1 U14512 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14513 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11523) );
  NAND4_X1 U14514 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n11532) );
  INV_X2 U14515 ( .A(n10200), .ZN(n17195) );
  AOI22_X1 U14516 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14517 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14518 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14519 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11527) );
  NAND4_X1 U14520 ( .A1(n11530), .A2(n11529), .A3(n11528), .A4(n11527), .ZN(
        n11531) );
  INV_X1 U14521 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18973) );
  INV_X1 U14522 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18921) );
  NAND2_X1 U14523 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18921), .ZN(n18805) );
  NOR2_X1 U14524 ( .A1(n18973), .A2(n18805), .ZN(n18955) );
  AOI22_X1 U14525 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18579), .B2(n18934), .ZN(
        n11645) );
  NAND2_X1 U14526 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20991), .ZN(
        n11540) );
  NOR2_X1 U14527 ( .A1(n11645), .A2(n11540), .ZN(n11533) );
  AOI21_X1 U14528 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18579), .A(
        n11533), .ZN(n11535) );
  INV_X1 U14529 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U14530 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18298), .B2(n11534), .ZN(
        n11536) );
  XOR2_X1 U14531 ( .A(n11535), .B(n11536), .Z(n11544) );
  INV_X1 U14532 ( .A(n11544), .ZN(n11549) );
  INV_X1 U14533 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21096) );
  OR2_X1 U14534 ( .A1(n11536), .A2(n11535), .ZN(n11537) );
  OAI21_X1 U14535 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n11534), .A(
        n11537), .ZN(n11538) );
  OAI22_X1 U14536 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21096), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11538), .ZN(n11542) );
  NOR2_X1 U14537 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21096), .ZN(
        n11539) );
  NAND2_X1 U14538 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11538), .ZN(
        n11541) );
  AOI22_X1 U14539 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11542), .B1(
        n11539), .B2(n11541), .ZN(n11545) );
  OAI211_X1 U14540 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20991), .A(
        n11545), .B(n11540), .ZN(n11644) );
  XOR2_X1 U14541 ( .A(n11645), .B(n11540), .Z(n11548) );
  INV_X1 U14542 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16966) );
  AND2_X1 U14543 ( .A1(n11541), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11543) );
  OAI22_X1 U14544 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16966), .B1(
        n11543), .B2(n11542), .ZN(n11547) );
  AOI21_X1 U14545 ( .B1(n11545), .B2(n11544), .A(n11547), .ZN(n11643) );
  INV_X1 U14546 ( .A(n11643), .ZN(n11546) );
  OAI21_X1 U14547 ( .B1(n11549), .B2(n11644), .A(n18746), .ZN(n18753) );
  AOI22_X1 U14548 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14549 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14550 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14551 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11550) );
  NAND4_X1 U14552 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11559) );
  AOI22_X1 U14553 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14554 ( .A1(n15869), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14555 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14556 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11554) );
  NAND4_X1 U14557 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n11558) );
  AOI22_X1 U14558 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14559 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14560 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14561 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U14562 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11569) );
  AOI22_X1 U14563 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14564 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14565 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14566 ( .A1(n15869), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11564) );
  NAND4_X1 U14567 ( .A1(n11567), .A2(n11566), .A3(n11565), .A4(n11564), .ZN(
        n11568) );
  AOI22_X1 U14568 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14569 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14570 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14571 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11570) );
  NAND4_X1 U14572 ( .A1(n11573), .A2(n11572), .A3(n11571), .A4(n11570), .ZN(
        n11579) );
  AOI22_X1 U14573 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14574 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14575 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14576 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11574) );
  NAND4_X1 U14577 ( .A1(n11577), .A2(n11576), .A3(n11575), .A4(n11574), .ZN(
        n11578) );
  NOR2_X1 U14578 ( .A1(n18331), .A2(n18336), .ZN(n11634) );
  AOI22_X1 U14579 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14580 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11588) );
  INV_X1 U14581 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18310) );
  AOI22_X1 U14582 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11580) );
  OAI21_X1 U14583 ( .B1(n11591), .B2(n18310), .A(n11580), .ZN(n11586) );
  AOI22_X1 U14584 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14585 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14586 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14587 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11581) );
  NAND4_X1 U14588 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11585) );
  AOI22_X1 U14589 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14590 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11599) );
  INV_X1 U14591 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U14592 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11590) );
  OAI21_X1 U14593 ( .B1(n11591), .B2(n18329), .A(n11590), .ZN(n11597) );
  AOI22_X1 U14594 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14595 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14596 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14597 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14598 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11596) );
  AOI211_X1 U14599 ( .C1(n17259), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n11597), .B(n11596), .ZN(n11598) );
  NAND3_X1 U14600 ( .A1(n11600), .A2(n11599), .A3(n11598), .ZN(n13000) );
  NOR2_X1 U14601 ( .A1(n17492), .A2(n13000), .ZN(n12993) );
  AOI22_X1 U14602 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17275), .ZN(n11612) );
  AOI22_X1 U14603 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17270), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11611) );
  INV_X1 U14604 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n21066) );
  INV_X2 U14605 ( .A(n9850), .ZN(n17268) );
  AOI22_X1 U14606 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17268), .ZN(n11601) );
  OAI21_X1 U14607 ( .B1(n21066), .B2(n11602), .A(n11601), .ZN(n11603) );
  INV_X1 U14608 ( .A(n11603), .ZN(n11605) );
  AOI22_X1 U14609 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17195), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14610 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17295), .ZN(n11609) );
  AOI22_X1 U14611 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17294), .ZN(n11608) );
  AOI22_X1 U14612 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17252), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n11606), .ZN(n11607) );
  NAND4_X1 U14613 ( .A1(n18321), .A2(n11634), .A3(n12993), .A4(n17459), .ZN(
        n11635) );
  AOI22_X1 U14614 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14615 ( .A1(n15826), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11621) );
  INV_X1 U14616 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n21233) );
  AOI22_X1 U14617 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11613) );
  OAI21_X1 U14618 ( .B1(n9822), .B2(n21233), .A(n11613), .ZN(n11619) );
  AOI22_X1 U14619 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14620 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14621 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14622 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11614) );
  NAND4_X1 U14623 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11618) );
  AOI211_X1 U14624 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n11619), .B(n11618), .ZN(n11620) );
  NAND3_X1 U14625 ( .A1(n11622), .A2(n11621), .A3(n11620), .ZN(n12988) );
  NAND2_X1 U14626 ( .A1(n18315), .A2(n18321), .ZN(n18758) );
  INV_X1 U14627 ( .A(n18758), .ZN(n11623) );
  NOR2_X1 U14628 ( .A1(n18336), .A2(n17343), .ZN(n12992) );
  NAND2_X1 U14629 ( .A1(n11623), .A2(n12992), .ZN(n15885) );
  NOR2_X1 U14630 ( .A1(n15915), .A2(n17492), .ZN(n16010) );
  NAND2_X1 U14631 ( .A1(n16010), .A2(n17459), .ZN(n11626) );
  OAI21_X2 U14632 ( .B1(n15885), .B2(n11626), .A(n18748), .ZN(n11642) );
  INV_X1 U14633 ( .A(n18336), .ZN(n11624) );
  NOR2_X1 U14634 ( .A1(n18331), .A2(n11624), .ZN(n16014) );
  INV_X1 U14635 ( .A(n16014), .ZN(n18768) );
  OAI211_X1 U14636 ( .C1(n13000), .C2(n18768), .A(n11637), .B(n18315), .ZN(
        n11625) );
  INV_X1 U14637 ( .A(n11625), .ZN(n12995) );
  AND2_X1 U14638 ( .A1(n11637), .A2(n11626), .ZN(n11630) );
  NAND2_X1 U14639 ( .A1(n18315), .A2(n17343), .ZN(n12990) );
  NAND2_X1 U14640 ( .A1(n18961), .A2(n17492), .ZN(n11636) );
  NOR2_X1 U14641 ( .A1(n16013), .A2(n11636), .ZN(n12996) );
  AOI21_X1 U14642 ( .B1(n12990), .B2(n11631), .A(n12996), .ZN(n11628) );
  OAI21_X1 U14643 ( .B1(n18343), .B2(n11634), .A(n13000), .ZN(n11627) );
  OAI21_X1 U14644 ( .B1(n11628), .B2(n18321), .A(n11627), .ZN(n11629) );
  INV_X1 U14645 ( .A(n11631), .ZN(n11632) );
  NOR2_X1 U14646 ( .A1(n18336), .A2(n12990), .ZN(n13001) );
  OAI21_X1 U14647 ( .B1(n11632), .B2(n13001), .A(n18307), .ZN(n11633) );
  INV_X1 U14648 ( .A(n11642), .ZN(n11640) );
  INV_X4 U14649 ( .A(n18771), .ZN(n18763) );
  NAND2_X1 U14650 ( .A1(n11637), .A2(n11636), .ZN(n18975) );
  INV_X1 U14651 ( .A(n18975), .ZN(n18964) );
  NAND2_X1 U14652 ( .A1(n18336), .A2(n13000), .ZN(n18759) );
  NOR3_X1 U14653 ( .A1(n12991), .A2(n12990), .A3(n18759), .ZN(n15883) );
  NOR2_X1 U14654 ( .A1(n18961), .A2(n11638), .ZN(n11641) );
  AOI21_X1 U14655 ( .B1(n11641), .B2(n11640), .A(n11639), .ZN(n18757) );
  XOR2_X1 U14656 ( .A(n18961), .B(n18315), .Z(n12989) );
  OAI21_X1 U14657 ( .B1(n11645), .B2(n11644), .A(n11643), .ZN(n12999) );
  NAND2_X2 U14658 ( .A1(n18961), .A2(n18230), .ZN(n18750) );
  INV_X1 U14659 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18010) );
  NOR2_X1 U14660 ( .A1(n18023), .A2(n18010), .ZN(n17971) );
  NAND2_X1 U14661 ( .A1(n18018), .A2(n17971), .ZN(n17968) );
  INV_X1 U14662 ( .A(n11646), .ZN(n17479) );
  NOR2_X1 U14663 ( .A1(n17475), .A2(n11651), .ZN(n11662) );
  AND2_X1 U14664 ( .A1(n11647), .A2(n11662), .ZN(n11649) );
  NAND2_X1 U14665 ( .A1(n11649), .A2(n11648), .ZN(n11665) );
  NOR2_X1 U14666 ( .A1(n17465), .A2(n11665), .ZN(n11669) );
  NAND2_X1 U14667 ( .A1(n11669), .A2(n16534), .ZN(n11670) );
  XNOR2_X1 U14668 ( .A(n17468), .B(n11649), .ZN(n11650) );
  AND2_X1 U14669 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11650), .ZN(
        n11664) );
  XNOR2_X1 U14670 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11650), .ZN(
        n17908) );
  XNOR2_X1 U14671 ( .A(n17475), .B(n11651), .ZN(n11660) );
  NOR2_X1 U14672 ( .A1(n18246), .A2(n11660), .ZN(n11661) );
  XOR2_X1 U14673 ( .A(n17479), .B(n11652), .Z(n11657) );
  NOR2_X1 U14674 ( .A1(n11657), .A2(n18278), .ZN(n11659) );
  INV_X1 U14675 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18938) );
  NOR2_X1 U14676 ( .A1(n11654), .A2(n18938), .ZN(n11656) );
  INV_X1 U14677 ( .A(n17959), .ZN(n11655) );
  NAND3_X1 U14678 ( .A1(n11655), .A2(n11654), .A3(n18938), .ZN(n11653) );
  OAI221_X1 U14679 ( .B1(n11656), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n11655), .C2(n11654), .A(n11653), .ZN(n17944) );
  XNOR2_X1 U14680 ( .A(n18278), .B(n11657), .ZN(n17943) );
  NOR2_X1 U14681 ( .A1(n17944), .A2(n17943), .ZN(n11658) );
  NOR2_X1 U14682 ( .A1(n11659), .A2(n11658), .ZN(n17933) );
  XNOR2_X1 U14683 ( .A(n18246), .B(n11660), .ZN(n17932) );
  NOR2_X1 U14684 ( .A1(n17933), .A2(n17932), .ZN(n17931) );
  XOR2_X1 U14685 ( .A(n17471), .B(n11662), .Z(n17916) );
  NOR2_X1 U14686 ( .A1(n17915), .A2(n17916), .ZN(n11663) );
  NAND2_X1 U14687 ( .A1(n17915), .A2(n17916), .ZN(n17914) );
  OAI21_X1 U14688 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n11663), .A(
        n17914), .ZN(n17907) );
  XNOR2_X1 U14689 ( .A(n17465), .B(n11665), .ZN(n11667) );
  NOR2_X1 U14690 ( .A1(n11666), .A2(n11667), .ZN(n11668) );
  INV_X1 U14691 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18238) );
  XNOR2_X1 U14692 ( .A(n11667), .B(n11666), .ZN(n17894) );
  NOR2_X1 U14693 ( .A1(n11668), .A2(n17893), .ZN(n11671) );
  XNOR2_X1 U14694 ( .A(n16534), .B(n11669), .ZN(n11672) );
  NAND2_X1 U14695 ( .A1(n11671), .A2(n11672), .ZN(n17879) );
  NAND2_X1 U14696 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17879), .ZN(
        n11674) );
  NOR2_X1 U14697 ( .A1(n11670), .A2(n11674), .ZN(n11676) );
  INV_X1 U14698 ( .A(n11670), .ZN(n11675) );
  OR2_X1 U14699 ( .A1(n11672), .A2(n11671), .ZN(n17880) );
  OAI21_X1 U14700 ( .B1(n11675), .B2(n11674), .A(n17880), .ZN(n11673) );
  AOI21_X1 U14701 ( .B1(n11675), .B2(n11674), .A(n11673), .ZN(n17871) );
  NOR2_X2 U14702 ( .A1(n15915), .A2(n16654), .ZN(n17950) );
  OAI22_X2 U14703 ( .A1(n17827), .A2(n17965), .B1(n17878), .B2(n18170), .ZN(
        n17856) );
  NOR3_X1 U14704 ( .A1(n17996), .A2(n17968), .A3(n17771), .ZN(n17631) );
  NAND2_X1 U14705 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17631), .ZN(
        n17621) );
  INV_X1 U14706 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U14707 ( .A1(n11684), .A2(n15983), .ZN(n15990) );
  NOR2_X1 U14708 ( .A1(n17621), .A2(n15990), .ZN(n11689) );
  NOR2_X1 U14709 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18974) );
  INV_X1 U14710 ( .A(n18974), .ZN(n18913) );
  NAND2_X1 U14711 ( .A1(n18973), .A2(n18910), .ZN(n16650) );
  AND2_X1 U14712 ( .A1(n18913), .A2(n16650), .ZN(n20992) );
  NAND2_X1 U14713 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17864) );
  INV_X1 U14714 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17653) );
  INV_X1 U14715 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17825) );
  NOR2_X2 U14716 ( .A1(n17822), .A2(n17825), .ZN(n17810) );
  INV_X1 U14717 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17787) );
  INV_X1 U14718 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17750) );
  INV_X1 U14719 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17018) );
  NOR2_X2 U14720 ( .A1(n17711), .A2(n17018), .ZN(n13414) );
  NAND2_X1 U14721 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n13414), .ZN(
        n13412) );
  INV_X1 U14722 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17696) );
  INV_X1 U14723 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17694) );
  NOR2_X1 U14724 ( .A1(n17696), .A2(n17694), .ZN(n17683) );
  INV_X1 U14725 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17628) );
  NOR2_X2 U14726 ( .A1(n17598), .A2(n17628), .ZN(n16670) );
  NAND2_X1 U14727 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17600) );
  INV_X1 U14728 ( .A(n17600), .ZN(n11677) );
  INV_X1 U14729 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20999) );
  XOR2_X1 U14730 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16519), .Z(
        n16684) );
  INV_X1 U14731 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17710) );
  NOR2_X1 U14732 ( .A1(n17711), .A2(n17710), .ZN(n17682) );
  NAND3_X1 U14733 ( .A1(n17682), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17664) );
  INV_X1 U14734 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17666) );
  NOR2_X1 U14735 ( .A1(n17664), .A2(n17666), .ZN(n17640) );
  NAND3_X1 U14736 ( .A1(n17640), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17627) );
  NOR2_X1 U14737 ( .A1(n17628), .A2(n17627), .ZN(n17599) );
  NAND3_X1 U14738 ( .A1(n17599), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16516) );
  NOR2_X1 U14739 ( .A1(n20999), .A2(n16516), .ZN(n11678) );
  NOR2_X1 U14740 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18973), .ZN(n17680) );
  NOR2_X1 U14741 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18910), .ZN(
        n18936) );
  AOI221_X1 U14742 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18973), .C1(n18921), 
        .C2(P3_STATE2_REG_2__SCAN_IN), .A(n18936), .ZN(n18306) );
  NOR2_X1 U14743 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18306), .ZN(n18661) );
  INV_X1 U14744 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18960) );
  NOR3_X1 U14745 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18960), .ZN(n18601) );
  NAND2_X1 U14746 ( .A1(n18661), .A2(n18601), .ZN(n18411) );
  NAND2_X1 U14747 ( .A1(n11678), .A2(n17809), .ZN(n13028) );
  NOR2_X1 U14748 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17678), .ZN(
        n16520) );
  INV_X1 U14749 ( .A(n16673), .ZN(n11680) );
  INV_X1 U14750 ( .A(n17680), .ZN(n17961) );
  OR2_X1 U14751 ( .A1(n18411), .A2(n11678), .ZN(n11679) );
  OAI211_X1 U14752 ( .C1(n11680), .C2(n17961), .A(n17960), .B(n11679), .ZN(
        n16526) );
  NOR2_X1 U14753 ( .A1(n16520), .A2(n16526), .ZN(n13026) );
  INV_X1 U14754 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20997) );
  NAND2_X1 U14755 ( .A1(n9768), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n15988) );
  OAI221_X1 U14756 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n13028), .C1(
        n9912), .C2(n13026), .A(n15988), .ZN(n11681) );
  AOI21_X1 U14757 ( .B1(n17812), .B2(n16684), .A(n11681), .ZN(n11687) );
  NAND2_X1 U14758 ( .A1(n16536), .A2(n18074), .ZN(n18027) );
  INV_X1 U14759 ( .A(n18027), .ZN(n18107) );
  NAND2_X1 U14760 ( .A1(n18107), .A2(n17650), .ZN(n17655) );
  INV_X1 U14761 ( .A(n17655), .ZN(n18005) );
  NAND2_X1 U14762 ( .A1(n18005), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17646) );
  NOR2_X1 U14763 ( .A1(n17996), .A2(n17646), .ZN(n17645) );
  NAND2_X1 U14764 ( .A1(n17645), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17974) );
  NOR2_X2 U14765 ( .A1(n17827), .A2(n16538), .ZN(n18026) );
  NAND2_X1 U14766 ( .A1(n17650), .A2(n18026), .ZN(n18007) );
  NAND2_X1 U14767 ( .A1(n11684), .A2(n17976), .ZN(n16528) );
  INV_X1 U14768 ( .A(n16528), .ZN(n13009) );
  OAI22_X1 U14769 ( .A1(n16517), .A2(n17878), .B1(n13009), .B2(n17965), .ZN(
        n11685) );
  NAND2_X1 U14770 ( .A1(n11685), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11686) );
  NAND2_X1 U14771 ( .A1(n11687), .A2(n11686), .ZN(n11688) );
  NAND2_X1 U14772 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n13684), .ZN(
        n11692) );
  INV_X1 U14773 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11697) );
  NOR2_X4 U14774 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14775 ( .A1(n11946), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11696) );
  AND2_X2 U14776 ( .A1(n11707), .A2(n13621), .ZN(n11847) );
  NAND2_X1 U14777 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11695) );
  OAI211_X1 U14778 ( .C1(n11945), .C2(n11697), .A(n11696), .B(n11695), .ZN(
        n11698) );
  INV_X1 U14779 ( .A(n11698), .ZN(n11703) );
  AOI22_X1 U14781 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14783 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10222), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11701) );
  AND2_X4 U14784 ( .A1(n11699), .A2(n13655), .ZN(n11896) );
  NAND2_X1 U14785 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11700) );
  NAND4_X1 U14786 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(
        n11715) );
  AOI22_X1 U14787 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12001), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14788 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11854), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11712) );
  AND2_X2 U14789 ( .A1(n11706), .A2(n13621), .ZN(n12427) );
  AOI22_X1 U14790 ( .A1(n12427), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14791 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11710) );
  NAND4_X1 U14792 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11714) );
  AOI22_X1 U14793 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12001), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14794 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11854), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14795 ( .A1(n12427), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14796 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11716) );
  INV_X1 U14797 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U14798 ( .A1(n11946), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14799 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11720) );
  OAI211_X1 U14800 ( .C1(n11945), .C2(n11722), .A(n11721), .B(n11720), .ZN(
        n11723) );
  INV_X1 U14801 ( .A(n11723), .ZN(n11727) );
  AOI22_X1 U14802 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14803 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10222), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U14804 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11724) );
  NAND2_X4 U14805 ( .A1(n10223), .A2(n9799), .ZN(n11827) );
  AOI22_X1 U14806 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11735) );
  INV_X1 U14807 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11730) );
  NAND2_X1 U14808 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U14809 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11728) );
  OAI211_X1 U14810 ( .C1(n11945), .C2(n11730), .A(n11729), .B(n11728), .ZN(
        n11731) );
  INV_X1 U14811 ( .A(n11731), .ZN(n11733) );
  NAND2_X1 U14812 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11732) );
  AOI22_X1 U14813 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11854), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14814 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10222), .B1(
        n12427), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14815 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11946), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14816 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14817 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11854), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14818 ( .A1(n12427), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14819 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U14820 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11753) );
  AOI22_X1 U14821 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10222), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14822 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11750) );
  INV_X1 U14823 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11746) );
  NAND2_X1 U14824 ( .A1(n11946), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14825 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11744) );
  OAI211_X1 U14826 ( .C1(n11945), .C2(n11746), .A(n11745), .B(n11744), .ZN(
        n11747) );
  INV_X1 U14827 ( .A(n11747), .ZN(n11749) );
  NAND2_X1 U14828 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11748) );
  NAND4_X1 U14829 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11752) );
  AOI22_X1 U14831 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12001), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14832 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11854), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14833 ( .A1(n12427), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11755) );
  INV_X1 U14834 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14835 ( .A1(n11946), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U14836 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11758) );
  OAI211_X1 U14837 ( .C1(n11945), .C2(n11760), .A(n11759), .B(n11758), .ZN(
        n11761) );
  INV_X1 U14838 ( .A(n11761), .ZN(n11765) );
  AOI22_X1 U14839 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14840 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10222), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11763) );
  NAND2_X1 U14841 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11762) );
  AOI22_X1 U14842 ( .A1(n12001), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12427), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14843 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14844 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11854), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14845 ( .A1(n11946), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11768) );
  INV_X1 U14846 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11774) );
  NAND2_X1 U14847 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U14848 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11772) );
  OAI211_X1 U14849 ( .C1(n11945), .C2(n11774), .A(n11773), .B(n11772), .ZN(
        n11775) );
  INV_X1 U14850 ( .A(n11775), .ZN(n11780) );
  AOI22_X1 U14851 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U14852 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11777) );
  AOI22_X1 U14853 ( .A1(n10222), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11955), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U14855 ( .A1(n12691), .A2(n11782), .ZN(n11784) );
  OAI21_X1 U14856 ( .B1(n11788), .B2(n12691), .A(n11784), .ZN(n11785) );
  INV_X1 U14857 ( .A(n11785), .ZN(n11786) );
  AOI22_X1 U14858 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12001), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14859 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11854), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14860 ( .A1(n12427), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14861 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11789) );
  NAND4_X1 U14862 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11802) );
  INV_X1 U14863 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11795) );
  NAND2_X1 U14864 ( .A1(n11946), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U14865 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11793) );
  OAI211_X1 U14866 ( .C1(n11945), .C2(n11795), .A(n11794), .B(n11793), .ZN(
        n11796) );
  INV_X1 U14867 ( .A(n11796), .ZN(n11800) );
  AOI22_X1 U14868 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14869 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10222), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U14870 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11797) );
  NAND4_X1 U14871 ( .A1(n11800), .A2(n11799), .A3(n11798), .A4(n11797), .ZN(
        n11801) );
  NAND2_X1 U14872 ( .A1(n12624), .A2(n14197), .ZN(n11803) );
  INV_X1 U14873 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11806) );
  NAND2_X1 U14874 ( .A1(n12001), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U14875 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11804) );
  OAI211_X1 U14876 ( .C1(n11945), .C2(n11806), .A(n11805), .B(n11804), .ZN(
        n11807) );
  INV_X1 U14877 ( .A(n11807), .ZN(n11811) );
  AOI22_X1 U14878 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11955), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14879 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11809) );
  NAND2_X1 U14880 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11808) );
  NAND4_X1 U14881 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11818) );
  AOI22_X1 U14882 ( .A1(n11946), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12427), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14883 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11853), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14884 ( .A1(n10222), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14885 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11862), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11813) );
  NAND4_X1 U14886 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11817) );
  NAND2_X1 U14887 ( .A1(n12831), .A2(n11824), .ZN(n13616) );
  AND2_X2 U14888 ( .A1(n13469), .A2(n11820), .ZN(n12824) );
  NAND2_X1 U14889 ( .A1(n13616), .A2(n14125), .ZN(n12842) );
  XNOR2_X1 U14890 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12821) );
  NAND3_X1 U14891 ( .A1(n13732), .A2(n11767), .A3(n13480), .ZN(n13612) );
  OAI21_X1 U14892 ( .B1(n12842), .B2(n11822), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11918) );
  NAND2_X1 U14893 ( .A1(n12624), .A2(n9817), .ZN(n13611) );
  NAND2_X1 U14894 ( .A1(n20261), .A2(n20278), .ZN(n12948) );
  OAI211_X1 U14895 ( .C1(n12847), .C2(n20982), .A(n13611), .B(n12948), .ZN(
        n11842) );
  NAND2_X1 U14896 ( .A1(n9771), .A2(n20261), .ZN(n12853) );
  NOR2_X1 U14897 ( .A1(n11842), .A2(n12950), .ZN(n11834) );
  NAND2_X1 U14898 ( .A1(n9801), .A2(n12847), .ZN(n11829) );
  NAND2_X1 U14899 ( .A1(n12835), .A2(n15030), .ZN(n11837) );
  INV_X1 U14900 ( .A(n13732), .ZN(n12951) );
  NAND2_X1 U14901 ( .A1(n12951), .A2(n11824), .ZN(n11832) );
  OAI21_X1 U14902 ( .B1(n11831), .B2(n11832), .A(n14197), .ZN(n11833) );
  NAND3_X1 U14903 ( .A1(n11834), .A2(n11837), .A3(n11833), .ZN(n12943) );
  NAND2_X1 U14904 ( .A1(n12943), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11835) );
  NOR2_X1 U14905 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13683) );
  NAND2_X1 U14906 ( .A1(n13683), .A2(n20885), .ZN(n12683) );
  MUX2_X1 U14907 ( .A(n12683), .B(n15963), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11836) );
  NAND2_X1 U14908 ( .A1(n11837), .A2(n20261), .ZN(n11838) );
  NAND2_X1 U14909 ( .A1(n11838), .A2(n20272), .ZN(n11846) );
  INV_X1 U14910 ( .A(n9801), .ZN(n14134) );
  INV_X1 U14911 ( .A(n13480), .ZN(n14650) );
  NAND3_X1 U14912 ( .A1(n14134), .A2(n20284), .A3(n14650), .ZN(n11844) );
  INV_X1 U14913 ( .A(n13683), .ZN(n16312) );
  NOR2_X1 U14914 ( .A1(n16312), .A2(n20885), .ZN(n11839) );
  NAND2_X1 U14915 ( .A1(n13732), .A2(n11819), .ZN(n12958) );
  OAI211_X1 U14916 ( .C1(n11840), .C2(n20982), .A(n11839), .B(n12958), .ZN(
        n11841) );
  AOI21_X1 U14917 ( .B1(n11831), .B2(n11844), .A(n11843), .ZN(n11845) );
  NAND2_X1 U14918 ( .A1(n11982), .A2(n20885), .ZN(n11886) );
  INV_X1 U14919 ( .A(n12759), .ZN(n11927) );
  BUF_X2 U14920 ( .A(n11945), .Z(n12600) );
  INV_X1 U14921 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U14922 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11849) );
  NAND2_X1 U14923 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11848) );
  OAI211_X1 U14924 ( .C1(n12600), .C2(n11850), .A(n11849), .B(n11848), .ZN(
        n11851) );
  INV_X1 U14925 ( .A(n11851), .ZN(n11859) );
  INV_X1 U14926 ( .A(n11852), .ZN(n11895) );
  AOI22_X1 U14927 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11858) );
  INV_X1 U14928 ( .A(n11853), .ZN(n12559) );
  INV_X2 U14929 ( .A(n12559), .ZN(n12578) );
  INV_X1 U14930 ( .A(n11854), .ZN(n11855) );
  INV_X2 U14931 ( .A(n11855), .ZN(n12565) );
  AOI22_X1 U14932 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U14933 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11856) );
  NAND4_X1 U14934 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11868) );
  INV_X1 U14935 ( .A(n10222), .ZN(n12589) );
  AOI22_X1 U14936 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11866) );
  INV_X1 U14937 ( .A(n12427), .ZN(n13627) );
  AOI22_X1 U14938 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11865) );
  INV_X1 U14939 ( .A(n11861), .ZN(n12002) );
  AOI22_X1 U14940 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14941 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11863) );
  NAND4_X1 U14942 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11867) );
  INV_X1 U14943 ( .A(n12690), .ZN(n11883) );
  INV_X1 U14944 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11871) );
  NAND2_X1 U14945 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U14946 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11869) );
  OAI211_X1 U14947 ( .C1(n12600), .C2(n11871), .A(n11870), .B(n11869), .ZN(
        n11872) );
  INV_X1 U14948 ( .A(n11872), .ZN(n11876) );
  AOI22_X1 U14949 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14950 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U14952 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11873) );
  NAND4_X1 U14953 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11882) );
  AOI22_X1 U14954 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14955 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14956 ( .A1(n12427), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14957 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U14958 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11881) );
  XNOR2_X1 U14959 ( .A(n11883), .B(n12763), .ZN(n11884) );
  NAND2_X1 U14960 ( .A1(n11927), .A2(n11884), .ZN(n11885) );
  INV_X1 U14961 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20271) );
  AOI21_X1 U14962 ( .B1(n14197), .B2(n12690), .A(n20885), .ZN(n11888) );
  NAND2_X1 U14963 ( .A1(n12847), .A2(n12763), .ZN(n11887) );
  OAI211_X1 U14964 ( .C1(n12661), .C2(n20271), .A(n11888), .B(n11887), .ZN(
        n11978) );
  NAND2_X1 U14965 ( .A1(n11980), .A2(n11978), .ZN(n11890) );
  NAND2_X1 U14966 ( .A1(n11927), .A2(n12763), .ZN(n11889) );
  INV_X1 U14967 ( .A(n11992), .ZN(n11908) );
  INV_X1 U14968 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U14969 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U14970 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11891) );
  OAI211_X1 U14971 ( .C1(n12600), .C2(n11893), .A(n11892), .B(n11891), .ZN(
        n11894) );
  INV_X1 U14972 ( .A(n11894), .ZN(n11900) );
  INV_X2 U14973 ( .A(n11895), .ZN(n12553) );
  AOI22_X1 U14974 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12582), .ZN(n11899) );
  AOI22_X1 U14975 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U14976 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11897) );
  NAND4_X1 U14977 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n11907) );
  INV_X1 U14978 ( .A(n9751), .ZN(n12555) );
  INV_X2 U14979 ( .A(n12555), .ZN(n12583) );
  AOI22_X1 U14980 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11905) );
  INV_X2 U14981 ( .A(n13627), .ZN(n12579) );
  AOI22_X1 U14982 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14983 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14985 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12577), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11902) );
  NAND4_X1 U14986 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11906) );
  NAND2_X1 U14987 ( .A1(n11908), .A2(n12689), .ZN(n11910) );
  NAND2_X1 U14988 ( .A1(n12669), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11909) );
  OAI211_X1 U14989 ( .C1(n12759), .C2(n12763), .A(n11910), .B(n11909), .ZN(
        n11911) );
  NAND2_X1 U14990 ( .A1(n11912), .A2(n11911), .ZN(n11913) );
  NAND2_X1 U14991 ( .A1(n11933), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U14992 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11936) );
  OAI21_X1 U14993 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11936), .ZN(n20608) );
  INV_X1 U14994 ( .A(n15963), .ZN(n11914) );
  NAND2_X1 U14995 ( .A1(n11914), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11930) );
  OAI21_X1 U14996 ( .B1(n12683), .B2(n20608), .A(n11930), .ZN(n11915) );
  INV_X1 U14997 ( .A(n11915), .ZN(n11916) );
  XNOR2_X2 U14998 ( .A(n11920), .B(n11919), .ZN(n20390) );
  INV_X1 U14999 ( .A(n11921), .ZN(n11922) );
  NAND2_X2 U15000 ( .A1(n20390), .A2(n11924), .ZN(n11943) );
  INV_X1 U15001 ( .A(n20390), .ZN(n11926) );
  NAND2_X1 U15002 ( .A1(n11926), .A2(n11925), .ZN(n20321) );
  NAND2_X1 U15004 ( .A1(n11927), .A2(n12689), .ZN(n11928) );
  NAND2_X1 U15005 ( .A1(n11930), .A2(n10119), .ZN(n11931) );
  NOR2_X1 U15006 ( .A1(n15963), .A2(n20611), .ZN(n11934) );
  INV_X1 U15007 ( .A(n12683), .ZN(n11989) );
  INV_X1 U15008 ( .A(n11936), .ZN(n11935) );
  NAND2_X1 U15009 ( .A1(n11935), .A2(n20611), .ZN(n20653) );
  NAND2_X1 U15010 ( .A1(n11936), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U15011 ( .A1(n20653), .A2(n11937), .ZN(n20265) );
  NAND2_X1 U15012 ( .A1(n11989), .A2(n20265), .ZN(n11940) );
  NAND2_X2 U15013 ( .A1(n11939), .A2(n11938), .ZN(n13819) );
  NAND4_X1 U15014 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11944) );
  INV_X1 U15015 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11949) );
  NAND2_X1 U15016 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U15017 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11947) );
  OAI211_X1 U15018 ( .C1(n12600), .C2(n11949), .A(n11948), .B(n11947), .ZN(
        n11950) );
  INV_X1 U15019 ( .A(n11950), .ZN(n11954) );
  INV_X1 U15020 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n21011) );
  AOI22_X1 U15021 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11953) );
  INV_X2 U15022 ( .A(n12589), .ZN(n12538) );
  AOI22_X1 U15023 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U15024 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11951) );
  NAND4_X1 U15025 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11961) );
  AOI22_X1 U15026 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15027 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15028 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15029 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U15030 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  INV_X1 U15031 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20283) );
  OAI22_X1 U15032 ( .A1(n12706), .A2(n11992), .B1(n12661), .B2(n20283), .ZN(
        n11962) );
  INV_X1 U15033 ( .A(n11962), .ZN(n11963) );
  NAND2_X1 U15034 ( .A1(n11819), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12120) );
  NAND2_X1 U15036 ( .A1(n9777), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12042) );
  NOR2_X1 U15037 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11985) );
  XNOR2_X1 U15038 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14676) );
  INV_X2 U15039 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20888) );
  AND2_X1 U15040 ( .A1(n20888), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12614) );
  AOI21_X1 U15041 ( .B1(n11985), .B2(n14676), .A(n12614), .ZN(n11968) );
  INV_X2 U15042 ( .A(n10208), .ZN(n12615) );
  NAND2_X1 U15043 ( .A1(n12615), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11967) );
  OAI211_X1 U15044 ( .C1(n12042), .C2(n13655), .A(n11968), .B(n11967), .ZN(
        n11969) );
  INV_X1 U15045 ( .A(n11969), .ZN(n11970) );
  NAND2_X1 U15046 ( .A1(n12614), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11987) );
  XNOR2_X2 U15047 ( .A(n9807), .B(n12695), .ZN(n13831) );
  NAND2_X1 U15048 ( .A1(n13831), .A2(n12247), .ZN(n11977) );
  NAND2_X1 U15049 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20888), .ZN(
        n11974) );
  NAND2_X1 U15050 ( .A1(n12615), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n11973) );
  OAI211_X1 U15051 ( .C1(n12042), .C2(n9784), .A(n11974), .B(n11973), .ZN(
        n11975) );
  INV_X1 U15052 ( .A(n11975), .ZN(n11976) );
  NAND2_X1 U15053 ( .A1(n11977), .A2(n11976), .ZN(n13784) );
  INV_X1 U15054 ( .A(n11978), .ZN(n11979) );
  INV_X1 U15055 ( .A(n12686), .ZN(n20349) );
  NAND2_X1 U15056 ( .A1(n20349), .A2(n11819), .ZN(n11981) );
  NAND2_X1 U15057 ( .A1(n11981), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13739) );
  AOI22_X1 U15058 ( .A1(n12615), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20888), .ZN(n11983) );
  OAI21_X1 U15059 ( .B1(n13684), .B2(n12042), .A(n11983), .ZN(n11984) );
  AOI21_X1 U15060 ( .B1(n9785), .B2(n12247), .A(n11984), .ZN(n13740) );
  INV_X1 U15061 ( .A(n11985), .ZN(n12609) );
  NAND2_X1 U15062 ( .A1(n13740), .A2(n11985), .ZN(n11986) );
  NAND2_X1 U15063 ( .A1(n13737), .A2(n11986), .ZN(n13783) );
  NAND2_X1 U15064 ( .A1(n11933), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11991) );
  NOR3_X1 U15065 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20611), .A3(
        n20693), .ZN(n20526) );
  NAND2_X1 U15066 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20526), .ZN(
        n20519) );
  NAND3_X1 U15067 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20821) );
  NOR2_X1 U15068 ( .A1(n20755), .A2(n20821), .ZN(n20873) );
  AOI21_X1 U15069 ( .B1(n20519), .B2(n20652), .A(n20873), .ZN(n20551) );
  NOR2_X1 U15070 ( .A1(n15963), .A2(n20652), .ZN(n11988) );
  AOI21_X1 U15071 ( .B1(n20551), .B2(n11989), .A(n11988), .ZN(n11990) );
  XNOR2_X2 U15072 ( .A(n13819), .B(n20427), .ZN(n20549) );
  INV_X1 U15073 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11995) );
  NAND2_X1 U15074 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11994) );
  NAND2_X1 U15075 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11993) );
  OAI211_X1 U15076 ( .C1(n12600), .C2(n11995), .A(n11994), .B(n11993), .ZN(
        n11996) );
  INV_X1 U15077 ( .A(n11996), .ZN(n12000) );
  AOI22_X1 U15078 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15079 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U15080 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11997) );
  NAND4_X1 U15081 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12008) );
  AOI22_X1 U15082 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15083 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12005) );
  INV_X2 U15084 ( .A(n12002), .ZN(n12590) );
  AOI22_X1 U15085 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15086 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12003) );
  NAND4_X1 U15087 ( .A1(n12006), .A2(n12005), .A3(n12004), .A4(n12003), .ZN(
        n12007) );
  AOI22_X1 U15088 ( .A1(n12640), .A2(n12716), .B1(n12669), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12009) );
  INV_X1 U15089 ( .A(n13829), .ZN(n13830) );
  NAND2_X1 U15090 ( .A1(n9752), .A2(n12247), .ZN(n12020) );
  INV_X1 U15091 ( .A(n12609), .ZN(n14192) );
  INV_X1 U15092 ( .A(n12013), .ZN(n12015) );
  INV_X1 U15093 ( .A(n12039), .ZN(n12014) );
  OAI21_X1 U15094 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12015), .A(
        n12014), .ZN(n14665) );
  AOI22_X1 U15095 ( .A1(n14192), .A2(n14665), .B1(n12614), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U15096 ( .A1(n12615), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12016) );
  OAI211_X1 U15097 ( .C1(n12042), .C2(n12011), .A(n12017), .B(n12016), .ZN(
        n12018) );
  INV_X1 U15098 ( .A(n12018), .ZN(n12019) );
  NAND2_X1 U15099 ( .A1(n12020), .A2(n12019), .ZN(n13921) );
  NAND2_X1 U15100 ( .A1(n13922), .A2(n13921), .ZN(n13920) );
  INV_X1 U15101 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12507) );
  NAND2_X1 U15102 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12022) );
  NAND2_X1 U15103 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12021) );
  OAI211_X1 U15104 ( .C1(n12600), .C2(n12507), .A(n12022), .B(n12021), .ZN(
        n12023) );
  INV_X1 U15105 ( .A(n12023), .ZN(n12027) );
  AOI22_X1 U15106 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15107 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12025) );
  NAND2_X1 U15108 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12024) );
  NAND4_X1 U15109 ( .A1(n12027), .A2(n12026), .A3(n12025), .A4(n12024), .ZN(
        n12033) );
  AOI22_X1 U15110 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15111 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15112 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15113 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12028) );
  NAND4_X1 U15114 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12032) );
  NAND2_X1 U15115 ( .A1(n12640), .A2(n12723), .ZN(n12035) );
  NAND2_X1 U15116 ( .A1(n12669), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12034) );
  NAND2_X1 U15117 ( .A1(n12035), .A2(n12034), .ZN(n12036) );
  OR2_X1 U15118 ( .A1(n12037), .A2(n12036), .ZN(n12038) );
  NAND2_X1 U15119 ( .A1(n12064), .A2(n12038), .ZN(n12714) );
  OAI21_X1 U15120 ( .B1(n12039), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12066), .ZN(n20178) );
  INV_X1 U15121 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16315) );
  INV_X1 U15122 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20092) );
  AOI21_X1 U15123 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20092), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12040) );
  AOI21_X1 U15124 ( .B1(n12615), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12040), .ZN(
        n12041) );
  OAI21_X1 U15125 ( .B1(n12042), .B2(n16315), .A(n12041), .ZN(n12043) );
  OAI21_X1 U15126 ( .B1(n20178), .B2(n12609), .A(n12043), .ZN(n12044) );
  NOR2_X2 U15127 ( .A1(n13920), .A2(n14139), .ZN(n13988) );
  INV_X1 U15128 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U15129 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U15130 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12047) );
  OAI211_X1 U15131 ( .C1(n12600), .C2(n12049), .A(n12048), .B(n12047), .ZN(
        n12050) );
  INV_X1 U15132 ( .A(n12050), .ZN(n12054) );
  AOI22_X1 U15133 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15134 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12052) );
  NAND2_X1 U15135 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12051) );
  NAND4_X1 U15136 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n12060) );
  AOI22_X1 U15137 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15138 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15139 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15140 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12055) );
  NAND4_X1 U15141 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12059) );
  AOI22_X1 U15142 ( .A1(n12640), .A2(n12733), .B1(n12669), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12063) );
  NAND2_X1 U15143 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  NAND2_X1 U15144 ( .A1(n12092), .A2(n12065), .ZN(n12722) );
  INV_X1 U15145 ( .A(n12614), .ZN(n12161) );
  NAND2_X1 U15146 ( .A1(n12066), .A2(n20073), .ZN(n12067) );
  INV_X1 U15147 ( .A(n12085), .ZN(n12086) );
  NAND2_X1 U15148 ( .A1(n12067), .A2(n12086), .ZN(n20084) );
  NAND2_X1 U15149 ( .A1(n20084), .A2(n11985), .ZN(n12068) );
  OAI21_X1 U15150 ( .B1(n20073), .B2(n12161), .A(n12068), .ZN(n12069) );
  AOI21_X1 U15151 ( .B1(n12615), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12069), .ZN(
        n12070) );
  INV_X1 U15152 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12554) );
  NAND2_X1 U15153 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12073) );
  NAND2_X1 U15154 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12072) );
  OAI211_X1 U15155 ( .C1(n12600), .C2(n12554), .A(n12073), .B(n12072), .ZN(
        n12074) );
  INV_X1 U15156 ( .A(n12074), .ZN(n12078) );
  AOI22_X1 U15157 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15158 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12076) );
  NAND2_X1 U15159 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12075) );
  NAND4_X1 U15160 ( .A1(n12078), .A2(n12077), .A3(n12076), .A4(n12075), .ZN(
        n12084) );
  AOI22_X1 U15161 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15162 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11955), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15163 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15164 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12079) );
  NAND4_X1 U15165 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        n12083) );
  OR2_X1 U15166 ( .A1(n12084), .A2(n12083), .ZN(n12744) );
  AOI22_X1 U15167 ( .A1(n12640), .A2(n12744), .B1(n12669), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12093) );
  INV_X1 U15168 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14235) );
  INV_X1 U15169 ( .A(n12097), .ZN(n12098) );
  INV_X1 U15170 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20063) );
  NAND2_X1 U15171 ( .A1(n20063), .A2(n12086), .ZN(n12087) );
  NAND2_X1 U15172 ( .A1(n12098), .A2(n12087), .ZN(n20070) );
  AOI22_X1 U15173 ( .A1(n20070), .A2(n11985), .B1(n12614), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12088) );
  OAI21_X1 U15174 ( .B1(n10208), .B2(n14235), .A(n12088), .ZN(n12089) );
  INV_X1 U15175 ( .A(n14234), .ZN(n12090) );
  NAND2_X1 U15176 ( .A1(n12091), .A2(n12090), .ZN(n14162) );
  NAND2_X1 U15177 ( .A1(n12640), .A2(n12763), .ZN(n12095) );
  NAND2_X1 U15178 ( .A1(n12669), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12094) );
  NAND2_X1 U15179 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  INV_X1 U15180 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12102) );
  INV_X1 U15181 ( .A(n12121), .ZN(n12100) );
  INV_X1 U15182 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16149) );
  NAND2_X1 U15183 ( .A1(n12098), .A2(n16149), .ZN(n12099) );
  NAND2_X1 U15184 ( .A1(n12100), .A2(n12099), .ZN(n20059) );
  AOI22_X1 U15185 ( .A1(n20059), .A2(n11985), .B1(n12614), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12101) );
  OAI21_X1 U15186 ( .B1(n10208), .B2(n12102), .A(n12101), .ZN(n12103) );
  AOI21_X1 U15187 ( .B1(n12743), .B2(n12247), .A(n12103), .ZN(n14161) );
  NAND2_X1 U15188 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12105) );
  NAND2_X1 U15189 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12104) );
  OAI211_X1 U15190 ( .C1(n12600), .C2(n20271), .A(n12105), .B(n12104), .ZN(
        n12106) );
  INV_X1 U15191 ( .A(n12106), .ZN(n12110) );
  AOI22_X1 U15192 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11955), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15193 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U15194 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12107) );
  NAND4_X1 U15195 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12116) );
  AOI22_X1 U15196 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15197 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15198 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15199 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12111) );
  NAND4_X1 U15200 ( .A1(n12114), .A2(n12113), .A3(n12112), .A4(n12111), .ZN(
        n12115) );
  NOR2_X1 U15201 ( .A1(n12116), .A2(n12115), .ZN(n12119) );
  XNOR2_X1 U15202 ( .A(n12121), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14272) );
  AOI22_X1 U15203 ( .A1(n14272), .A2(n11985), .B1(n12614), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U15204 ( .A1(n12615), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12117) );
  OAI211_X1 U15205 ( .C1(n12120), .C2(n12119), .A(n12118), .B(n12117), .ZN(
        n14171) );
  XNOR2_X1 U15206 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12140), .ZN(
        n20038) );
  INV_X1 U15207 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U15208 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12123) );
  NAND2_X1 U15209 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12122) );
  OAI211_X1 U15210 ( .C1(n12600), .C2(n12124), .A(n12123), .B(n12122), .ZN(
        n12125) );
  INV_X1 U15211 ( .A(n12125), .ZN(n12129) );
  AOI22_X1 U15212 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12582), .ZN(n12128) );
  AOI22_X1 U15213 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11955), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U15214 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12126) );
  NAND4_X1 U15215 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12135) );
  AOI22_X1 U15216 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12578), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15217 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11901), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15218 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15219 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12130) );
  NAND4_X1 U15220 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12134) );
  OR2_X1 U15221 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  AOI22_X1 U15222 ( .A1(n12247), .A2(n12136), .B1(n12614), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U15223 ( .A1(n12615), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12137) );
  OAI211_X1 U15224 ( .C1(n20038), .C2(n12609), .A(n12138), .B(n12137), .ZN(
        n14238) );
  INV_X1 U15225 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12139) );
  XNOR2_X1 U15226 ( .A(n12158), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14970) );
  AOI22_X1 U15227 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15228 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15229 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15230 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12141) );
  NAND4_X1 U15231 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .ZN(
        n12153) );
  NAND2_X1 U15232 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U15233 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12145) );
  OAI211_X1 U15234 ( .C1(n12600), .C2(n20283), .A(n12146), .B(n12145), .ZN(
        n12147) );
  INV_X1 U15235 ( .A(n12147), .ZN(n12151) );
  AOI22_X1 U15236 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15237 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12149) );
  NAND2_X1 U15238 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12148) );
  NAND4_X1 U15239 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n12152) );
  OAI21_X1 U15240 ( .B1(n12153), .B2(n12152), .A(n12247), .ZN(n12156) );
  NAND2_X1 U15241 ( .A1(n12615), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12155) );
  NAND2_X1 U15242 ( .A1(n12614), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12154) );
  NAND3_X1 U15243 ( .A1(n12156), .A2(n12155), .A3(n12154), .ZN(n12157) );
  AOI21_X1 U15244 ( .B1(n14970), .B2(n14192), .A(n12157), .ZN(n14635) );
  INV_X1 U15245 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12162) );
  OAI21_X1 U15246 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12159), .A(
        n12210), .ZN(n16142) );
  NAND2_X1 U15247 ( .A1(n16142), .A2(n11985), .ZN(n12160) );
  OAI21_X1 U15248 ( .B1(n12162), .B2(n12161), .A(n12160), .ZN(n12163) );
  AOI21_X1 U15249 ( .B1(n12615), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12163), .ZN(
        n14621) );
  INV_X1 U15250 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12167) );
  NAND2_X1 U15251 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15252 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12165) );
  OAI211_X1 U15253 ( .C1(n12600), .C2(n12167), .A(n12166), .B(n12165), .ZN(
        n12168) );
  INV_X1 U15254 ( .A(n12168), .ZN(n12172) );
  AOI22_X1 U15255 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15256 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12170) );
  NAND2_X1 U15257 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12169) );
  NAND4_X1 U15258 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12178) );
  AOI22_X1 U15259 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15260 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15261 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15262 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12173) );
  NAND4_X1 U15263 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12177) );
  OR2_X1 U15264 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  NAND2_X1 U15265 ( .A1(n12247), .A2(n12179), .ZN(n14858) );
  INV_X1 U15266 ( .A(n14858), .ZN(n12180) );
  INV_X1 U15267 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16061) );
  XOR2_X1 U15268 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12214), .Z(
        n14963) );
  INV_X1 U15269 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20304) );
  NAND2_X1 U15270 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12182) );
  NAND2_X1 U15271 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12181) );
  OAI211_X1 U15272 ( .C1(n12600), .C2(n20304), .A(n12182), .B(n12181), .ZN(
        n12183) );
  INV_X1 U15273 ( .A(n12183), .ZN(n12187) );
  AOI22_X1 U15274 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15275 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12185) );
  NAND2_X1 U15276 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12184) );
  NAND4_X1 U15277 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12193) );
  AOI22_X1 U15278 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15279 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15280 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15281 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15282 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12192) );
  OR2_X1 U15283 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  AOI22_X1 U15284 ( .A1(n12247), .A2(n12194), .B1(n12614), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U15285 ( .A1(n12615), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12195) );
  OAI211_X1 U15286 ( .C1(n14963), .C2(n12609), .A(n12196), .B(n12195), .ZN(
        n14624) );
  INV_X1 U15287 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U15288 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15289 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15290 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15291 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15292 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12209) );
  INV_X1 U15293 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20295) );
  NAND2_X1 U15294 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12202) );
  NAND2_X1 U15295 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12201) );
  OAI211_X1 U15296 ( .C1(n12600), .C2(n20295), .A(n12202), .B(n12201), .ZN(
        n12203) );
  INV_X1 U15297 ( .A(n12203), .ZN(n12207) );
  AOI22_X1 U15298 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15299 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12205) );
  NAND2_X1 U15300 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12204) );
  NAND4_X1 U15301 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12208) );
  OAI21_X1 U15302 ( .B1(n12209), .B2(n12208), .A(n12247), .ZN(n12213) );
  XNOR2_X1 U15303 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12210), .ZN(
        n16129) );
  INV_X1 U15304 ( .A(n16129), .ZN(n12211) );
  AOI22_X1 U15305 ( .A1(n12614), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n14192), .B2(n12211), .ZN(n12212) );
  OAI211_X1 U15306 ( .C1(n10208), .C2(n14855), .A(n12213), .B(n12212), .ZN(
        n14851) );
  INV_X1 U15307 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21015) );
  NAND2_X1 U15308 ( .A1(n12215), .A2(n21015), .ZN(n12217) );
  INV_X1 U15309 ( .A(n12273), .ZN(n12216) );
  NAND2_X1 U15310 ( .A1(n12217), .A2(n12216), .ZN(n14949) );
  NAND2_X1 U15311 ( .A1(n14949), .A2(n11985), .ZN(n12235) );
  AOI22_X1 U15312 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15313 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15314 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15315 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12218) );
  NAND4_X1 U15316 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12218), .ZN(
        n12230) );
  INV_X1 U15317 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20309) );
  NAND2_X1 U15318 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12223) );
  NAND2_X1 U15319 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12222) );
  OAI211_X1 U15320 ( .C1(n12600), .C2(n20309), .A(n12223), .B(n12222), .ZN(
        n12224) );
  INV_X1 U15321 ( .A(n12224), .ZN(n12228) );
  AOI22_X1 U15322 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15323 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U15324 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12225) );
  NAND4_X1 U15325 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12229) );
  OAI21_X1 U15326 ( .B1(n12230), .B2(n12229), .A(n12247), .ZN(n12233) );
  NAND2_X1 U15327 ( .A1(n12615), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12232) );
  NAND2_X1 U15328 ( .A1(n12614), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12231) );
  AND3_X1 U15329 ( .A1(n12233), .A2(n12232), .A3(n12231), .ZN(n12234) );
  NAND2_X1 U15330 ( .A1(n12235), .A2(n12234), .ZN(n14606) );
  NAND2_X1 U15331 ( .A1(n14607), .A2(n14606), .ZN(n14608) );
  INV_X1 U15332 ( .A(n14608), .ZN(n12255) );
  AOI22_X1 U15333 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15334 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15335 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15336 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12236) );
  NAND4_X1 U15337 ( .A1(n12239), .A2(n12238), .A3(n12237), .A4(n12236), .ZN(
        n12249) );
  INV_X1 U15338 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U15339 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12241) );
  NAND2_X1 U15340 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12240) );
  OAI211_X1 U15341 ( .C1(n11945), .C2(n12591), .A(n12241), .B(n12240), .ZN(
        n12242) );
  INV_X1 U15342 ( .A(n12242), .ZN(n12246) );
  AOI22_X1 U15343 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15344 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U15345 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12243) );
  NAND4_X1 U15346 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12248) );
  OAI21_X1 U15347 ( .B1(n12249), .B2(n12248), .A(n12247), .ZN(n12253) );
  XOR2_X1 U15348 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12273), .Z(
        n16124) );
  INV_X1 U15349 ( .A(n16124), .ZN(n12250) );
  AOI22_X1 U15350 ( .A1(n12614), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n14192), .B2(n12250), .ZN(n12252) );
  NAND2_X1 U15351 ( .A1(n12615), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12251) );
  AND3_X1 U15352 ( .A1(n12253), .A2(n12252), .A3(n12251), .ZN(n14755) );
  NAND2_X1 U15353 ( .A1(n12255), .A2(n12254), .ZN(n14591) );
  INV_X1 U15354 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U15355 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12257) );
  NAND2_X1 U15356 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12256) );
  OAI211_X1 U15357 ( .C1(n11945), .C2(n12258), .A(n12257), .B(n12256), .ZN(
        n12259) );
  INV_X1 U15358 ( .A(n12259), .ZN(n12263) );
  AOI22_X1 U15359 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15360 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U15361 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12260) );
  NAND4_X1 U15362 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12269) );
  AOI22_X1 U15363 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15364 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15365 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15366 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U15367 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12268) );
  NOR2_X1 U15368 ( .A1(n12269), .A2(n12268), .ZN(n12272) );
  INV_X1 U15369 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12276) );
  AOI21_X1 U15370 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n12276), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12270) );
  AOI21_X1 U15371 ( .B1(n12615), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12270), .ZN(
        n12271) );
  OAI21_X1 U15372 ( .B1(n12574), .B2(n12272), .A(n12271), .ZN(n12275) );
  XNOR2_X1 U15373 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B(n12277), .ZN(
        n14934) );
  NAND2_X1 U15374 ( .A1(n14192), .A2(n14934), .ZN(n12274) );
  NAND2_X1 U15375 ( .A1(n12275), .A2(n12274), .ZN(n14594) );
  XNOR2_X1 U15376 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12294), .ZN(
        n16114) );
  AOI22_X1 U15377 ( .A1(n12615), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12614), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15378 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15379 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12577), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15380 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11901), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15381 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U15382 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12291) );
  INV_X1 U15383 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12284) );
  NAND2_X1 U15384 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12283) );
  NAND2_X1 U15385 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12282) );
  OAI211_X1 U15386 ( .C1(n11945), .C2(n12284), .A(n12283), .B(n12282), .ZN(
        n12285) );
  INV_X1 U15387 ( .A(n12285), .ZN(n12289) );
  AOI22_X1 U15388 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15389 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12287) );
  NAND2_X1 U15390 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12286) );
  NAND4_X1 U15391 ( .A1(n12289), .A2(n12288), .A3(n12287), .A4(n12286), .ZN(
        n12290) );
  INV_X1 U15392 ( .A(n12574), .ZN(n12605) );
  OAI21_X1 U15393 ( .B1(n12291), .B2(n12290), .A(n12605), .ZN(n12292) );
  OAI211_X1 U15394 ( .C1(n16114), .C2(n12609), .A(n12293), .B(n12292), .ZN(
        n14742) );
  INV_X1 U15395 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16044) );
  INV_X1 U15396 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12295) );
  XNOR2_X1 U15397 ( .A(n12330), .B(n12295), .ZN(n14922) );
  AOI22_X1 U15398 ( .A1(n12615), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20888), .ZN(n12311) );
  AOI22_X1 U15399 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15400 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15401 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15402 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15403 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12309) );
  AOI22_X1 U15404 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12307) );
  INV_X1 U15405 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U15406 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12301) );
  NAND2_X1 U15407 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12300) );
  OAI211_X1 U15408 ( .C1(n12600), .C2(n12302), .A(n12301), .B(n12300), .ZN(
        n12303) );
  INV_X1 U15409 ( .A(n12303), .ZN(n12306) );
  AOI21_X1 U15410 ( .B1(n12538), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n14192), .ZN(n12305) );
  AOI22_X1 U15411 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12304) );
  NAND4_X1 U15412 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12304), .ZN(
        n12308) );
  NAND2_X1 U15413 ( .A1(n12574), .A2(n12609), .ZN(n12384) );
  OAI21_X1 U15414 ( .B1(n12309), .B2(n12308), .A(n12384), .ZN(n12310) );
  AOI22_X1 U15415 ( .A1(n14922), .A2(n11985), .B1(n12311), .B2(n12310), .ZN(
        n14579) );
  INV_X1 U15416 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12314) );
  NAND2_X1 U15417 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12313) );
  NAND2_X1 U15418 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12312) );
  OAI211_X1 U15419 ( .C1(n11945), .C2(n12314), .A(n12313), .B(n12312), .ZN(
        n12315) );
  INV_X1 U15420 ( .A(n12315), .ZN(n12319) );
  AOI22_X1 U15421 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15422 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U15423 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12316) );
  NAND4_X1 U15424 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12325) );
  AOI22_X1 U15425 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15426 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15427 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15428 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12320) );
  NAND4_X1 U15429 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12324) );
  NOR2_X1 U15430 ( .A1(n12325), .A2(n12324), .ZN(n12329) );
  NAND2_X1 U15431 ( .A1(n20888), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12326) );
  NAND2_X1 U15432 ( .A1(n12609), .A2(n12326), .ZN(n12327) );
  AOI21_X1 U15433 ( .B1(n12615), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12327), .ZN(
        n12328) );
  OAI21_X1 U15434 ( .B1(n12574), .B2(n12329), .A(n12328), .ZN(n12333) );
  OAI21_X1 U15435 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12331), .A(
        n12369), .ZN(n16108) );
  OR2_X1 U15436 ( .A1(n12609), .A2(n16108), .ZN(n12332) );
  NAND2_X1 U15437 ( .A1(n12333), .A2(n12332), .ZN(n14563) );
  AOI22_X1 U15438 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15439 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15440 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15441 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12334) );
  NAND4_X1 U15442 ( .A1(n12337), .A2(n12336), .A3(n12335), .A4(n12334), .ZN(
        n12346) );
  AOI22_X1 U15443 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12344) );
  INV_X1 U15444 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12508) );
  NAND2_X1 U15445 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12339) );
  NAND2_X1 U15446 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12338) );
  OAI211_X1 U15447 ( .C1(n12600), .C2(n12508), .A(n12339), .B(n12338), .ZN(
        n12340) );
  INV_X1 U15448 ( .A(n12340), .ZN(n12343) );
  AOI21_X1 U15449 ( .B1(n12596), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n14192), .ZN(n12342) );
  AOI22_X1 U15450 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12341) );
  NAND4_X1 U15451 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .ZN(
        n12345) );
  OAI21_X1 U15452 ( .B1(n12346), .B2(n12345), .A(n12384), .ZN(n12348) );
  AOI22_X1 U15453 ( .A1(n12615), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20888), .ZN(n12347) );
  NAND2_X1 U15454 ( .A1(n12348), .A2(n12347), .ZN(n12350) );
  XNOR2_X1 U15455 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12369), .ZN(
        n14916) );
  NAND2_X1 U15456 ( .A1(n14192), .A2(n14916), .ZN(n12349) );
  NAND2_X1 U15457 ( .A1(n12350), .A2(n12349), .ZN(n14552) );
  INV_X1 U15458 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12353) );
  NAND2_X1 U15459 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12352) );
  NAND2_X1 U15460 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12351) );
  OAI211_X1 U15461 ( .C1(n11945), .C2(n12353), .A(n12352), .B(n12351), .ZN(
        n12354) );
  INV_X1 U15462 ( .A(n12354), .ZN(n12358) );
  AOI22_X1 U15463 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15464 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12356) );
  NAND2_X1 U15465 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12355) );
  NAND4_X1 U15466 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12364) );
  AOI22_X1 U15467 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15468 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12427), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15469 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15470 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12359) );
  NAND4_X1 U15471 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12363) );
  NOR2_X1 U15472 ( .A1(n12364), .A2(n12363), .ZN(n12368) );
  INV_X1 U15473 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20789) );
  OAI21_X1 U15474 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20789), .A(
        n20888), .ZN(n12365) );
  INV_X1 U15475 ( .A(n12365), .ZN(n12366) );
  AOI21_X1 U15476 ( .B1(n12615), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12366), .ZN(
        n12367) );
  OAI21_X1 U15477 ( .B1(n12574), .B2(n12368), .A(n12367), .ZN(n12372) );
  INV_X1 U15478 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14914) );
  OAI21_X1 U15479 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12370), .A(
        n12440), .ZN(n16101) );
  OR2_X1 U15480 ( .A1(n12609), .A2(n16101), .ZN(n12371) );
  INV_X1 U15481 ( .A(n14532), .ZN(n12392) );
  AOI22_X1 U15482 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15483 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15484 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15485 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U15486 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12386) );
  AOI22_X1 U15487 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11896), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12383) );
  INV_X1 U15488 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12557) );
  NAND2_X1 U15489 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12378) );
  NAND2_X1 U15490 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12377) );
  OAI211_X1 U15491 ( .C1(n11945), .C2(n12557), .A(n12378), .B(n12377), .ZN(
        n12379) );
  INV_X1 U15492 ( .A(n12379), .ZN(n12382) );
  AOI21_X1 U15493 ( .B1(n12565), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n14192), .ZN(n12381) );
  AOI22_X1 U15494 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15495 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12385) );
  OAI21_X1 U15496 ( .B1(n12386), .B2(n12385), .A(n12384), .ZN(n12388) );
  AOI22_X1 U15497 ( .A1(n12615), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20888), .ZN(n12387) );
  NAND2_X1 U15498 ( .A1(n12388), .A2(n12387), .ZN(n12390) );
  XNOR2_X1 U15499 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12440), .ZN(
        n14531) );
  NAND2_X1 U15500 ( .A1(n14192), .A2(n14531), .ZN(n12389) );
  NAND2_X1 U15501 ( .A1(n12390), .A2(n12389), .ZN(n14534) );
  NAND2_X1 U15502 ( .A1(n12392), .A2(n12391), .ZN(n14520) );
  INV_X1 U15503 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12588) );
  NAND2_X1 U15504 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12394) );
  NAND2_X1 U15505 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12393) );
  OAI211_X1 U15506 ( .C1(n12600), .C2(n12588), .A(n12394), .B(n12393), .ZN(
        n12395) );
  INV_X1 U15507 ( .A(n12395), .ZN(n12399) );
  AOI22_X1 U15508 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15509 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12397) );
  NAND2_X1 U15510 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12396) );
  NAND4_X1 U15511 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12405) );
  AOI22_X1 U15512 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15513 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15514 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15515 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12400) );
  NAND4_X1 U15516 ( .A1(n12403), .A2(n12402), .A3(n12401), .A4(n12400), .ZN(
        n12404) );
  OR2_X1 U15517 ( .A1(n12405), .A2(n12404), .ZN(n12443) );
  INV_X1 U15518 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U15519 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12407) );
  NAND2_X1 U15520 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12406) );
  OAI211_X1 U15521 ( .C1(n12600), .C2(n12408), .A(n12407), .B(n12406), .ZN(
        n12409) );
  INV_X1 U15522 ( .A(n12409), .ZN(n12413) );
  AOI22_X1 U15523 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15524 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12411) );
  NAND2_X1 U15525 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12410) );
  NAND4_X1 U15526 ( .A1(n12413), .A2(n12412), .A3(n12411), .A4(n12410), .ZN(
        n12419) );
  AOI22_X1 U15527 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15528 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15529 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15530 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12414) );
  NAND4_X1 U15531 ( .A1(n12417), .A2(n12416), .A3(n12415), .A4(n12414), .ZN(
        n12418) );
  OR2_X1 U15532 ( .A1(n12419), .A2(n12418), .ZN(n12444) );
  NAND2_X1 U15533 ( .A1(n12443), .A2(n12444), .ZN(n12456) );
  INV_X1 U15534 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15535 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12596), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12421) );
  NAND2_X1 U15536 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12420) );
  OAI211_X1 U15537 ( .C1(n12422), .C2(n12600), .A(n12421), .B(n12420), .ZN(
        n12423) );
  INV_X1 U15538 ( .A(n12423), .ZN(n12426) );
  AOI22_X1 U15539 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11901), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15540 ( .A1(n12565), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12424) );
  NAND3_X1 U15541 ( .A1(n12426), .A2(n12425), .A3(n12424), .ZN(n12433) );
  AOI22_X1 U15542 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15543 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12427), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U15544 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15545 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12590), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12428) );
  NAND4_X1 U15546 ( .A1(n12431), .A2(n12430), .A3(n12429), .A4(n12428), .ZN(
        n12432) );
  NOR2_X1 U15547 ( .A1(n12433), .A2(n12432), .ZN(n12457) );
  XOR2_X1 U15548 ( .A(n12456), .B(n12457), .Z(n12434) );
  NAND2_X1 U15549 ( .A1(n12434), .A2(n12605), .ZN(n12438) );
  INV_X1 U15550 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12435) );
  AOI21_X1 U15551 ( .B1(n12435), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12436) );
  AOI21_X1 U15552 ( .B1(n12615), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12436), .ZN(
        n12437) );
  NAND2_X1 U15553 ( .A1(n12438), .A2(n12437), .ZN(n12442) );
  INV_X1 U15554 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12439) );
  XNOR2_X1 U15555 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12453), .ZN(
        n14895) );
  NAND2_X1 U15556 ( .A1(n14192), .A2(n14895), .ZN(n12441) );
  NAND2_X1 U15557 ( .A1(n12442), .A2(n12441), .ZN(n14523) );
  XNOR2_X1 U15558 ( .A(n12444), .B(n12443), .ZN(n12448) );
  NAND2_X1 U15559 ( .A1(n20888), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12445) );
  NAND2_X1 U15560 ( .A1(n12609), .A2(n12445), .ZN(n12446) );
  AOI21_X1 U15561 ( .B1(n12615), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12446), .ZN(
        n12447) );
  OAI21_X1 U15562 ( .B1(n12574), .B2(n12448), .A(n12447), .ZN(n12451) );
  OAI21_X1 U15563 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n12449), .A(
        n12453), .ZN(n16096) );
  OR2_X1 U15564 ( .A1(n12609), .A2(n16096), .ZN(n12450) );
  NAND2_X1 U15565 ( .A1(n12451), .A2(n12450), .ZN(n14714) );
  OR2_X1 U15566 ( .A1(n12454), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12455) );
  NAND2_X1 U15567 ( .A1(n12479), .A2(n12455), .ZN(n16088) );
  NOR2_X1 U15568 ( .A1(n12457), .A2(n12456), .ZN(n12482) );
  INV_X1 U15569 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U15570 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12459) );
  NAND2_X1 U15571 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12458) );
  OAI211_X1 U15572 ( .C1(n12600), .C2(n12460), .A(n12459), .B(n12458), .ZN(
        n12461) );
  INV_X1 U15573 ( .A(n12461), .ZN(n12465) );
  AOI22_X1 U15574 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15575 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12463) );
  NAND2_X1 U15576 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12462) );
  NAND4_X1 U15577 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n12471) );
  AOI22_X1 U15578 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15579 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U15580 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15581 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12466) );
  NAND4_X1 U15582 ( .A1(n12469), .A2(n12468), .A3(n12467), .A4(n12466), .ZN(
        n12470) );
  OR2_X1 U15583 ( .A1(n12471), .A2(n12470), .ZN(n12481) );
  XNOR2_X1 U15584 ( .A(n12482), .B(n12481), .ZN(n12475) );
  INV_X1 U15585 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12472) );
  AOI21_X1 U15586 ( .B1(n12472), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12473) );
  AOI21_X1 U15587 ( .B1(n12615), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12473), .ZN(
        n12474) );
  OAI21_X1 U15588 ( .B1(n12475), .B2(n12574), .A(n12474), .ZN(n12476) );
  OAI21_X1 U15589 ( .B1(n16088), .B2(n12609), .A(n12476), .ZN(n12477) );
  INV_X1 U15590 ( .A(n12477), .ZN(n14703) );
  INV_X1 U15591 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U15592 ( .A1(n12479), .A2(n14889), .ZN(n12480) );
  AND2_X1 U15593 ( .A1(n12503), .A2(n12480), .ZN(n14891) );
  NAND2_X1 U15594 ( .A1(n12482), .A2(n12481), .ZN(n12505) );
  INV_X1 U15595 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15596 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12484) );
  NAND2_X1 U15597 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12483) );
  OAI211_X1 U15598 ( .C1(n12485), .C2(n12600), .A(n12484), .B(n12483), .ZN(
        n12486) );
  INV_X1 U15599 ( .A(n12486), .ZN(n12489) );
  AOI22_X1 U15600 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15601 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12487) );
  NAND3_X1 U15602 ( .A1(n12489), .A2(n12488), .A3(n12487), .ZN(n12496) );
  AOI22_X1 U15603 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15604 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15605 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15606 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12491) );
  NAND4_X1 U15607 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12495) );
  NOR2_X1 U15608 ( .A1(n12496), .A2(n12495), .ZN(n12506) );
  XOR2_X1 U15609 ( .A(n12505), .B(n12506), .Z(n12499) );
  INV_X1 U15610 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14796) );
  NAND2_X1 U15611 ( .A1(n20888), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12497) );
  OAI211_X1 U15612 ( .C1(n10208), .C2(n14796), .A(n12609), .B(n12497), .ZN(
        n12498) );
  AOI21_X1 U15613 ( .B1(n12499), .B2(n12605), .A(n12498), .ZN(n12500) );
  AOI21_X1 U15614 ( .B1(n14891), .B2(n14192), .A(n12500), .ZN(n14508) );
  INV_X1 U15615 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U15616 ( .A1(n12503), .A2(n12502), .ZN(n12504) );
  NAND2_X1 U15617 ( .A1(n12526), .A2(n12504), .ZN(n14880) );
  NOR2_X1 U15618 ( .A1(n12506), .A2(n12505), .ZN(n12529) );
  INV_X1 U15619 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12514) );
  INV_X1 U15620 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21046) );
  OAI22_X1 U15621 ( .A1(n11895), .A2(n21046), .B1(n12555), .B2(n12507), .ZN(
        n12511) );
  INV_X1 U15622 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12509) );
  OAI22_X1 U15623 ( .A1(n12559), .A2(n12509), .B1(n12589), .B2(n12508), .ZN(
        n12510) );
  AOI211_X1 U15624 ( .C1(n12490), .C2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n12511), .B(n12510), .ZN(n12513) );
  AOI22_X1 U15625 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12512) );
  OAI211_X1 U15626 ( .C1(n11945), .C2(n12514), .A(n12513), .B(n12512), .ZN(
        n12520) );
  AOI22_X1 U15627 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15628 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15629 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U15630 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12515) );
  NAND4_X1 U15631 ( .A1(n12518), .A2(n12517), .A3(n12516), .A4(n12515), .ZN(
        n12519) );
  OR2_X1 U15632 ( .A1(n12520), .A2(n12519), .ZN(n12528) );
  XNOR2_X1 U15633 ( .A(n12529), .B(n12528), .ZN(n12523) );
  OAI21_X1 U15634 ( .B1(n20789), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n20888), .ZN(n12522) );
  NAND2_X1 U15635 ( .A1(n12615), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12521) );
  OAI211_X1 U15636 ( .C1(n12523), .C2(n12574), .A(n12522), .B(n12521), .ZN(
        n12524) );
  OAI21_X1 U15637 ( .B1(n14880), .B2(n12609), .A(n12524), .ZN(n14496) );
  INV_X1 U15638 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13046) );
  INV_X1 U15639 ( .A(n12526), .ZN(n12525) );
  AOI21_X1 U15640 ( .B1(n13046), .B2(n12526), .A(n12547), .ZN(n14490) );
  NOR2_X1 U15641 ( .A1(n13046), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12527) );
  AOI211_X1 U15642 ( .C1(n12615), .C2(P1_EAX_REG_28__SCAN_IN), .A(n14192), .B(
        n12527), .ZN(n12546) );
  NAND2_X1 U15643 ( .A1(n12529), .A2(n12528), .ZN(n12551) );
  AOI22_X1 U15644 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15645 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15646 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15647 ( .A1(n12590), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12530) );
  NAND4_X1 U15648 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        n12543) );
  INV_X1 U15649 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15650 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U15651 ( .A1(n12553), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12534) );
  OAI211_X1 U15652 ( .C1(n12536), .C2(n12600), .A(n12535), .B(n12534), .ZN(
        n12537) );
  INV_X1 U15653 ( .A(n12537), .ZN(n12541) );
  AOI22_X1 U15654 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15655 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12539) );
  NAND3_X1 U15656 ( .A1(n12541), .A2(n12540), .A3(n12539), .ZN(n12542) );
  NOR2_X1 U15657 ( .A1(n12543), .A2(n12542), .ZN(n12552) );
  XOR2_X1 U15658 ( .A(n12551), .B(n12552), .Z(n12544) );
  NAND2_X1 U15659 ( .A1(n12544), .A2(n12605), .ZN(n12545) );
  INV_X1 U15660 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12548) );
  NAND2_X1 U15661 ( .A1(n12549), .A2(n12548), .ZN(n12550) );
  NAND2_X1 U15662 ( .A1(n12619), .A2(n12550), .ZN(n14871) );
  NOR2_X1 U15663 ( .A1(n12552), .A2(n12551), .ZN(n12604) );
  INV_X1 U15664 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12564) );
  INV_X1 U15665 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12556) );
  OAI22_X1 U15666 ( .A1(n11895), .A2(n12556), .B1(n12555), .B2(n12554), .ZN(
        n12561) );
  INV_X1 U15667 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12558) );
  OAI22_X1 U15668 ( .A1(n12559), .A2(n12558), .B1(n12589), .B2(n12557), .ZN(
        n12560) );
  AOI22_X1 U15669 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12562) );
  OAI211_X1 U15670 ( .C1(n12600), .C2(n12564), .A(n12563), .B(n12562), .ZN(
        n12571) );
  AOI22_X1 U15671 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15672 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12565), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15673 ( .A1(n12579), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12590), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15674 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12566) );
  NAND4_X1 U15675 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        n12570) );
  OR2_X1 U15676 ( .A1(n12571), .A2(n12570), .ZN(n12603) );
  XNOR2_X1 U15677 ( .A(n12604), .B(n12603), .ZN(n12575) );
  AOI21_X1 U15678 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20888), .A(
        n14192), .ZN(n12573) );
  NAND2_X1 U15679 ( .A1(n12615), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12572) );
  OAI211_X1 U15680 ( .C1(n12575), .C2(n12574), .A(n12573), .B(n12572), .ZN(
        n12576) );
  OAI21_X1 U15681 ( .B1(n14871), .B2(n12609), .A(n12576), .ZN(n14467) );
  XNOR2_X1 U15682 ( .A(n12619), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14459) );
  AOI22_X1 U15683 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15684 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12579), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15685 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15686 ( .A1(n12583), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12584) );
  NAND4_X1 U15687 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n12602) );
  INV_X1 U15688 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12599) );
  INV_X1 U15689 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21197) );
  OAI22_X1 U15690 ( .A1(n12589), .A2(n12588), .B1(n11855), .B2(n21197), .ZN(
        n12594) );
  INV_X1 U15691 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12592) );
  OAI22_X1 U15692 ( .A1(n11895), .A2(n12592), .B1(n12002), .B2(n12591), .ZN(
        n12593) );
  AOI22_X1 U15693 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12597) );
  OAI211_X1 U15694 ( .C1(n12600), .C2(n12599), .A(n12598), .B(n12597), .ZN(
        n12601) );
  NOR2_X1 U15695 ( .A1(n12602), .A2(n12601), .ZN(n12608) );
  NAND2_X1 U15696 ( .A1(n12604), .A2(n12603), .ZN(n12607) );
  OAI21_X1 U15697 ( .B1(n12608), .B2(n12607), .A(n12605), .ZN(n12606) );
  AOI21_X1 U15698 ( .B1(n12608), .B2(n12607), .A(n12606), .ZN(n12612) );
  INV_X1 U15699 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14773) );
  NAND2_X1 U15700 ( .A1(n20888), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12610) );
  OAI211_X1 U15701 ( .C1(n10208), .C2(n14773), .A(n12610), .B(n12609), .ZN(
        n12611) );
  NOR2_X1 U15702 ( .A1(n12612), .A2(n12611), .ZN(n12613) );
  NAND2_X1 U15703 ( .A1(n14466), .A2(n12804), .ZN(n12618) );
  AOI22_X1 U15704 ( .A1(n12615), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12614), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12616) );
  INV_X1 U15705 ( .A(n12616), .ZN(n12617) );
  NAND2_X1 U15706 ( .A1(n20885), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16318) );
  NAND2_X1 U15707 ( .A1(n20888), .A2(n20701), .ZN(n20822) );
  NAND2_X1 U15708 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20829), .ZN(n13840) );
  INV_X1 U15709 ( .A(n20258), .ZN(n20194) );
  INV_X1 U15710 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12806) );
  INV_X1 U15711 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12620) );
  INV_X1 U15712 ( .A(n12622), .ZN(n13468) );
  NAND2_X1 U15713 ( .A1(n15030), .A2(n14197), .ZN(n12623) );
  NAND3_X1 U15714 ( .A1(n12952), .A2(n13468), .A3(n12623), .ZN(n12844) );
  NAND2_X1 U15715 ( .A1(n15963), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20012) );
  INV_X1 U15716 ( .A(n20012), .ZN(n14132) );
  NAND2_X1 U15717 ( .A1(n12624), .A2(n14132), .ZN(n12625) );
  NOR2_X1 U15718 ( .A1(n12844), .A2(n12625), .ZN(n12678) );
  XNOR2_X1 U15719 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12637) );
  NAND2_X1 U15720 ( .A1(n20755), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12641) );
  INV_X1 U15721 ( .A(n12641), .ZN(n12636) );
  NAND2_X1 U15722 ( .A1(n12637), .A2(n12636), .ZN(n12627) );
  NAND2_X1 U15723 ( .A1(n20693), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12626) );
  NAND2_X1 U15724 ( .A1(n12627), .A2(n12626), .ZN(n12652) );
  XNOR2_X1 U15725 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12651) );
  NAND2_X1 U15726 ( .A1(n12652), .A2(n12651), .ZN(n12629) );
  NAND2_X1 U15727 ( .A1(n20611), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12628) );
  NAND2_X1 U15728 ( .A1(n12629), .A2(n12628), .ZN(n12635) );
  XNOR2_X1 U15729 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12634) );
  NAND2_X1 U15730 ( .A1(n12635), .A2(n12634), .ZN(n12631) );
  NAND2_X1 U15731 ( .A1(n20652), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12630) );
  NAND2_X1 U15732 ( .A1(n12631), .A2(n12630), .ZN(n12665) );
  NOR2_X1 U15733 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16315), .ZN(
        n12632) );
  OR2_X1 U15734 ( .A1(n12665), .A2(n12632), .ZN(n12633) );
  INV_X1 U15735 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20250) );
  OR2_X1 U15736 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20250), .ZN(
        n12664) );
  NAND2_X1 U15737 ( .A1(n12663), .A2(n12820), .ZN(n12677) );
  NAND2_X1 U15738 ( .A1(n12820), .A2(n12640), .ZN(n12675) );
  XNOR2_X1 U15739 ( .A(n12635), .B(n12634), .ZN(n12815) );
  XNOR2_X1 U15740 ( .A(n12637), .B(n12636), .ZN(n12817) );
  NAND2_X1 U15741 ( .A1(n12640), .A2(n20272), .ZN(n12639) );
  NAND2_X1 U15742 ( .A1(n11767), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12638) );
  NOR2_X1 U15743 ( .A1(n12817), .A2(n12648), .ZN(n12647) );
  OAI21_X1 U15744 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20755), .A(
        n12641), .ZN(n12643) );
  NOR2_X1 U15745 ( .A1(n12658), .A2(n12643), .ZN(n12646) );
  INV_X1 U15746 ( .A(n12624), .ZN(n12843) );
  NAND2_X1 U15747 ( .A1(n11767), .A2(n20261), .ZN(n12642) );
  NAND2_X1 U15748 ( .A1(n12642), .A2(n11824), .ZN(n12657) );
  INV_X1 U15749 ( .A(n12643), .ZN(n12644) );
  OAI211_X1 U15750 ( .C1(n14197), .C2(n12843), .A(n12657), .B(n12644), .ZN(
        n12645) );
  OAI21_X1 U15751 ( .B1(n12663), .B2(n12646), .A(n12645), .ZN(n12649) );
  NAND2_X1 U15752 ( .A1(n12647), .A2(n12649), .ZN(n12656) );
  INV_X1 U15753 ( .A(n12648), .ZN(n12650) );
  OAI211_X1 U15754 ( .C1(n12650), .C2(n12649), .A(n12817), .B(n12667), .ZN(
        n12655) );
  XNOR2_X1 U15755 ( .A(n12652), .B(n12651), .ZN(n12816) );
  NAND2_X1 U15756 ( .A1(n12669), .A2(n12816), .ZN(n12653) );
  OAI211_X1 U15757 ( .C1(n12658), .C2(n12816), .A(n12653), .B(n12657), .ZN(
        n12654) );
  NAND3_X1 U15758 ( .A1(n12656), .A2(n12655), .A3(n12654), .ZN(n12660) );
  AOI22_X1 U15759 ( .A1(n12661), .A2(n12815), .B1(n12660), .B2(n12659), .ZN(
        n12662) );
  AOI21_X1 U15760 ( .B1(n12663), .B2(n12815), .A(n12662), .ZN(n12672) );
  NOR2_X1 U15761 ( .A1(n12665), .A2(n12664), .ZN(n12818) );
  INV_X1 U15762 ( .A(n12818), .ZN(n12666) );
  NOR2_X1 U15763 ( .A1(n12669), .A2(n12666), .ZN(n12671) );
  INV_X1 U15764 ( .A(n12667), .ZN(n12668) );
  NAND3_X1 U15765 ( .A1(n12669), .A2(n12668), .A3(n12818), .ZN(n12670) );
  OAI21_X1 U15766 ( .B1(n12672), .B2(n12671), .A(n12670), .ZN(n12673) );
  AOI21_X1 U15767 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20885), .A(
        n12673), .ZN(n12674) );
  NAND2_X1 U15768 ( .A1(n12675), .A2(n12674), .ZN(n12676) );
  NAND2_X1 U15769 ( .A1(n12683), .A2(n20822), .ZN(n20977) );
  AND2_X1 U15770 ( .A1(n20977), .A2(n20885), .ZN(n12679) );
  NAND2_X1 U15771 ( .A1(n20885), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12681) );
  NAND2_X1 U15772 ( .A1(n20789), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12680) );
  AND2_X1 U15773 ( .A1(n12681), .A2(n12680), .ZN(n20191) );
  INV_X1 U15774 ( .A(n20191), .ZN(n12682) );
  INV_X2 U15775 ( .A(n20190), .ZN(n20180) );
  OR2_X1 U15776 ( .A1(n12683), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16230) );
  INV_X1 U15777 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20951) );
  NOR2_X1 U15778 ( .A1(n16230), .A2(n20951), .ZN(n14285) );
  AOI21_X1 U15779 ( .B1(n20180), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14285), .ZN(n12684) );
  OAI21_X1 U15780 ( .B1(n14215), .B2(n20179), .A(n12684), .ZN(n12685) );
  AOI21_X1 U15781 ( .B1(n14439), .B2(n20194), .A(n12685), .ZN(n12796) );
  INV_X1 U15782 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12775) );
  INV_X1 U15783 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12914) );
  INV_X1 U15784 ( .A(n12758), .ZN(n12742) );
  NAND2_X1 U15785 ( .A1(n14197), .A2(n20284), .ZN(n12700) );
  OAI21_X1 U15786 ( .B1(n20982), .B2(n12690), .A(n12700), .ZN(n12687) );
  INV_X1 U15787 ( .A(n12687), .ZN(n12688) );
  NAND2_X1 U15788 ( .A1(n12689), .A2(n12690), .ZN(n12707) );
  OAI21_X1 U15789 ( .B1(n12690), .B2(n12689), .A(n12707), .ZN(n12692) );
  INV_X1 U15790 ( .A(n12693), .ZN(n12694) );
  NAND2_X1 U15791 ( .A1(n20182), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20181) );
  INV_X1 U15792 ( .A(n12696), .ZN(n12698) );
  NAND2_X1 U15793 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  NAND2_X1 U15794 ( .A1(n20181), .A2(n12699), .ZN(n12704) );
  INV_X1 U15795 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21112) );
  XNOR2_X1 U15796 ( .A(n12704), .B(n21112), .ZN(n13792) );
  XNOR2_X1 U15797 ( .A(n12707), .B(n12706), .ZN(n12702) );
  INV_X1 U15798 ( .A(n20982), .ZN(n12749) );
  INV_X1 U15799 ( .A(n12700), .ZN(n12701) );
  AOI21_X1 U15800 ( .B1(n12702), .B2(n12749), .A(n12701), .ZN(n12703) );
  OAI21_X1 U15801 ( .B1(n13828), .B2(n12758), .A(n12703), .ZN(n13793) );
  NAND2_X1 U15802 ( .A1(n13793), .A2(n13792), .ZN(n13794) );
  NAND2_X1 U15803 ( .A1(n12704), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12705) );
  INV_X1 U15804 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20200) );
  XNOR2_X1 U15805 ( .A(n12712), .B(n20200), .ZN(n13954) );
  NAND2_X1 U15806 ( .A1(n9752), .A2(n12742), .ZN(n12711) );
  NAND2_X1 U15807 ( .A1(n12707), .A2(n12706), .ZN(n12715) );
  INV_X1 U15808 ( .A(n12716), .ZN(n12708) );
  XNOR2_X1 U15809 ( .A(n12715), .B(n12708), .ZN(n12709) );
  NAND2_X1 U15810 ( .A1(n12709), .A2(n12749), .ZN(n12710) );
  NAND2_X1 U15811 ( .A1(n12711), .A2(n12710), .ZN(n13953) );
  NAND2_X1 U15812 ( .A1(n13954), .A2(n13953), .ZN(n13952) );
  NAND2_X1 U15813 ( .A1(n12712), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12713) );
  OR2_X1 U15814 ( .A1(n12714), .A2(n12758), .ZN(n12719) );
  NAND2_X1 U15815 ( .A1(n12716), .A2(n12715), .ZN(n12724) );
  XNOR2_X1 U15816 ( .A(n12723), .B(n12724), .ZN(n12717) );
  NAND2_X1 U15817 ( .A1(n12749), .A2(n12717), .ZN(n12718) );
  NAND2_X1 U15818 ( .A1(n12719), .A2(n12718), .ZN(n12720) );
  INV_X1 U15819 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20201) );
  XNOR2_X1 U15820 ( .A(n12720), .B(n20201), .ZN(n20172) );
  NAND2_X1 U15821 ( .A1(n20173), .A2(n20172), .ZN(n20171) );
  NAND2_X1 U15822 ( .A1(n12720), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12721) );
  OR2_X1 U15823 ( .A1(n12722), .A2(n12758), .ZN(n12729) );
  INV_X1 U15824 ( .A(n12723), .ZN(n12725) );
  NOR2_X1 U15825 ( .A1(n12725), .A2(n12724), .ZN(n12734) );
  INV_X1 U15826 ( .A(n12734), .ZN(n12726) );
  XNOR2_X1 U15827 ( .A(n12733), .B(n12726), .ZN(n12727) );
  NAND2_X1 U15828 ( .A1(n12749), .A2(n12727), .ZN(n12728) );
  NAND2_X1 U15829 ( .A1(n12729), .A2(n12728), .ZN(n12730) );
  INV_X1 U15830 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16279) );
  XNOR2_X1 U15831 ( .A(n12730), .B(n16279), .ZN(n16157) );
  NAND2_X1 U15832 ( .A1(n12730), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12731) );
  NAND3_X1 U15833 ( .A1(n12761), .A2(n12742), .A3(n12732), .ZN(n12737) );
  NAND2_X1 U15834 ( .A1(n12734), .A2(n12733), .ZN(n12745) );
  XNOR2_X1 U15835 ( .A(n12744), .B(n12745), .ZN(n12735) );
  NAND2_X1 U15836 ( .A1(n12749), .A2(n12735), .ZN(n12736) );
  INV_X1 U15837 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16150) );
  NAND2_X1 U15838 ( .A1(n16151), .A2(n16150), .ZN(n12738) );
  INV_X1 U15839 ( .A(n16151), .ZN(n12739) );
  NAND2_X1 U15840 ( .A1(n12739), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12740) );
  NAND2_X1 U15841 ( .A1(n12741), .A2(n12740), .ZN(n16144) );
  NAND2_X1 U15842 ( .A1(n12743), .A2(n12742), .ZN(n12751) );
  INV_X1 U15843 ( .A(n12744), .ZN(n12746) );
  NOR2_X1 U15844 ( .A1(n12746), .A2(n12745), .ZN(n12762) );
  INV_X1 U15845 ( .A(n12762), .ZN(n12747) );
  XNOR2_X1 U15846 ( .A(n12763), .B(n12747), .ZN(n12748) );
  NAND2_X1 U15847 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  NAND2_X1 U15848 ( .A1(n12751), .A2(n12750), .ZN(n12753) );
  XNOR2_X1 U15849 ( .A(n12753), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16145) );
  INV_X1 U15850 ( .A(n16145), .ZN(n12752) );
  INV_X1 U15851 ( .A(n12753), .ZN(n12755) );
  INV_X1 U15852 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12754) );
  NAND2_X1 U15853 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  INV_X1 U15854 ( .A(n12763), .ZN(n12757) );
  NOR3_X1 U15855 ( .A1(n12759), .A2(n12758), .A3(n12757), .ZN(n12760) );
  NAND2_X1 U15856 ( .A1(n12763), .A2(n12762), .ZN(n12764) );
  NOR2_X1 U15857 ( .A1(n20982), .A2(n12764), .ZN(n12765) );
  INV_X1 U15858 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12766) );
  INV_X1 U15859 ( .A(n12767), .ZN(n12768) );
  OR2_X2 U15860 ( .A1(n14974), .A2(n12769), .ZN(n14967) );
  INV_X1 U15861 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16275) );
  BUF_X4 U15862 ( .A(n12771), .Z(n16121) );
  NOR2_X1 U15863 ( .A1(n12771), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14958) );
  AOI21_X1 U15864 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n12771), .ZN(n14954) );
  NAND2_X1 U15865 ( .A1(n12771), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14943) );
  INV_X1 U15866 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14945) );
  NAND2_X1 U15867 ( .A1(n16134), .A2(n14945), .ZN(n12772) );
  NAND2_X1 U15868 ( .A1(n16121), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12773) );
  NAND2_X1 U15869 ( .A1(n16121), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12774) );
  MUX2_X1 U15870 ( .A(n12775), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .S(
        n16121), .Z(n14932) );
  NOR2_X1 U15871 ( .A1(n14932), .A2(n16120), .ZN(n12776) );
  NAND2_X1 U15872 ( .A1(n12777), .A2(n12776), .ZN(n16109) );
  INV_X1 U15873 ( .A(n14931), .ZN(n12780) );
  NAND2_X1 U15874 ( .A1(n16121), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14956) );
  INV_X1 U15875 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12778) );
  INV_X1 U15876 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16137) );
  NAND2_X1 U15877 ( .A1(n12778), .A2(n16137), .ZN(n12779) );
  NAND2_X1 U15878 ( .A1(n16121), .A2(n12779), .ZN(n14953) );
  NAND2_X1 U15879 ( .A1(n14956), .A2(n14953), .ZN(n14941) );
  INV_X1 U15880 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16208) );
  XNOR2_X1 U15881 ( .A(n16121), .B(n16208), .ZN(n14921) );
  AND2_X1 U15882 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U15883 ( .A1(n15995), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12781) );
  OAI21_X2 U15884 ( .B1(n14911), .B2(n12781), .A(n16134), .ZN(n14903) );
  INV_X1 U15885 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12783) );
  INV_X1 U15886 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16102) );
  INV_X1 U15887 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15980) );
  NAND4_X1 U15888 ( .A1(n12783), .A2(n16102), .A3(n15980), .A4(n16208), .ZN(
        n12784) );
  INV_X1 U15889 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16089) );
  INV_X1 U15890 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16083) );
  INV_X1 U15891 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U15892 ( .A1(n16083), .A2(n12813), .ZN(n13037) );
  OAI21_X1 U15893 ( .B1(n16080), .B2(n13037), .A(n16121), .ZN(n14887) );
  NAND3_X1 U15894 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14885) );
  INV_X1 U15895 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14282) );
  AOI21_X1 U15896 ( .B1(n12785), .B2(n14885), .A(n14282), .ZN(n14875) );
  NAND2_X1 U15897 ( .A1(n12786), .A2(n16134), .ZN(n12811) );
  NAND2_X1 U15898 ( .A1(n14875), .A2(n12811), .ZN(n12787) );
  NAND2_X1 U15899 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14988) );
  NOR2_X2 U15900 ( .A1(n9842), .A2(n14988), .ZN(n12799) );
  INV_X1 U15901 ( .A(n12799), .ZN(n12791) );
  NOR2_X1 U15902 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15003) );
  NAND2_X1 U15903 ( .A1(n9842), .A2(n15003), .ZN(n12797) );
  INV_X1 U15904 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12789) );
  NAND2_X1 U15905 ( .A1(n14867), .A2(n12789), .ZN(n12793) );
  XOR2_X1 U15906 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n16121), .Z(
        n14869) );
  OAI21_X1 U15907 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12789), .A(
        n14869), .ZN(n12790) );
  NAND2_X1 U15908 ( .A1(n12793), .A2(n12792), .ZN(n12795) );
  NOR2_X1 U15909 ( .A1(n12797), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U15910 ( .A1(n12798), .A2(n16121), .ZN(n12802) );
  AND2_X1 U15911 ( .A1(n12799), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12800) );
  INV_X1 U15912 ( .A(n12804), .ZN(n12805) );
  XNOR2_X1 U15913 ( .A(n14466), .B(n12805), .ZN(n14450) );
  INV_X1 U15914 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21043) );
  NOR2_X1 U15915 ( .A1(n16230), .A2(n21043), .ZN(n14981) );
  NOR2_X1 U15916 ( .A1(n20190), .A2(n12806), .ZN(n12807) );
  AOI211_X1 U15917 ( .C1(n14459), .C2(n20185), .A(n14981), .B(n12807), .ZN(
        n12808) );
  INV_X1 U15918 ( .A(n12808), .ZN(n12809) );
  AOI21_X1 U15919 ( .B1(n14450), .B2(n20194), .A(n12809), .ZN(n12810) );
  OAI21_X1 U15920 ( .B1(n14987), .B2(n20198), .A(n12810), .ZN(P1_U2969) );
  NAND2_X1 U15921 ( .A1(n12811), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16082) );
  NAND2_X1 U15922 ( .A1(n16082), .A2(n14884), .ZN(n12812) );
  MUX2_X1 U15923 ( .A(n12812), .B(n16082), .S(n16134), .Z(n12814) );
  XNOR2_X1 U15924 ( .A(n12814), .B(n12813), .ZN(n14901) );
  INV_X1 U15925 ( .A(n14901), .ZN(n12849) );
  NOR4_X1 U15926 ( .A1(n12818), .A2(n12817), .A3(n12816), .A4(n12815), .ZN(
        n12819) );
  NOR2_X1 U15927 ( .A1(n12820), .A2(n12819), .ZN(n13472) );
  NAND2_X1 U15928 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20978) );
  NAND2_X1 U15929 ( .A1(n13472), .A2(n20978), .ZN(n13638) );
  INV_X1 U15930 ( .A(n12821), .ZN(n12822) );
  INV_X1 U15931 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20897) );
  NAND2_X1 U15932 ( .A1(n12822), .A2(n20897), .ZN(n15993) );
  AND2_X1 U15933 ( .A1(n20272), .A2(n15993), .ZN(n12823) );
  OR2_X1 U15934 ( .A1(n13638), .A2(n12823), .ZN(n12830) );
  AOI21_X1 U15935 ( .B1(n12824), .B2(n20978), .A(n14197), .ZN(n12827) );
  INV_X1 U15936 ( .A(n15993), .ZN(n15960) );
  NOR2_X1 U15937 ( .A1(n20982), .A2(n15960), .ZN(n12826) );
  OAI21_X1 U15938 ( .B1(n12827), .B2(n12826), .A(n12825), .ZN(n12828) );
  NAND2_X1 U15939 ( .A1(n12828), .A2(n14128), .ZN(n12829) );
  MUX2_X1 U15940 ( .A(n12830), .B(n12829), .S(n12691), .Z(n12840) );
  INV_X1 U15941 ( .A(n12844), .ZN(n12833) );
  OR2_X1 U15942 ( .A1(n12832), .A2(n12833), .ZN(n12836) );
  NAND2_X1 U15943 ( .A1(n9801), .A2(n20272), .ZN(n12944) );
  AND2_X1 U15944 ( .A1(n12944), .A2(n20261), .ZN(n12834) );
  NAND2_X1 U15945 ( .A1(n12835), .A2(n12834), .ZN(n12955) );
  NAND2_X1 U15946 ( .A1(n12836), .A2(n12955), .ZN(n13643) );
  INV_X1 U15947 ( .A(n13643), .ZN(n12839) );
  INV_X1 U15948 ( .A(n15030), .ZN(n12837) );
  NAND3_X1 U15949 ( .A1(n13646), .A2(n12837), .A3(n20272), .ZN(n12838) );
  NAND3_X1 U15950 ( .A1(n12840), .A2(n12839), .A3(n12838), .ZN(n12841) );
  INV_X1 U15951 ( .A(n12842), .ZN(n12846) );
  NOR2_X1 U15952 ( .A1(n12844), .A2(n14650), .ZN(n13639) );
  NOR2_X1 U15953 ( .A1(n12844), .A2(n12843), .ZN(n15951) );
  OR2_X1 U15954 ( .A1(n13639), .A2(n15951), .ZN(n13471) );
  INV_X1 U15955 ( .A(n13471), .ZN(n12845) );
  OAI211_X1 U15956 ( .C1(n12847), .C2(n9853), .A(n12846), .B(n12845), .ZN(
        n12848) );
  NAND2_X1 U15957 ( .A1(n12963), .A2(n12848), .ZN(n16291) );
  MUX2_X1 U15958 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12852) );
  OR2_X1 U15959 ( .A1(n9815), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12851) );
  NAND2_X1 U15960 ( .A1(n12852), .A2(n12851), .ZN(n12854) );
  INV_X1 U15961 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14686) );
  OAI22_X1 U15962 ( .A1(n14296), .A2(n14686), .B1(n14291), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13730) );
  XNOR2_X1 U15963 ( .A(n12854), .B(n13730), .ZN(n14678) );
  INV_X1 U15964 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21194) );
  NAND2_X1 U15965 ( .A1(n12875), .A2(n21194), .ZN(n12858) );
  NAND2_X1 U15966 ( .A1(n9818), .A2(n21194), .ZN(n12856) );
  NAND2_X1 U15967 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12855) );
  NAND3_X1 U15968 ( .A1(n12856), .A2(n14296), .A3(n12855), .ZN(n12857) );
  AND2_X2 U15969 ( .A1(n13798), .A2(n13797), .ZN(n20086) );
  INV_X1 U15970 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21063) );
  NAND2_X1 U15971 ( .A1(n12875), .A2(n21063), .ZN(n12862) );
  NAND2_X1 U15972 ( .A1(n9818), .A2(n21063), .ZN(n12860) );
  NAND2_X1 U15973 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12859) );
  NAND3_X1 U15974 ( .A1(n12860), .A2(n14296), .A3(n12859), .ZN(n12861) );
  AND2_X1 U15975 ( .A1(n12862), .A2(n12861), .ZN(n20087) );
  INV_X1 U15976 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12864) );
  NAND2_X1 U15977 ( .A1(n14295), .A2(n12864), .ZN(n12868) );
  NAND2_X1 U15978 ( .A1(n14296), .A2(n20200), .ZN(n12866) );
  NAND2_X1 U15979 ( .A1(n9818), .A2(n12864), .ZN(n12865) );
  NAND3_X1 U15980 ( .A1(n12866), .A2(n14291), .A3(n12865), .ZN(n12867) );
  NAND2_X1 U15981 ( .A1(n12868), .A2(n12867), .ZN(n20085) );
  NAND2_X1 U15982 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U15983 ( .A1(n14296), .A2(n12870), .ZN(n12873) );
  INV_X1 U15984 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12871) );
  NAND2_X1 U15985 ( .A1(n9818), .A2(n12871), .ZN(n12872) );
  NAND2_X1 U15986 ( .A1(n12873), .A2(n12872), .ZN(n12874) );
  OAI21_X1 U15987 ( .B1(n14306), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12874), .ZN(
        n16298) );
  INV_X1 U15988 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20111) );
  NAND2_X1 U15989 ( .A1(n12875), .A2(n20111), .ZN(n12879) );
  NAND2_X1 U15990 ( .A1(n9818), .A2(n20111), .ZN(n12877) );
  NAND2_X1 U15991 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12876) );
  NAND3_X1 U15992 ( .A1(n12877), .A2(n14296), .A3(n12876), .ZN(n12878) );
  NAND2_X1 U15993 ( .A1(n16298), .A2(n16297), .ZN(n12880) );
  NOR2_X2 U15994 ( .A1(n13990), .A2(n12880), .ZN(n16300) );
  NAND2_X1 U15995 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12881) );
  NAND2_X1 U15996 ( .A1(n14296), .A2(n12881), .ZN(n12883) );
  INV_X1 U15997 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U15998 ( .A1(n9818), .A2(n14165), .ZN(n12882) );
  NAND2_X1 U15999 ( .A1(n12883), .A2(n12882), .ZN(n12884) );
  OAI21_X1 U16000 ( .B1(n14306), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12884), .ZN(
        n14159) );
  INV_X1 U16001 ( .A(n14176), .ZN(n12889) );
  INV_X1 U16002 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14208) );
  NAND2_X1 U16003 ( .A1(n9818), .A2(n14208), .ZN(n12886) );
  NAND2_X1 U16004 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12885) );
  NAND3_X1 U16005 ( .A1(n12886), .A2(n14296), .A3(n12885), .ZN(n12887) );
  OAI21_X1 U16006 ( .B1(n14301), .B2(P1_EBX_REG_8__SCAN_IN), .A(n12887), .ZN(
        n14177) );
  INV_X1 U16007 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14243) );
  NAND2_X1 U16008 ( .A1(n9818), .A2(n14243), .ZN(n12892) );
  NAND2_X1 U16009 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12890) );
  NAND2_X1 U16010 ( .A1(n14296), .A2(n12890), .ZN(n12891) );
  AOI22_X1 U16011 ( .A1(n14295), .A2(n14243), .B1(n12892), .B2(n12891), .ZN(
        n14242) );
  MUX2_X1 U16012 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12893) );
  INV_X1 U16013 ( .A(n12893), .ZN(n12895) );
  NOR2_X1 U16014 ( .A1(n9815), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12894) );
  NOR2_X1 U16015 ( .A1(n12895), .A2(n12894), .ZN(n14639) );
  INV_X1 U16016 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U16017 ( .A1(n14295), .A2(n16079), .ZN(n12899) );
  NAND2_X1 U16018 ( .A1(n14296), .A2(n16137), .ZN(n12897) );
  NAND2_X1 U16019 ( .A1(n9818), .A2(n16079), .ZN(n12896) );
  NAND3_X1 U16020 ( .A1(n12897), .A2(n14291), .A3(n12896), .ZN(n12898) );
  INV_X1 U16021 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16077) );
  NAND2_X1 U16022 ( .A1(n9818), .A2(n16077), .ZN(n12901) );
  NAND2_X1 U16023 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12900) );
  NAND3_X1 U16024 ( .A1(n12901), .A2(n14296), .A3(n12900), .ZN(n12902) );
  OAI21_X1 U16025 ( .B1(n14301), .B2(P1_EBX_REG_12__SCAN_IN), .A(n12902), .ZN(
        n15013) );
  INV_X1 U16026 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U16027 ( .A1(n14295), .A2(n14764), .ZN(n12907) );
  INV_X1 U16028 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12903) );
  NAND2_X1 U16029 ( .A1(n14296), .A2(n12903), .ZN(n12905) );
  NAND2_X1 U16030 ( .A1(n9818), .A2(n14764), .ZN(n12904) );
  NAND3_X1 U16031 ( .A1(n12905), .A2(n14291), .A3(n12904), .ZN(n12906) );
  AND2_X1 U16032 ( .A1(n12907), .A2(n12906), .ZN(n14628) );
  MUX2_X1 U16033 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12908) );
  OAI21_X1 U16034 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n9815), .A(
        n12908), .ZN(n14612) );
  INV_X1 U16035 ( .A(n14612), .ZN(n12909) );
  AND2_X2 U16036 ( .A1(n14629), .A2(n12909), .ZN(n14757) );
  INV_X1 U16037 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16224) );
  NAND2_X1 U16038 ( .A1(n14296), .A2(n16224), .ZN(n12911) );
  INV_X1 U16039 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n16053) );
  NAND2_X1 U16040 ( .A1(n9818), .A2(n16053), .ZN(n12910) );
  NAND3_X1 U16041 ( .A1(n12911), .A2(n14291), .A3(n12910), .ZN(n12912) );
  OAI21_X1 U16042 ( .B1(n14306), .B2(P1_EBX_REG_15__SCAN_IN), .A(n12912), .ZN(
        n14756) );
  MUX2_X1 U16043 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12913) );
  OAI21_X1 U16044 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n9815), .A(
        n12913), .ZN(n14595) );
  INV_X1 U16045 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16045) );
  NAND2_X1 U16046 ( .A1(n14295), .A2(n16045), .ZN(n12918) );
  NAND2_X1 U16047 ( .A1(n14296), .A2(n12914), .ZN(n12916) );
  NAND2_X1 U16048 ( .A1(n9818), .A2(n16045), .ZN(n12915) );
  NAND3_X1 U16049 ( .A1(n12916), .A2(n14291), .A3(n12915), .ZN(n12917) );
  AND2_X1 U16050 ( .A1(n12918), .A2(n12917), .ZN(n14745) );
  INV_X1 U16051 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14585) );
  NAND2_X1 U16052 ( .A1(n9818), .A2(n14585), .ZN(n12920) );
  NAND2_X1 U16053 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12919) );
  NAND3_X1 U16054 ( .A1(n12920), .A2(n14296), .A3(n12919), .ZN(n12921) );
  OAI21_X1 U16055 ( .B1(n14301), .B2(P1_EBX_REG_18__SCAN_IN), .A(n12921), .ZN(
        n14581) );
  NAND2_X1 U16056 ( .A1(n14296), .A2(n16102), .ZN(n12923) );
  INV_X1 U16057 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14737) );
  NAND2_X1 U16058 ( .A1(n9818), .A2(n14737), .ZN(n12922) );
  NAND3_X1 U16059 ( .A1(n12923), .A2(n14291), .A3(n12922), .ZN(n12924) );
  OAI21_X1 U16060 ( .B1(n14306), .B2(P1_EBX_REG_19__SCAN_IN), .A(n12924), .ZN(
        n14564) );
  INV_X1 U16061 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U16062 ( .A1(n9818), .A2(n14734), .ZN(n12926) );
  NAND2_X1 U16063 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12925) );
  NAND3_X1 U16064 ( .A1(n12926), .A2(n14296), .A3(n12925), .ZN(n12927) );
  OAI21_X1 U16065 ( .B1(n14301), .B2(P1_EBX_REG_20__SCAN_IN), .A(n12927), .ZN(
        n14554) );
  INV_X1 U16066 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14731) );
  NAND2_X1 U16067 ( .A1(n14295), .A2(n14731), .ZN(n12931) );
  NAND2_X1 U16068 ( .A1(n14296), .A2(n15980), .ZN(n12929) );
  NAND2_X1 U16069 ( .A1(n9818), .A2(n14731), .ZN(n12928) );
  NAND3_X1 U16070 ( .A1(n12929), .A2(n14291), .A3(n12928), .ZN(n12930) );
  AND2_X1 U16071 ( .A1(n12931), .A2(n12930), .ZN(n14728) );
  MUX2_X1 U16072 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12932) );
  OAI21_X1 U16073 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n9815), .A(
        n12932), .ZN(n12933) );
  INV_X1 U16074 ( .A(n12933), .ZN(n14535) );
  NAND2_X1 U16075 ( .A1(n14296), .A2(n16089), .ZN(n12935) );
  INV_X1 U16076 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14721) );
  NAND3_X1 U16077 ( .A1(n12935), .A2(n14291), .A3(n12934), .ZN(n12936) );
  OAI21_X1 U16078 ( .B1(n14306), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12936), .ZN(
        n14717) );
  MUX2_X1 U16079 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12937) );
  OAI21_X1 U16080 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n9815), .A(
        n12937), .ZN(n12938) );
  AND2_X1 U16081 ( .A1(n14720), .A2(n12938), .ZN(n12939) );
  OR2_X1 U16082 ( .A1(n14706), .A2(n12939), .ZN(n14712) );
  INV_X1 U16083 ( .A(n14712), .ZN(n12978) );
  INV_X1 U16084 ( .A(n12940), .ZN(n12941) );
  NAND2_X1 U16085 ( .A1(n12941), .A2(n11824), .ZN(n15965) );
  OAI21_X1 U16086 ( .B1(n9853), .B2(n11823), .A(n15965), .ZN(n12942) );
  INV_X1 U16087 ( .A(n12943), .ZN(n12946) );
  INV_X1 U16088 ( .A(n12944), .ZN(n12945) );
  NAND2_X1 U16089 ( .A1(n12946), .A2(n12945), .ZN(n13637) );
  INV_X1 U16090 ( .A(n13637), .ZN(n12947) );
  AND2_X1 U16091 ( .A1(n12832), .A2(n20272), .ZN(n15940) );
  NAND2_X1 U16092 ( .A1(n11831), .A2(n13480), .ZN(n12957) );
  INV_X1 U16093 ( .A(n12948), .ZN(n12949) );
  NOR2_X1 U16094 ( .A1(n12950), .A2(n12949), .ZN(n12956) );
  OAI211_X1 U16095 ( .C1(n12624), .C2(n20261), .A(n12952), .B(n12951), .ZN(
        n12953) );
  NAND2_X1 U16096 ( .A1(n12953), .A2(n20272), .ZN(n12954) );
  NAND4_X1 U16097 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n13615) );
  INV_X1 U16098 ( .A(n13615), .ZN(n12959) );
  OAI211_X1 U16099 ( .C1(n13611), .C2(n20261), .A(n12959), .B(n12958), .ZN(
        n12960) );
  INV_X1 U16100 ( .A(n13801), .ZN(n12961) );
  NAND2_X1 U16101 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16194) );
  NOR2_X1 U16102 ( .A1(n15999), .A2(n14277), .ZN(n16283) );
  INV_X1 U16103 ( .A(n16283), .ZN(n20219) );
  NAND2_X1 U16104 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16280) );
  NOR2_X1 U16105 ( .A1(n20201), .A2(n20200), .ZN(n20199) );
  NAND2_X1 U16106 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20199), .ZN(
        n15019) );
  NOR2_X1 U16107 ( .A1(n16280), .A2(n15019), .ZN(n16261) );
  NAND3_X1 U16108 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16262) );
  NOR3_X1 U16109 ( .A1(n12778), .A2(n16275), .A3(n16262), .ZN(n16238) );
  NAND2_X1 U16110 ( .A1(n16261), .A2(n16238), .ZN(n15016) );
  NAND2_X1 U16111 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16239) );
  NOR2_X1 U16112 ( .A1(n15016), .A2(n16239), .ZN(n12971) );
  NAND4_X1 U16113 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16215) );
  NOR2_X1 U16114 ( .A1(n16208), .A2(n16215), .ZN(n12972) );
  NAND3_X1 U16115 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12971), .A3(
        n12972), .ZN(n12965) );
  INV_X1 U16116 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20241) );
  INV_X1 U16117 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20247) );
  OAI21_X1 U16118 ( .B1(n20241), .B2(n20247), .A(n21112), .ZN(n20223) );
  INV_X1 U16119 ( .A(n20223), .ZN(n12962) );
  NOR2_X1 U16120 ( .A1(n12962), .A2(n15019), .ZN(n16281) );
  NAND4_X1 U16121 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n16238), .A4(n16281), .ZN(
        n12970) );
  NOR2_X1 U16122 ( .A1(n12903), .A2(n12970), .ZN(n16207) );
  AOI21_X1 U16123 ( .B1(n12972), .B2(n16207), .A(n20205), .ZN(n12964) );
  INV_X1 U16124 ( .A(n14277), .ZN(n12967) );
  OAI22_X1 U16125 ( .A1(n20236), .A2(n12963), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n12967), .ZN(n20218) );
  AOI211_X1 U16126 ( .C1(n20219), .C2(n12965), .A(n12964), .B(n20218), .ZN(
        n15996) );
  NOR2_X1 U16127 ( .A1(n16263), .A2(n20218), .ZN(n12966) );
  AOI21_X1 U16128 ( .B1(n15995), .B2(n15996), .A(n12966), .ZN(n16191) );
  OAI21_X1 U16130 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20205), .A(
        n16185), .ZN(n14281) );
  INV_X1 U16131 ( .A(n15999), .ZN(n20240) );
  OAI21_X1 U16132 ( .B1(n20241), .B2(n12967), .A(n20240), .ZN(n20217) );
  OAI221_X1 U16133 ( .B1(n14281), .B2(n20217), .C1(n14281), .C2(n16089), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12976) );
  INV_X1 U16134 ( .A(n12971), .ZN(n12969) );
  NAND2_X1 U16135 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14277), .ZN(
        n12968) );
  OAI22_X1 U16136 ( .A1(n20205), .A2(n12970), .B1(n12969), .B2(n12968), .ZN(
        n15997) );
  AOI21_X1 U16137 ( .B1(n15999), .B2(n12971), .A(n15997), .ZN(n16250) );
  INV_X1 U16138 ( .A(n16195), .ZN(n12973) );
  NOR2_X1 U16139 ( .A1(n16194), .A2(n12973), .ZN(n14284) );
  NAND3_X1 U16140 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14284), .A3(
        n12813), .ZN(n12975) );
  NAND2_X1 U16141 ( .A1(n20236), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n12974) );
  NAND3_X1 U16142 ( .A1(n12976), .A2(n12975), .A3(n12974), .ZN(n12977) );
  NOR2_X1 U16143 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17873), .ZN(
        n12981) );
  NAND2_X1 U16144 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17873), .ZN(
        n12987) );
  OAI22_X1 U16145 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17873), .B1(
        n12987), .B2(n15983), .ZN(n12986) );
  OAI211_X1 U16146 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n15983), .A(
        n12984), .B(n12983), .ZN(n12985) );
  NOR4_X1 U16147 ( .A1(n18961), .A2(n18336), .A3(n18753), .A4(n12988), .ZN(
        n13005) );
  INV_X1 U16148 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18830) );
  NAND2_X1 U16149 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18830), .ZN(n18970) );
  INV_X1 U16150 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18833) );
  NOR2_X1 U16151 ( .A1(n18970), .A2(n18833), .ZN(n18832) );
  NOR2_X1 U16152 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18816) );
  NOR3_X1 U16153 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18832), .A3(n18816), 
        .ZN(n18822) );
  NAND2_X1 U16154 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18962) );
  OAI21_X1 U16155 ( .B1(n18822), .B2(n12989), .A(n18962), .ZN(n16652) );
  NAND2_X1 U16156 ( .A1(n18746), .A2(n12990), .ZN(n13003) );
  NOR3_X1 U16157 ( .A1(n12993), .A2(n12992), .A3(n12991), .ZN(n12994) );
  OAI211_X1 U16158 ( .C1(n18326), .C2(n16014), .A(n12995), .B(n12994), .ZN(
        n12997) );
  AOI21_X1 U16159 ( .B1(n12998), .B2(n12997), .A(n12996), .ZN(n15918) );
  INV_X1 U16160 ( .A(n12999), .ZN(n18749) );
  OAI21_X1 U16161 ( .B1(n13001), .B2(n13000), .A(n18749), .ZN(n13002) );
  OAI211_X1 U16162 ( .C1(n16652), .C2(n13003), .A(n15918), .B(n13002), .ZN(
        n13004) );
  NAND2_X1 U16163 ( .A1(n13025), .A2(n9895), .ZN(n13024) );
  NAND2_X1 U16164 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16517), .ZN(
        n13006) );
  XOR2_X1 U16165 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13006), .Z(
        n13031) );
  INV_X1 U16166 ( .A(n13031), .ZN(n13008) );
  INV_X1 U16167 ( .A(n18781), .ZN(n18268) );
  INV_X1 U16168 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21099) );
  NOR3_X1 U16169 ( .A1(n21099), .A2(n18246), .A3(n10115), .ZN(n18232) );
  NAND2_X1 U16170 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18232), .ZN(
        n18221) );
  OR2_X1 U16171 ( .A1(n18222), .A2(n18221), .ZN(n18202) );
  NOR2_X1 U16172 ( .A1(n18193), .A2(n18202), .ZN(n18072) );
  OAI21_X1 U16173 ( .B1(n18923), .B2(n18938), .A(n18278), .ZN(n18208) );
  NAND2_X1 U16174 ( .A1(n18072), .A2(n18208), .ZN(n18097) );
  NOR2_X1 U16175 ( .A1(n16538), .A2(n18097), .ZN(n13011) );
  INV_X1 U16176 ( .A(n18192), .ZN(n18769) );
  OAI21_X1 U16177 ( .B1(n18769), .B2(n18938), .A(n18763), .ZN(n18269) );
  NAND2_X1 U16178 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18206) );
  NOR2_X1 U16179 ( .A1(n18206), .A2(n18202), .ZN(n18196) );
  NAND2_X1 U16180 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18196), .ZN(
        n18171) );
  NOR2_X1 U16181 ( .A1(n16538), .A2(n18171), .ZN(n18025) );
  AOI22_X1 U16182 ( .A1(n18268), .A2(n13011), .B1(n18269), .B2(n18025), .ZN(
        n16537) );
  NOR2_X1 U16183 ( .A1(n16537), .A2(n17968), .ZN(n17993) );
  NAND2_X1 U16184 ( .A1(n17972), .A2(n17993), .ZN(n15931) );
  NOR4_X1 U16185 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13017), .A3(
        n15983), .A4(n15931), .ZN(n13007) );
  AOI21_X1 U16186 ( .B1(n18204), .B2(n13008), .A(n13007), .ZN(n13021) );
  NAND2_X1 U16187 ( .A1(n13009), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13010) );
  XNOR2_X1 U16188 ( .A(n13010), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13034) );
  NOR2_X2 U16189 ( .A1(n18750), .A2(n18217), .ZN(n18292) );
  NAND2_X1 U16190 ( .A1(n13034), .A2(n18292), .ZN(n13020) );
  INV_X1 U16191 ( .A(n18230), .ZN(n18209) );
  NAND2_X1 U16192 ( .A1(n18288), .A2(n18209), .ZN(n18210) );
  INV_X1 U16193 ( .A(n18210), .ZN(n18283) );
  INV_X1 U16194 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18041) );
  NAND2_X1 U16195 ( .A1(n17972), .A2(n17971), .ZN(n13014) );
  NOR3_X1 U16196 ( .A1(n18041), .A2(n17622), .A3(n13014), .ZN(n16539) );
  INV_X1 U16197 ( .A(n17743), .ZN(n18081) );
  INV_X1 U16198 ( .A(n13011), .ZN(n17969) );
  NOR2_X1 U16199 ( .A1(n18081), .A2(n17969), .ZN(n18075) );
  AOI21_X1 U16200 ( .B1(n13012), .B2(n18075), .A(n18781), .ZN(n18009) );
  AOI211_X1 U16201 ( .C1(n18268), .C2(n13014), .A(n18254), .B(n18009), .ZN(
        n13016) );
  NAND2_X1 U16202 ( .A1(n18018), .A2(n18025), .ZN(n17967) );
  INV_X1 U16203 ( .A(n18171), .ZN(n18098) );
  NAND2_X1 U16204 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18098), .ZN(
        n18191) );
  NOR2_X1 U16205 ( .A1(n16538), .A2(n18191), .ZN(n18100) );
  INV_X1 U16206 ( .A(n13013), .ZN(n18033) );
  NOR2_X1 U16207 ( .A1(n18043), .A2(n18033), .ZN(n16535) );
  AOI21_X1 U16208 ( .B1(n18100), .B2(n16535), .A(n18769), .ZN(n18032) );
  AOI221_X1 U16209 ( .B1(n13014), .B2(n18771), .C1(n17967), .C2(n18771), .A(
        n18032), .ZN(n13015) );
  OAI211_X1 U16210 ( .C1(n18769), .C2(n16539), .A(n13016), .B(n13015), .ZN(
        n15927) );
  AOI22_X1 U16211 ( .A1(n18283), .A2(n13017), .B1(n18289), .B2(n15927), .ZN(
        n15985) );
  OAI21_X1 U16212 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18210), .A(
        n15985), .ZN(n13018) );
  INV_X1 U16213 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18892) );
  NOR2_X1 U16214 ( .A1(n18892), .A2(n18289), .ZN(n13030) );
  AOI21_X1 U16215 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13018), .A(
        n13030), .ZN(n13019) );
  INV_X1 U16216 ( .A(n13022), .ZN(n13023) );
  NAND2_X1 U16217 ( .A1(n13024), .A2(n13023), .ZN(P3_U2831) );
  XOR2_X1 U16218 ( .A(n9910), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(n13027) );
  OAI22_X1 U16219 ( .A1(n13028), .A2(n13027), .B1(n13026), .B2(n9910), .ZN(
        n13029) );
  AOI211_X1 U16220 ( .C1(n17812), .C2(n9921), .A(n13030), .B(n13029), .ZN(
        n13032) );
  NAND2_X1 U16221 ( .A1(n13036), .A2(n13035), .ZN(P3_U2799) );
  INV_X1 U16222 ( .A(n13040), .ZN(n13039) );
  NOR4_X1 U16223 ( .A1(n13037), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16224 ( .A1(n13039), .A2(n13038), .ZN(n13042) );
  NAND3_X1 U16225 ( .A1(n13040), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13041) );
  XNOR2_X1 U16226 ( .A(n13043), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15009) );
  NAND2_X1 U16227 ( .A1(n15009), .A2(n20186), .ZN(n13051) );
  OAI21_X2 U16228 ( .B1(n13044), .B2(n13045), .A(n9844), .ZN(n14790) );
  INV_X1 U16229 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20948) );
  NOR2_X1 U16230 ( .A1(n16230), .A2(n20948), .ZN(n15000) );
  NOR2_X1 U16231 ( .A1(n20190), .A2(n13046), .ZN(n13047) );
  AOI211_X1 U16232 ( .C1(n14490), .C2(n20185), .A(n15000), .B(n13047), .ZN(
        n13048) );
  NAND2_X1 U16233 ( .A1(n13051), .A2(n13050), .ZN(P1_U2971) );
  INV_X1 U16234 ( .A(n13069), .ZN(n13059) );
  NAND2_X1 U16235 ( .A1(n10392), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13052) );
  NAND2_X1 U16236 ( .A1(n13052), .A2(n20000), .ZN(n13072) );
  AOI22_X1 U16237 ( .A1(n13072), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19942), .B2(n19976), .ZN(n13053) );
  NOR2_X1 U16238 ( .A1(n10392), .A2(n16509), .ZN(n13054) );
  NAND2_X1 U16239 ( .A1(n13054), .A2(n9772), .ZN(n13083) );
  OR2_X1 U16240 ( .A1(n13083), .A2(n13055), .ZN(n13060) );
  NAND2_X1 U16241 ( .A1(n13072), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13057) );
  NAND2_X1 U16242 ( .A1(n19968), .A2(n19976), .ZN(n13056) );
  NAND2_X1 U16243 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19661) );
  AND2_X1 U16244 ( .A1(n13056), .A2(n19661), .ZN(n19452) );
  NAND2_X1 U16245 ( .A1(n19452), .A2(n19942), .ZN(n19634) );
  NAND2_X1 U16246 ( .A1(n13057), .A2(n19634), .ZN(n13058) );
  NAND2_X1 U16247 ( .A1(n13558), .A2(n13557), .ZN(n13560) );
  INV_X1 U16248 ( .A(n15775), .ZN(n13544) );
  NAND2_X1 U16249 ( .A1(n13544), .A2(n13060), .ZN(n13061) );
  NAND2_X1 U16250 ( .A1(n19661), .A2(n19958), .ZN(n13062) );
  NOR2_X1 U16251 ( .A1(n19958), .A2(n19968), .ZN(n14089) );
  NAND2_X1 U16252 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14089), .ZN(
        n14090) );
  AND2_X1 U16253 ( .A1(n13062), .A2(n14090), .ZN(n19453) );
  AND2_X1 U16254 ( .A1(n19453), .A2(n19942), .ZN(n19698) );
  AOI21_X1 U16255 ( .B1(n13072), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19698), .ZN(n13063) );
  INV_X1 U16256 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13064) );
  OR2_X1 U16257 ( .A1(n13083), .A2(n13064), .ZN(n13065) );
  NAND2_X1 U16258 ( .A1(n13667), .A2(n13666), .ZN(n13665) );
  INV_X1 U16259 ( .A(n13065), .ZN(n13066) );
  NAND2_X1 U16260 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  NOR2_X1 U16261 ( .A1(n13726), .A2(n13069), .ZN(n13075) );
  NAND2_X1 U16262 ( .A1(n14090), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13071) );
  NAND2_X1 U16263 ( .A1(n14089), .A2(n19950), .ZN(n19544) );
  INV_X1 U16264 ( .A(n19544), .ZN(n13070) );
  NAND2_X1 U16265 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13070), .ZN(
        n19574) );
  NAND2_X1 U16266 ( .A1(n13071), .A2(n19574), .ZN(n19696) );
  AOI22_X1 U16267 ( .A1(n13072), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19942), .B2(n19696), .ZN(n13073) );
  INV_X1 U16268 ( .A(n13073), .ZN(n13074) );
  INV_X1 U16269 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13076) );
  OR2_X1 U16270 ( .A1(n13083), .A2(n13076), .ZN(n13077) );
  NAND2_X1 U16271 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  NAND2_X1 U16272 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10392), .ZN(
        n13080) );
  INV_X1 U16273 ( .A(n13083), .ZN(n13302) );
  INV_X1 U16274 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13084) );
  INV_X1 U16275 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U16276 ( .A1(n13963), .A2(n13962), .ZN(n13961) );
  AOI22_X1 U16277 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16278 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16279 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16280 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13089) );
  NAND4_X1 U16281 ( .A1(n13092), .A2(n13091), .A3(n13090), .A4(n13089), .ZN(
        n13098) );
  AOI22_X1 U16282 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16283 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13175), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16284 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16285 ( .A1(n13173), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13093) );
  NAND4_X1 U16286 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13093), .ZN(
        n13097) );
  OR2_X1 U16287 ( .A1(n13098), .A2(n13097), .ZN(n15151) );
  AOI22_X1 U16288 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U16289 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16290 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16291 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10680), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13099) );
  NAND4_X1 U16292 ( .A1(n13102), .A2(n13101), .A3(n13100), .A4(n13099), .ZN(
        n13108) );
  AOI22_X1 U16293 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16294 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n13175), .ZN(n13105) );
  AOI22_X1 U16295 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U16296 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13173), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13103) );
  NAND4_X1 U16297 ( .A1(n13106), .A2(n13105), .A3(n13104), .A4(n13103), .ZN(
        n13107) );
  NOR2_X1 U16298 ( .A1(n13108), .A2(n13107), .ZN(n15159) );
  AOI22_X1 U16299 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U16300 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16301 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U16302 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10680), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13109) );
  NAND4_X1 U16303 ( .A1(n13112), .A2(n13111), .A3(n13110), .A4(n13109), .ZN(
        n13118) );
  AOI22_X1 U16304 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16305 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n13175), .ZN(n13115) );
  AOI22_X1 U16306 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16307 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13173), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13113) );
  NAND4_X1 U16308 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        n13117) );
  NOR2_X1 U16309 ( .A1(n13118), .A2(n13117), .ZN(n15167) );
  AOI22_X1 U16310 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16311 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16312 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16313 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10680), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13119) );
  NAND4_X1 U16314 ( .A1(n13122), .A2(n13121), .A3(n13120), .A4(n13119), .ZN(
        n13128) );
  AOI22_X1 U16315 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13126) );
  AOI22_X1 U16316 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n13175), .ZN(n13125) );
  AOI22_X1 U16317 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16318 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13173), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13123) );
  NAND4_X1 U16319 ( .A1(n13126), .A2(n13125), .A3(n13124), .A4(n13123), .ZN(
        n13127) );
  NOR2_X1 U16320 ( .A1(n13128), .A2(n13127), .ZN(n15170) );
  OR2_X1 U16321 ( .A1(n15167), .A2(n15170), .ZN(n15157) );
  NOR2_X1 U16322 ( .A1(n15159), .A2(n15157), .ZN(n15149) );
  AND2_X1 U16323 ( .A1(n15151), .A2(n15149), .ZN(n13139) );
  AOI22_X1 U16324 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U16325 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16326 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U16327 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10680), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13129) );
  NAND4_X1 U16328 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13138) );
  AOI22_X1 U16329 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16330 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13175), .ZN(n13135) );
  AOI22_X1 U16331 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U16332 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13173), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13133) );
  NAND4_X1 U16333 ( .A1(n13136), .A2(n13135), .A3(n13134), .A4(n13133), .ZN(
        n13137) );
  OR2_X1 U16334 ( .A1(n13138), .A2(n13137), .ZN(n15182) );
  AND2_X1 U16335 ( .A1(n13139), .A2(n15182), .ZN(n15144) );
  AOI22_X1 U16336 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U16337 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U16338 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U16339 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10680), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13140) );
  NAND4_X1 U16340 ( .A1(n13143), .A2(n13142), .A3(n13141), .A4(n13140), .ZN(
        n13149) );
  AOI22_X1 U16341 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10730), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U16342 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n13175), .ZN(n13146) );
  AOI22_X1 U16343 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U16344 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13173), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13144) );
  NAND4_X1 U16345 ( .A1(n13147), .A2(n13146), .A3(n13145), .A4(n13144), .ZN(
        n13148) );
  NOR2_X1 U16346 ( .A1(n13149), .A2(n13148), .ZN(n15146) );
  INV_X1 U16347 ( .A(n15146), .ZN(n13150) );
  AND2_X1 U16348 ( .A1(n15144), .A2(n13150), .ZN(n13161) );
  AOI22_X1 U16349 ( .A1(n13164), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U16350 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U16351 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13152) );
  AOI22_X1 U16352 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13151) );
  NAND4_X1 U16353 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13160) );
  AOI22_X1 U16354 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13171), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16355 ( .A1(n10725), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13175), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16356 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16357 ( .A1(n13173), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13155) );
  NAND4_X1 U16358 ( .A1(n13158), .A2(n13157), .A3(n13156), .A4(n13155), .ZN(
        n13159) );
  OR2_X1 U16359 ( .A1(n13160), .A2(n13159), .ZN(n15191) );
  NAND2_X1 U16360 ( .A1(n13161), .A2(n15191), .ZN(n13162) );
  NOR2_X1 U16361 ( .A1(n15197), .A2(n13162), .ZN(n13163) );
  AOI22_X1 U16362 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13164), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U16363 ( .A1(n13165), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13169) );
  AOI22_X1 U16364 ( .A1(n13166), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10603), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U16365 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10680), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13167) );
  NAND4_X1 U16366 ( .A1(n13170), .A2(n13169), .A3(n13168), .A4(n13167), .ZN(
        n13181) );
  AOI22_X1 U16367 ( .A1(n13171), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10725), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U16368 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U16369 ( .A1(n13174), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13173), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U16370 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13175), .ZN(n13176) );
  NAND4_X1 U16371 ( .A1(n13179), .A2(n13178), .A3(n13177), .A4(n13176), .ZN(
        n13180) );
  NOR2_X1 U16372 ( .A1(n13181), .A2(n13180), .ZN(n13222) );
  AOI22_X1 U16373 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13191) );
  INV_X1 U16374 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13182) );
  OR2_X1 U16375 ( .A1(n10588), .A2(n13182), .ZN(n13187) );
  NAND2_X1 U16376 ( .A1(n9756), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13186) );
  NAND2_X1 U16377 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13185) );
  NAND2_X1 U16378 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13184) );
  AND4_X1 U16379 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13190) );
  AOI22_X1 U16380 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13189) );
  XNOR2_X1 U16381 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13353) );
  NAND4_X1 U16382 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13353), .ZN(
        n13200) );
  AOI22_X1 U16383 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10589), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16384 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13194) );
  NAND2_X1 U16385 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13193) );
  NAND2_X1 U16386 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13192) );
  AND4_X1 U16387 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13197) );
  INV_X1 U16388 ( .A(n13353), .ZN(n13358) );
  AOI22_X1 U16389 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13196) );
  NAND4_X1 U16390 ( .A1(n13198), .A2(n13197), .A3(n13358), .A4(n13196), .ZN(
        n13199) );
  NAND2_X1 U16391 ( .A1(n13200), .A2(n13199), .ZN(n13227) );
  NOR2_X1 U16392 ( .A1(n10625), .A2(n13227), .ZN(n13201) );
  XOR2_X1 U16393 ( .A(n13222), .B(n13201), .Z(n13228) );
  INV_X1 U16394 ( .A(n13227), .ZN(n13223) );
  NAND2_X1 U16395 ( .A1(n10625), .A2(n13223), .ZN(n15140) );
  INV_X1 U16396 ( .A(n13228), .ZN(n13203) );
  AOI22_X1 U16397 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9767), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13211) );
  OR2_X1 U16398 ( .A1(n10588), .A2(n13204), .ZN(n13208) );
  NAND2_X1 U16399 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13207) );
  NAND2_X1 U16400 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13206) );
  NAND2_X1 U16401 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13205) );
  AND4_X1 U16402 ( .A1(n13208), .A2(n13207), .A3(n13206), .A4(n13205), .ZN(
        n13210) );
  AOI22_X1 U16403 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9762), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13209) );
  NAND4_X1 U16404 ( .A1(n13211), .A2(n13210), .A3(n13209), .A4(n13353), .ZN(
        n13221) );
  AOI22_X1 U16405 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9767), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13219) );
  INV_X1 U16406 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13212) );
  OR2_X1 U16407 ( .A1(n10588), .A2(n13212), .ZN(n13216) );
  NAND2_X1 U16408 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13215) );
  NAND2_X1 U16409 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13214) );
  NAND2_X1 U16410 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13213) );
  AND4_X1 U16411 ( .A1(n13216), .A2(n13215), .A3(n13214), .A4(n13213), .ZN(
        n13218) );
  AOI22_X1 U16412 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13217) );
  NAND4_X1 U16413 ( .A1(n13219), .A2(n13218), .A3(n13358), .A4(n13217), .ZN(
        n13220) );
  NAND2_X1 U16414 ( .A1(n13221), .A2(n13220), .ZN(n13230) );
  INV_X1 U16415 ( .A(n13222), .ZN(n13224) );
  NAND2_X1 U16416 ( .A1(n13224), .A2(n13223), .ZN(n13231) );
  XOR2_X1 U16417 ( .A(n13230), .B(n13231), .Z(n13225) );
  NAND2_X1 U16418 ( .A1(n13225), .A2(n13302), .ZN(n15130) );
  INV_X1 U16419 ( .A(n13230), .ZN(n13226) );
  NAND2_X1 U16420 ( .A1(n10625), .A2(n13226), .ZN(n15132) );
  NOR3_X1 U16421 ( .A1(n13228), .A2(n13227), .A3(n15132), .ZN(n13229) );
  NOR2_X1 U16422 ( .A1(n13231), .A2(n13230), .ZN(n13250) );
  AOI22_X1 U16423 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13239) );
  INV_X1 U16424 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13232) );
  OR2_X1 U16425 ( .A1(n10588), .A2(n13232), .ZN(n13236) );
  NAND2_X1 U16426 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U16427 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13234) );
  NAND2_X1 U16428 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13233) );
  AND4_X1 U16429 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13238) );
  AOI22_X1 U16430 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13237) );
  NAND4_X1 U16431 ( .A1(n13239), .A2(n13238), .A3(n13237), .A4(n13353), .ZN(
        n13249) );
  AOI22_X1 U16432 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13247) );
  INV_X1 U16433 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13240) );
  OR2_X1 U16434 ( .A1(n10588), .A2(n13240), .ZN(n13244) );
  NAND2_X1 U16435 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13243) );
  NAND2_X1 U16436 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13242) );
  NAND2_X1 U16437 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13241) );
  AND4_X1 U16438 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13246) );
  AOI22_X1 U16439 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9762), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13245) );
  NAND4_X1 U16440 ( .A1(n13247), .A2(n13246), .A3(n13358), .A4(n13245), .ZN(
        n13248) );
  AND2_X1 U16441 ( .A1(n13249), .A2(n13248), .ZN(n13251) );
  NAND2_X1 U16442 ( .A1(n13250), .A2(n13251), .ZN(n13299) );
  OAI211_X1 U16443 ( .C1(n13250), .C2(n13251), .A(n13302), .B(n13299), .ZN(
        n13254) );
  INV_X1 U16444 ( .A(n13251), .ZN(n13252) );
  NOR2_X1 U16445 ( .A1(n19990), .A2(n13252), .ZN(n14315) );
  AOI22_X1 U16446 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13264) );
  INV_X1 U16447 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13257) );
  OR2_X1 U16448 ( .A1(n10588), .A2(n13257), .ZN(n13261) );
  NAND2_X1 U16449 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13260) );
  NAND2_X1 U16450 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13259) );
  NAND2_X1 U16451 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13258) );
  AND4_X1 U16452 ( .A1(n13261), .A2(n13260), .A3(n13259), .A4(n13258), .ZN(
        n13263) );
  AOI22_X1 U16453 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13262) );
  NAND4_X1 U16454 ( .A1(n13264), .A2(n13263), .A3(n13262), .A4(n13353), .ZN(
        n13274) );
  AOI22_X1 U16455 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9767), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13272) );
  INV_X1 U16456 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13265) );
  OR2_X1 U16457 ( .A1(n10588), .A2(n13265), .ZN(n13269) );
  NAND2_X1 U16458 ( .A1(n9756), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13268) );
  NAND2_X1 U16459 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13267) );
  NAND2_X1 U16460 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13266) );
  AND4_X1 U16461 ( .A1(n13269), .A2(n13268), .A3(n13267), .A4(n13266), .ZN(
        n13271) );
  AOI22_X1 U16462 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9762), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13270) );
  NAND4_X1 U16463 ( .A1(n13272), .A2(n13271), .A3(n13358), .A4(n13270), .ZN(
        n13273) );
  AND2_X1 U16464 ( .A1(n13274), .A2(n13273), .ZN(n13297) );
  XNOR2_X1 U16465 ( .A(n13299), .B(n13297), .ZN(n13275) );
  NAND2_X1 U16466 ( .A1(n10625), .A2(n13297), .ZN(n15121) );
  INV_X1 U16467 ( .A(n15120), .ZN(n13278) );
  NAND2_X1 U16468 ( .A1(n13276), .A2(n10219), .ZN(n13277) );
  AOI22_X1 U16469 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13286) );
  INV_X1 U16470 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13279) );
  OR2_X1 U16471 ( .A1(n10588), .A2(n13279), .ZN(n13283) );
  NAND2_X1 U16472 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13282) );
  NAND2_X1 U16473 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13281) );
  NAND2_X1 U16474 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13280) );
  AND4_X1 U16475 ( .A1(n13283), .A2(n13282), .A3(n13281), .A4(n13280), .ZN(
        n13285) );
  AOI22_X1 U16476 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13284) );
  NAND4_X1 U16477 ( .A1(n13286), .A2(n13285), .A3(n13284), .A4(n13353), .ZN(
        n13296) );
  AOI22_X1 U16478 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13294) );
  INV_X1 U16479 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13287) );
  OR2_X1 U16480 ( .A1(n10588), .A2(n13287), .ZN(n13291) );
  NAND2_X1 U16481 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13290) );
  NAND2_X1 U16482 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13289) );
  NAND2_X1 U16483 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13288) );
  AND4_X1 U16484 ( .A1(n13291), .A2(n13290), .A3(n13289), .A4(n13288), .ZN(
        n13293) );
  AOI22_X1 U16485 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13292) );
  NAND4_X1 U16486 ( .A1(n13294), .A2(n13293), .A3(n13358), .A4(n13292), .ZN(
        n13295) );
  NAND2_X1 U16487 ( .A1(n13296), .A2(n13295), .ZN(n13300) );
  INV_X1 U16488 ( .A(n13300), .ZN(n13308) );
  INV_X1 U16489 ( .A(n13297), .ZN(n13298) );
  OR2_X1 U16490 ( .A1(n13299), .A2(n13298), .ZN(n13301) );
  INV_X1 U16491 ( .A(n13301), .ZN(n13303) );
  OR2_X1 U16492 ( .A1(n13301), .A2(n13300), .ZN(n15108) );
  OAI211_X1 U16493 ( .C1(n13308), .C2(n13303), .A(n15108), .B(n13302), .ZN(
        n13305) );
  NAND2_X1 U16494 ( .A1(n13306), .A2(n13305), .ZN(n13307) );
  NAND2_X1 U16495 ( .A1(n10625), .A2(n13308), .ZN(n15115) );
  INV_X1 U16496 ( .A(n15109), .ZN(n13327) );
  AOI22_X1 U16497 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13316) );
  INV_X1 U16498 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13309) );
  OR2_X1 U16499 ( .A1(n10588), .A2(n13309), .ZN(n13313) );
  NAND2_X1 U16500 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13312) );
  NAND2_X1 U16501 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13311) );
  NAND2_X1 U16502 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13310) );
  AND4_X1 U16503 ( .A1(n13313), .A2(n13312), .A3(n13311), .A4(n13310), .ZN(
        n13315) );
  AOI22_X1 U16504 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9762), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13314) );
  NAND4_X1 U16505 ( .A1(n13316), .A2(n13315), .A3(n13314), .A4(n13353), .ZN(
        n13326) );
  AOI22_X1 U16506 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9767), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13324) );
  INV_X1 U16507 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13317) );
  OR2_X1 U16508 ( .A1(n10588), .A2(n13317), .ZN(n13321) );
  NAND2_X1 U16509 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13320) );
  NAND2_X1 U16510 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13319) );
  NAND2_X1 U16511 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n13318) );
  AND4_X1 U16512 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n13323) );
  AOI22_X1 U16513 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13322) );
  NAND4_X1 U16514 ( .A1(n13324), .A2(n13323), .A3(n13358), .A4(n13322), .ZN(
        n13325) );
  AND2_X1 U16515 ( .A1(n13326), .A2(n13325), .ZN(n15110) );
  NAND2_X1 U16516 ( .A1(n9772), .A2(n15110), .ZN(n13328) );
  NOR2_X1 U16517 ( .A1(n15108), .A2(n13328), .ZN(n13347) );
  AOI22_X1 U16518 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13356), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13335) );
  INV_X1 U16519 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n21029) );
  OR2_X1 U16520 ( .A1(n10588), .A2(n21029), .ZN(n13332) );
  NAND2_X1 U16521 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13331) );
  NAND2_X1 U16522 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n13330) );
  INV_X1 U16523 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21142) );
  NAND2_X1 U16524 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13329) );
  AND4_X1 U16525 ( .A1(n13332), .A2(n13331), .A3(n13330), .A4(n13329), .ZN(
        n13334) );
  AOI22_X1 U16526 ( .A1(n9756), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13352), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13333) );
  NAND4_X1 U16527 ( .A1(n13335), .A2(n13334), .A3(n13333), .A4(n13353), .ZN(
        n13345) );
  AOI22_X1 U16528 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9767), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13343) );
  INV_X1 U16529 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13336) );
  OR2_X1 U16530 ( .A1(n10588), .A2(n13336), .ZN(n13340) );
  NAND2_X1 U16531 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13339) );
  INV_X1 U16532 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n19770) );
  NAND2_X1 U16533 ( .A1(n13352), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13338) );
  NAND2_X1 U16534 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n13337) );
  AND4_X1 U16535 ( .A1(n13340), .A2(n13339), .A3(n13338), .A4(n13337), .ZN(
        n13342) );
  AOI22_X1 U16536 ( .A1(n10589), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13341) );
  NAND4_X1 U16537 ( .A1(n13343), .A2(n13342), .A3(n13358), .A4(n13341), .ZN(
        n13344) );
  AND2_X1 U16538 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  NAND2_X1 U16539 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  OAI21_X1 U16540 ( .B1(n13347), .B2(n13346), .A(n13348), .ZN(n14410) );
  INV_X1 U16541 ( .A(n13348), .ZN(n13349) );
  AOI22_X1 U16542 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10589), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13351) );
  AOI22_X1 U16543 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9762), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U16544 ( .A1(n13351), .A2(n13350), .ZN(n13365) );
  AOI22_X1 U16545 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13352), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13355) );
  AOI22_X1 U16546 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9757), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13354) );
  NAND3_X1 U16547 ( .A1(n13355), .A2(n13354), .A3(n13353), .ZN(n13364) );
  AOI22_X1 U16548 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13352), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13359) );
  AOI22_X1 U16549 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13357) );
  NAND3_X1 U16550 ( .A1(n13359), .A2(n13358), .A3(n13357), .ZN(n13363) );
  AOI22_X1 U16551 ( .A1(n10587), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10589), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U16552 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U16553 ( .A1(n13361), .A2(n13360), .ZN(n13362) );
  OAI22_X1 U16554 ( .A1(n13365), .A2(n13364), .B1(n13363), .B2(n13362), .ZN(
        n13366) );
  XNOR2_X1 U16555 ( .A(n13367), .B(n13366), .ZN(n14408) );
  NAND2_X1 U16556 ( .A1(n11015), .A2(n20001), .ZN(n14050) );
  NOR2_X1 U16557 ( .A1(n14052), .A2(n14050), .ZN(n13368) );
  AOI21_X1 U16558 ( .B1(n14093), .B2(n14041), .A(n13368), .ZN(n14009) );
  NAND2_X1 U16559 ( .A1(n13370), .A2(n13369), .ZN(n13371) );
  NAND2_X1 U16560 ( .A1(n14009), .A2(n13371), .ZN(n13372) );
  NAND2_X1 U16561 ( .A1(n19249), .A2(n13373), .ZN(n15282) );
  NOR4_X1 U16562 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n13378) );
  NOR4_X1 U16563 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13377) );
  NOR4_X1 U16564 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n13376) );
  NOR4_X1 U16565 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13375) );
  NAND4_X1 U16566 ( .A1(n13378), .A2(n13377), .A3(n13376), .A4(n13375), .ZN(
        n13383) );
  NOR4_X1 U16567 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_0__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13381) );
  NOR4_X1 U16568 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13380) );
  NOR4_X1 U16569 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13379) );
  INV_X1 U16570 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19888) );
  NAND4_X1 U16571 ( .A1(n13381), .A2(n13380), .A3(n13379), .A4(n19888), .ZN(
        n13382) );
  OAI21_X1 U16572 ( .B1(n13383), .B2(n13382), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13574) );
  NOR2_X1 U16573 ( .A1(n10402), .A2(n13574), .ZN(n13384) );
  INV_X1 U16574 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13385) );
  NOR2_X1 U16575 ( .A1(n19249), .A2(n13385), .ZN(n13386) );
  AOI21_X1 U16576 ( .B1(n19223), .B2(BUF1_REG_30__SCAN_IN), .A(n13386), .ZN(
        n13387) );
  INV_X1 U16577 ( .A(n13387), .ZN(n13388) );
  INV_X1 U16578 ( .A(n13574), .ZN(n14106) );
  AND2_X1 U16579 ( .A1(n10904), .A2(n13564), .ZN(n13390) );
  MUX2_X1 U16580 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n14104), .Z(n19230) );
  AOI22_X1 U16581 ( .A1(n19222), .A2(BUF2_REG_30__SCAN_IN), .B1(n19221), .B2(
        n19230), .ZN(n13391) );
  AND2_X1 U16582 ( .A1(n13392), .A2(n13391), .ZN(n13393) );
  OAI21_X1 U16583 ( .B1(n14408), .B2(n15282), .A(n13393), .ZN(P2_U2889) );
  NOR4_X1 U16584 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13397) );
  NOR4_X1 U16585 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13396) );
  NOR4_X1 U16586 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13395) );
  NOR4_X1 U16587 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13394) );
  AND4_X1 U16588 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13402) );
  NOR4_X1 U16589 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13400) );
  NOR4_X1 U16590 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13399) );
  NOR4_X1 U16591 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13398) );
  INV_X1 U16592 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20909) );
  AND4_X1 U16593 ( .A1(n13400), .A2(n13399), .A3(n13398), .A4(n20909), .ZN(
        n13401) );
  NAND2_X1 U16594 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  INV_X1 U16595 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20975) );
  NOR3_X1 U16596 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20975), .ZN(n13405) );
  NOR4_X1 U16597 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13404) );
  NAND4_X1 U16598 ( .A1(n20259), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13405), .A4(
        n13404), .ZN(U214) );
  NOR2_X1 U16599 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13407) );
  NOR4_X1 U16600 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13406) );
  NAND4_X1 U16601 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13407), .A4(n13406), .ZN(n13408) );
  NOR2_X1 U16602 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13408), .ZN(n16638)
         );
  NOR2_X1 U16603 ( .A1(n14104), .A2(n13408), .ZN(n16559) );
  NAND2_X1 U16604 ( .A1(n16559), .A2(U214), .ZN(U212) );
  NOR3_X1 U16605 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16994) );
  INV_X1 U16606 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17320) );
  NAND2_X1 U16607 ( .A1(n16994), .A2(n17320), .ZN(n16978) );
  NOR2_X1 U16608 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16978), .ZN(n16965) );
  INV_X1 U16609 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17312) );
  NAND2_X1 U16610 ( .A1(n16965), .A2(n17312), .ZN(n16956) );
  NOR2_X1 U16611 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16956), .ZN(n16937) );
  INV_X1 U16612 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17306) );
  NAND2_X1 U16613 ( .A1(n16937), .A2(n17306), .ZN(n16928) );
  NOR2_X1 U16614 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16928), .ZN(n16913) );
  INV_X1 U16615 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17263) );
  NAND2_X1 U16616 ( .A1(n16913), .A2(n17263), .ZN(n16900) );
  NOR2_X1 U16617 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16900), .ZN(n16887) );
  INV_X1 U16618 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16883) );
  NAND2_X1 U16619 ( .A1(n16887), .A2(n16883), .ZN(n16882) );
  NOR2_X1 U16620 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16882), .ZN(n16867) );
  INV_X1 U16621 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17215) );
  NAND2_X1 U16622 ( .A1(n16867), .A2(n17215), .ZN(n16854) );
  NOR2_X1 U16623 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16854), .ZN(n16840) );
  INV_X1 U16624 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16834) );
  NAND2_X1 U16625 ( .A1(n16840), .A2(n16834), .ZN(n16833) );
  NOR2_X1 U16626 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16833), .ZN(n16819) );
  INV_X1 U16627 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21210) );
  NAND2_X1 U16628 ( .A1(n16819), .A2(n21210), .ZN(n16809) );
  NOR2_X1 U16629 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16809), .ZN(n16795) );
  INV_X1 U16630 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16788) );
  NAND2_X1 U16631 ( .A1(n16795), .A2(n16788), .ZN(n16786) );
  NOR2_X1 U16632 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16786), .ZN(n16775) );
  INV_X1 U16633 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U16634 ( .A1(n16775), .A2(n16767), .ZN(n16766) );
  NOR2_X1 U16635 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16766), .ZN(n16755) );
  INV_X1 U16636 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16748) );
  NAND2_X1 U16637 ( .A1(n16755), .A2(n16748), .ZN(n16747) );
  NOR2_X1 U16638 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16747), .ZN(n16723) );
  INV_X1 U16639 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17031) );
  NAND2_X1 U16640 ( .A1(n16723), .A2(n17031), .ZN(n13410) );
  NOR2_X1 U16641 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n13410), .ZN(n16719) );
  NAND2_X1 U16642 ( .A1(n18955), .A2(n18746), .ZN(n17530) );
  NAND2_X1 U16643 ( .A1(n18976), .A2(n17492), .ZN(n13423) );
  NAND2_X1 U16644 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n15915), .ZN(n13409) );
  AOI211_X4 U16645 ( .C1(n18960), .C2(n18962), .A(n13423), .B(n13409), .ZN(
        n16977) );
  AOI211_X1 U16646 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n13410), .A(n16719), .B(
        n17022), .ZN(n13427) );
  INV_X1 U16647 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18880) );
  INV_X1 U16648 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18882) );
  OAI211_X1 U16649 ( .C1(n15915), .C2(n18822), .A(n18962), .B(n18960), .ZN(
        n13422) );
  NOR2_X2 U16650 ( .A1(n13422), .A2(n13423), .ZN(n17001) );
  INV_X1 U16651 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18878) );
  INV_X1 U16652 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21048) );
  INV_X1 U16653 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18859) );
  INV_X1 U16654 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18853) );
  INV_X1 U16655 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18845) );
  INV_X1 U16656 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18841) );
  INV_X1 U16657 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18837) );
  NAND2_X1 U16658 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17002) );
  NOR2_X1 U16659 ( .A1(n18837), .A2(n17002), .ZN(n16961) );
  NAND2_X1 U16660 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16961), .ZN(n16949) );
  NOR2_X1 U16661 ( .A1(n18841), .A2(n16949), .ZN(n16925) );
  NAND2_X1 U16662 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16925), .ZN(n16926) );
  NOR2_X1 U16663 ( .A1(n18845), .A2(n16926), .ZN(n16914) );
  NAND2_X1 U16664 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16914), .ZN(n16886) );
  NAND2_X1 U16665 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16888) );
  NOR3_X1 U16666 ( .A1(n18853), .A2(n16886), .A3(n16888), .ZN(n16869) );
  NAND2_X1 U16667 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16869), .ZN(n16852) );
  NOR3_X1 U16668 ( .A1(n21048), .A2(n18859), .A3(n16852), .ZN(n16823) );
  INV_X1 U16669 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18871) );
  INV_X1 U16670 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18865) );
  NAND2_X1 U16671 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16812) );
  NOR2_X1 U16672 ( .A1(n18865), .A2(n16812), .ZN(n16791) );
  NAND3_X1 U16673 ( .A1(n16791), .A2(P3_REIP_REG_19__SCAN_IN), .A3(
        P3_REIP_REG_18__SCAN_IN), .ZN(n16772) );
  NOR2_X1 U16674 ( .A1(n18871), .A2(n16772), .ZN(n16754) );
  INV_X1 U16675 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18874) );
  INV_X1 U16676 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18872) );
  NOR2_X1 U16677 ( .A1(n18874), .A2(n18872), .ZN(n16752) );
  NAND4_X1 U16678 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16823), .A3(n16754), 
        .A4(n16752), .ZN(n16741) );
  NOR2_X1 U16679 ( .A1(n18878), .A2(n16741), .ZN(n13411) );
  NAND2_X1 U16680 ( .A1(n17001), .A2(n13411), .ZN(n16726) );
  NAND3_X1 U16681 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n13411), .ZN(n16675) );
  NAND3_X1 U16682 ( .A1(n18973), .A2(n20997), .A3(n18960), .ZN(n18813) );
  NAND2_X1 U16683 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18973), .ZN(n18806) );
  NOR2_X1 U16684 ( .A1(n18805), .A2(n18806), .ZN(n18801) );
  NOR4_X2 U16685 ( .A1(n9768), .A2(n18976), .A3(n16987), .A4(n18801), .ZN(
        n17012) );
  AOI21_X1 U16686 ( .B1(n17001), .B2(n16675), .A(n17012), .ZN(n16722) );
  AOI221_X1 U16687 ( .B1(n18880), .B2(n18882), .C1(n16726), .C2(n18882), .A(
        n16722), .ZN(n13426) );
  AOI21_X1 U16688 ( .B1(n17628), .B2(n17598), .A(n16670), .ZN(n17630) );
  AOI22_X1 U16689 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13415), .B1(
        n13412), .B2(n17696), .ZN(n17699) );
  INV_X1 U16690 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17726) );
  INV_X1 U16691 ( .A(n17724), .ZN(n17722) );
  NOR2_X1 U16692 ( .A1(n17018), .A2(n17722), .ZN(n17723) );
  INV_X1 U16693 ( .A(n17810), .ZN(n17799) );
  NOR2_X1 U16694 ( .A1(n17018), .A2(n17799), .ZN(n17801) );
  NAND3_X1 U16695 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A3(n17801), .ZN(n16850) );
  NOR2_X1 U16696 ( .A1(n17787), .A2(n16850), .ZN(n17764) );
  NAND2_X1 U16697 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17764), .ZN(
        n16828) );
  NOR2_X1 U16698 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16828), .ZN(
        n16818) );
  NAND2_X1 U16699 ( .A1(n17723), .A2(n16818), .ZN(n16798) );
  NOR2_X1 U16700 ( .A1(n17726), .A2(n16798), .ZN(n16783) );
  AND2_X1 U16701 ( .A1(n16783), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13413) );
  INV_X1 U16702 ( .A(n13414), .ZN(n17679) );
  AOI21_X1 U16703 ( .B1(n17710), .B2(n17679), .A(n13415), .ZN(n17713) );
  NOR2_X1 U16704 ( .A1(n16774), .A2(n9920), .ZN(n16763) );
  NAND2_X1 U16706 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13415), .ZN(
        n13416) );
  AOI21_X1 U16707 ( .B1(n17694), .B2(n13416), .A(n17638), .ZN(n17685) );
  OAI21_X1 U16708 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17638), .A(
        n13419), .ZN(n13417) );
  INV_X1 U16709 ( .A(n13417), .ZN(n17669) );
  AOI21_X1 U16710 ( .B1(n17653), .B2(n13419), .A(n13420), .ZN(n17660) );
  OAI21_X1 U16711 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13420), .A(
        n17598), .ZN(n17642) );
  INV_X1 U16712 ( .A(n17642), .ZN(n16725) );
  INV_X1 U16713 ( .A(n16987), .ZN(n18811) );
  AOI211_X1 U16714 ( .C1(n17630), .C2(n13421), .A(n16672), .B(n18811), .ZN(
        n13425) );
  INV_X1 U16715 ( .A(n13422), .ZN(n18797) );
  AOI211_X4 U16716 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n15915), .A(n18797), .B(
        n13423), .ZN(n17006) );
  INV_X1 U16717 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17032) );
  OAI22_X1 U16718 ( .A1(n17628), .A2(n17013), .B1(n17023), .B2(n17032), .ZN(
        n13424) );
  OR4_X1 U16719 ( .A1(n13427), .A2(n13426), .A3(n13425), .A4(n13424), .ZN(
        P3_U2645) );
  AOI211_X1 U16720 ( .C1(n15309), .C2(n13429), .A(n13428), .B(n19216), .ZN(
        n13442) );
  OAI22_X1 U16721 ( .A1(n15307), .A2(n19178), .B1(n19919), .B2(n19204), .ZN(
        n13441) );
  INV_X1 U16722 ( .A(n13430), .ZN(n13432) );
  INV_X1 U16723 ( .A(n19207), .ZN(n19188) );
  INV_X1 U16724 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13431) );
  OAI22_X1 U16725 ( .A1(n13432), .A2(n19201), .B1(n19188), .B2(n13431), .ZN(
        n13440) );
  NAND2_X1 U16726 ( .A1(n13433), .A2(n13434), .ZN(n13435) );
  NAND2_X1 U16727 ( .A1(n9841), .A2(n13435), .ZN(n15491) );
  OR2_X1 U16728 ( .A1(n15231), .A2(n13437), .ZN(n13438) );
  NAND2_X1 U16729 ( .A1(n13436), .A2(n13438), .ZN(n15494) );
  OAI22_X1 U16730 ( .A1(n15491), .A2(n19209), .B1(n15494), .B2(n19203), .ZN(
        n13439) );
  OR4_X1 U16731 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        P2_U2828) );
  AOI211_X1 U16732 ( .C1(n16415), .C2(n13443), .A(n19102), .B(n9883), .ZN(
        n13459) );
  OAI21_X1 U16733 ( .B1(n13446), .B2(n13444), .A(n13445), .ZN(n15677) );
  AOI22_X1 U16734 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19167), .ZN(n13447) );
  OAI211_X1 U16735 ( .C1(n15677), .C2(n19203), .A(n13447), .B(n19151), .ZN(
        n13458) );
  INV_X1 U16736 ( .A(n13448), .ZN(n13449) );
  OAI22_X1 U16737 ( .A1(n13449), .A2(n19201), .B1(n10918), .B2(n19188), .ZN(
        n13457) );
  INV_X1 U16738 ( .A(n13450), .ZN(n13452) );
  NAND2_X1 U16739 ( .A1(n13452), .A2(n13451), .ZN(n13453) );
  AND2_X1 U16740 ( .A1(n13453), .A2(n14245), .ZN(n16419) );
  INV_X1 U16741 ( .A(n16419), .ZN(n13455) );
  INV_X1 U16742 ( .A(n16415), .ZN(n13454) );
  NAND2_X1 U16743 ( .A1(n19192), .A2(n19174), .ZN(n19091) );
  OAI22_X1 U16744 ( .A1(n13455), .A2(n19209), .B1(n13454), .B2(n19091), .ZN(
        n13456) );
  OR4_X1 U16745 ( .A1(n13459), .A2(n13458), .A3(n13457), .A4(n13456), .ZN(
        P2_U2844) );
  NOR2_X1 U16746 ( .A1(n13646), .A2(n20012), .ZN(n13460) );
  NAND2_X1 U16747 ( .A1(n15940), .A2(n13460), .ZN(n13463) );
  NOR2_X1 U16748 ( .A1(n12940), .A2(n20012), .ZN(n13461) );
  OR2_X1 U16749 ( .A1(n14437), .A2(n20272), .ZN(n13462) );
  NAND2_X1 U16750 ( .A1(n13463), .A2(n13462), .ZN(n13464) );
  NOR2_X1 U16751 ( .A1(n20888), .A2(n20884), .ZN(n16324) );
  INV_X1 U16752 ( .A(n16324), .ZN(n16326) );
  OR2_X1 U16753 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16326), .ZN(n20117) );
  INV_X2 U16754 ( .A(n20117), .ZN(n20979) );
  AND2_X1 U16755 ( .A1(n20132), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U16756 ( .A(n10983), .ZN(n14054) );
  NAND2_X1 U16757 ( .A1(n14054), .A2(n16503), .ZN(n13465) );
  NOR2_X1 U16758 ( .A1(n14043), .A2(n13465), .ZN(n19211) );
  INV_X1 U16759 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n21020) );
  INV_X1 U16760 ( .A(n14372), .ZN(n13466) );
  OAI211_X1 U16761 ( .C1(n19211), .C2(n21020), .A(n13483), .B(n13466), .ZN(
        P2_U2814) );
  NAND2_X1 U16762 ( .A1(n12832), .A2(n13472), .ZN(n13479) );
  AOI22_X1 U16763 ( .A1(n13479), .A2(n12940), .B1(n13646), .B2(n14650), .ZN(
        n20011) );
  INV_X1 U16764 ( .A(n9818), .ZN(n14307) );
  NAND2_X1 U16765 ( .A1(n14307), .A2(n15993), .ZN(n13644) );
  OAI21_X1 U16766 ( .B1(n13644), .B2(n13480), .A(n20978), .ZN(n20980) );
  AND2_X1 U16767 ( .A1(n20011), .A2(n20980), .ZN(n15952) );
  NOR2_X1 U16768 ( .A1(n15952), .A2(n20012), .ZN(n20019) );
  INV_X1 U16769 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21078) );
  AND3_X1 U16770 ( .A1(n13469), .A2(n13468), .A3(n20261), .ZN(n13470) );
  OAI21_X1 U16771 ( .B1(n13471), .B2(n13470), .A(n13646), .ZN(n13475) );
  INV_X1 U16772 ( .A(n13472), .ZN(n13473) );
  NAND2_X1 U16773 ( .A1(n12832), .A2(n13473), .ZN(n13474) );
  OAI211_X1 U16774 ( .C1(n13637), .C2(n13646), .A(n13475), .B(n13474), .ZN(
        n13476) );
  NAND2_X1 U16775 ( .A1(n13476), .A2(n11827), .ZN(n15954) );
  INV_X1 U16776 ( .A(n15954), .ZN(n13477) );
  NAND2_X1 U16777 ( .A1(n20019), .A2(n13477), .ZN(n13478) );
  OAI21_X1 U16778 ( .B1(n20019), .B2(n21078), .A(n13478), .ZN(P1_U3484) );
  NOR2_X1 U16779 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20822), .ZN(n14436) );
  OR2_X1 U16780 ( .A1(n13479), .A2(n20012), .ZN(n14435) );
  OAI21_X1 U16781 ( .B1(n14436), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14196), 
        .ZN(n13482) );
  OAI21_X1 U16782 ( .B1(n13480), .B2(n9817), .A(n20976), .ZN(n13481) );
  NAND2_X1 U16783 ( .A1(n13482), .A2(n13481), .ZN(P1_U3487) );
  INV_X1 U16784 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13486) );
  INV_X1 U16785 ( .A(n13589), .ZN(n13530) );
  AOI22_X1 U16786 ( .A1(n14106), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14104), .ZN(n19370) );
  NOR2_X1 U16787 ( .A1(n13530), .A2(n19370), .ZN(n13500) );
  AOI21_X1 U16788 ( .B1(n13523), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13500), .ZN(
        n13485) );
  OAI21_X1 U16789 ( .B1(n13484), .B2(n13486), .A(n13485), .ZN(P2_U2974) );
  INV_X1 U16790 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U16791 ( .A1(n14106), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13574), .ZN(n19345) );
  NOR2_X1 U16792 ( .A1(n13530), .A2(n19345), .ZN(n13497) );
  AOI21_X1 U16793 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n13523), .A(n13497), .ZN(
        n13487) );
  OAI21_X1 U16794 ( .B1(n13484), .B2(n13488), .A(n13487), .ZN(P2_U2968) );
  INV_X1 U16795 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13490) );
  AOI22_X1 U16796 ( .A1(n14106), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14104), .ZN(n19348) );
  NOR2_X1 U16797 ( .A1(n13530), .A2(n19348), .ZN(n13509) );
  AOI21_X1 U16798 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n13523), .A(n13509), .ZN(
        n13489) );
  OAI21_X1 U16799 ( .B1(n13484), .B2(n13490), .A(n13489), .ZN(P2_U2969) );
  INV_X1 U16800 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13492) );
  OAI22_X1 U16801 ( .A1(n13574), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14106), .ZN(n19362) );
  NOR2_X1 U16802 ( .A1(n13530), .A2(n19362), .ZN(n13506) );
  AOI21_X1 U16803 ( .B1(n13523), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13506), .ZN(
        n13491) );
  OAI21_X1 U16804 ( .B1(n13484), .B2(n13492), .A(n13491), .ZN(P2_U2958) );
  INV_X1 U16805 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13494) );
  AOI22_X1 U16806 ( .A1(n14106), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13574), .ZN(n19352) );
  NOR2_X1 U16807 ( .A1(n13530), .A2(n19352), .ZN(n13503) );
  AOI21_X1 U16808 ( .B1(n13523), .B2(P2_EAX_REG_3__SCAN_IN), .A(n13503), .ZN(
        n13493) );
  OAI21_X1 U16809 ( .B1(n13484), .B2(n13494), .A(n13493), .ZN(P2_U2970) );
  INV_X1 U16810 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13496) );
  AOI22_X1 U16811 ( .A1(n14106), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14104), .ZN(n19359) );
  NOR2_X1 U16812 ( .A1(n13530), .A2(n19359), .ZN(n13512) );
  AOI21_X1 U16813 ( .B1(n13523), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13512), .ZN(
        n13495) );
  OAI21_X1 U16814 ( .B1(n13484), .B2(n13496), .A(n13495), .ZN(P2_U2957) );
  INV_X1 U16815 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13499) );
  AOI21_X1 U16816 ( .B1(n13523), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13497), .ZN(
        n13498) );
  OAI21_X1 U16817 ( .B1(n13484), .B2(n13499), .A(n13498), .ZN(P2_U2953) );
  INV_X1 U16818 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13502) );
  AOI21_X1 U16819 ( .B1(n13523), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13500), .ZN(
        n13501) );
  OAI21_X1 U16820 ( .B1(n13484), .B2(n13502), .A(n13501), .ZN(P2_U2959) );
  INV_X1 U16821 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13505) );
  AOI21_X1 U16822 ( .B1(n13523), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13503), .ZN(
        n13504) );
  OAI21_X1 U16823 ( .B1(n13484), .B2(n13505), .A(n13504), .ZN(P2_U2955) );
  INV_X1 U16824 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13508) );
  AOI21_X1 U16825 ( .B1(n13523), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13506), .ZN(
        n13507) );
  OAI21_X1 U16826 ( .B1(n13484), .B2(n13508), .A(n13507), .ZN(P2_U2973) );
  INV_X1 U16827 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13511) );
  AOI21_X1 U16828 ( .B1(n13523), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13509), .ZN(
        n13510) );
  OAI21_X1 U16829 ( .B1(n13484), .B2(n13511), .A(n13510), .ZN(P2_U2954) );
  INV_X1 U16830 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13514) );
  AOI21_X1 U16831 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n13523), .A(n13512), .ZN(
        n13513) );
  OAI21_X1 U16832 ( .B1(n13484), .B2(n13514), .A(n13513), .ZN(P2_U2972) );
  INV_X1 U16833 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n13519) );
  INV_X1 U16834 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13700) );
  OR2_X1 U16835 ( .A1(n13574), .A2(n13700), .ZN(n13516) );
  NAND2_X1 U16836 ( .A1(n13574), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13515) );
  AND2_X1 U16837 ( .A1(n13516), .A2(n13515), .ZN(n15225) );
  INV_X1 U16838 ( .A(n15225), .ZN(n13517) );
  NAND2_X1 U16839 ( .A1(n13589), .A2(n13517), .ZN(n13580) );
  NAND2_X1 U16840 ( .A1(n13523), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n13518) );
  OAI211_X1 U16841 ( .C1(n13484), .C2(n13519), .A(n13580), .B(n13518), .ZN(
        P2_U2978) );
  INV_X1 U16842 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13525) );
  INV_X1 U16843 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13520) );
  OR2_X1 U16844 ( .A1(n14104), .A2(n13520), .ZN(n13522) );
  NAND2_X1 U16845 ( .A1(n14104), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13521) );
  NAND2_X1 U16846 ( .A1(n13522), .A2(n13521), .ZN(n14412) );
  NAND2_X1 U16847 ( .A1(n13589), .A2(n14412), .ZN(n13572) );
  NAND2_X1 U16848 ( .A1(n13523), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13524) );
  OAI211_X1 U16849 ( .C1(n13484), .C2(n13525), .A(n13572), .B(n13524), .ZN(
        P2_U2980) );
  INV_X1 U16850 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U16851 ( .A1(n14106), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14104), .ZN(n14147) );
  INV_X1 U16852 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13526) );
  OAI222_X1 U16853 ( .A1(n13484), .A2(n13527), .B1(n13530), .B2(n14147), .C1(
        n13526), .C2(n13597), .ZN(P2_U2982) );
  INV_X1 U16854 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13528) );
  INV_X1 U16855 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13759) );
  INV_X1 U16856 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16609) );
  INV_X1 U16857 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18304) );
  AOI22_X1 U16858 ( .A1(n14106), .A2(n16609), .B1(n18304), .B2(n13574), .ZN(
        n19220) );
  INV_X1 U16859 ( .A(n19220), .ZN(n14101) );
  OAI222_X1 U16860 ( .A1(n13528), .A2(n13484), .B1(n13597), .B2(n13759), .C1(
        n13530), .C2(n14101), .ZN(P2_U2952) );
  INV_X1 U16861 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13531) );
  INV_X1 U16862 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13529) );
  OAI222_X1 U16863 ( .A1(n13531), .A2(n13484), .B1(n13530), .B2(n14101), .C1(
        n13529), .C2(n13597), .ZN(P2_U2967) );
  OAI21_X1 U16864 ( .B1(n15089), .B2(n13673), .A(n13532), .ZN(n13533) );
  XNOR2_X1 U16865 ( .A(n13533), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15767) );
  AOI22_X1 U16866 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19296), .B1(
        n19283), .B2(n15767), .ZN(n13536) );
  INV_X1 U16867 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14261) );
  XNOR2_X1 U16868 ( .A(n13534), .B(n14261), .ZN(n15763) );
  AND2_X1 U16869 ( .A1(n15730), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15765) );
  AOI21_X1 U16870 ( .B1(n19300), .B2(n15763), .A(n15765), .ZN(n13535) );
  OAI211_X1 U16871 ( .C1(n19294), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13536), .B(n13535), .ZN(n13537) );
  AOI21_X1 U16872 ( .B1(n19302), .B2(n15764), .A(n13537), .ZN(n13538) );
  INV_X1 U16873 ( .A(n13538), .ZN(P2_U3013) );
  AND2_X1 U16874 ( .A1(n13539), .A2(n13564), .ZN(n13540) );
  NAND2_X1 U16875 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13542) );
  NAND4_X1 U16876 ( .A1(n13541), .A2(n13542), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20000), .ZN(n13543) );
  INV_X1 U16877 ( .A(n10650), .ZN(n13550) );
  INV_X1 U16878 ( .A(n13545), .ZN(n13548) );
  INV_X1 U16879 ( .A(n13546), .ZN(n13547) );
  NAND2_X1 U16880 ( .A1(n13548), .A2(n13547), .ZN(n13549) );
  NAND2_X1 U16881 ( .A1(n13550), .A2(n13549), .ZN(n19202) );
  INV_X1 U16882 ( .A(n19202), .ZN(n13552) );
  NOR2_X1 U16883 ( .A1(n19971), .A2(n19202), .ZN(n13718) );
  INV_X1 U16884 ( .A(n13718), .ZN(n13551) );
  INV_X1 U16885 ( .A(n15282), .ZN(n19225) );
  OAI211_X1 U16886 ( .C1(n19212), .C2(n13552), .A(n13551), .B(n19225), .ZN(
        n13554) );
  AOI22_X1 U16887 ( .A1(n13389), .A2(n13552), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19239), .ZN(n13553) );
  OAI211_X1 U16888 ( .C1(n14148), .C2(n14101), .A(n13554), .B(n13553), .ZN(
        P2_U2919) );
  XNOR2_X1 U16889 ( .A(n13555), .B(n13556), .ZN(n19163) );
  INV_X1 U16890 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19269) );
  OAI222_X1 U16891 ( .A1(n14148), .A2(n19362), .B1(n19163), .B2(n19243), .C1(
        n19269), .C2(n19249), .ZN(P2_U2913) );
  OR2_X1 U16892 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  INV_X1 U16893 ( .A(n14093), .ZN(n13562) );
  INV_X1 U16894 ( .A(n13561), .ZN(n14044) );
  NAND2_X1 U16895 ( .A1(n13562), .A2(n14044), .ZN(n14008) );
  INV_X1 U16896 ( .A(n11022), .ZN(n13996) );
  NAND2_X1 U16897 ( .A1(n14008), .A2(n13996), .ZN(n13563) );
  NAND2_X1 U16898 ( .A1(n15205), .A2(n13564), .ZN(n15178) );
  INV_X1 U16899 ( .A(n15764), .ZN(n15092) );
  MUX2_X1 U16900 ( .A(n15092), .B(n15094), .S(n9750), .Z(n13565) );
  OAI21_X1 U16901 ( .B1(n19961), .B2(n15178), .A(n13565), .ZN(P2_U2886) );
  INV_X1 U16902 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19265) );
  NAND2_X1 U16903 ( .A1(n13591), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13566) );
  MUX2_X1 U16904 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n14104), .Z(n19244) );
  NAND2_X1 U16905 ( .A1(n13589), .A2(n19244), .ZN(n13582) );
  OAI211_X1 U16906 ( .C1(n19265), .C2(n13597), .A(n13566), .B(n13582), .ZN(
        P2_U2975) );
  INV_X1 U16907 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19263) );
  NAND2_X1 U16908 ( .A1(n13591), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13568) );
  INV_X1 U16909 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16592) );
  NOR2_X1 U16910 ( .A1(n13574), .A2(n16592), .ZN(n13567) );
  AOI21_X1 U16911 ( .B1(n14104), .B2(BUF2_REG_9__SCAN_IN), .A(n13567), .ZN(
        n14321) );
  INV_X1 U16912 ( .A(n14321), .ZN(n19240) );
  NAND2_X1 U16913 ( .A1(n13589), .A2(n19240), .ZN(n13570) );
  OAI211_X1 U16914 ( .C1(n19263), .C2(n13597), .A(n13568), .B(n13570), .ZN(
        P2_U2976) );
  INV_X1 U16915 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19261) );
  NAND2_X1 U16916 ( .A1(n13591), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13569) );
  MUX2_X1 U16917 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n14104), .Z(n19236) );
  NAND2_X1 U16918 ( .A1(n13589), .A2(n19236), .ZN(n13584) );
  OAI211_X1 U16919 ( .C1(n19261), .C2(n13597), .A(n13569), .B(n13584), .ZN(
        P2_U2977) );
  INV_X1 U16920 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14319) );
  NAND2_X1 U16921 ( .A1(n13591), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13571) );
  OAI211_X1 U16922 ( .C1(n13597), .C2(n14319), .A(n13571), .B(n13570), .ZN(
        P2_U2961) );
  INV_X1 U16923 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n21179) );
  NAND2_X1 U16924 ( .A1(n13591), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13573) );
  OAI211_X1 U16925 ( .C1(n13597), .C2(n21179), .A(n13573), .B(n13572), .ZN(
        P2_U2965) );
  INV_X1 U16926 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n13576) );
  NAND2_X1 U16927 ( .A1(n13591), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n13575) );
  OAI22_X1 U16928 ( .A1(n13574), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14106), .ZN(n19356) );
  INV_X1 U16929 ( .A(n19356), .ZN(n16397) );
  NAND2_X1 U16930 ( .A1(n13589), .A2(n16397), .ZN(n13586) );
  OAI211_X1 U16931 ( .C1(n13597), .C2(n13576), .A(n13575), .B(n13586), .ZN(
        P2_U2971) );
  INV_X1 U16932 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19257) );
  NAND2_X1 U16933 ( .A1(n13591), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13577) );
  MUX2_X1 U16934 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n14104), .Z(n19233) );
  NAND2_X1 U16935 ( .A1(n13589), .A2(n19233), .ZN(n13578) );
  OAI211_X1 U16936 ( .C1(n19257), .C2(n13597), .A(n13577), .B(n13578), .ZN(
        P2_U2979) );
  INV_X1 U16937 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13604) );
  NAND2_X1 U16938 ( .A1(n13591), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13579) );
  OAI211_X1 U16939 ( .C1(n13604), .C2(n13597), .A(n13579), .B(n13578), .ZN(
        P2_U2964) );
  INV_X1 U16940 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15223) );
  NAND2_X1 U16941 ( .A1(n13591), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13581) );
  OAI211_X1 U16942 ( .C1(n13597), .C2(n15223), .A(n13581), .B(n13580), .ZN(
        P2_U2963) );
  INV_X1 U16943 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U16944 ( .A1(n13591), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13583) );
  OAI211_X1 U16945 ( .C1(n13608), .C2(n13597), .A(n13583), .B(n13582), .ZN(
        P2_U2960) );
  INV_X1 U16946 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13602) );
  NAND2_X1 U16947 ( .A1(n13591), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13585) );
  OAI211_X1 U16948 ( .C1(n13602), .C2(n13597), .A(n13585), .B(n13584), .ZN(
        P2_U2962) );
  INV_X1 U16949 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U16950 ( .A1(n13591), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13587) );
  OAI211_X1 U16951 ( .C1(n13597), .C2(n13588), .A(n13587), .B(n13586), .ZN(
        P2_U2956) );
  INV_X1 U16952 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19253) );
  NAND2_X1 U16953 ( .A1(n13591), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U16954 ( .A1(n13589), .A2(n19230), .ZN(n13592) );
  OAI211_X1 U16955 ( .C1(n19253), .C2(n13597), .A(n13590), .B(n13592), .ZN(
        P2_U2981) );
  NAND2_X1 U16956 ( .A1(n13591), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13593) );
  OAI211_X1 U16957 ( .C1(n13385), .C2(n13597), .A(n13593), .B(n13592), .ZN(
        P2_U2966) );
  NOR2_X1 U16958 ( .A1(n9750), .A2(n10072), .ZN(n13594) );
  AOI21_X1 U16959 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n9769), .A(n13594), .ZN(
        n13595) );
  OAI21_X1 U16960 ( .B1(n15178), .B2(n19971), .A(n13595), .ZN(P2_U2887) );
  NOR2_X1 U16961 ( .A1(n13596), .A2(n10983), .ZN(n14006) );
  NAND2_X1 U16962 ( .A1(n14006), .A2(n16503), .ZN(n13598) );
  NAND2_X1 U16963 ( .A1(n13598), .A2(n13597), .ZN(n13599) );
  INV_X1 U16964 ( .A(n19875), .ZN(n19989) );
  NAND2_X1 U16965 ( .A1(n19250), .A2(n13600), .ZN(n13768) );
  NAND2_X1 U16966 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14094) );
  NOR2_X1 U16967 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14094), .ZN(n19280) );
  AOI22_X1 U16968 ( .A1(n20002), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13601) );
  OAI21_X1 U16969 ( .B1(n13602), .B2(n13768), .A(n13601), .ZN(P2_U2925) );
  AOI22_X1 U16970 ( .A1(n20002), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13603) );
  OAI21_X1 U16971 ( .B1(n13604), .B2(n13768), .A(n13603), .ZN(P2_U2923) );
  AOI22_X1 U16972 ( .A1(n20002), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13605) );
  OAI21_X1 U16973 ( .B1(n13385), .B2(n13768), .A(n13605), .ZN(P2_U2921) );
  AOI22_X1 U16974 ( .A1(n20002), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13606) );
  OAI21_X1 U16975 ( .B1(n15223), .B2(n13768), .A(n13606), .ZN(P2_U2924) );
  AOI22_X1 U16976 ( .A1(n20002), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13607) );
  OAI21_X1 U16977 ( .B1(n13608), .B2(n13768), .A(n13607), .ZN(P2_U2927) );
  AOI22_X1 U16978 ( .A1(n20002), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13609) );
  OAI21_X1 U16979 ( .B1(n14319), .B2(n13768), .A(n13609), .ZN(P2_U2926) );
  AOI22_X1 U16980 ( .A1(n20002), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13610) );
  OAI21_X1 U16981 ( .B1(n21179), .B2(n13768), .A(n13610), .ZN(P2_U2922) );
  INV_X1 U16982 ( .A(n12824), .ZN(n13613) );
  NAND3_X1 U16983 ( .A1(n13613), .A2(n13612), .A3(n13611), .ZN(n13614) );
  NOR2_X1 U16984 ( .A1(n13615), .A2(n13614), .ZN(n13618) );
  AND2_X1 U16985 ( .A1(n13618), .A2(n13617), .ZN(n15031) );
  INV_X1 U16986 ( .A(n15031), .ZN(n13619) );
  NAND2_X1 U16987 ( .A1(n20549), .A2(n13619), .ZN(n13635) );
  INV_X1 U16988 ( .A(n13639), .ZN(n13620) );
  NAND2_X1 U16989 ( .A1(n13637), .A2(n13620), .ZN(n13659) );
  INV_X1 U16990 ( .A(n13621), .ZN(n15037) );
  OAI21_X1 U16991 ( .B1(n13621), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12011), .ZN(n13622) );
  NAND2_X1 U16992 ( .A1(n13623), .A2(n13622), .ZN(n13624) );
  NAND2_X1 U16993 ( .A1(n13659), .A2(n13624), .ZN(n13633) );
  NOR2_X1 U16994 ( .A1(n13621), .A2(n12011), .ZN(n13625) );
  NAND2_X1 U16995 ( .A1(n13627), .A2(n13626), .ZN(n13636) );
  NAND3_X1 U16996 ( .A1(n15031), .A2(n13732), .A3(n13636), .ZN(n13632) );
  OR2_X1 U16997 ( .A1(n11694), .A2(n9784), .ZN(n13630) );
  NAND2_X1 U16998 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13628) );
  NAND2_X1 U16999 ( .A1(n12011), .A2(n13628), .ZN(n13629) );
  NAND3_X1 U17000 ( .A1(n15940), .A2(n13630), .A3(n13629), .ZN(n13631) );
  AND3_X1 U17001 ( .A1(n13633), .A2(n13632), .A3(n13631), .ZN(n13634) );
  NAND2_X1 U17002 ( .A1(n13635), .A2(n13634), .ZN(n13815) );
  AOI22_X1 U17003 ( .A1(n13815), .A2(n13683), .B1(n15038), .B2(n13636), .ZN(
        n13652) );
  OR2_X1 U17004 ( .A1(n13617), .A2(n13638), .ZN(n13641) );
  NAND2_X1 U17005 ( .A1(n13639), .A2(n14128), .ZN(n13640) );
  NAND2_X1 U17006 ( .A1(n14197), .A2(n20272), .ZN(n14657) );
  NOR2_X1 U17007 ( .A1(n14657), .A2(n20278), .ZN(n13642) );
  NOR2_X1 U17008 ( .A1(n13643), .A2(n13642), .ZN(n13649) );
  NAND2_X1 U17009 ( .A1(n13644), .A2(n20978), .ZN(n13645) );
  NOR2_X1 U17010 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  OAI21_X1 U17011 ( .B1(n15940), .B2(n12824), .A(n13647), .ZN(n13648) );
  NAND4_X1 U17012 ( .A1(n13735), .A2(n14131), .A3(n13649), .A4(n13648), .ZN(
        n13821) );
  NOR2_X1 U17013 ( .A1(n20885), .A2(n16326), .ZN(n13826) );
  AND2_X1 U17014 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13826), .ZN(n13650) );
  AOI21_X1 U17015 ( .B1(n13821), .B2(n14132), .A(n13650), .ZN(n16313) );
  NAND2_X1 U17016 ( .A1(n20885), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13651) );
  NAND2_X1 U17017 ( .A1(n16313), .A2(n13651), .ZN(n16316) );
  MUX2_X1 U17018 ( .A(n12011), .B(n13652), .S(n16316), .Z(n13653) );
  INV_X1 U17019 ( .A(n13653), .ZN(P1_U3469) );
  XNOR2_X1 U17020 ( .A(n13621), .B(n13655), .ZN(n13662) );
  AND2_X1 U17021 ( .A1(n13732), .A2(n13662), .ZN(n13657) );
  XNOR2_X1 U17022 ( .A(n10119), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13656) );
  AOI22_X1 U17023 ( .A1(n15031), .A2(n13657), .B1(n15940), .B2(n13656), .ZN(
        n13661) );
  INV_X1 U17024 ( .A(n13662), .ZN(n13658) );
  NAND2_X1 U17025 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  OAI211_X1 U17026 ( .C1(n20690), .C2(n15031), .A(n13661), .B(n13660), .ZN(
        n13816) );
  NOR2_X1 U17027 ( .A1(n20884), .A2(n20241), .ZN(n15036) );
  AOI22_X1 U17028 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20247), .B2(n12794), .ZN(
        n15034) );
  AOI222_X1 U17029 ( .A1(n13816), .A2(n13683), .B1(n15036), .B2(n15034), .C1(
        n13662), .C2(n15038), .ZN(n13664) );
  INV_X1 U17030 ( .A(n16316), .ZN(n13686) );
  NAND2_X1 U17031 ( .A1(n13686), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13663) );
  OAI21_X1 U17032 ( .B1(n13664), .B2(n13686), .A(n13663), .ZN(P1_U3472) );
  MUX2_X1 U17033 ( .A(n13670), .B(n10411), .S(n9769), .Z(n13671) );
  OAI21_X1 U17034 ( .B1(n19953), .B2(n15178), .A(n13671), .ZN(P2_U2885) );
  MUX2_X1 U17035 ( .A(n15616), .B(n13672), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13681) );
  OAI21_X1 U17036 ( .B1(n19199), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13673), .ZN(n19306) );
  INV_X1 U17037 ( .A(n19317), .ZN(n16486) );
  NAND2_X1 U17038 ( .A1(n16486), .A2(n19301), .ZN(n13674) );
  NAND2_X1 U17039 ( .A1(n15730), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19297) );
  OAI211_X1 U17040 ( .C1(n19306), .C2(n15761), .A(n13674), .B(n19297), .ZN(
        n13679) );
  AOI21_X1 U17041 ( .B1(n10031), .B2(n13676), .A(n13675), .ZN(n19299) );
  NAND2_X1 U17042 ( .A1(n19319), .A2(n19299), .ZN(n13677) );
  OAI21_X1 U17043 ( .B1(n19202), .B2(n16466), .A(n13677), .ZN(n13678) );
  NOR2_X1 U17044 ( .A1(n13679), .A2(n13678), .ZN(n13680) );
  NAND2_X1 U17045 ( .A1(n13681), .A2(n13680), .ZN(P2_U3046) );
  INV_X1 U17046 ( .A(n11982), .ZN(n13847) );
  OAI22_X1 U17047 ( .A1(n13847), .A2(n15031), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15030), .ZN(n15939) );
  OAI22_X1 U17048 ( .A1(n20884), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15967), .ZN(n13682) );
  AOI21_X1 U17049 ( .B1(n15939), .B2(n13683), .A(n13682), .ZN(n13687) );
  AOI21_X1 U17050 ( .B1(n15940), .B2(n13683), .A(n13686), .ZN(n13685) );
  OAI22_X1 U17051 ( .A1(n13687), .A2(n13686), .B1(n13685), .B2(n13684), .ZN(
        P1_U3474) );
  OR2_X1 U17052 ( .A1(n13689), .A2(n13688), .ZN(n13691) );
  NAND2_X1 U17053 ( .A1(n13691), .A2(n13690), .ZN(n19146) );
  INV_X1 U17054 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19267) );
  OAI222_X1 U17055 ( .A1(n14148), .A2(n19370), .B1(n19146), .B2(n19243), .C1(
        n19267), .C2(n19249), .ZN(P2_U2912) );
  INV_X1 U17056 ( .A(n20978), .ZN(n20890) );
  AND2_X1 U17057 ( .A1(n20982), .A2(n20890), .ZN(n13692) );
  OR2_X1 U17058 ( .A1(n20144), .A2(n20272), .ZN(n13850) );
  NAND2_X1 U17059 ( .A1(n20144), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13696) );
  NOR2_X2 U17060 ( .A1(n20144), .A2(n11824), .ZN(n20155) );
  INV_X1 U17061 ( .A(DATAI_10_), .ZN(n13694) );
  INV_X1 U17062 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n13693) );
  MUX2_X1 U17063 ( .A(n13694), .B(n13693), .S(n20259), .Z(n14863) );
  INV_X1 U17064 ( .A(n14863), .ZN(n13695) );
  NAND2_X1 U17065 ( .A1(n20155), .A2(n13695), .ZN(n20161) );
  OAI211_X1 U17066 ( .C1(n13850), .C2(n14796), .A(n13696), .B(n20161), .ZN(
        P1_U2947) );
  INV_X1 U17067 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14843) );
  INV_X1 U17068 ( .A(n20155), .ZN(n13699) );
  INV_X1 U17069 ( .A(n20259), .ZN(n20257) );
  INV_X1 U17070 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13697) );
  NOR2_X1 U17071 ( .A1(n20257), .A2(n13697), .ZN(n13698) );
  AOI21_X1 U17072 ( .B1(DATAI_15_), .B2(n20257), .A(n13698), .ZN(n14842) );
  INV_X1 U17073 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20118) );
  OAI222_X1 U17074 ( .A1(n13850), .A2(n14843), .B1(n13699), .B2(n14842), .C1(
        n13859), .C2(n20118), .ZN(P1_U2967) );
  INV_X1 U17075 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n21189) );
  NAND2_X1 U17076 ( .A1(n20144), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13703) );
  INV_X1 U17077 ( .A(DATAI_11_), .ZN(n13701) );
  MUX2_X1 U17078 ( .A(n13701), .B(n13700), .S(n20259), .Z(n14859) );
  INV_X1 U17079 ( .A(n14859), .ZN(n13702) );
  NAND2_X1 U17080 ( .A1(n20155), .A2(n13702), .ZN(n13885) );
  OAI211_X1 U17081 ( .C1(n13850), .C2(n21189), .A(n13703), .B(n13885), .ZN(
        P1_U2963) );
  INV_X1 U17082 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13705) );
  NAND2_X1 U17083 ( .A1(n20119), .A2(n20261), .ZN(n13950) );
  AOI22_X1 U17084 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13704) );
  OAI21_X1 U17085 ( .B1(n13705), .B2(n13950), .A(n13704), .ZN(P1_U2912) );
  INV_X1 U17086 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13707) );
  AOI22_X1 U17087 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13706) );
  OAI21_X1 U17088 ( .B1(n13707), .B2(n13950), .A(n13706), .ZN(P1_U2907) );
  INV_X1 U17089 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21190) );
  AOI22_X1 U17090 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U17091 ( .B1(n21190), .B2(n13950), .A(n13708), .ZN(P1_U2911) );
  INV_X1 U17092 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13710) );
  AOI22_X1 U17093 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13709) );
  OAI21_X1 U17094 ( .B1(n13710), .B2(n13950), .A(n13709), .ZN(P1_U2908) );
  AOI22_X1 U17095 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13711) );
  OAI21_X1 U17096 ( .B1(n14796), .B2(n13950), .A(n13711), .ZN(P1_U2910) );
  AOI22_X1 U17097 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13712) );
  OAI21_X1 U17098 ( .B1(n14773), .B2(n13950), .A(n13712), .ZN(P1_U2906) );
  INV_X1 U17099 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14791) );
  AOI22_X1 U17100 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13713) );
  OAI21_X1 U17101 ( .B1(n14791), .B2(n13950), .A(n13713), .ZN(P1_U2909) );
  XNOR2_X1 U17102 ( .A(n13714), .B(n13715), .ZN(n19966) );
  INV_X1 U17103 ( .A(n19966), .ZN(n13716) );
  NAND2_X1 U17104 ( .A1(n19961), .A2(n13716), .ZN(n13770) );
  OAI21_X1 U17105 ( .B1(n19961), .B2(n13716), .A(n13770), .ZN(n13717) );
  NOR2_X1 U17106 ( .A1(n13717), .A2(n13718), .ZN(n13772) );
  AOI21_X1 U17107 ( .B1(n13718), .B2(n13717), .A(n13772), .ZN(n13721) );
  INV_X1 U17108 ( .A(n19345), .ZN(n15288) );
  AOI22_X1 U17109 ( .A1(n19245), .A2(n15288), .B1(n19239), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U17110 ( .A1(n13389), .A2(n19966), .ZN(n13719) );
  OAI211_X1 U17111 ( .C1(n13721), .C2(n15282), .A(n13720), .B(n13719), .ZN(
        P2_U2918) );
  NOR2_X1 U17112 ( .A1(n13727), .A2(n9750), .ZN(n13728) );
  AOI21_X1 U17113 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n9750), .A(n13728), .ZN(
        n13729) );
  OAI21_X1 U17114 ( .B1(n19944), .B2(n15178), .A(n13729), .ZN(P2_U2884) );
  NOR2_X1 U17115 ( .A1(n9815), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13731) );
  OR2_X1 U17116 ( .A1(n13731), .A2(n13730), .ZN(n14687) );
  NAND4_X1 U17117 ( .A1(n13733), .A2(n13732), .A3(n11828), .A4(n11826), .ZN(
        n14126) );
  OR2_X1 U17118 ( .A1(n14126), .A2(n14307), .ZN(n13734) );
  NAND2_X1 U17119 ( .A1(n13735), .A2(n13734), .ZN(n13736) );
  INV_X1 U17120 ( .A(n13737), .ZN(n13738) );
  AOI21_X1 U17121 ( .B1(n13740), .B2(n13739), .A(n13738), .ZN(n20193) );
  INV_X1 U17122 ( .A(n20193), .ZN(n14693) );
  NAND2_X1 U17123 ( .A1(n20115), .A2(n11827), .ZN(n14767) );
  OAI222_X1 U17124 ( .A1(n14687), .A2(n14769), .B1(n14686), .B2(n20115), .C1(
        n14693), .C2(n14767), .ZN(P1_U2872) );
  XOR2_X1 U17125 ( .A(n13741), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13745)
         );
  AND2_X1 U17126 ( .A1(n13752), .A2(n13742), .ZN(n13743) );
  OR2_X1 U17127 ( .A1(n13743), .A2(n13808), .ZN(n16454) );
  MUX2_X1 U17128 ( .A(n16454), .B(n10916), .S(n9769), .Z(n13744) );
  OAI21_X1 U17129 ( .B1(n13745), .B2(n15178), .A(n13744), .ZN(P2_U2882) );
  OR2_X1 U17130 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  AND2_X1 U17131 ( .A1(n13741), .A2(n13748), .ZN(n19190) );
  INV_X1 U17132 ( .A(n19190), .ZN(n13974) );
  NAND2_X1 U17133 ( .A1(n13750), .A2(n13749), .ZN(n13751) );
  NAND2_X1 U17134 ( .A1(n13752), .A2(n13751), .ZN(n19288) );
  NOR2_X1 U17135 ( .A1(n19288), .A2(n9769), .ZN(n13753) );
  AOI21_X1 U17136 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n9769), .A(n13753), .ZN(
        n13754) );
  OAI21_X1 U17137 ( .B1(n13974), .B2(n15178), .A(n13754), .ZN(P2_U2883) );
  INV_X1 U17138 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U17139 ( .A1(n20002), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13755) );
  OAI21_X1 U17140 ( .B1(n13756), .B2(n13768), .A(n13755), .ZN(P2_U2932) );
  INV_X1 U17141 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U17142 ( .A1(n20002), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13757) );
  OAI21_X1 U17143 ( .B1(n15273), .B2(n13768), .A(n13757), .ZN(P2_U2933) );
  AOI22_X1 U17144 ( .A1(n20002), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13758) );
  OAI21_X1 U17145 ( .B1(n13759), .B2(n13768), .A(n13758), .ZN(P2_U2935) );
  INV_X1 U17146 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U17147 ( .A1(n20002), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13760) );
  OAI21_X1 U17148 ( .B1(n13761), .B2(n13768), .A(n13760), .ZN(P2_U2929) );
  INV_X1 U17149 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U17150 ( .A1(n20002), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13762) );
  OAI21_X1 U17151 ( .B1(n13763), .B2(n13768), .A(n13762), .ZN(P2_U2934) );
  AOI22_X1 U17152 ( .A1(n20002), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13764) );
  OAI21_X1 U17153 ( .B1(n13588), .B2(n13768), .A(n13764), .ZN(P2_U2931) );
  INV_X1 U17154 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13766) );
  AOI22_X1 U17155 ( .A1(n20002), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13765) );
  OAI21_X1 U17156 ( .B1(n13766), .B2(n13768), .A(n13765), .ZN(P2_U2928) );
  INV_X1 U17157 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U17158 ( .A1(n20002), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13767) );
  OAI21_X1 U17159 ( .B1(n13769), .B2(n13768), .A(n13767), .ZN(P2_U2930) );
  INV_X1 U17160 ( .A(n13770), .ZN(n13771) );
  NOR2_X1 U17161 ( .A1(n13772), .A2(n13771), .ZN(n13778) );
  NAND2_X1 U17162 ( .A1(n13774), .A2(n13773), .ZN(n13776) );
  AND2_X1 U17163 ( .A1(n13776), .A2(n9770), .ZN(n19951) );
  NAND2_X1 U17164 ( .A1(n19953), .A2(n19951), .ZN(n13925) );
  OAI21_X1 U17165 ( .B1(n19953), .B2(n19951), .A(n13925), .ZN(n13777) );
  NOR2_X1 U17166 ( .A1(n13778), .A2(n13777), .ZN(n13927) );
  AOI21_X1 U17167 ( .B1(n13778), .B2(n13777), .A(n13927), .ZN(n13781) );
  INV_X1 U17168 ( .A(n19348), .ZN(n15271) );
  AOI22_X1 U17169 ( .A1(n19245), .A2(n15271), .B1(n19239), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13780) );
  INV_X1 U17170 ( .A(n19951), .ZN(n19327) );
  NAND2_X1 U17171 ( .A1(n19327), .A2(n13389), .ZN(n13779) );
  OAI211_X1 U17172 ( .C1(n13781), .C2(n15282), .A(n13780), .B(n13779), .ZN(
        P2_U2917) );
  XNOR2_X1 U17173 ( .A(n14678), .B(n14307), .ZN(n20235) );
  INV_X1 U17174 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13786) );
  OR2_X1 U17175 ( .A1(n13784), .A2(n13783), .ZN(n13785) );
  NAND2_X1 U17176 ( .A1(n13782), .A2(n13785), .ZN(n20189) );
  OAI222_X1 U17177 ( .A1(n20235), .A2(n14769), .B1(n13786), .B2(n20115), .C1(
        n20189), .C2(n14753), .ZN(P1_U2871) );
  NAND2_X1 U17178 ( .A1(n13787), .A2(n13782), .ZN(n13788) );
  AND2_X1 U17179 ( .A1(n13789), .A2(n13788), .ZN(n14666) );
  AOI22_X1 U17180 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13790) );
  OAI21_X1 U17181 ( .B1(n20179), .B2(n14676), .A(n13790), .ZN(n13791) );
  AOI21_X1 U17182 ( .B1(n14666), .B2(n20194), .A(n13791), .ZN(n13796) );
  OR2_X1 U17183 ( .A1(n13793), .A2(n13792), .ZN(n20221) );
  NAND3_X1 U17184 ( .A1(n20221), .A2(n13794), .A3(n20186), .ZN(n13795) );
  NAND2_X1 U17185 ( .A1(n13796), .A2(n13795), .ZN(P1_U2997) );
  INV_X1 U17186 ( .A(n14666), .ZN(n14136) );
  NOR2_X1 U17187 ( .A1(n13798), .A2(n13797), .ZN(n13799) );
  NOR2_X1 U17188 ( .A1(n20086), .A2(n13799), .ZN(n20220) );
  INV_X1 U17189 ( .A(n20115), .ZN(n14740) );
  AOI22_X1 U17190 ( .A1(n20112), .A2(n20220), .B1(n14740), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13800) );
  OAI21_X1 U17191 ( .B1(n14136), .B2(n14767), .A(n13800), .ZN(P1_U2870) );
  AOI21_X1 U17192 ( .B1(n20226), .B2(n20241), .A(n20218), .ZN(n20248) );
  AOI22_X1 U17193 ( .A1(n20248), .A2(n20240), .B1(n13801), .B2(n20241), .ZN(
        n13806) );
  OAI21_X1 U17194 ( .B1(n13802), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12696), .ZN(n20197) );
  NOR2_X1 U17195 ( .A1(n20197), .A2(n16291), .ZN(n13805) );
  INV_X1 U17196 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13803) );
  OR2_X1 U17197 ( .A1(n16230), .A2(n13803), .ZN(n20195) );
  OAI21_X1 U17198 ( .B1(n20230), .B2(n14687), .A(n20195), .ZN(n13804) );
  OR3_X1 U17199 ( .A1(n13806), .A2(n13805), .A3(n13804), .ZN(P1_U3031) );
  OR2_X1 U17200 ( .A1(n13808), .A2(n13807), .ZN(n13809) );
  AND2_X1 U17201 ( .A1(n13809), .A2(n13905), .ZN(n19159) );
  INV_X1 U17202 ( .A(n19159), .ZN(n13814) );
  NOR2_X1 U17203 ( .A1(n13741), .A2(n13810), .ZN(n13811) );
  OAI211_X1 U17204 ( .C1(n13811), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15212), .B(n13904), .ZN(n13813) );
  NAND2_X1 U17205 ( .A1(n9769), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13812) );
  OAI211_X1 U17206 ( .C1(n13814), .C2(n9769), .A(n13813), .B(n13812), .ZN(
        P2_U2881) );
  MUX2_X1 U17207 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13815), .S(
        n13821), .Z(n15947) );
  NOR2_X1 U17208 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20884), .ZN(n13822) );
  AOI22_X1 U17209 ( .A1(n15947), .A2(n20884), .B1(n13822), .B2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13818) );
  MUX2_X1 U17210 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13816), .S(
        n13821), .Z(n15945) );
  AOI22_X1 U17211 ( .A1(n13822), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15945), .B2(n20884), .ZN(n13817) );
  NOR2_X1 U17212 ( .A1(n13818), .A2(n13817), .ZN(n15958) );
  INV_X1 U17213 ( .A(n15958), .ZN(n13825) );
  INV_X1 U17214 ( .A(n20427), .ZN(n20689) );
  NOR2_X1 U17215 ( .A1(n13819), .A2(n20689), .ZN(n13820) );
  XNOR2_X1 U17216 ( .A(n13820), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20096) );
  OAI21_X1 U17217 ( .B1(n20096), .B2(n13617), .A(n13821), .ZN(n13824) );
  INV_X1 U17218 ( .A(n13821), .ZN(n15937) );
  AOI21_X1 U17219 ( .B1(n15937), .B2(n16315), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13823) );
  AOI22_X1 U17220 ( .A1(n13824), .A2(n13823), .B1(n13822), .B2(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15956) );
  OAI21_X1 U17221 ( .B1(n13825), .B2(n11708), .A(n15956), .ZN(n13846) );
  OAI21_X1 U17222 ( .B1(n13846), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13826), .ZN(
        n13827) );
  NOR2_X1 U17223 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20983) );
  NAND2_X1 U17224 ( .A1(n13827), .A2(n20432), .ZN(n20249) );
  OR2_X1 U17225 ( .A1(n13828), .A2(n13829), .ZN(n20759) );
  OR2_X1 U17226 ( .A1(n13828), .A2(n13830), .ZN(n20457) );
  MUX2_X1 U17227 ( .A(n20759), .B(n20457), .S(n13831), .Z(n13832) );
  NAND2_X1 U17228 ( .A1(n9752), .A2(n13828), .ZN(n20656) );
  AOI21_X1 U17229 ( .B1(n13832), .B2(n20656), .A(n13840), .ZN(n13835) );
  NOR2_X1 U17230 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20822), .ZN(n13838) );
  NAND2_X1 U17231 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20701), .ZN(n13837) );
  AOI22_X1 U17232 ( .A1(n9752), .A2(n13838), .B1(n13837), .B2(n20549), .ZN(
        n13833) );
  INV_X1 U17233 ( .A(n13833), .ZN(n13834) );
  OAI21_X1 U17234 ( .B1(n13835), .B2(n13834), .A(n20249), .ZN(n13836) );
  OAI21_X1 U17235 ( .B1(n20249), .B2(n20652), .A(n13836), .ZN(P1_U3475) );
  INV_X1 U17236 ( .A(n13837), .ZN(n15028) );
  NOR2_X1 U17237 ( .A1(n20690), .A2(n15028), .ZN(n13844) );
  OR2_X1 U17238 ( .A1(n13831), .A2(n20822), .ZN(n13839) );
  INV_X1 U17239 ( .A(n13838), .ZN(n20687) );
  NAND2_X1 U17240 ( .A1(n13839), .A2(n20687), .ZN(n20825) );
  INV_X1 U17241 ( .A(n13831), .ZN(n13841) );
  NOR2_X1 U17242 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  MUX2_X1 U17243 ( .A(n20825), .B(n13842), .S(n13828), .Z(n13843) );
  OAI21_X1 U17244 ( .B1(n13844), .B2(n13843), .A(n20249), .ZN(n13845) );
  OAI21_X1 U17245 ( .B1(n20249), .B2(n20611), .A(n13845), .ZN(P1_U3476) );
  NOR2_X1 U17246 ( .A1(n13846), .A2(n16326), .ZN(n15970) );
  OAI22_X1 U17247 ( .A1(n20349), .A2(n20822), .B1(n13847), .B2(n15028), .ZN(
        n13848) );
  OAI21_X1 U17248 ( .B1(n15970), .B2(n13848), .A(n20249), .ZN(n13849) );
  OAI21_X1 U17249 ( .B1(n20249), .B2(n20755), .A(n13849), .ZN(P1_U3478) );
  INV_X1 U17250 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19259) );
  OAI222_X1 U17251 ( .A1(n14148), .A2(n15225), .B1(n15677), .B2(n19243), .C1(
        n19259), .C2(n19249), .ZN(P2_U2908) );
  INV_X2 U17252 ( .A(n13850), .ZN(n20168) );
  AOI22_X1 U17253 ( .A1(n20168), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20167), .ZN(n13854) );
  NAND2_X1 U17254 ( .A1(n20257), .A2(DATAI_0_), .ZN(n13852) );
  NAND2_X1 U17255 ( .A1(n20259), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13851) );
  AND2_X1 U17256 ( .A1(n13852), .A2(n13851), .ZN(n20264) );
  INV_X1 U17257 ( .A(n20264), .ZN(n13853) );
  NAND2_X1 U17258 ( .A1(n20155), .A2(n13853), .ZN(n13891) );
  NAND2_X1 U17259 ( .A1(n13854), .A2(n13891), .ZN(P1_U2952) );
  AOI22_X1 U17260 ( .A1(n20168), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20167), .ZN(n13858) );
  NAND2_X1 U17261 ( .A1(n20257), .A2(DATAI_3_), .ZN(n13856) );
  NAND2_X1 U17262 ( .A1(n20259), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13855) );
  AND2_X1 U17263 ( .A1(n13856), .A2(n13855), .ZN(n20286) );
  INV_X1 U17264 ( .A(n20286), .ZN(n13857) );
  NAND2_X1 U17265 ( .A1(n20155), .A2(n13857), .ZN(n13860) );
  NAND2_X1 U17266 ( .A1(n13858), .A2(n13860), .ZN(P1_U2940) );
  INV_X1 U17267 ( .A(n13859), .ZN(n20167) );
  AOI22_X1 U17268 ( .A1(n20168), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20167), .ZN(n13861) );
  NAND2_X1 U17269 ( .A1(n13861), .A2(n13860), .ZN(P1_U2955) );
  AOI22_X1 U17270 ( .A1(n20168), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20167), .ZN(n13865) );
  NAND2_X1 U17271 ( .A1(n20257), .A2(DATAI_4_), .ZN(n13863) );
  NAND2_X1 U17272 ( .A1(n20259), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13862) );
  AND2_X1 U17273 ( .A1(n13863), .A2(n13862), .ZN(n20292) );
  INV_X1 U17274 ( .A(n20292), .ZN(n13864) );
  NAND2_X1 U17275 ( .A1(n20155), .A2(n13864), .ZN(n13881) );
  NAND2_X1 U17276 ( .A1(n13865), .A2(n13881), .ZN(P1_U2956) );
  AOI22_X1 U17277 ( .A1(n20168), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20167), .ZN(n13869) );
  NAND2_X1 U17278 ( .A1(n20257), .A2(DATAI_5_), .ZN(n13867) );
  NAND2_X1 U17279 ( .A1(n20259), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13866) );
  AND2_X1 U17280 ( .A1(n13867), .A2(n13866), .ZN(n20297) );
  INV_X1 U17281 ( .A(n20297), .ZN(n13868) );
  NAND2_X1 U17282 ( .A1(n20155), .A2(n13868), .ZN(n13897) );
  NAND2_X1 U17283 ( .A1(n13869), .A2(n13897), .ZN(P1_U2942) );
  AOI22_X1 U17284 ( .A1(n20168), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20167), .ZN(n13873) );
  NAND2_X1 U17285 ( .A1(n20257), .A2(DATAI_2_), .ZN(n13871) );
  NAND2_X1 U17286 ( .A1(n20259), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13870) );
  AND2_X1 U17287 ( .A1(n13871), .A2(n13870), .ZN(n20280) );
  INV_X1 U17288 ( .A(n20280), .ZN(n13872) );
  NAND2_X1 U17289 ( .A1(n20155), .A2(n13872), .ZN(n13899) );
  NAND2_X1 U17290 ( .A1(n13873), .A2(n13899), .ZN(P1_U2954) );
  AOI22_X1 U17291 ( .A1(n20168), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20167), .ZN(n13877) );
  NAND2_X1 U17292 ( .A1(n20257), .A2(DATAI_1_), .ZN(n13875) );
  NAND2_X1 U17293 ( .A1(n20259), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13874) );
  AND2_X1 U17294 ( .A1(n13875), .A2(n13874), .ZN(n20274) );
  INV_X1 U17295 ( .A(n20274), .ZN(n13876) );
  NAND2_X1 U17296 ( .A1(n20155), .A2(n13876), .ZN(n13895) );
  NAND2_X1 U17297 ( .A1(n13877), .A2(n13895), .ZN(P1_U2938) );
  AOI22_X1 U17298 ( .A1(n20168), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20167), .ZN(n13880) );
  INV_X1 U17299 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16595) );
  NAND2_X1 U17300 ( .A1(n20259), .A2(n16595), .ZN(n13878) );
  OAI21_X1 U17301 ( .B1(n20259), .B2(DATAI_7_), .A(n13878), .ZN(n20316) );
  INV_X1 U17302 ( .A(n20316), .ZN(n13879) );
  NAND2_X1 U17303 ( .A1(n20155), .A2(n13879), .ZN(n13883) );
  NAND2_X1 U17304 ( .A1(n13880), .A2(n13883), .ZN(P1_U2944) );
  AOI22_X1 U17305 ( .A1(n20168), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20167), .ZN(n13882) );
  NAND2_X1 U17306 ( .A1(n13882), .A2(n13881), .ZN(P1_U2941) );
  AOI22_X1 U17307 ( .A1(n20168), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20167), .ZN(n13884) );
  NAND2_X1 U17308 ( .A1(n13884), .A2(n13883), .ZN(P1_U2959) );
  AOI22_X1 U17309 ( .A1(n20168), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20167), .ZN(n13886) );
  NAND2_X1 U17310 ( .A1(n13886), .A2(n13885), .ZN(P1_U2948) );
  AOI22_X1 U17311 ( .A1(n20168), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20167), .ZN(n13890) );
  NAND2_X1 U17312 ( .A1(n20257), .A2(DATAI_6_), .ZN(n13888) );
  NAND2_X1 U17313 ( .A1(n20259), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13887) );
  AND2_X1 U17314 ( .A1(n13888), .A2(n13887), .ZN(n20306) );
  INV_X1 U17315 ( .A(n20306), .ZN(n13889) );
  NAND2_X1 U17316 ( .A1(n20155), .A2(n13889), .ZN(n13893) );
  NAND2_X1 U17317 ( .A1(n13890), .A2(n13893), .ZN(P1_U2943) );
  AOI22_X1 U17318 ( .A1(n20168), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20167), .ZN(n13892) );
  NAND2_X1 U17319 ( .A1(n13892), .A2(n13891), .ZN(P1_U2937) );
  AOI22_X1 U17320 ( .A1(n20168), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20167), .ZN(n13894) );
  NAND2_X1 U17321 ( .A1(n13894), .A2(n13893), .ZN(P1_U2958) );
  AOI22_X1 U17322 ( .A1(n20168), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20167), .ZN(n13896) );
  NAND2_X1 U17323 ( .A1(n13896), .A2(n13895), .ZN(P1_U2953) );
  AOI22_X1 U17324 ( .A1(n20168), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20167), .ZN(n13898) );
  NAND2_X1 U17325 ( .A1(n13898), .A2(n13897), .ZN(P1_U2957) );
  AOI22_X1 U17326 ( .A1(n20168), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20167), .ZN(n13900) );
  NAND2_X1 U17327 ( .A1(n13900), .A2(n13899), .ZN(P1_U2939) );
  AOI22_X1 U17328 ( .A1(n20168), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20167), .ZN(n13903) );
  INV_X1 U17329 ( .A(DATAI_9_), .ZN(n13901) );
  MUX2_X1 U17330 ( .A(n13901), .B(n16592), .S(n20259), .Z(n14800) );
  INV_X1 U17331 ( .A(n14800), .ZN(n13902) );
  NAND2_X1 U17332 ( .A1(n20155), .A2(n13902), .ZN(n20159) );
  NAND2_X1 U17333 ( .A1(n13903), .A2(n20159), .ZN(P1_U2946) );
  XOR2_X1 U17334 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13904), .Z(n13911)
         );
  NAND2_X1 U17335 ( .A1(n13906), .A2(n13905), .ZN(n13908) );
  INV_X1 U17336 ( .A(n13960), .ZN(n13907) );
  NAND2_X1 U17337 ( .A1(n13908), .A2(n13907), .ZN(n19145) );
  INV_X1 U17338 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13909) );
  MUX2_X1 U17339 ( .A(n19145), .B(n13909), .S(n9750), .Z(n13910) );
  OAI21_X1 U17340 ( .B1(n13911), .B2(n15178), .A(n13910), .ZN(P2_U2880) );
  INV_X1 U17341 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n13919) );
  AOI21_X1 U17342 ( .B1(n13914), .B2(n13912), .A(n13913), .ZN(n19183) );
  NAND2_X1 U17343 ( .A1(n19190), .A2(n19183), .ZN(n13975) );
  INV_X1 U17344 ( .A(n13975), .ZN(n13917) );
  OAI21_X1 U17345 ( .B1(n13913), .B2(n13916), .A(n13915), .ZN(n19177) );
  INV_X1 U17346 ( .A(n19177), .ZN(n15753) );
  AOI21_X1 U17347 ( .B1(n13917), .B2(n19225), .A(n15753), .ZN(n13918) );
  OAI222_X1 U17348 ( .A1(n13919), .A2(n19249), .B1(n14148), .B2(n19359), .C1(
        n19243), .C2(n13918), .ZN(P2_U2914) );
  OR2_X1 U17349 ( .A1(n13922), .A2(n13921), .ZN(n13923) );
  AND2_X1 U17350 ( .A1(n13920), .A2(n13923), .ZN(n14651) );
  INV_X1 U17351 ( .A(n14651), .ZN(n14138) );
  XOR2_X1 U17352 ( .A(n20085), .B(n20086), .Z(n20210) );
  AOI22_X1 U17353 ( .A1(n20210), .A2(n20112), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14740), .ZN(n13924) );
  OAI21_X1 U17354 ( .B1(n14138), .B2(n14753), .A(n13924), .ZN(P1_U2869) );
  INV_X1 U17355 ( .A(n13925), .ZN(n13926) );
  NOR2_X1 U17356 ( .A1(n13927), .A2(n13926), .ZN(n13932) );
  OR2_X1 U17357 ( .A1(n13929), .A2(n13928), .ZN(n13930) );
  NAND2_X1 U17358 ( .A1(n13930), .A2(n13912), .ZN(n13972) );
  XNOR2_X1 U17359 ( .A(n19944), .B(n13972), .ZN(n13931) );
  NOR2_X1 U17360 ( .A1(n13932), .A2(n13931), .ZN(n13971) );
  AOI21_X1 U17361 ( .B1(n13932), .B2(n13931), .A(n13971), .ZN(n13935) );
  INV_X1 U17362 ( .A(n19352), .ZN(n15266) );
  AOI22_X1 U17363 ( .A1(n19245), .A2(n15266), .B1(n19239), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n13934) );
  INV_X1 U17364 ( .A(n13972), .ZN(n19948) );
  NAND2_X1 U17365 ( .A1(n19948), .A2(n13389), .ZN(n13933) );
  OAI211_X1 U17366 ( .C1(n13935), .C2(n15282), .A(n13934), .B(n13933), .ZN(
        P2_U2916) );
  INV_X1 U17367 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U17368 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13936) );
  OAI21_X1 U17369 ( .B1(n13937), .B2(n13950), .A(n13936), .ZN(P1_U2920) );
  INV_X1 U17370 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17371 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13938) );
  OAI21_X1 U17372 ( .B1(n13939), .B2(n13950), .A(n13938), .ZN(P1_U2914) );
  INV_X1 U17373 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13941) );
  AOI22_X1 U17374 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13940) );
  OAI21_X1 U17375 ( .B1(n13941), .B2(n13950), .A(n13940), .ZN(P1_U2913) );
  INV_X1 U17376 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U17377 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13942) );
  OAI21_X1 U17378 ( .B1(n13943), .B2(n13950), .A(n13942), .ZN(P1_U2918) );
  INV_X1 U17379 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13945) );
  AOI22_X1 U17380 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13944) );
  OAI21_X1 U17381 ( .B1(n13945), .B2(n13950), .A(n13944), .ZN(P1_U2917) );
  INV_X1 U17382 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U17383 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13946) );
  OAI21_X1 U17384 ( .B1(n13947), .B2(n13950), .A(n13946), .ZN(P1_U2916) );
  INV_X1 U17385 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14816) );
  AOI22_X1 U17386 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13948) );
  OAI21_X1 U17387 ( .B1(n14816), .B2(n13950), .A(n13948), .ZN(P1_U2915) );
  INV_X1 U17388 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U17389 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13949) );
  OAI21_X1 U17390 ( .B1(n13951), .B2(n13950), .A(n13949), .ZN(P1_U2919) );
  OAI21_X1 U17391 ( .B1(n13954), .B2(n13953), .A(n13952), .ZN(n20211) );
  AOI22_X1 U17392 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13955) );
  OAI21_X1 U17393 ( .B1(n20179), .B2(n14665), .A(n13955), .ZN(n13956) );
  AOI21_X1 U17394 ( .B1(n14651), .B2(n20194), .A(n13956), .ZN(n13957) );
  OAI21_X1 U17395 ( .B1(n20211), .B2(n20198), .A(n13957), .ZN(P1_U2996) );
  INV_X1 U17396 ( .A(n13967), .ZN(n13958) );
  OAI21_X1 U17397 ( .B1(n13960), .B2(n13959), .A(n13958), .ZN(n19139) );
  OAI211_X1 U17398 ( .C1(n13963), .C2(n13962), .A(n13961), .B(n15212), .ZN(
        n13965) );
  NAND2_X1 U17399 ( .A1(n9769), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13964) );
  OAI211_X1 U17400 ( .C1(n19139), .C2(n9769), .A(n13965), .B(n13964), .ZN(
        P2_U2879) );
  XNOR2_X1 U17401 ( .A(n13961), .B(n14080), .ZN(n13970) );
  NOR2_X1 U17402 ( .A1(n13967), .A2(n13966), .ZN(n13968) );
  OR2_X1 U17403 ( .A1(n14084), .A2(n13968), .ZN(n15702) );
  MUX2_X1 U17404 ( .A(n15702), .B(n10917), .S(n9750), .Z(n13969) );
  OAI21_X1 U17405 ( .B1(n13970), .B2(n15178), .A(n13969), .ZN(P2_U2878) );
  AOI21_X1 U17406 ( .B1(n13972), .B2(n19944), .A(n13971), .ZN(n13977) );
  INV_X1 U17407 ( .A(n19183), .ZN(n13973) );
  NAND2_X1 U17408 ( .A1(n13974), .A2(n13973), .ZN(n13976) );
  OAI211_X1 U17409 ( .C1(n13977), .C2(n13976), .A(n19225), .B(n13975), .ZN(
        n13979) );
  AOI22_X1 U17410 ( .A1(n13389), .A2(n19183), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19239), .ZN(n13978) );
  OAI211_X1 U17411 ( .C1(n19356), .C2(n14148), .A(n13979), .B(n13978), .ZN(
        P2_U2915) );
  INV_X1 U17412 ( .A(n14412), .ZN(n13985) );
  INV_X1 U17413 ( .A(n13980), .ZN(n13984) );
  INV_X1 U17414 ( .A(n13981), .ZN(n13982) );
  NAND2_X1 U17415 ( .A1(n13982), .A2(n9866), .ZN(n13983) );
  NAND2_X1 U17416 ( .A1(n13984), .A2(n13983), .ZN(n19097) );
  INV_X1 U17417 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19255) );
  OAI222_X1 U17418 ( .A1(n14148), .A2(n13985), .B1(n19097), .B2(n19243), .C1(
        n19255), .C2(n19249), .ZN(P2_U2906) );
  OR2_X1 U17419 ( .A1(n13988), .A2(n13987), .ZN(n13989) );
  AND2_X1 U17420 ( .A1(n13986), .A2(n13989), .ZN(n20082) );
  INV_X1 U17421 ( .A(n20082), .ZN(n14137) );
  XNOR2_X1 U17422 ( .A(n13990), .B(n16298), .ZN(n20079) );
  AOI22_X1 U17423 ( .A1(n20112), .A2(n20079), .B1(n14740), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13991) );
  OAI21_X1 U17424 ( .B1(n14137), .B2(n14767), .A(n13991), .ZN(P1_U2867) );
  INV_X1 U17425 ( .A(n14021), .ZN(n14028) );
  OR2_X1 U17426 ( .A1(n13727), .A2(n14028), .ZN(n14005) );
  NOR2_X1 U17427 ( .A1(n14041), .A2(n14044), .ZN(n14027) );
  NOR2_X1 U17428 ( .A1(n13992), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14024) );
  NAND2_X1 U17429 ( .A1(n13993), .A2(n10371), .ZN(n13994) );
  AOI21_X1 U17430 ( .B1(n11005), .B2(n13998), .A(n13994), .ZN(n13995) );
  OAI21_X1 U17431 ( .B1(n14027), .B2(n14024), .A(n13995), .ZN(n14003) );
  NAND2_X1 U17432 ( .A1(n10436), .A2(n13996), .ZN(n14031) );
  OAI21_X1 U17433 ( .B1(n14031), .B2(n10371), .A(n13997), .ZN(n14001) );
  INV_X1 U17434 ( .A(n13998), .ZN(n13999) );
  NAND2_X1 U17435 ( .A1(n11005), .A2(n13999), .ZN(n14026) );
  INV_X1 U17436 ( .A(n14024), .ZN(n14000) );
  NAND3_X1 U17437 ( .A1(n14001), .A2(n14026), .A3(n14000), .ZN(n14002) );
  NAND2_X1 U17438 ( .A1(n14003), .A2(n14002), .ZN(n14004) );
  AND2_X1 U17439 ( .A1(n14005), .A2(n14004), .ZN(n15785) );
  NAND2_X1 U17440 ( .A1(n14006), .A2(n14048), .ZN(n14011) );
  AND3_X1 U17441 ( .A1(n14009), .A2(n14008), .A3(n14007), .ZN(n14010) );
  NAND2_X1 U17442 ( .A1(n15785), .A2(n14264), .ZN(n14013) );
  NAND2_X1 U17443 ( .A1(n14040), .A2(n10371), .ZN(n14012) );
  INV_X1 U17444 ( .A(n14014), .ZN(n14015) );
  OR2_X1 U17445 ( .A1(n11000), .A2(n14015), .ZN(n14019) );
  NOR2_X1 U17446 ( .A1(n14016), .A2(n13992), .ZN(n14017) );
  AOI22_X1 U17447 ( .A1(n10563), .A2(n11005), .B1(n14019), .B2(n14017), .ZN(
        n14018) );
  OAI21_X1 U17448 ( .B1(n15092), .B2(n14028), .A(n14018), .ZN(n15781) );
  INV_X1 U17449 ( .A(n15781), .ZN(n14022) );
  MUX2_X1 U17450 ( .A(n14019), .B(n11005), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14020) );
  AOI21_X1 U17451 ( .B1(n19301), .B2(n14021), .A(n14020), .ZN(n15774) );
  OAI211_X1 U17452 ( .C1(n14022), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15774), .ZN(n14023) );
  OAI211_X1 U17453 ( .C1(n19968), .C2(n15781), .A(n14023), .B(n14264), .ZN(
        n14036) );
  NOR2_X1 U17454 ( .A1(n14024), .A2(n9767), .ZN(n14032) );
  OAI22_X1 U17455 ( .A1(n14027), .A2(n14032), .B1(n14025), .B2(n14026), .ZN(
        n14030) );
  NOR2_X1 U17456 ( .A1(n13670), .A2(n14028), .ZN(n14029) );
  AOI211_X1 U17457 ( .C1(n14032), .C2(n14031), .A(n14030), .B(n14029), .ZN(
        n14033) );
  INV_X1 U17458 ( .A(n14033), .ZN(n14263) );
  AOI22_X1 U17459 ( .A1(n14040), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n14263), .B2(n14264), .ZN(n14039) );
  OR2_X1 U17460 ( .A1(n14039), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14035) );
  OAI21_X1 U17461 ( .B1(n19950), .B2(n14064), .A(n19958), .ZN(n14034) );
  AOI222_X1 U17462 ( .A1(n14036), .A2(n14035), .B1(n14036), .B2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C1(n14035), .C2(n14034), .ZN(
        n14037) );
  AOI21_X1 U17463 ( .B1(n19950), .B2(n14064), .A(n14037), .ZN(n14038) );
  OR2_X1 U17464 ( .A1(n14038), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n14066) );
  INV_X1 U17465 ( .A(n14039), .ZN(n14063) );
  NAND2_X1 U17466 ( .A1(n14040), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14061) );
  INV_X1 U17467 ( .A(n14041), .ZN(n14047) );
  NAND2_X1 U17468 ( .A1(n14043), .A2(n14042), .ZN(n14046) );
  NAND2_X1 U17469 ( .A1(n14093), .A2(n14044), .ZN(n14045) );
  OAI211_X1 U17470 ( .C1(n14093), .C2(n14047), .A(n14046), .B(n14045), .ZN(
        n19984) );
  INV_X1 U17471 ( .A(n14048), .ZN(n14049) );
  NAND2_X1 U17472 ( .A1(n14050), .A2(n14049), .ZN(n14051) );
  NOR2_X1 U17473 ( .A1(n14052), .A2(n14051), .ZN(n18986) );
  OAI21_X1 U17474 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n18986), .ZN(n14056) );
  INV_X1 U17475 ( .A(n15788), .ZN(n14053) );
  NAND3_X1 U17476 ( .A1(n14054), .A2(n10625), .A3(n14053), .ZN(n14055) );
  OAI211_X1 U17477 ( .C1(n14058), .C2(n14057), .A(n14056), .B(n14055), .ZN(
        n14059) );
  NOR2_X1 U17478 ( .A1(n19984), .A2(n14059), .ZN(n14060) );
  NAND2_X1 U17479 ( .A1(n14061), .A2(n14060), .ZN(n14062) );
  AOI21_X1 U17480 ( .B1(n14064), .B2(n14063), .A(n14062), .ZN(n14065) );
  NAND2_X1 U17481 ( .A1(n16515), .A2(n10456), .ZN(n14072) );
  OR2_X1 U17482 ( .A1(n14067), .A2(n19995), .ZN(n19999) );
  INV_X1 U17483 ( .A(n19999), .ZN(n14068) );
  OAI21_X1 U17484 ( .B1(n14070), .B2(n14069), .A(n14068), .ZN(n14071) );
  AOI21_X1 U17485 ( .B1(n14072), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14071), 
        .ZN(n16510) );
  OAI21_X1 U17486 ( .B1(n16510), .B2(n16509), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14074) );
  NOR2_X1 U17487 ( .A1(n16509), .A2(n14094), .ZN(n16507) );
  INV_X1 U17488 ( .A(n16507), .ZN(n14073) );
  NAND2_X1 U17489 ( .A1(n14074), .A2(n14073), .ZN(P2_U3593) );
  OAI211_X1 U17490 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20001), .A(n14076), 
        .B(n14075), .ZN(n14078) );
  NOR2_X1 U17491 ( .A1(n16509), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n18982) );
  OAI211_X1 U17492 ( .C1(n16510), .C2(n18982), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n19996), .ZN(n14077) );
  OAI211_X1 U17493 ( .C1(n16510), .C2(n14078), .A(n14077), .B(n19216), .ZN(
        P2_U3177) );
  OAI21_X1 U17494 ( .B1(n13961), .B2(n14080), .A(n14079), .ZN(n14082) );
  NAND3_X1 U17495 ( .A1(n14082), .A2(n15212), .A3(n14081), .ZN(n14088) );
  OR2_X1 U17496 ( .A1(n14084), .A2(n14083), .ZN(n14085) );
  NAND2_X1 U17497 ( .A1(n14085), .A2(n13451), .ZN(n19119) );
  INV_X1 U17498 ( .A(n19119), .ZN(n14086) );
  NAND2_X1 U17499 ( .A1(n15205), .A2(n14086), .ZN(n14087) );
  OAI211_X1 U17500 ( .C1(n15205), .C2(n19111), .A(n14088), .B(n14087), .ZN(
        P2_U2877) );
  NOR2_X1 U17501 ( .A1(n19944), .A2(n19781), .ZN(n19732) );
  NAND2_X1 U17502 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14089), .ZN(
        n19778) );
  INV_X1 U17503 ( .A(n19778), .ZN(n14098) );
  AOI21_X1 U17504 ( .B1(n19732), .B2(n19545), .A(n14098), .ZN(n14097) );
  INV_X1 U17505 ( .A(n14090), .ZN(n14091) );
  AND2_X1 U17506 ( .A1(n14091), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19855) );
  OR2_X1 U17507 ( .A1(n19855), .A2(n19995), .ZN(n14092) );
  NOR2_X1 U17508 ( .A1(n11123), .A2(n14092), .ZN(n14100) );
  AOI21_X1 U17509 ( .B1(n10456), .B2(n19995), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19993) );
  NAND2_X1 U17510 ( .A1(n19993), .A2(n14094), .ZN(n14095) );
  OAI21_X1 U17511 ( .B1(n19855), .B2(n20000), .A(n19738), .ZN(n14096) );
  INV_X1 U17512 ( .A(n19849), .ZN(n19865) );
  INV_X1 U17513 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14112) );
  AOI21_X1 U17514 ( .B1(n20000), .B2(n14098), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14099) );
  NOR2_X1 U17515 ( .A1(n14100), .A2(n14099), .ZN(n19857) );
  NOR2_X2 U17516 ( .A1(n14101), .A2(n19784), .ZN(n19790) );
  INV_X1 U17517 ( .A(n19367), .ZN(n14102) );
  AND2_X1 U17518 ( .A1(n14103), .A2(n14102), .ZN(n19779) );
  INV_X1 U17519 ( .A(n19779), .ZN(n14109) );
  INV_X1 U17520 ( .A(n19855), .ZN(n14108) );
  AOI22_X1 U17521 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19365), .ZN(n19793) );
  NOR2_X2 U17522 ( .A1(n19744), .A2(n19937), .ZN(n19861) );
  AOI22_X1 U17523 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19365), .ZN(n19710) );
  INV_X1 U17524 ( .A(n19710), .ZN(n19780) );
  AOI22_X1 U17525 ( .A1(n19859), .A2(n19747), .B1(n19861), .B2(n19780), .ZN(
        n14107) );
  OAI21_X1 U17526 ( .B1(n14109), .B2(n14108), .A(n14107), .ZN(n14110) );
  AOI21_X1 U17527 ( .B1(n19857), .B2(n19790), .A(n14110), .ZN(n14111) );
  OAI21_X1 U17528 ( .B1(n19865), .B2(n14112), .A(n14111), .ZN(P2_U3168) );
  NAND2_X1 U17529 ( .A1(n14114), .A2(n14113), .ZN(n14116) );
  XNOR2_X1 U17530 ( .A(n14116), .B(n14115), .ZN(n16499) );
  XNOR2_X1 U17531 ( .A(n14117), .B(n14118), .ZN(n16497) );
  NAND2_X1 U17532 ( .A1(n15730), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16493) );
  OAI21_X1 U17533 ( .B1(n16462), .B2(n14185), .A(n16493), .ZN(n14119) );
  AOI21_X1 U17534 ( .B1(n16453), .B2(n14182), .A(n14119), .ZN(n14122) );
  NAND2_X1 U17535 ( .A1(n14120), .A2(n19302), .ZN(n14121) );
  OAI211_X1 U17536 ( .C1(n16497), .C2(n16456), .A(n14122), .B(n14121), .ZN(
        n14123) );
  AOI21_X1 U17537 ( .B1(n16499), .B2(n19283), .A(n14123), .ZN(n14124) );
  INV_X1 U17538 ( .A(n14124), .ZN(P2_U3011) );
  NOR2_X1 U17539 ( .A1(n14125), .A2(n20890), .ZN(n14129) );
  NOR2_X1 U17540 ( .A1(n14126), .A2(n14650), .ZN(n14127) );
  AOI21_X1 U17541 ( .B1(n14129), .B2(n14128), .A(n14127), .ZN(n14130) );
  NAND2_X1 U17542 ( .A1(n14131), .A2(n14130), .ZN(n14133) );
  NAND2_X1 U17543 ( .A1(n14134), .A2(n11827), .ZN(n14135) );
  INV_X1 U17544 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20137) );
  OAI222_X1 U17545 ( .A1(n14866), .A2(n14136), .B1(n14861), .B2(n20137), .C1(
        n14864), .C2(n20280), .ZN(P1_U2902) );
  INV_X1 U17546 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20131) );
  OAI222_X1 U17547 ( .A1(n14866), .A2(n14137), .B1(n14861), .B2(n20131), .C1(
        n14864), .C2(n20297), .ZN(P1_U2899) );
  INV_X1 U17548 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20135) );
  OAI222_X1 U17549 ( .A1(n14866), .A2(n14138), .B1(n14861), .B2(n20135), .C1(
        n14864), .C2(n20286), .ZN(P1_U2901) );
  INV_X1 U17550 ( .A(n14139), .ZN(n14140) );
  XNOR2_X1 U17551 ( .A(n13920), .B(n14140), .ZN(n20175) );
  INV_X1 U17552 ( .A(n20175), .ZN(n14142) );
  INV_X1 U17553 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n14141) );
  OAI222_X1 U17554 ( .A1(n14866), .A2(n14142), .B1(n14141), .B2(n14861), .C1(
        n14864), .C2(n20292), .ZN(P1_U2900) );
  INV_X1 U17555 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20139) );
  OAI222_X1 U17556 ( .A1(n14866), .A2(n20189), .B1(n14861), .B2(n20139), .C1(
        n14864), .C2(n20274), .ZN(P1_U2903) );
  INV_X1 U17557 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20143) );
  OAI222_X1 U17558 ( .A1(n14866), .A2(n14693), .B1(n14861), .B2(n20143), .C1(
        n14864), .C2(n20264), .ZN(P1_U2904) );
  AND2_X1 U17559 ( .A1(n14143), .A2(n14144), .ZN(n14146) );
  OR2_X1 U17560 ( .A1(n14146), .A2(n14145), .ZN(n19069) );
  OAI222_X1 U17561 ( .A1(n14148), .A2(n14147), .B1(n19069), .B2(n19243), .C1(
        n13526), .C2(n19249), .ZN(P2_U2904) );
  NAND2_X1 U17562 ( .A1(n14150), .A2(n14149), .ZN(n14151) );
  XNOR2_X1 U17563 ( .A(n14151), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19285) );
  INV_X1 U17564 ( .A(n19285), .ZN(n14158) );
  XNOR2_X1 U17565 ( .A(n14152), .B(n9882), .ZN(n19284) );
  AOI22_X1 U17566 ( .A1(n19326), .A2(n19183), .B1(n15730), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n14153) );
  OAI21_X1 U17567 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15748), .A(
        n14153), .ZN(n14156) );
  NAND2_X1 U17568 ( .A1(n14154), .A2(n16492), .ZN(n15756) );
  OAI22_X1 U17569 ( .A1(n15756), .A2(n15750), .B1(n19317), .B2(n19288), .ZN(
        n14155) );
  AOI211_X1 U17570 ( .C1(n19284), .C2(n19316), .A(n14156), .B(n14155), .ZN(
        n14157) );
  OAI21_X1 U17571 ( .B1(n16496), .B2(n14158), .A(n14157), .ZN(P2_U3042) );
  OR2_X1 U17572 ( .A1(n16300), .A2(n14159), .ZN(n14160) );
  NAND2_X1 U17573 ( .A1(n14176), .A2(n14160), .ZN(n20048) );
  AND2_X1 U17574 ( .A1(n14162), .A2(n14161), .ZN(n14164) );
  OR2_X1 U17575 ( .A1(n14164), .A2(n14163), .ZN(n20052) );
  OAI222_X1 U17576 ( .A1(n20048), .A2(n14769), .B1(n14165), .B2(n20115), .C1(
        n20052), .C2(n14767), .ZN(P1_U2865) );
  AOI211_X1 U17577 ( .C1(n14167), .C2(n14081), .A(n15178), .B(n14166), .ZN(
        n14168) );
  INV_X1 U17578 ( .A(n14168), .ZN(n14170) );
  NAND2_X1 U17579 ( .A1(n15205), .A2(n16419), .ZN(n14169) );
  OAI211_X1 U17580 ( .C1(n15205), .C2(n10918), .A(n14170), .B(n14169), .ZN(
        P2_U2876) );
  INV_X1 U17581 ( .A(n14171), .ZN(n14174) );
  INV_X1 U17582 ( .A(n14163), .ZN(n14173) );
  AOI21_X1 U17583 ( .B1(n14174), .B2(n14173), .A(n14172), .ZN(n14274) );
  INV_X1 U17584 ( .A(n14274), .ZN(n14233) );
  INV_X1 U17585 ( .A(n14241), .ZN(n14175) );
  AOI21_X1 U17586 ( .B1(n14177), .B2(n14176), .A(n14175), .ZN(n16278) );
  AOI22_X1 U17587 ( .A1(n16278), .A2(n20112), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14740), .ZN(n14178) );
  OAI21_X1 U17588 ( .B1(n14233), .B2(n14767), .A(n14178), .ZN(P1_U2864) );
  INV_X1 U17589 ( .A(n19211), .ZN(n14229) );
  NAND2_X1 U17590 ( .A1(n9977), .A2(n14180), .ZN(n14181) );
  XNOR2_X1 U17591 ( .A(n14182), .B(n14181), .ZN(n14183) );
  NAND2_X1 U17592 ( .A1(n14183), .A2(n19174), .ZN(n14191) );
  NOR2_X1 U17593 ( .A1(n19201), .A2(n14184), .ZN(n14187) );
  OAI22_X1 U17594 ( .A1(n14185), .A2(n19178), .B1(n10663), .B2(n19204), .ZN(
        n14186) );
  AOI211_X1 U17595 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19207), .A(n14187), .B(
        n14186), .ZN(n14188) );
  OAI21_X1 U17596 ( .B1(n13727), .B2(n19209), .A(n14188), .ZN(n14189) );
  AOI21_X1 U17597 ( .B1(n19182), .B2(n19948), .A(n14189), .ZN(n14190) );
  OAI211_X1 U17598 ( .C1(n14229), .C2(n19944), .A(n14191), .B(n14190), .ZN(
        P2_U2852) );
  NAND2_X1 U17599 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20983), .ZN(n16320) );
  NAND2_X1 U17600 ( .A1(n14192), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14193) );
  MUX2_X1 U17601 ( .A(n16320), .B(n14193), .S(n20885), .Z(n14194) );
  AND2_X1 U17602 ( .A1(n16230), .A2(n14194), .ZN(n14195) );
  NAND2_X1 U17603 ( .A1(n14636), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14213) );
  INV_X1 U17604 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20910) );
  NAND3_X1 U17605 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20100) );
  NOR2_X1 U17606 ( .A1(n20910), .A2(n20100), .ZN(n14440) );
  NAND2_X1 U17607 ( .A1(n14440), .A2(n14636), .ZN(n14199) );
  AND2_X1 U17608 ( .A1(n20978), .A2(n20789), .ZN(n15961) );
  OAI21_X1 U17609 ( .B1(n20272), .B2(n15960), .A(n15961), .ZN(n14204) );
  NOR2_X1 U17610 ( .A1(n14204), .A2(n14197), .ZN(n14198) );
  NAND2_X1 U17611 ( .A1(n20101), .A2(n14636), .ZN(n14685) );
  AND2_X1 U17612 ( .A1(n14199), .A2(n14685), .ZN(n20103) );
  INV_X1 U17613 ( .A(n20103), .ZN(n20045) );
  INV_X1 U17614 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20917) );
  NAND3_X1 U17615 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .ZN(n14203) );
  NOR2_X1 U17616 ( .A1(n20917), .A2(n14203), .ZN(n20041) );
  INV_X1 U17617 ( .A(n20041), .ZN(n14200) );
  NAND2_X1 U17618 ( .A1(n14685), .A2(n14200), .ZN(n14201) );
  NAND2_X1 U17619 ( .A1(n20045), .A2(n14201), .ZN(n20033) );
  INV_X1 U17620 ( .A(n16278), .ZN(n14212) );
  NAND2_X1 U17621 ( .A1(n9818), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14205) );
  NOR2_X1 U17622 ( .A1(n14205), .A2(n15961), .ZN(n14202) );
  NOR3_X1 U17623 ( .A1(n20101), .A2(n20100), .A3(n20910), .ZN(n20074) );
  NOR2_X1 U17624 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14203), .ZN(n14210) );
  AND3_X1 U17625 ( .A1(n14205), .A2(n20261), .A3(n14204), .ZN(n14206) );
  INV_X1 U17626 ( .A(n20071), .ZN(n20094) );
  NAND2_X1 U17627 ( .A1(n14636), .A2(n14436), .ZN(n20091) );
  INV_X1 U17628 ( .A(n20091), .ZN(n20050) );
  AOI21_X1 U17629 ( .B1(n20051), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20050), .ZN(n14207) );
  OAI21_X1 U17630 ( .B1(n20094), .B2(n14208), .A(n14207), .ZN(n14209) );
  AOI21_X1 U17631 ( .B1(n20074), .B2(n14210), .A(n14209), .ZN(n14211) );
  OAI21_X1 U17632 ( .B1(n14212), .B2(n20061), .A(n14211), .ZN(n14217) );
  INV_X1 U17633 ( .A(n14213), .ZN(n14214) );
  NOR2_X1 U17634 ( .A1(n20107), .A2(n14272), .ZN(n14216) );
  AOI211_X1 U17635 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n20033), .A(n14217), .B(
        n14216), .ZN(n14218) );
  OAI21_X1 U17636 ( .B1(n14233), .B2(n14648), .A(n14218), .ZN(P1_U2832) );
  NOR2_X1 U17637 ( .A1(n19192), .A2(n14219), .ZN(n14258) );
  XNOR2_X1 U17638 ( .A(n14258), .B(n14427), .ZN(n14220) );
  NAND2_X1 U17639 ( .A1(n14220), .A2(n19174), .ZN(n14228) );
  OAI22_X1 U17640 ( .A1(n19188), .A2(n10411), .B1(n19951), .B2(n19203), .ZN(
        n14224) );
  NOR2_X1 U17641 ( .A1(n19201), .A2(n14222), .ZN(n14223) );
  AOI211_X1 U17642 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19213), .A(
        n14224), .B(n14223), .ZN(n14225) );
  OAI21_X1 U17643 ( .B1(n19885), .B2(n19204), .A(n14225), .ZN(n14226) );
  AOI21_X1 U17644 ( .B1(n14221), .B2(n19172), .A(n14226), .ZN(n14227) );
  OAI211_X1 U17645 ( .C1(n14229), .C2(n19953), .A(n14228), .B(n14227), .ZN(
        P2_U2853) );
  INV_X1 U17646 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14232) );
  INV_X1 U17647 ( .A(DATAI_8_), .ZN(n14231) );
  INV_X1 U17648 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n14230) );
  MUX2_X1 U17649 ( .A(n14231), .B(n14230), .S(n20259), .Z(n20145) );
  OAI222_X1 U17650 ( .A1(n14233), .A2(n14866), .B1(n14232), .B2(n14861), .C1(
        n14864), .C2(n20145), .ZN(P1_U2896) );
  XOR2_X1 U17651 ( .A(n13986), .B(n14234), .Z(n20109) );
  INV_X1 U17652 ( .A(n20109), .ZN(n14236) );
  OAI222_X1 U17653 ( .A1(n14864), .A2(n20306), .B1(n14866), .B2(n14236), .C1(
        n14235), .C2(n14861), .ZN(P1_U2898) );
  OR2_X1 U17654 ( .A1(n14172), .A2(n14238), .ZN(n14239) );
  NAND2_X1 U17655 ( .A1(n14237), .A2(n14239), .ZN(n20037) );
  INV_X1 U17656 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14240) );
  OAI222_X1 U17657 ( .A1(n20037), .A2(n14866), .B1(n14240), .B2(n14861), .C1(
        n14864), .C2(n14800), .ZN(P1_U2895) );
  AOI21_X1 U17658 ( .B1(n14242), .B2(n14241), .A(n14640), .ZN(n16271) );
  INV_X1 U17659 ( .A(n16271), .ZN(n20035) );
  OAI222_X1 U17660 ( .A1(n20037), .A2(n14753), .B1(n14243), .B2(n20115), .C1(
        n20035), .C2(n14769), .ZN(P1_U2863) );
  AOI21_X1 U17661 ( .B1(n14246), .B2(n14245), .A(n14244), .ZN(n16470) );
  INV_X1 U17662 ( .A(n16470), .ZN(n19108) );
  INV_X1 U17663 ( .A(n14247), .ZN(n14248) );
  OAI211_X1 U17664 ( .C1(n14166), .C2(n14249), .A(n14248), .B(n15212), .ZN(
        n14251) );
  NAND2_X1 U17665 ( .A1(n9750), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14250) );
  OAI211_X1 U17666 ( .C1(n19108), .C2(n9750), .A(n14251), .B(n14250), .ZN(
        P2_U2875) );
  OAI222_X1 U17667 ( .A1(n14864), .A2(n20316), .B1(n14861), .B2(n12102), .C1(
        n20052), .C2(n14866), .ZN(P1_U2897) );
  OAI211_X1 U17668 ( .C1(n14247), .C2(n14253), .A(n14252), .B(n15212), .ZN(
        n14257) );
  NOR2_X1 U17669 ( .A1(n14244), .A2(n14254), .ZN(n14255) );
  OR2_X1 U17670 ( .A1(n15207), .A2(n14255), .ZN(n15660) );
  INV_X1 U17671 ( .A(n15660), .ZN(n19094) );
  NAND2_X1 U17672 ( .A1(n15205), .A2(n19094), .ZN(n14256) );
  OAI211_X1 U17673 ( .C1(n15205), .C2(n10919), .A(n14257), .B(n14256), .ZN(
        P2_U2874) );
  OAI21_X1 U17674 ( .B1(n14260), .B2(n14259), .A(n14258), .ZN(n15098) );
  OAI21_X1 U17675 ( .B1(n9977), .B2(n14261), .A(n15098), .ZN(n15777) );
  AOI22_X1 U17676 ( .A1(n19192), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19198), .B2(n9977), .ZN(n15772) );
  NOR2_X1 U17677 ( .A1(n15772), .A2(n10456), .ZN(n15778) );
  INV_X1 U17678 ( .A(n16508), .ZN(n15780) );
  INV_X1 U17679 ( .A(n19953), .ZN(n14262) );
  AOI222_X1 U17680 ( .A1(n14263), .A2(n19941), .B1(n15777), .B2(n15778), .C1(
        n15780), .C2(n14262), .ZN(n14267) );
  AOI22_X1 U17681 ( .A1(n14264), .A2(n16503), .B1(P2_FLUSH_REG_SCAN_IN), .B2(
        n16507), .ZN(n14265) );
  OAI21_X1 U17682 ( .B1(n20000), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14265), 
        .ZN(n15789) );
  INV_X1 U17683 ( .A(n15789), .ZN(n15784) );
  NAND2_X1 U17684 ( .A1(n15784), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14266) );
  OAI21_X1 U17685 ( .B1(n14267), .B2(n15784), .A(n14266), .ZN(P2_U3599) );
  NOR2_X1 U17686 ( .A1(n9870), .A2(n14268), .ZN(n14269) );
  XNOR2_X1 U17687 ( .A(n14270), .B(n14269), .ZN(n16285) );
  INV_X1 U17688 ( .A(n16285), .ZN(n14276) );
  AOI22_X1 U17689 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14271) );
  OAI21_X1 U17690 ( .B1(n20179), .B2(n14272), .A(n14271), .ZN(n14273) );
  AOI21_X1 U17691 ( .B1(n14274), .B2(n20194), .A(n14273), .ZN(n14275) );
  OAI21_X1 U17692 ( .B1(n14276), .B2(n20198), .A(n14275), .ZN(P1_U2991) );
  NAND2_X1 U17693 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16172) );
  AOI22_X1 U17694 ( .A1(n16172), .A2(n14277), .B1(n12813), .B2(n20226), .ZN(
        n14279) );
  NAND2_X1 U17695 ( .A1(n15999), .A2(n14885), .ZN(n14278) );
  NAND2_X1 U17696 ( .A1(n14279), .A2(n14278), .ZN(n14280) );
  NOR2_X1 U17697 ( .A1(n14282), .A2(n16179), .ZN(n16173) );
  NAND2_X1 U17698 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n16173), .ZN(
        n14997) );
  INV_X1 U17699 ( .A(n16179), .ZN(n14283) );
  NAND2_X1 U17700 ( .A1(n14283), .A2(n20239), .ZN(n14998) );
  OAI211_X1 U17702 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n20239), .A(
        n14993), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14983) );
  AND3_X1 U17703 ( .A1(n14983), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14998), .ZN(n14287) );
  INV_X1 U17704 ( .A(n14284), .ZN(n16186) );
  NOR2_X1 U17705 ( .A1(n14885), .A2(n16186), .ZN(n16175) );
  NAND2_X1 U17706 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16175), .ZN(
        n14989) );
  INV_X1 U17707 ( .A(n14989), .ZN(n16163) );
  INV_X1 U17708 ( .A(n14988), .ZN(n15002) );
  NAND3_X1 U17709 ( .A1(n16163), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15002), .ZN(n14980) );
  NOR3_X1 U17710 ( .A1(n14980), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12789), .ZN(n14286) );
  NOR3_X1 U17711 ( .A1(n14287), .A2(n14286), .A3(n14285), .ZN(n14312) );
  NAND2_X1 U17712 ( .A1(n9815), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14289) );
  NAND2_X1 U17713 ( .A1(n14307), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14288) );
  NAND2_X1 U17714 ( .A1(n14289), .A2(n14288), .ZN(n14456) );
  NAND2_X1 U17715 ( .A1(n14296), .A2(n16083), .ZN(n14292) );
  INV_X1 U17716 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14709) );
  NAND2_X1 U17717 ( .A1(n9818), .A2(n14709), .ZN(n14290) );
  NAND3_X1 U17718 ( .A1(n14292), .A2(n14291), .A3(n14290), .ZN(n14293) );
  OAI21_X1 U17719 ( .B1(n14306), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14293), .ZN(
        n14705) );
  MUX2_X1 U17720 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14294) );
  OAI21_X1 U17721 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n9815), .A(
        n14294), .ZN(n14515) );
  INV_X1 U17722 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14701) );
  NAND2_X1 U17723 ( .A1(n14295), .A2(n14701), .ZN(n14300) );
  NAND2_X1 U17724 ( .A1(n14296), .A2(n9809), .ZN(n14298) );
  NAND2_X1 U17725 ( .A1(n9818), .A2(n14701), .ZN(n14297) );
  NAND3_X1 U17726 ( .A1(n14298), .A2(n14291), .A3(n14297), .ZN(n14299) );
  AND2_X1 U17727 ( .A1(n14300), .A2(n14299), .ZN(n14492) );
  MUX2_X1 U17728 ( .A(n14301), .B(n14291), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14302) );
  OAI21_X1 U17729 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n9815), .A(
        n14302), .ZN(n14485) );
  OR2_X1 U17730 ( .A1(n9815), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14305) );
  INV_X1 U17731 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14303) );
  NAND2_X1 U17732 ( .A1(n14305), .A2(n14304), .ZN(n14452) );
  OAI22_X1 U17733 ( .A1(n14452), .A2(n9817), .B1(P1_EBX_REG_29__SCAN_IN), .B2(
        n14306), .ZN(n14468) );
  AOI22_X1 U17734 ( .A1(n9815), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14307), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14309) );
  XNOR2_X2 U17735 ( .A(n14310), .B(n14309), .ZN(n14695) );
  NAND2_X1 U17736 ( .A1(n14695), .A2(n20238), .ZN(n14311) );
  OAI211_X1 U17737 ( .C1(n14313), .C2(n16291), .A(n14312), .B(n14311), .ZN(
        P1_U3000) );
  OAI21_X1 U17738 ( .B1(n14316), .B2(n14315), .A(n14314), .ZN(n14331) );
  INV_X1 U17739 ( .A(n14317), .ZN(n14318) );
  XNOR2_X1 U17740 ( .A(n15240), .B(n14318), .ZN(n16376) );
  INV_X1 U17741 ( .A(n16376), .ZN(n14320) );
  OAI22_X1 U17742 ( .A1(n15276), .A2(n14320), .B1(n19249), .B2(n14319), .ZN(
        n14324) );
  INV_X1 U17743 ( .A(n19222), .ZN(n15278) );
  INV_X1 U17744 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n14322) );
  INV_X1 U17745 ( .A(n19221), .ZN(n15224) );
  OAI22_X1 U17746 ( .A1(n15278), .A2(n14322), .B1(n14321), .B2(n15224), .ZN(
        n14323) );
  AOI211_X1 U17747 ( .C1(n19223), .C2(BUF1_REG_25__SCAN_IN), .A(n14324), .B(
        n14323), .ZN(n14325) );
  OAI21_X1 U17748 ( .B1(n14331), .B2(n15282), .A(n14325), .ZN(P2_U2894) );
  NOR2_X1 U17749 ( .A1(n14326), .A2(n14327), .ZN(n14328) );
  OR2_X1 U17750 ( .A1(n15125), .A2(n14328), .ZN(n16380) );
  MUX2_X1 U17751 ( .A(n16380), .B(n14329), .S(n9769), .Z(n14330) );
  OAI21_X1 U17752 ( .B1(n14331), .B2(n15178), .A(n14330), .ZN(P2_U2862) );
  NOR2_X1 U17753 ( .A1(n14332), .A2(n11342), .ZN(n14333) );
  INV_X1 U17754 ( .A(n15293), .ZN(n14335) );
  NOR2_X1 U17755 ( .A1(n14338), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14339) );
  MUX2_X1 U17756 ( .A(n14340), .B(n14339), .S(n10904), .Z(n16328) );
  NAND2_X1 U17757 ( .A1(n16328), .A2(n10137), .ZN(n14341) );
  XNOR2_X1 U17758 ( .A(n14341), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14342) );
  XNOR2_X1 U17759 ( .A(n14343), .B(n14342), .ZN(n14371) );
  NAND2_X1 U17760 ( .A1(n15298), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14344) );
  NAND2_X1 U17762 ( .A1(n14357), .A2(n19300), .ZN(n14356) );
  AOI22_X1 U17763 ( .A1(n10511), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14348) );
  NAND2_X1 U17764 ( .A1(n14346), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14347) );
  OAI211_X1 U17765 ( .C1(n14349), .C2(n14363), .A(n14348), .B(n14347), .ZN(
        n14350) );
  XNOR2_X1 U17766 ( .A(n14351), .B(n14350), .ZN(n16336) );
  INV_X1 U17767 ( .A(n16336), .ZN(n15099) );
  NAND2_X1 U17768 ( .A1(n15730), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14365) );
  NAND2_X1 U17769 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14352) );
  OAI211_X1 U17770 ( .C1(n19294), .C2(n14353), .A(n14365), .B(n14352), .ZN(
        n14354) );
  AOI21_X1 U17771 ( .B1(n15099), .B2(n19302), .A(n14354), .ZN(n14355) );
  OAI211_X1 U17772 ( .C1(n14371), .C2(n19305), .A(n14356), .B(n14355), .ZN(
        P2_U2983) );
  NAND2_X1 U17773 ( .A1(n14357), .A2(n19319), .ZN(n14370) );
  OAI21_X1 U17774 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15616), .A(
        n14358), .ZN(n14359) );
  INV_X1 U17775 ( .A(n14359), .ZN(n14367) );
  AOI222_X1 U17776 ( .A1(n14361), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14360), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10657), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14362) );
  OAI211_X1 U17777 ( .C1(n14367), .C2(n14363), .A(n10195), .B(n14366), .ZN(
        n14368) );
  INV_X1 U17778 ( .A(n14368), .ZN(n14369) );
  OAI211_X1 U17779 ( .C1(n14371), .C2(n15761), .A(n14370), .B(n14369), .ZN(
        P2_U3015) );
  OAI21_X1 U17780 ( .B1(n14372), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20003), 
        .ZN(n14373) );
  OAI21_X1 U17781 ( .B1(n19991), .B2(n20003), .A(n14373), .ZN(P2_U3612) );
  NAND2_X1 U17782 ( .A1(n14375), .A2(n14374), .ZN(n14377) );
  INV_X1 U17783 ( .A(n14377), .ZN(n14379) );
  XNOR2_X1 U17784 ( .A(n14380), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14381) );
  INV_X1 U17785 ( .A(n15497), .ZN(n14382) );
  NAND2_X1 U17786 ( .A1(n15481), .A2(n15479), .ZN(n15492) );
  NAND2_X1 U17787 ( .A1(n14382), .A2(n15492), .ZN(n15486) );
  AND2_X1 U17788 ( .A1(n9841), .A2(n14383), .ZN(n14384) );
  INV_X1 U17789 ( .A(n14415), .ZN(n14385) );
  AOI21_X1 U17790 ( .B1(n14386), .B2(n13436), .A(n14385), .ZN(n16356) );
  NAND2_X1 U17791 ( .A1(n15730), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14400) );
  OAI21_X1 U17792 ( .B1(n14387), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14400), .ZN(n14388) );
  AOI21_X1 U17793 ( .B1(n16356), .B2(n19326), .A(n14388), .ZN(n14389) );
  OAI21_X1 U17794 ( .B1(n16358), .B2(n19317), .A(n14389), .ZN(n14392) );
  OR2_X1 U17795 ( .A1(n15306), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14390) );
  NOR2_X1 U17796 ( .A1(n14402), .A2(n16496), .ZN(n14391) );
  OAI21_X1 U17797 ( .B1(n14405), .B2(n15761), .A(n14393), .ZN(P2_U3018) );
  NAND2_X1 U17798 ( .A1(n14861), .A2(n9777), .ZN(n14396) );
  INV_X1 U17799 ( .A(n14396), .ZN(n14395) );
  NAND2_X1 U17800 ( .A1(n14395), .A2(n20259), .ZN(n14782) );
  INV_X1 U17801 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16560) );
  NAND3_X1 U17802 ( .A1(n14439), .A2(n11828), .A3(n14861), .ZN(n14399) );
  AOI22_X1 U17803 ( .A1(n14397), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14847), .ZN(n14398) );
  OAI211_X1 U17804 ( .C1(n14782), .C2(n16560), .A(n14399), .B(n14398), .ZN(
        P1_U2873) );
  INV_X1 U17805 ( .A(n16358), .ZN(n14404) );
  NAND2_X1 U17806 ( .A1(n16453), .A2(n10206), .ZN(n14401) );
  OAI211_X1 U17807 ( .C1(n16462), .C2(n9973), .A(n14401), .B(n14400), .ZN(
        n14403) );
  NOR2_X1 U17808 ( .A1(n11028), .A2(n9750), .ZN(n14406) );
  AOI21_X1 U17809 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n9769), .A(n14406), .ZN(
        n14407) );
  OAI21_X1 U17810 ( .B1(n14408), .B2(n15178), .A(n14407), .ZN(P2_U2857) );
  NAND2_X1 U17811 ( .A1(n14411), .A2(n14410), .ZN(n15105) );
  NAND2_X1 U17812 ( .A1(n15105), .A2(n19225), .ZN(n14421) );
  AOI22_X1 U17813 ( .A1(n19222), .A2(BUF2_REG_29__SCAN_IN), .B1(n19221), .B2(
        n14412), .ZN(n14420) );
  INV_X1 U17814 ( .A(n14413), .ZN(n14417) );
  NAND2_X1 U17815 ( .A1(n14415), .A2(n14414), .ZN(n14416) );
  NAND2_X1 U17816 ( .A1(n14417), .A2(n14416), .ZN(n16340) );
  OAI22_X1 U17817 ( .A1(n16340), .A2(n15276), .B1(n19249), .B2(n21179), .ZN(
        n14418) );
  AOI21_X1 U17818 ( .B1(n19223), .B2(BUF1_REG_29__SCAN_IN), .A(n14418), .ZN(
        n14419) );
  OAI211_X1 U17819 ( .C1(n14409), .C2(n14421), .A(n14420), .B(n14419), .ZN(
        P2_U2890) );
  NAND2_X1 U17820 ( .A1(n14423), .A2(n14422), .ZN(n14424) );
  AND2_X1 U17821 ( .A1(n14425), .A2(n14424), .ZN(n19315) );
  INV_X1 U17822 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14426) );
  NAND2_X1 U17823 ( .A1(n15730), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19321) );
  OAI21_X1 U17824 ( .B1(n16462), .B2(n14426), .A(n19321), .ZN(n14429) );
  NOR2_X1 U17825 ( .A1(n19294), .A2(n14427), .ZN(n14428) );
  AOI211_X1 U17826 ( .C1(n19315), .C2(n19283), .A(n14429), .B(n14428), .ZN(
        n14434) );
  INV_X1 U17827 ( .A(n14430), .ZN(n14431) );
  XNOR2_X1 U17828 ( .A(n14432), .B(n14431), .ZN(n19318) );
  NAND2_X1 U17829 ( .A1(n19318), .A2(n19300), .ZN(n14433) );
  OAI211_X1 U17830 ( .C1(n19289), .C2(n13670), .A(n14434), .B(n14433), .ZN(
        P2_U3012) );
  NAND2_X1 U17831 ( .A1(n14435), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14438)
         );
  INV_X1 U17832 ( .A(n14436), .ZN(n20015) );
  NAND3_X1 U17833 ( .A1(n14438), .A2(n20015), .A3(n14437), .ZN(P1_U2801) );
  INV_X1 U17834 ( .A(n14439), .ZN(n14449) );
  INV_X1 U17835 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20944) );
  INV_X1 U17836 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14441) );
  NAND3_X1 U17837 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n14440), .A3(n20041), 
        .ZN(n14643) );
  NOR2_X1 U17838 ( .A1(n14441), .A2(n14643), .ZN(n14638) );
  NAND3_X1 U17839 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(n14638), .ZN(n14627) );
  NAND2_X1 U17840 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14599) );
  NOR2_X1 U17841 ( .A1(n14627), .A2(n14599), .ZN(n14600) );
  NAND4_X1 U17842 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14600), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U17843 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14571) );
  NOR2_X1 U17844 ( .A1(n14570), .A2(n14571), .ZN(n14540) );
  INV_X1 U17845 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21230) );
  NAND2_X1 U17846 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14543) );
  NOR2_X1 U17847 ( .A1(n21230), .A2(n14543), .ZN(n16027) );
  AND3_X1 U17848 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14540), .A3(n16027), 
        .ZN(n14525) );
  AND2_X1 U17849 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14525), .ZN(n16020) );
  NAND2_X1 U17850 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n16020), .ZN(n14513) );
  NOR2_X1 U17851 ( .A1(n20944), .A2(n14513), .ZN(n14499) );
  NAND2_X1 U17852 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14499), .ZN(n14484) );
  NOR2_X1 U17853 ( .A1(n20948), .A2(n14484), .ZN(n14473) );
  NAND2_X1 U17854 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14473), .ZN(n14443) );
  INV_X1 U17855 ( .A(n14443), .ZN(n14458) );
  NAND2_X1 U17856 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n14458), .ZN(n14442) );
  INV_X1 U17857 ( .A(n14636), .ZN(n14679) );
  AOI21_X1 U17858 ( .B1(n16021), .B2(n14442), .A(n14679), .ZN(n14463) );
  NOR4_X1 U17859 ( .A1(n20101), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14443), 
        .A4(n21043), .ZN(n14444) );
  AOI21_X1 U17860 ( .B1(n20051), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14444), .ZN(n14446) );
  NAND2_X1 U17861 ( .A1(n20071), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14445) );
  OAI211_X1 U17862 ( .C1(n14463), .C2(n20951), .A(n14446), .B(n14445), .ZN(
        n14447) );
  OAI21_X1 U17863 ( .B1(n14449), .B2(n14648), .A(n14448), .ZN(P1_U2809) );
  INV_X1 U17864 ( .A(n14450), .ZN(n14777) );
  NAND2_X1 U17865 ( .A1(n14451), .A2(n9817), .ZN(n14453) );
  NAND2_X1 U17866 ( .A1(n14453), .A2(n14452), .ZN(n14455) );
  OR2_X1 U17867 ( .A1(n14487), .A2(n9817), .ZN(n14454) );
  NAND2_X1 U17868 ( .A1(n14455), .A2(n14454), .ZN(n14457) );
  AOI21_X1 U17869 ( .B1(n16021), .B2(n14458), .A(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14462) );
  NAND2_X1 U17870 ( .A1(n20039), .A2(n14459), .ZN(n14461) );
  AOI22_X1 U17871 ( .A1(n20071), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20051), .ZN(n14460) );
  OAI211_X1 U17872 ( .C1(n14463), .C2(n14462), .A(n14461), .B(n14460), .ZN(
        n14464) );
  AOI21_X1 U17873 ( .B1(n14984), .B2(n20099), .A(n14464), .ZN(n14465) );
  OAI21_X1 U17874 ( .B1(n14777), .B2(n14648), .A(n14465), .ZN(P1_U2810) );
  AOI21_X1 U17875 ( .B1(n14467), .B2(n9844), .A(n14466), .ZN(n14873) );
  INV_X1 U17876 ( .A(n14873), .ZN(n14785) );
  INV_X1 U17877 ( .A(n14468), .ZN(n14469) );
  XNOR2_X1 U17878 ( .A(n14487), .B(n14469), .ZN(n14992) );
  INV_X1 U17879 ( .A(n14871), .ZN(n14470) );
  NAND2_X1 U17880 ( .A1(n20039), .A2(n14470), .ZN(n14477) );
  INV_X1 U17881 ( .A(n14473), .ZN(n14471) );
  NOR2_X1 U17882 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14471), .ZN(n14472) );
  AOI22_X1 U17883 ( .A1(n16021), .A2(n14472), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20051), .ZN(n14476) );
  OR2_X1 U17884 ( .A1(n20101), .A2(n14473), .ZN(n14483) );
  NAND2_X1 U17885 ( .A1(n14483), .A2(n14636), .ZN(n14480) );
  NAND2_X1 U17886 ( .A1(n14480), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14475) );
  NAND2_X1 U17887 ( .A1(n20071), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14474) );
  NAND4_X1 U17888 ( .A1(n14477), .A2(n14476), .A3(n14475), .A4(n14474), .ZN(
        n14478) );
  AOI21_X1 U17889 ( .B1(n14992), .B2(n20099), .A(n14478), .ZN(n14479) );
  OAI21_X1 U17890 ( .B1(n14785), .B2(n14648), .A(n14479), .ZN(P1_U2811) );
  NAND2_X1 U17891 ( .A1(n14480), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U17892 ( .A1(n20071), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20051), .ZN(n14481) );
  OAI211_X1 U17893 ( .C1(n14484), .C2(n14483), .A(n14482), .B(n14481), .ZN(
        n14489) );
  AND2_X1 U17894 ( .A1(n14494), .A2(n14485), .ZN(n14486) );
  NOR2_X1 U17895 ( .A1(n14999), .A2(n20061), .ZN(n14488) );
  AOI211_X1 U17896 ( .C1(n20039), .C2(n14490), .A(n14489), .B(n14488), .ZN(
        n14491) );
  OAI21_X1 U17897 ( .B1(n14790), .B2(n14648), .A(n14491), .ZN(P1_U2812) );
  NAND2_X1 U17898 ( .A1(n14517), .A2(n14492), .ZN(n14493) );
  NAND2_X1 U17899 ( .A1(n14494), .A2(n14493), .ZN(n16169) );
  AOI21_X1 U17900 ( .B1(n14496), .B2(n14495), .A(n13044), .ZN(n14882) );
  NAND2_X1 U17901 ( .A1(n14882), .A2(n20066), .ZN(n14505) );
  INV_X1 U17902 ( .A(n14880), .ZN(n14503) );
  INV_X1 U17903 ( .A(n14499), .ZN(n14497) );
  NOR2_X1 U17904 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14497), .ZN(n14498) );
  AOI22_X1 U17905 ( .A1(n16021), .A2(n14498), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20051), .ZN(n14501) );
  OR2_X1 U17906 ( .A1(n20101), .A2(n14499), .ZN(n14512) );
  NAND2_X1 U17907 ( .A1(n14512), .A2(n14636), .ZN(n14509) );
  NAND2_X1 U17908 ( .A1(n14509), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14500) );
  OAI211_X1 U17909 ( .C1(n14701), .C2(n20094), .A(n14501), .B(n14500), .ZN(
        n14502) );
  AOI21_X1 U17910 ( .B1(n20039), .B2(n14503), .A(n14502), .ZN(n14504) );
  OAI211_X1 U17911 ( .C1(n16169), .C2(n20061), .A(n14505), .B(n14504), .ZN(
        P1_U2813) );
  OAI21_X1 U17912 ( .B1(n14507), .B2(n14508), .A(n14495), .ZN(n14894) );
  NAND2_X1 U17913 ( .A1(n14509), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U17914 ( .A1(n20071), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20051), .ZN(n14510) );
  OAI211_X1 U17915 ( .C1(n14513), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14514) );
  AOI21_X1 U17916 ( .B1(n20039), .B2(n14891), .A(n14514), .ZN(n14519) );
  NAND2_X1 U17917 ( .A1(n14708), .A2(n14515), .ZN(n14516) );
  AND2_X1 U17918 ( .A1(n14517), .A2(n14516), .ZN(n16170) );
  NAND2_X1 U17919 ( .A1(n16170), .A2(n20099), .ZN(n14518) );
  OAI211_X1 U17920 ( .C1(n14894), .C2(n14648), .A(n14519), .B(n14518), .ZN(
        P1_U2814) );
  OR2_X1 U17921 ( .A1(n14520), .A2(n14714), .ZN(n14716) );
  AOI21_X1 U17922 ( .B1(n14523), .B2(n14716), .A(n14522), .ZN(n14899) );
  INV_X1 U17923 ( .A(n14899), .ZN(n14807) );
  NOR2_X1 U17924 ( .A1(n20101), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U17925 ( .A1(n16019), .A2(n14525), .B1(n20071), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14524) );
  OAI21_X1 U17926 ( .B1(n12435), .B2(n20093), .A(n14524), .ZN(n14529) );
  OR2_X1 U17927 ( .A1(n20101), .A2(n14525), .ZN(n14526) );
  NAND2_X1 U17928 ( .A1(n14526), .A2(n14636), .ZN(n16018) );
  INV_X1 U17929 ( .A(n16018), .ZN(n16032) );
  INV_X1 U17930 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14527) );
  OAI22_X1 U17931 ( .A1(n14712), .A2(n20061), .B1(n16032), .B2(n14527), .ZN(
        n14528) );
  AOI211_X1 U17932 ( .C1(n20039), .C2(n14895), .A(n14529), .B(n14528), .ZN(
        n14530) );
  OAI21_X1 U17933 ( .B1(n14807), .B2(n14648), .A(n14530), .ZN(P1_U2816) );
  INV_X1 U17934 ( .A(n14531), .ZN(n14906) );
  INV_X1 U17935 ( .A(n14520), .ZN(n14533) );
  AOI21_X1 U17936 ( .B1(n14534), .B2(n14532), .A(n14533), .ZN(n14908) );
  NAND2_X1 U17937 ( .A1(n14908), .A2(n20066), .ZN(n14549) );
  NOR2_X1 U17938 ( .A1(n14729), .A2(n14535), .ZN(n14536) );
  OR2_X1 U17939 ( .A1(n14718), .A2(n14536), .ZN(n14724) );
  INV_X1 U17940 ( .A(n14724), .ZN(n16192) );
  INV_X1 U17941 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14725) );
  NAND2_X1 U17942 ( .A1(n14540), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16033) );
  INV_X1 U17943 ( .A(n16033), .ZN(n14537) );
  NAND2_X1 U17944 ( .A1(n14636), .A2(n14537), .ZN(n14538) );
  NAND2_X1 U17945 ( .A1(n14685), .A2(n14538), .ZN(n16034) );
  OAI21_X1 U17946 ( .B1(n20101), .B2(P1_REIP_REG_21__SCAN_IN), .A(n16034), 
        .ZN(n14539) );
  NAND2_X1 U17947 ( .A1(n14539), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14546) );
  INV_X1 U17948 ( .A(n14540), .ZN(n14541) );
  NOR2_X1 U17949 ( .A1(n20101), .A2(n14541), .ZN(n16026) );
  NAND2_X1 U17950 ( .A1(n16026), .A2(n21230), .ZN(n14542) );
  NOR2_X1 U17951 ( .A1(n14543), .A2(n14542), .ZN(n14544) );
  AOI21_X1 U17952 ( .B1(n20051), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14544), .ZN(n14545) );
  OAI211_X1 U17953 ( .C1(n14725), .C2(n20094), .A(n14546), .B(n14545), .ZN(
        n14547) );
  AOI21_X1 U17954 ( .B1(n16192), .B2(n20099), .A(n14547), .ZN(n14548) );
  OAI211_X1 U17955 ( .C1(n14906), .C2(n20107), .A(n14549), .B(n14548), .ZN(
        P1_U2818) );
  AOI21_X1 U17956 ( .B1(n14552), .B2(n10168), .A(n14551), .ZN(n14553) );
  INV_X1 U17957 ( .A(n14553), .ZN(n14919) );
  NAND2_X1 U17958 ( .A1(n14566), .A2(n14554), .ZN(n14555) );
  AND2_X1 U17959 ( .A1(n9874), .A2(n14555), .ZN(n16000) );
  INV_X1 U17960 ( .A(n16000), .ZN(n14559) );
  AOI22_X1 U17961 ( .A1(n20071), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n20051), 
        .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14558) );
  INV_X1 U17962 ( .A(n16034), .ZN(n14556) );
  OAI21_X1 U17963 ( .B1(n16026), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14556), 
        .ZN(n14557) );
  OAI211_X1 U17964 ( .C1(n14559), .C2(n20061), .A(n14558), .B(n14557), .ZN(
        n14560) );
  AOI21_X1 U17965 ( .B1(n20039), .B2(n14916), .A(n14560), .ZN(n14561) );
  OAI21_X1 U17966 ( .B1(n14919), .B2(n14648), .A(n14561), .ZN(P1_U2820) );
  AOI21_X1 U17967 ( .B1(n14563), .B2(n14562), .A(n14550), .ZN(n16105) );
  INV_X1 U17968 ( .A(n16105), .ZN(n14827) );
  INV_X1 U17969 ( .A(n16108), .ZN(n14576) );
  OR2_X1 U17970 ( .A1(n14580), .A2(n14564), .ZN(n14565) );
  NAND2_X1 U17971 ( .A1(n14566), .A2(n14565), .ZN(n16204) );
  INV_X1 U17972 ( .A(n14570), .ZN(n14567) );
  OR2_X1 U17973 ( .A1(n20101), .A2(n14567), .ZN(n14568) );
  NAND2_X1 U17974 ( .A1(n14568), .A2(n14636), .ZN(n16048) );
  AOI22_X1 U17975 ( .A1(n16048), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n20071), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n14569) );
  OAI21_X1 U17976 ( .B1(n16204), .B2(n20061), .A(n14569), .ZN(n14575) );
  INV_X1 U17977 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14573) );
  NOR2_X1 U17978 ( .A1(n20101), .A2(n14570), .ZN(n14582) );
  OAI211_X1 U17979 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14582), .B(n14571), .ZN(n14572) );
  OAI211_X1 U17980 ( .C1(n20093), .C2(n14573), .A(n14572), .B(n20091), .ZN(
        n14574) );
  AOI211_X1 U17981 ( .C1(n20039), .C2(n14576), .A(n14575), .B(n14574), .ZN(
        n14577) );
  OAI21_X1 U17982 ( .B1(n14827), .B2(n14648), .A(n14577), .ZN(P1_U2821) );
  XOR2_X1 U17983 ( .A(n14579), .B(n14578), .Z(n14926) );
  INV_X1 U17984 ( .A(n14926), .ZN(n14831) );
  AOI21_X1 U17985 ( .B1(n14581), .B2(n14748), .A(n14580), .ZN(n16211) );
  INV_X1 U17986 ( .A(n16211), .ZN(n14588) );
  INV_X1 U17987 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20932) );
  NAND2_X1 U17988 ( .A1(n14582), .A2(n20932), .ZN(n14584) );
  AOI21_X1 U17989 ( .B1(n20051), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20050), .ZN(n14583) );
  OAI211_X1 U17990 ( .C1(n14585), .C2(n20094), .A(n14584), .B(n14583), .ZN(
        n14586) );
  AOI21_X1 U17991 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n16048), .A(n14586), 
        .ZN(n14587) );
  OAI21_X1 U17992 ( .B1(n14588), .B2(n20061), .A(n14587), .ZN(n14589) );
  AOI21_X1 U17993 ( .B1(n14922), .B2(n20039), .A(n14589), .ZN(n14590) );
  OAI21_X1 U17994 ( .B1(n14831), .B2(n14648), .A(n14590), .ZN(P1_U2822) );
  AOI21_X1 U17995 ( .B1(n14594), .B2(n14592), .A(n14593), .ZN(n14938) );
  INV_X1 U17996 ( .A(n14938), .ZN(n14841) );
  NAND2_X1 U17997 ( .A1(n14759), .A2(n14595), .ZN(n14596) );
  AND2_X1 U17998 ( .A1(n14746), .A2(n14596), .ZN(n16225) );
  INV_X1 U17999 ( .A(n16225), .ZN(n14751) );
  AOI21_X1 U18000 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20051), .A(
        n20050), .ZN(n14597) );
  OAI21_X1 U18001 ( .B1(n14751), .B2(n20061), .A(n14597), .ZN(n14604) );
  INV_X1 U18002 ( .A(n14627), .ZN(n14598) );
  NAND2_X1 U18003 ( .A1(n16021), .A2(n14598), .ZN(n14626) );
  OR2_X1 U18004 ( .A1(n14626), .A2(n14599), .ZN(n16054) );
  NAND2_X1 U18005 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n16047) );
  OAI21_X1 U18006 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n16047), .ZN(n14602) );
  OAI21_X1 U18007 ( .B1(n20101), .B2(n14600), .A(n14636), .ZN(n16057) );
  AOI22_X1 U18008 ( .A1(n16057), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n20071), 
        .B2(P1_EBX_REG_16__SCAN_IN), .ZN(n14601) );
  OAI21_X1 U18009 ( .B1(n16054), .B2(n14602), .A(n14601), .ZN(n14603) );
  AOI211_X1 U18010 ( .C1(n20039), .C2(n14934), .A(n14604), .B(n14603), .ZN(
        n14605) );
  OAI21_X1 U18011 ( .B1(n14841), .B2(n14648), .A(n14605), .ZN(P1_U2824) );
  INV_X1 U18012 ( .A(n14606), .ZN(n14610) );
  INV_X1 U18013 ( .A(n14607), .ZN(n14623) );
  NAND2_X1 U18014 ( .A1(n14951), .A2(n20066), .ZN(n14618) );
  INV_X1 U18015 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20923) );
  INV_X1 U18016 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20924) );
  OAI21_X1 U18017 ( .B1(n20923), .B2(n14626), .A(n20924), .ZN(n14616) );
  INV_X1 U18018 ( .A(n14629), .ZN(n14611) );
  AOI21_X1 U18019 ( .B1(n14612), .B2(n14611), .A(n14757), .ZN(n16243) );
  INV_X1 U18020 ( .A(n16243), .ZN(n14762) );
  NOR2_X1 U18021 ( .A1(n14762), .A2(n20061), .ZN(n14615) );
  NAND2_X1 U18022 ( .A1(n20071), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n14613) );
  OAI211_X1 U18023 ( .C1(n20093), .C2(n21015), .A(n14613), .B(n20091), .ZN(
        n14614) );
  AOI211_X1 U18024 ( .C1(n14616), .C2(n16057), .A(n14615), .B(n14614), .ZN(
        n14617) );
  OAI211_X1 U18025 ( .C1(n20107), .C2(n14949), .A(n14618), .B(n14617), .ZN(
        P1_U2826) );
  NAND2_X1 U18026 ( .A1(n14634), .A2(n14621), .ZN(n14622) );
  NAND2_X1 U18027 ( .A1(n14619), .A2(n14622), .ZN(n14857) );
  OAI21_X1 U18028 ( .B1(n14857), .B2(n14858), .A(n14619), .ZN(n14850) );
  AOI22_X1 U18029 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n20051), .B1(
        n20071), .B2(P1_EBX_REG_13__SCAN_IN), .ZN(n14625) );
  OAI211_X1 U18030 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n14626), .A(n14625), 
        .B(n20091), .ZN(n14632) );
  OAI21_X1 U18031 ( .B1(n14679), .B2(n14627), .A(n14685), .ZN(n16066) );
  AND2_X1 U18032 ( .A1(n15014), .A2(n14628), .ZN(n14630) );
  OR2_X1 U18033 ( .A1(n14630), .A2(n14629), .ZN(n16254) );
  OAI22_X1 U18034 ( .A1(n16066), .A2(n20923), .B1(n20061), .B2(n16254), .ZN(
        n14631) );
  AOI211_X1 U18035 ( .C1(n14963), .C2(n20039), .A(n14632), .B(n14631), .ZN(
        n14633) );
  OAI21_X1 U18036 ( .B1(n14966), .B2(n14648), .A(n14633), .ZN(P1_U2827) );
  AOI21_X1 U18037 ( .B1(n14635), .B2(n14237), .A(n14620), .ZN(n14972) );
  NAND2_X1 U18038 ( .A1(n14972), .A2(n20066), .ZN(n14647) );
  OAI21_X1 U18039 ( .B1(n20101), .B2(n14638), .A(n14636), .ZN(n16070) );
  INV_X1 U18040 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14637) );
  OAI21_X1 U18041 ( .B1(n20093), .B2(n14637), .A(n20091), .ZN(n14645) );
  INV_X1 U18042 ( .A(n14638), .ZN(n16060) );
  NAND2_X1 U18043 ( .A1(n16021), .A2(n16060), .ZN(n14642) );
  OAI21_X1 U18044 ( .B1(n14640), .B2(n14639), .A(n16068), .ZN(n14770) );
  INV_X1 U18045 ( .A(n14770), .ZN(n16265) );
  AOI22_X1 U18046 ( .A1(n16265), .A2(n20099), .B1(n20071), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14641) );
  OAI21_X1 U18047 ( .B1(n14643), .B2(n14642), .A(n14641), .ZN(n14644) );
  AOI211_X1 U18048 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n16070), .A(n14645), 
        .B(n14644), .ZN(n14646) );
  OAI211_X1 U18049 ( .C1(n20107), .C2(n14970), .A(n14647), .B(n14646), .ZN(
        P1_U2830) );
  INV_X1 U18050 ( .A(n14659), .ZN(n14649) );
  OAI21_X1 U18051 ( .B1(n14650), .B2(n14649), .A(n14648), .ZN(n20104) );
  NAND2_X1 U18052 ( .A1(n20104), .A2(n14651), .ZN(n14664) );
  NAND2_X1 U18053 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n14668) );
  AOI21_X1 U18054 ( .B1(n16021), .B2(n14668), .A(n14679), .ZN(n14656) );
  INV_X1 U18055 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14655) );
  AOI22_X1 U18056 ( .A1(n20071), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20051), .ZN(n14654) );
  INV_X1 U18057 ( .A(n14668), .ZN(n14652) );
  NAND3_X1 U18058 ( .A1(n16021), .A2(n14652), .A3(n14655), .ZN(n14653) );
  OAI211_X1 U18059 ( .C1(n14656), .C2(n14655), .A(n14654), .B(n14653), .ZN(
        n14662) );
  INV_X1 U18060 ( .A(n20549), .ZN(n14660) );
  INV_X1 U18061 ( .A(n14657), .ZN(n14658) );
  NAND2_X1 U18062 ( .A1(n14659), .A2(n14658), .ZN(n20095) );
  NOR2_X1 U18063 ( .A1(n14660), .A2(n20095), .ZN(n14661) );
  AOI211_X1 U18064 ( .C1(n20099), .C2(n20210), .A(n14662), .B(n14661), .ZN(
        n14663) );
  OAI211_X1 U18065 ( .C1(n20107), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        P1_U2837) );
  NAND2_X1 U18066 ( .A1(n20104), .A2(n14666), .ZN(n14675) );
  INV_X1 U18067 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20908) );
  INV_X1 U18068 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20966) );
  NAND2_X1 U18069 ( .A1(n20908), .A2(n20966), .ZN(n14667) );
  NAND2_X1 U18070 ( .A1(n14668), .A2(n14667), .ZN(n14671) );
  NAND2_X1 U18071 ( .A1(n20071), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14670) );
  AOI22_X1 U18072 ( .A1(n20051), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n14679), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14669) );
  OAI211_X1 U18073 ( .C1(n14671), .C2(n20101), .A(n14670), .B(n14669), .ZN(
        n14673) );
  NOR2_X1 U18074 ( .A1(n20690), .A2(n20095), .ZN(n14672) );
  AOI211_X1 U18075 ( .C1(n20220), .C2(n20099), .A(n14673), .B(n14672), .ZN(
        n14674) );
  OAI211_X1 U18076 ( .C1(n20107), .C2(n14676), .A(n14675), .B(n14674), .ZN(
        P1_U2838) );
  INV_X1 U18077 ( .A(n20104), .ZN(n14694) );
  INV_X1 U18078 ( .A(n20095), .ZN(n14690) );
  INV_X1 U18079 ( .A(n20550), .ZN(n20791) );
  AOI22_X1 U18080 ( .A1(n20099), .A2(n14678), .B1(n20071), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U18081 ( .A1(n20051), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14679), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14680) );
  OAI211_X1 U18082 ( .C1(P1_REIP_REG_1__SCAN_IN), .C2(n20101), .A(n14681), .B(
        n14680), .ZN(n14683) );
  NOR2_X1 U18083 ( .A1(n20107), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14682) );
  AOI211_X1 U18084 ( .C1(n14690), .C2(n20791), .A(n14683), .B(n14682), .ZN(
        n14684) );
  OAI21_X1 U18085 ( .B1(n14694), .B2(n20189), .A(n14684), .ZN(P1_U2839) );
  INV_X1 U18086 ( .A(n14685), .ZN(n20046) );
  NOR2_X1 U18087 ( .A1(n20046), .A2(n13803), .ZN(n14689) );
  OAI22_X1 U18088 ( .A1(n20061), .A2(n14687), .B1(n20094), .B2(n14686), .ZN(
        n14688) );
  AOI211_X1 U18089 ( .C1(n14690), .C2(n9785), .A(n14689), .B(n14688), .ZN(
        n14692) );
  OAI21_X1 U18090 ( .B1(n20039), .B2(n20051), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14691) );
  OAI211_X1 U18091 ( .C1(n14694), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        P1_U2840) );
  INV_X1 U18092 ( .A(n14695), .ZN(n14697) );
  INV_X1 U18093 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14696) );
  OAI22_X1 U18094 ( .A1(n14697), .A2(n14769), .B1(n20115), .B2(n14696), .ZN(
        P1_U2841) );
  AOI22_X1 U18095 ( .A1(n14984), .A2(n20112), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14740), .ZN(n14698) );
  OAI21_X1 U18096 ( .B1(n14777), .B2(n14767), .A(n14698), .ZN(P1_U2842) );
  AOI22_X1 U18097 ( .A1(n14992), .A2(n20112), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14740), .ZN(n14699) );
  OAI21_X1 U18098 ( .B1(n14785), .B2(n14753), .A(n14699), .ZN(P1_U2843) );
  INV_X1 U18099 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14700) );
  OAI222_X1 U18100 ( .A1(n14767), .A2(n14790), .B1(n14700), .B2(n20115), .C1(
        n14999), .C2(n14769), .ZN(P1_U2844) );
  INV_X1 U18101 ( .A(n14882), .ZN(n14795) );
  OAI222_X1 U18102 ( .A1(n16169), .A2(n14769), .B1(n14701), .B2(n20115), .C1(
        n14795), .C2(n14767), .ZN(P1_U2845) );
  AOI22_X1 U18103 ( .A1(n16170), .A2(n20112), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14740), .ZN(n14702) );
  OAI21_X1 U18104 ( .B1(n14894), .B2(n14767), .A(n14702), .ZN(P1_U2846) );
  NOR2_X1 U18105 ( .A1(n14522), .A2(n14703), .ZN(n14704) );
  OR2_X1 U18106 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  NAND2_X1 U18107 ( .A1(n14708), .A2(n14707), .ZN(n16183) );
  OAI22_X1 U18108 ( .A1(n16183), .A2(n14769), .B1(n14709), .B2(n20115), .ZN(
        n14710) );
  INV_X1 U18109 ( .A(n14710), .ZN(n14711) );
  OAI21_X1 U18110 ( .B1(n16016), .B2(n14767), .A(n14711), .ZN(P1_U2847) );
  INV_X1 U18111 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14713) );
  OAI222_X1 U18112 ( .A1(n14767), .A2(n14807), .B1(n14713), .B2(n20115), .C1(
        n14712), .C2(n14769), .ZN(P1_U2848) );
  NAND2_X1 U18113 ( .A1(n14520), .A2(n14714), .ZN(n14715) );
  OR2_X1 U18114 ( .A1(n14718), .A2(n14717), .ZN(n14719) );
  NAND2_X1 U18115 ( .A1(n14720), .A2(n14719), .ZN(n16190) );
  OAI22_X1 U18116 ( .A1(n16190), .A2(n14769), .B1(n14721), .B2(n20115), .ZN(
        n14722) );
  INV_X1 U18117 ( .A(n14722), .ZN(n14723) );
  OAI21_X1 U18118 ( .B1(n14811), .B2(n14767), .A(n14723), .ZN(P1_U2849) );
  INV_X1 U18119 ( .A(n14908), .ZN(n14815) );
  OAI222_X1 U18120 ( .A1(n14753), .A2(n14815), .B1(n14725), .B2(n20115), .C1(
        n14724), .C2(n14769), .ZN(P1_U2850) );
  OR2_X1 U18121 ( .A1(n14551), .A2(n14726), .ZN(n14727) );
  AND2_X1 U18122 ( .A1(n14532), .A2(n14727), .ZN(n16097) );
  INV_X1 U18123 ( .A(n16097), .ZN(n14820) );
  AND2_X1 U18124 ( .A1(n9874), .A2(n14728), .ZN(n14730) );
  OR2_X1 U18125 ( .A1(n14730), .A2(n14729), .ZN(n16039) );
  OAI22_X1 U18126 ( .A1(n16039), .A2(n14769), .B1(n14731), .B2(n20115), .ZN(
        n14732) );
  INV_X1 U18127 ( .A(n14732), .ZN(n14733) );
  OAI21_X1 U18128 ( .B1(n14820), .B2(n14767), .A(n14733), .ZN(P1_U2851) );
  NOR2_X1 U18129 ( .A1(n20115), .A2(n14734), .ZN(n14735) );
  AOI21_X1 U18130 ( .B1(n16000), .B2(n20112), .A(n14735), .ZN(n14736) );
  OAI21_X1 U18131 ( .B1(n14919), .B2(n14767), .A(n14736), .ZN(P1_U2852) );
  OAI22_X1 U18132 ( .A1(n16204), .A2(n14769), .B1(n14737), .B2(n20115), .ZN(
        n14738) );
  INV_X1 U18133 ( .A(n14738), .ZN(n14739) );
  OAI21_X1 U18134 ( .B1(n14827), .B2(n14767), .A(n14739), .ZN(P1_U2853) );
  AOI22_X1 U18135 ( .A1(n16211), .A2(n20112), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n14740), .ZN(n14741) );
  OAI21_X1 U18136 ( .B1(n14831), .B2(n14753), .A(n14741), .ZN(P1_U2854) );
  INV_X1 U18137 ( .A(n14742), .ZN(n14744) );
  INV_X1 U18138 ( .A(n14593), .ZN(n14743) );
  AOI21_X1 U18139 ( .B1(n14744), .B2(n14743), .A(n14578), .ZN(n16115) );
  INV_X1 U18140 ( .A(n16115), .ZN(n14835) );
  NAND2_X1 U18141 ( .A1(n14746), .A2(n14745), .ZN(n14747) );
  NAND2_X1 U18142 ( .A1(n14748), .A2(n14747), .ZN(n16217) );
  OAI22_X1 U18143 ( .A1(n16217), .A2(n14769), .B1(n16045), .B2(n20115), .ZN(
        n14749) );
  INV_X1 U18144 ( .A(n14749), .ZN(n14750) );
  OAI21_X1 U18145 ( .B1(n14835), .B2(n14767), .A(n14750), .ZN(P1_U2855) );
  INV_X1 U18146 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14752) );
  OAI222_X1 U18147 ( .A1(n14841), .A2(n14753), .B1(n14752), .B2(n20115), .C1(
        n14751), .C2(n14769), .ZN(P1_U2856) );
  INV_X1 U18148 ( .A(n14592), .ZN(n14754) );
  AOI21_X1 U18149 ( .B1(n14755), .B2(n14609), .A(n14754), .ZN(n16125) );
  INV_X1 U18150 ( .A(n14767), .ZN(n20113) );
  OR2_X1 U18151 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  NAND2_X1 U18152 ( .A1(n14759), .A2(n14758), .ZN(n16231) );
  OAI22_X1 U18153 ( .A1(n16231), .A2(n14769), .B1(n16053), .B2(n20115), .ZN(
        n14760) );
  AOI21_X1 U18154 ( .B1(n16125), .B2(n20113), .A(n14760), .ZN(n14761) );
  INV_X1 U18155 ( .A(n14761), .ZN(P1_U2857) );
  INV_X1 U18156 ( .A(n14951), .ZN(n14846) );
  INV_X1 U18157 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14763) );
  OAI222_X1 U18158 ( .A1(n14846), .A2(n14767), .B1(n20115), .B2(n14763), .C1(
        n14762), .C2(n14769), .ZN(P1_U2858) );
  OAI22_X1 U18159 ( .A1(n16254), .A2(n14769), .B1(n14764), .B2(n20115), .ZN(
        n14765) );
  INV_X1 U18160 ( .A(n14765), .ZN(n14766) );
  OAI21_X1 U18161 ( .B1(n14966), .B2(n14767), .A(n14766), .ZN(P1_U2859) );
  INV_X1 U18162 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14768) );
  INV_X1 U18163 ( .A(n14972), .ZN(n14865) );
  OAI222_X1 U18164 ( .A1(n14770), .A2(n14769), .B1(n14768), .B2(n20115), .C1(
        n14865), .C2(n14767), .ZN(P1_U2862) );
  NAND3_X1 U18165 ( .A1(n14861), .A2(n11767), .A3(n11827), .ZN(n14836) );
  INV_X1 U18166 ( .A(DATAI_14_), .ZN(n14772) );
  INV_X1 U18167 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14771) );
  MUX2_X1 U18168 ( .A(n14772), .B(n14771), .S(n20259), .Z(n20153) );
  OAI22_X1 U18169 ( .A1(n14836), .A2(n20153), .B1(n14861), .B2(n14773), .ZN(
        n14774) );
  AOI21_X1 U18170 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14838), .A(n14774), .ZN(
        n14776) );
  NAND2_X1 U18171 ( .A1(n14397), .A2(DATAI_30_), .ZN(n14775) );
  OAI211_X1 U18172 ( .C1(n14777), .C2(n14866), .A(n14776), .B(n14775), .ZN(
        P1_U2874) );
  INV_X1 U18173 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16564) );
  INV_X1 U18174 ( .A(n14836), .ZN(n14780) );
  INV_X1 U18175 ( .A(DATAI_13_), .ZN(n14779) );
  NAND2_X1 U18176 ( .A1(n20259), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14778) );
  OAI21_X1 U18177 ( .B1(n20259), .B2(n14779), .A(n14778), .ZN(n20151) );
  AOI22_X1 U18178 ( .A1(n14780), .A2(n20151), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n14847), .ZN(n14781) );
  OAI21_X1 U18179 ( .B1(n16564), .B2(n14782), .A(n14781), .ZN(n14783) );
  AOI21_X1 U18180 ( .B1(n14397), .B2(DATAI_29_), .A(n14783), .ZN(n14784) );
  OAI21_X1 U18181 ( .B1(n14785), .B2(n14866), .A(n14784), .ZN(P1_U2875) );
  INV_X1 U18182 ( .A(DATAI_12_), .ZN(n14786) );
  INV_X1 U18183 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16589) );
  MUX2_X1 U18184 ( .A(n14786), .B(n16589), .S(n20259), .Z(n20148) );
  OAI22_X1 U18185 ( .A1(n14836), .A2(n20148), .B1(n14861), .B2(n13710), .ZN(
        n14787) );
  AOI21_X1 U18186 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14838), .A(n14787), .ZN(
        n14789) );
  NAND2_X1 U18187 ( .A1(n14397), .A2(DATAI_28_), .ZN(n14788) );
  OAI211_X1 U18188 ( .C1(n14790), .C2(n14866), .A(n14789), .B(n14788), .ZN(
        P1_U2876) );
  OAI22_X1 U18189 ( .A1(n14836), .A2(n14859), .B1(n14861), .B2(n14791), .ZN(
        n14792) );
  AOI21_X1 U18190 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14838), .A(n14792), .ZN(
        n14794) );
  NAND2_X1 U18191 ( .A1(n14397), .A2(DATAI_27_), .ZN(n14793) );
  OAI211_X1 U18192 ( .C1(n14795), .C2(n14866), .A(n14794), .B(n14793), .ZN(
        P1_U2877) );
  OAI22_X1 U18193 ( .A1(n14836), .A2(n14863), .B1(n14861), .B2(n14796), .ZN(
        n14797) );
  AOI21_X1 U18194 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14838), .A(n14797), .ZN(
        n14799) );
  NAND2_X1 U18195 ( .A1(n14397), .A2(DATAI_26_), .ZN(n14798) );
  OAI211_X1 U18196 ( .C1(n14894), .C2(n14866), .A(n14799), .B(n14798), .ZN(
        P1_U2878) );
  OAI22_X1 U18197 ( .A1(n14836), .A2(n14800), .B1(n14861), .B2(n21190), .ZN(
        n14801) );
  AOI21_X1 U18198 ( .B1(n14838), .B2(BUF1_REG_25__SCAN_IN), .A(n14801), .ZN(
        n14803) );
  NAND2_X1 U18199 ( .A1(n14397), .A2(DATAI_25_), .ZN(n14802) );
  OAI211_X1 U18200 ( .C1(n16016), .C2(n14866), .A(n14803), .B(n14802), .ZN(
        P1_U2879) );
  OAI22_X1 U18201 ( .A1(n14836), .A2(n20145), .B1(n14861), .B2(n13705), .ZN(
        n14804) );
  AOI21_X1 U18202 ( .B1(n14838), .B2(BUF1_REG_24__SCAN_IN), .A(n14804), .ZN(
        n14806) );
  NAND2_X1 U18203 ( .A1(n14397), .A2(DATAI_24_), .ZN(n14805) );
  OAI211_X1 U18204 ( .C1(n14807), .C2(n14866), .A(n14806), .B(n14805), .ZN(
        P1_U2880) );
  OAI22_X1 U18205 ( .A1(n14836), .A2(n20316), .B1(n14861), .B2(n13941), .ZN(
        n14808) );
  AOI21_X1 U18206 ( .B1(n14838), .B2(BUF1_REG_23__SCAN_IN), .A(n14808), .ZN(
        n14810) );
  NAND2_X1 U18207 ( .A1(n14397), .A2(DATAI_23_), .ZN(n14809) );
  OAI211_X1 U18208 ( .C1(n14811), .C2(n14866), .A(n14810), .B(n14809), .ZN(
        P1_U2881) );
  OAI22_X1 U18209 ( .A1(n14836), .A2(n20306), .B1(n14861), .B2(n13939), .ZN(
        n14812) );
  AOI21_X1 U18210 ( .B1(n14838), .B2(BUF1_REG_22__SCAN_IN), .A(n14812), .ZN(
        n14814) );
  NAND2_X1 U18211 ( .A1(n14397), .A2(DATAI_22_), .ZN(n14813) );
  OAI211_X1 U18212 ( .C1(n14815), .C2(n14866), .A(n14814), .B(n14813), .ZN(
        P1_U2882) );
  OAI22_X1 U18213 ( .A1(n14836), .A2(n20297), .B1(n14861), .B2(n14816), .ZN(
        n14817) );
  AOI21_X1 U18214 ( .B1(n14838), .B2(BUF1_REG_21__SCAN_IN), .A(n14817), .ZN(
        n14819) );
  NAND2_X1 U18215 ( .A1(n14397), .A2(DATAI_21_), .ZN(n14818) );
  OAI211_X1 U18216 ( .C1(n14820), .C2(n14866), .A(n14819), .B(n14818), .ZN(
        P1_U2883) );
  OAI22_X1 U18217 ( .A1(n14836), .A2(n20292), .B1(n14861), .B2(n13947), .ZN(
        n14821) );
  AOI21_X1 U18218 ( .B1(n14838), .B2(BUF1_REG_20__SCAN_IN), .A(n14821), .ZN(
        n14823) );
  NAND2_X1 U18219 ( .A1(n14397), .A2(DATAI_20_), .ZN(n14822) );
  OAI211_X1 U18220 ( .C1(n14919), .C2(n14866), .A(n14823), .B(n14822), .ZN(
        P1_U2884) );
  OAI22_X1 U18221 ( .A1(n14836), .A2(n20286), .B1(n14861), .B2(n13945), .ZN(
        n14824) );
  AOI21_X1 U18222 ( .B1(n14838), .B2(BUF1_REG_19__SCAN_IN), .A(n14824), .ZN(
        n14826) );
  NAND2_X1 U18223 ( .A1(n14397), .A2(DATAI_19_), .ZN(n14825) );
  OAI211_X1 U18224 ( .C1(n14827), .C2(n14866), .A(n14826), .B(n14825), .ZN(
        P1_U2885) );
  OAI22_X1 U18225 ( .A1(n14836), .A2(n20280), .B1(n14861), .B2(n13943), .ZN(
        n14828) );
  AOI21_X1 U18226 ( .B1(n14838), .B2(BUF1_REG_18__SCAN_IN), .A(n14828), .ZN(
        n14830) );
  NAND2_X1 U18227 ( .A1(n14397), .A2(DATAI_18_), .ZN(n14829) );
  OAI211_X1 U18228 ( .C1(n14831), .C2(n14866), .A(n14830), .B(n14829), .ZN(
        P1_U2886) );
  OAI22_X1 U18229 ( .A1(n14836), .A2(n20274), .B1(n14861), .B2(n13951), .ZN(
        n14832) );
  AOI21_X1 U18230 ( .B1(n14838), .B2(BUF1_REG_17__SCAN_IN), .A(n14832), .ZN(
        n14834) );
  NAND2_X1 U18231 ( .A1(n14397), .A2(DATAI_17_), .ZN(n14833) );
  OAI211_X1 U18232 ( .C1(n14835), .C2(n14866), .A(n14834), .B(n14833), .ZN(
        P1_U2887) );
  OAI22_X1 U18233 ( .A1(n14836), .A2(n20264), .B1(n14861), .B2(n13937), .ZN(
        n14837) );
  AOI21_X1 U18234 ( .B1(n14838), .B2(BUF1_REG_16__SCAN_IN), .A(n14837), .ZN(
        n14840) );
  NAND2_X1 U18235 ( .A1(n14397), .A2(DATAI_16_), .ZN(n14839) );
  OAI211_X1 U18236 ( .C1(n14841), .C2(n14866), .A(n14840), .B(n14839), .ZN(
        P1_U2888) );
  INV_X1 U18237 ( .A(n16125), .ZN(n14844) );
  OAI222_X1 U18238 ( .A1(n14866), .A2(n14844), .B1(n14861), .B2(n14843), .C1(
        n14864), .C2(n14842), .ZN(P1_U2889) );
  INV_X1 U18239 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14845) );
  OAI222_X1 U18240 ( .A1(n14846), .A2(n14866), .B1(n14845), .B2(n14861), .C1(
        n14864), .C2(n20153), .ZN(P1_U2890) );
  INV_X1 U18241 ( .A(n14864), .ZN(n14848) );
  AOI22_X1 U18242 ( .A1(n14848), .A2(n20151), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14847), .ZN(n14849) );
  OAI21_X1 U18243 ( .B1(n14966), .B2(n14866), .A(n14849), .ZN(P1_U2891) );
  INV_X1 U18244 ( .A(n14850), .ZN(n14854) );
  INV_X1 U18245 ( .A(n14851), .ZN(n14853) );
  INV_X1 U18246 ( .A(n16128), .ZN(n14856) );
  OAI222_X1 U18247 ( .A1(n14856), .A2(n14866), .B1(n14855), .B2(n14861), .C1(
        n14864), .C2(n20148), .ZN(P1_U2892) );
  INV_X1 U18248 ( .A(n16139), .ZN(n14860) );
  OAI222_X1 U18249 ( .A1(n14866), .A2(n14860), .B1(n14861), .B2(n21189), .C1(
        n14864), .C2(n14859), .ZN(P1_U2893) );
  INV_X1 U18250 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14862) );
  OAI222_X1 U18251 ( .A1(n14866), .A2(n14865), .B1(n14864), .B2(n14863), .C1(
        n14862), .C2(n14861), .ZN(P1_U2894) );
  INV_X1 U18252 ( .A(n14867), .ZN(n14868) );
  INV_X1 U18253 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21143) );
  NOR2_X1 U18254 ( .A1(n16230), .A2(n21143), .ZN(n14991) );
  AOI21_X1 U18255 ( .B1(n20180), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14991), .ZN(n14870) );
  OAI21_X1 U18256 ( .B1(n14871), .B2(n20179), .A(n14870), .ZN(n14872) );
  AOI21_X1 U18257 ( .B1(n14873), .B2(n20194), .A(n14872), .ZN(n14874) );
  OAI21_X1 U18258 ( .B1(n9847), .B2(n20198), .A(n14874), .ZN(P1_U2970) );
  INV_X1 U18259 ( .A(n14875), .ZN(n14876) );
  NOR2_X1 U18260 ( .A1(n14876), .A2(n12786), .ZN(n14877) );
  MUX2_X1 U18261 ( .A(n14877), .B(n9842), .S(n16121), .Z(n14878) );
  AOI22_X1 U18262 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n14879) );
  OAI21_X1 U18263 ( .B1(n14880), .B2(n20179), .A(n14879), .ZN(n14881) );
  AOI21_X1 U18264 ( .B1(n14882), .B2(n20194), .A(n14881), .ZN(n14883) );
  OAI21_X1 U18265 ( .B1(n16162), .B2(n20198), .A(n14883), .ZN(P1_U2972) );
  OAI21_X1 U18266 ( .B1(n14884), .B2(n14885), .A(n16134), .ZN(n14886) );
  NAND2_X1 U18267 ( .A1(n9779), .A2(n14886), .ZN(n14888) );
  XNOR2_X1 U18268 ( .A(n14888), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16171) );
  NAND2_X1 U18269 ( .A1(n16171), .A2(n20186), .ZN(n14893) );
  OAI22_X1 U18270 ( .A1(n20190), .A2(n14889), .B1(n16230), .B2(n20944), .ZN(
        n14890) );
  AOI21_X1 U18271 ( .B1(n14891), .B2(n20185), .A(n14890), .ZN(n14892) );
  OAI211_X1 U18272 ( .C1(n20258), .C2(n14894), .A(n14893), .B(n14892), .ZN(
        P1_U2973) );
  INV_X1 U18273 ( .A(n14895), .ZN(n14897) );
  AOI22_X1 U18274 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n14896) );
  OAI21_X1 U18275 ( .B1(n20179), .B2(n14897), .A(n14896), .ZN(n14898) );
  AOI21_X1 U18276 ( .B1(n14899), .B2(n20194), .A(n14898), .ZN(n14900) );
  OAI21_X1 U18277 ( .B1(n14901), .B2(n20198), .A(n14900), .ZN(P1_U2975) );
  NAND2_X1 U18278 ( .A1(n14903), .A2(n14902), .ZN(n14904) );
  XNOR2_X1 U18279 ( .A(n14904), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16193) );
  INV_X1 U18280 ( .A(n16193), .ZN(n14910) );
  AOI22_X1 U18281 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14905) );
  OAI21_X1 U18282 ( .B1(n20179), .B2(n14906), .A(n14905), .ZN(n14907) );
  AOI21_X1 U18283 ( .B1(n14908), .B2(n20194), .A(n14907), .ZN(n14909) );
  OAI21_X1 U18284 ( .B1(n20198), .B2(n14910), .A(n14909), .ZN(P1_U2977) );
  OAI21_X1 U18285 ( .B1(n16134), .B2(n16208), .A(n14920), .ZN(n16104) );
  NOR3_X1 U18286 ( .A1(n16104), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16134), .ZN(n14913) );
  NAND2_X1 U18287 ( .A1(n16134), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14912) );
  NOR2_X1 U18288 ( .A1(n14920), .A2(n14912), .ZN(n15978) );
  NOR2_X1 U18289 ( .A1(n14913), .A2(n15978), .ZN(n15976) );
  XNOR2_X1 U18290 ( .A(n15976), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16001) );
  NAND2_X1 U18291 ( .A1(n16001), .A2(n20186), .ZN(n14918) );
  NAND2_X1 U18292 ( .A1(n20236), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16002) );
  OAI21_X1 U18293 ( .B1(n20190), .B2(n14914), .A(n16002), .ZN(n14915) );
  AOI21_X1 U18294 ( .B1(n20185), .B2(n14916), .A(n14915), .ZN(n14917) );
  OAI211_X1 U18295 ( .C1(n20258), .C2(n14919), .A(n14918), .B(n14917), .ZN(
        P1_U2979) );
  OAI21_X1 U18296 ( .B1(n9776), .B2(n14921), .A(n14920), .ZN(n16209) );
  INV_X1 U18297 ( .A(n14922), .ZN(n14924) );
  AOI22_X1 U18298 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14923) );
  OAI21_X1 U18299 ( .B1(n14924), .B2(n20179), .A(n14923), .ZN(n14925) );
  AOI21_X1 U18300 ( .B1(n14926), .B2(n20194), .A(n14925), .ZN(n14927) );
  OAI21_X1 U18301 ( .B1(n16209), .B2(n20198), .A(n14927), .ZN(P1_U2981) );
  INV_X1 U18302 ( .A(n14928), .ZN(n14930) );
  INV_X1 U18303 ( .A(n16133), .ZN(n14942) );
  AOI21_X1 U18304 ( .B1(n14930), .B2(n14942), .A(n14941), .ZN(n16119) );
  AOI21_X1 U18305 ( .B1(n16119), .B2(n14931), .A(n16120), .ZN(n14933) );
  XNOR2_X1 U18306 ( .A(n14933), .B(n14932), .ZN(n16226) );
  INV_X1 U18307 ( .A(n16226), .ZN(n14940) );
  INV_X1 U18308 ( .A(n14934), .ZN(n14936) );
  AOI22_X1 U18309 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14935) );
  OAI21_X1 U18310 ( .B1(n20179), .B2(n14936), .A(n14935), .ZN(n14937) );
  AOI21_X1 U18311 ( .B1(n14938), .B2(n20194), .A(n14937), .ZN(n14939) );
  OAI21_X1 U18312 ( .B1(n14940), .B2(n20198), .A(n14939), .ZN(P1_U2983) );
  OAI21_X1 U18313 ( .B1(n14942), .B2(n14941), .A(n9876), .ZN(n14944) );
  NAND2_X1 U18314 ( .A1(n14944), .A2(n14943), .ZN(n14947) );
  MUX2_X1 U18315 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n14945), .S(
        n16121), .Z(n14946) );
  XNOR2_X1 U18316 ( .A(n14947), .B(n14946), .ZN(n16242) );
  AOI22_X1 U18317 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14948) );
  OAI21_X1 U18318 ( .B1(n20179), .B2(n14949), .A(n14948), .ZN(n14950) );
  AOI21_X1 U18319 ( .B1(n14951), .B2(n20194), .A(n14950), .ZN(n14952) );
  OAI21_X1 U18320 ( .B1(n16242), .B2(n20198), .A(n14952), .ZN(P1_U2985) );
  OAI21_X1 U18321 ( .B1(n16133), .B2(n14954), .A(n14953), .ZN(n15011) );
  INV_X1 U18322 ( .A(n14958), .ZN(n14955) );
  NAND2_X1 U18323 ( .A1(n14956), .A2(n14955), .ZN(n15012) );
  NOR2_X1 U18324 ( .A1(n15011), .A2(n15012), .ZN(n14957) );
  NOR2_X1 U18325 ( .A1(n14958), .A2(n14957), .ZN(n14960) );
  XNOR2_X1 U18326 ( .A(n14960), .B(n14959), .ZN(n16252) );
  NAND2_X1 U18327 ( .A1(n16252), .A2(n20186), .ZN(n14965) );
  INV_X1 U18328 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14961) );
  OAI22_X1 U18329 ( .A1(n20190), .A2(n14961), .B1(n16230), .B2(n20923), .ZN(
        n14962) );
  AOI21_X1 U18330 ( .B1(n20185), .B2(n14963), .A(n14962), .ZN(n14964) );
  OAI211_X1 U18331 ( .C1(n20258), .C2(n14966), .A(n14965), .B(n14964), .ZN(
        P1_U2986) );
  MUX2_X1 U18332 ( .A(n16133), .B(n14967), .S(n16121), .Z(n14968) );
  XNOR2_X1 U18333 ( .A(n14968), .B(n12778), .ZN(n16266) );
  AOI22_X1 U18334 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14969) );
  OAI21_X1 U18335 ( .B1(n20179), .B2(n14970), .A(n14969), .ZN(n14971) );
  AOI21_X1 U18336 ( .B1(n14972), .B2(n20194), .A(n14971), .ZN(n14973) );
  OAI21_X1 U18337 ( .B1(n16266), .B2(n20198), .A(n14973), .ZN(P1_U2989) );
  XNOR2_X1 U18338 ( .A(n12771), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14975) );
  XNOR2_X1 U18339 ( .A(n14974), .B(n14975), .ZN(n16272) );
  AOI22_X1 U18340 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14977) );
  NAND2_X1 U18341 ( .A1(n20185), .A2(n20038), .ZN(n14976) );
  OAI211_X1 U18342 ( .C1(n20037), .C2(n20258), .A(n14977), .B(n14976), .ZN(
        n14978) );
  AOI21_X1 U18343 ( .B1(n16272), .B2(n20186), .A(n14978), .ZN(n14979) );
  INV_X1 U18344 ( .A(n14979), .ZN(P1_U2990) );
  NAND2_X1 U18345 ( .A1(n12789), .A2(n14980), .ZN(n14982) );
  AOI21_X1 U18346 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(n14986) );
  NAND2_X1 U18347 ( .A1(n14984), .A2(n20238), .ZN(n14985) );
  OAI211_X1 U18348 ( .C1(n14987), .C2(n16291), .A(n14986), .B(n14985), .ZN(
        P1_U3001) );
  NOR3_X1 U18349 ( .A1(n14989), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14988), .ZN(n14990) );
  AOI211_X1 U18350 ( .C1(n20238), .C2(n14992), .A(n14991), .B(n14990), .ZN(
        n14996) );
  INV_X1 U18351 ( .A(n14993), .ZN(n14994) );
  NAND2_X1 U18352 ( .A1(n14994), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14995) );
  OAI211_X1 U18353 ( .C1(n9847), .C2(n16291), .A(n14996), .B(n14995), .ZN(
        P1_U3002) );
  NAND2_X1 U18354 ( .A1(n14998), .A2(n14997), .ZN(n16166) );
  INV_X1 U18355 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15007) );
  INV_X1 U18356 ( .A(n14999), .ZN(n15001) );
  AOI21_X1 U18357 ( .B1(n15001), .B2(n20238), .A(n15000), .ZN(n15006) );
  NOR2_X1 U18358 ( .A1(n15003), .A2(n15002), .ZN(n15004) );
  NAND2_X1 U18359 ( .A1(n16163), .A2(n15004), .ZN(n15005) );
  OAI211_X1 U18360 ( .C1(n16166), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        n15008) );
  AOI21_X1 U18361 ( .B1(n15009), .B2(n20243), .A(n15008), .ZN(n15010) );
  INV_X1 U18362 ( .A(n15010), .ZN(P1_U3003) );
  XOR2_X1 U18363 ( .A(n15012), .B(n15011), .Z(n16132) );
  OAI21_X1 U18364 ( .B1(n16068), .B2(n16069), .A(n15013), .ZN(n15015) );
  AND2_X1 U18365 ( .A1(n15015), .A2(n15014), .ZN(n16075) );
  AND2_X1 U18366 ( .A1(n20236), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15025) );
  AND2_X1 U18367 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16238), .ZN(
        n15020) );
  AND2_X1 U18368 ( .A1(n16281), .A2(n15020), .ZN(n15017) );
  AOI21_X1 U18369 ( .B1(n20219), .B2(n15016), .A(n20218), .ZN(n16206) );
  OAI21_X1 U18370 ( .B1(n15017), .B2(n20205), .A(n16206), .ZN(n16256) );
  AOI21_X1 U18371 ( .B1(n20217), .B2(n16137), .A(n16256), .ZN(n15023) );
  INV_X1 U18372 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15022) );
  INV_X1 U18373 ( .A(n16280), .ZN(n15018) );
  AOI22_X1 U18374 ( .A1(n20226), .A2(n20223), .B1(n15018), .B2(n20217), .ZN(
        n20216) );
  NOR2_X1 U18375 ( .A1(n20216), .A2(n15019), .ZN(n16302) );
  NAND3_X1 U18376 ( .A1(n15020), .A2(n16302), .A3(n15022), .ZN(n15021) );
  OAI21_X1 U18377 ( .B1(n15023), .B2(n15022), .A(n15021), .ZN(n15024) );
  AOI211_X1 U18378 ( .C1(n20238), .C2(n16075), .A(n15025), .B(n15024), .ZN(
        n15026) );
  OAI21_X1 U18379 ( .B1(n16132), .B2(n16291), .A(n15026), .ZN(P1_U3019) );
  OAI21_X1 U18380 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13831), .A(n20825), 
        .ZN(n15027) );
  OAI21_X1 U18381 ( .B1(n15028), .B2(n20550), .A(n15027), .ZN(n15029) );
  MUX2_X1 U18382 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15029), .S(
        n20249), .Z(P1_U3477) );
  NOR3_X1 U18383 ( .A1(n15030), .A2(n13621), .A3(n11708), .ZN(n15033) );
  NOR2_X1 U18384 ( .A1(n20550), .A2(n15031), .ZN(n15032) );
  AOI211_X1 U18385 ( .C1(n15940), .C2(n10119), .A(n15033), .B(n15032), .ZN(
        n15938) );
  INV_X1 U18386 ( .A(n15034), .ZN(n15035) );
  NAND2_X1 U18387 ( .A1(n15036), .A2(n15035), .ZN(n15041) );
  INV_X1 U18388 ( .A(n11708), .ZN(n15039) );
  NAND3_X1 U18389 ( .A1(n15039), .A2(n15038), .A3(n15037), .ZN(n15040) );
  OAI211_X1 U18390 ( .C1(n15938), .C2(n16312), .A(n15041), .B(n15040), .ZN(
        n15042) );
  MUX2_X1 U18391 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15042), .S(
        n16316), .Z(P1_U3473) );
  AOI211_X1 U18392 ( .C1(n15349), .C2(n15044), .A(n15043), .B(n19216), .ZN(
        n15046) );
  OAI22_X1 U18393 ( .A1(n15347), .A2(n19178), .B1(n19913), .B2(n19204), .ZN(
        n15045) );
  AOI211_X1 U18394 ( .C1(P2_EBX_REG_23__SCAN_IN), .C2(n19207), .A(n15046), .B(
        n15045), .ZN(n15055) );
  NAND2_X1 U18395 ( .A1(n15047), .A2(n15048), .ZN(n15049) );
  NAND2_X1 U18396 ( .A1(n15134), .A2(n15049), .ZN(n15534) );
  OR2_X1 U18397 ( .A1(n15067), .A2(n15051), .ZN(n15052) );
  NAND2_X1 U18398 ( .A1(n15050), .A2(n15052), .ZN(n15539) );
  OAI22_X1 U18399 ( .A1(n15534), .A2(n19209), .B1(n15539), .B2(n19203), .ZN(
        n15053) );
  INV_X1 U18400 ( .A(n15053), .ZN(n15054) );
  OAI211_X1 U18401 ( .C1(n15056), .C2(n19201), .A(n15055), .B(n15054), .ZN(
        P2_U2832) );
  INV_X1 U18402 ( .A(n15057), .ZN(n15071) );
  NOR2_X1 U18403 ( .A1(n19192), .A2(n15058), .ZN(n15059) );
  XOR2_X1 U18404 ( .A(n15362), .B(n15059), .Z(n15061) );
  AOI22_X1 U18405 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19167), .ZN(n15060) );
  OAI21_X1 U18406 ( .B1(n19216), .B2(n15061), .A(n15060), .ZN(n15062) );
  AOI21_X1 U18407 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n19207), .A(n15062), .ZN(
        n15070) );
  OR2_X1 U18408 ( .A1(n15079), .A2(n15063), .ZN(n15064) );
  NAND2_X1 U18409 ( .A1(n15047), .A2(n15064), .ZN(n15552) );
  INV_X1 U18410 ( .A(n15552), .ZN(n15068) );
  AND2_X1 U18411 ( .A1(n15083), .A2(n15065), .ZN(n15066) );
  NOR2_X1 U18412 ( .A1(n15067), .A2(n15066), .ZN(n16392) );
  AOI22_X1 U18413 ( .A1(n15068), .A2(n19172), .B1(n16392), .B2(n19182), .ZN(
        n15069) );
  OAI211_X1 U18414 ( .C1(n15071), .C2(n19201), .A(n15070), .B(n15069), .ZN(
        P2_U2833) );
  NAND2_X1 U18415 ( .A1(n9977), .A2(n15072), .ZN(n15073) );
  INV_X1 U18416 ( .A(n15073), .ZN(n19013) );
  INV_X1 U18417 ( .A(n15384), .ZN(n15074) );
  AOI221_X1 U18418 ( .B1(n15384), .B2(n19013), .C1(n15074), .C2(n15073), .A(
        n19216), .ZN(n15076) );
  OAI22_X1 U18419 ( .A1(n15382), .A2(n19178), .B1(n19910), .B2(n19204), .ZN(
        n15075) );
  AOI211_X1 U18420 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n19207), .A(n15076), .B(
        n15075), .ZN(n15088) );
  INV_X1 U18421 ( .A(n19201), .ZN(n19185) );
  NOR2_X1 U18422 ( .A1(n10218), .A2(n15077), .ZN(n15078) );
  OR2_X1 U18423 ( .A1(n15079), .A2(n15078), .ZN(n15559) );
  NAND2_X1 U18424 ( .A1(n15080), .A2(n15081), .ZN(n15082) );
  AND2_X1 U18425 ( .A1(n15083), .A2(n15082), .ZN(n15562) );
  INV_X1 U18426 ( .A(n15562), .ZN(n15084) );
  OAI22_X1 U18427 ( .A1(n15559), .A2(n19209), .B1(n15084), .B2(n19203), .ZN(
        n15085) );
  AOI21_X1 U18428 ( .B1(n15086), .B2(n19185), .A(n15085), .ZN(n15087) );
  NAND2_X1 U18429 ( .A1(n15088), .A2(n15087), .ZN(P2_U2834) );
  OAI22_X1 U18430 ( .A1(n19201), .A2(n15089), .B1(n19091), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15090) );
  AOI21_X1 U18431 ( .B1(n19182), .B2(n19966), .A(n15090), .ZN(n15091) );
  OAI21_X1 U18432 ( .B1(n15092), .B2(n19209), .A(n15091), .ZN(n15096) );
  AOI22_X1 U18433 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19167), .ZN(n15093) );
  OAI21_X1 U18434 ( .B1(n19188), .B2(n15094), .A(n15093), .ZN(n15095) );
  AOI211_X1 U18435 ( .C1(n19211), .C2(n19963), .A(n15096), .B(n15095), .ZN(
        n15097) );
  OAI21_X1 U18436 ( .B1(n15098), .B2(n19216), .A(n15097), .ZN(P2_U2854) );
  NAND2_X1 U18437 ( .A1(n15099), .A2(n15205), .ZN(n15100) );
  OAI21_X1 U18438 ( .B1(n15205), .B2(n16330), .A(n15100), .ZN(P2_U2856) );
  OR2_X1 U18439 ( .A1(n15102), .A2(n15101), .ZN(n15103) );
  NAND3_X1 U18440 ( .A1(n10062), .A2(n15212), .A3(n15105), .ZN(n15107) );
  NAND2_X1 U18441 ( .A1(n9750), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15106) );
  OAI211_X1 U18442 ( .C1(n9750), .C2(n16347), .A(n15107), .B(n15106), .ZN(
        P2_U2858) );
  NAND2_X1 U18443 ( .A1(n15109), .A2(n15108), .ZN(n15111) );
  XNOR2_X1 U18444 ( .A(n15111), .B(n15110), .ZN(n15222) );
  NOR2_X1 U18445 ( .A1(n16358), .A2(n9769), .ZN(n15112) );
  AOI21_X1 U18446 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n9750), .A(n15112), .ZN(
        n15113) );
  OAI21_X1 U18447 ( .B1(n15222), .B2(n15178), .A(n15113), .ZN(P2_U2859) );
  AOI21_X1 U18448 ( .B1(n15116), .B2(n15115), .A(n15114), .ZN(n15117) );
  INV_X1 U18449 ( .A(n15117), .ZN(n15230) );
  NOR2_X1 U18450 ( .A1(n15491), .A2(n9750), .ZN(n15118) );
  AOI21_X1 U18451 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n9769), .A(n15118), .ZN(
        n15119) );
  OAI21_X1 U18452 ( .B1(n15230), .B2(n15178), .A(n15119), .ZN(P2_U2860) );
  AOI21_X1 U18453 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15123) );
  INV_X1 U18454 ( .A(n15123), .ZN(n15239) );
  OR2_X1 U18455 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  NAND2_X1 U18456 ( .A1(n13433), .A2(n15126), .ZN(n16369) );
  NOR2_X1 U18457 ( .A1(n16369), .A2(n9769), .ZN(n15127) );
  AOI21_X1 U18458 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n9750), .A(n15127), .ZN(
        n15128) );
  OAI21_X1 U18459 ( .B1(n15239), .B2(n15178), .A(n15128), .ZN(P2_U2861) );
  AOI21_X1 U18460 ( .B1(n9869), .B2(n15130), .A(n15129), .ZN(n15131) );
  XOR2_X1 U18461 ( .A(n15132), .B(n15131), .Z(n15247) );
  AND2_X1 U18462 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  OR2_X1 U18463 ( .A1(n15135), .A2(n14326), .ZN(n16390) );
  MUX2_X1 U18464 ( .A(n16390), .B(n15136), .S(n9769), .Z(n15137) );
  OAI21_X1 U18465 ( .B1(n15247), .B2(n15178), .A(n15137), .ZN(P2_U2863) );
  AOI21_X1 U18466 ( .B1(n15138), .B2(n15140), .A(n15139), .ZN(n15248) );
  NAND2_X1 U18467 ( .A1(n15248), .A2(n15212), .ZN(n15142) );
  NAND2_X1 U18468 ( .A1(n9750), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15141) );
  OAI211_X1 U18469 ( .C1(n15534), .C2(n9750), .A(n15142), .B(n15141), .ZN(
        P2_U2864) );
  NAND2_X1 U18470 ( .A1(n15193), .A2(n15144), .ZN(n15150) );
  AOI21_X1 U18471 ( .B1(n15146), .B2(n15150), .A(n15145), .ZN(n16393) );
  NAND2_X1 U18472 ( .A1(n16393), .A2(n15212), .ZN(n15148) );
  NAND2_X1 U18473 ( .A1(n9769), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15147) );
  OAI211_X1 U18474 ( .C1(n15552), .C2(n9769), .A(n15148), .B(n15147), .ZN(
        P2_U2865) );
  NAND2_X1 U18475 ( .A1(n15193), .A2(n15182), .ZN(n15164) );
  INV_X1 U18476 ( .A(n15164), .ZN(n15183) );
  AND2_X1 U18477 ( .A1(n15183), .A2(n15149), .ZN(n15158) );
  OAI21_X1 U18478 ( .B1(n15158), .B2(n15151), .A(n15150), .ZN(n15260) );
  NOR2_X1 U18479 ( .A1(n15559), .A2(n9750), .ZN(n15152) );
  AOI21_X1 U18480 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n9769), .A(n15152), .ZN(
        n15153) );
  OAI21_X1 U18481 ( .B1(n15260), .B2(n15178), .A(n15153), .ZN(P2_U2866) );
  AND2_X1 U18482 ( .A1(n15162), .A2(n15155), .ZN(n15156) );
  OR2_X1 U18483 ( .A1(n15156), .A2(n10218), .ZN(n19010) );
  OR2_X1 U18484 ( .A1(n15164), .A2(n15157), .ZN(n15165) );
  AOI21_X1 U18485 ( .B1(n15159), .B2(n15165), .A(n15158), .ZN(n16398) );
  NAND2_X1 U18486 ( .A1(n16398), .A2(n15212), .ZN(n15161) );
  NAND2_X1 U18487 ( .A1(n9750), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15160) );
  OAI211_X1 U18488 ( .C1(n19010), .C2(n9750), .A(n15161), .B(n15160), .ZN(
        P2_U2867) );
  AOI21_X1 U18489 ( .B1(n15163), .B2(n15175), .A(n15154), .ZN(n19025) );
  INV_X1 U18490 ( .A(n19025), .ZN(n15588) );
  OR2_X1 U18491 ( .A1(n15164), .A2(n15170), .ZN(n15171) );
  INV_X1 U18492 ( .A(n15165), .ZN(n15166) );
  AOI21_X1 U18493 ( .B1(n15167), .B2(n15171), .A(n15166), .ZN(n15261) );
  NAND2_X1 U18494 ( .A1(n15261), .A2(n15212), .ZN(n15169) );
  NAND2_X1 U18495 ( .A1(n9769), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15168) );
  OAI211_X1 U18496 ( .C1(n15588), .C2(n9750), .A(n15169), .B(n15168), .ZN(
        P2_U2868) );
  INV_X1 U18497 ( .A(n15170), .ZN(n15172) );
  OAI21_X1 U18498 ( .B1(n15183), .B2(n15172), .A(n15171), .ZN(n15283) );
  OR2_X1 U18499 ( .A1(n15180), .A2(n15173), .ZN(n15174) );
  NAND2_X1 U18500 ( .A1(n15175), .A2(n15174), .ZN(n15595) );
  NOR2_X1 U18501 ( .A1(n15595), .A2(n9769), .ZN(n15176) );
  AOI21_X1 U18502 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n9750), .A(n15176), .ZN(
        n15177) );
  OAI21_X1 U18503 ( .B1(n15283), .B2(n15178), .A(n15177), .ZN(P2_U2869) );
  AND2_X1 U18504 ( .A1(n15190), .A2(n15179), .ZN(n15181) );
  OR2_X1 U18505 ( .A1(n15181), .A2(n15180), .ZN(n15608) );
  INV_X1 U18506 ( .A(n15182), .ZN(n15185) );
  INV_X1 U18507 ( .A(n15193), .ZN(n15184) );
  AOI21_X1 U18508 ( .B1(n15185), .B2(n15184), .A(n15183), .ZN(n15284) );
  NAND2_X1 U18509 ( .A1(n15284), .A2(n15212), .ZN(n15187) );
  NAND2_X1 U18510 ( .A1(n9769), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15186) );
  OAI211_X1 U18511 ( .C1(n15608), .C2(n9769), .A(n15187), .B(n15186), .ZN(
        P2_U2870) );
  NAND2_X1 U18512 ( .A1(n15201), .A2(n15188), .ZN(n15189) );
  NAND2_X1 U18513 ( .A1(n15190), .A2(n15189), .ZN(n19063) );
  INV_X1 U18514 ( .A(n15191), .ZN(n15194) );
  INV_X1 U18515 ( .A(n15192), .ZN(n15198) );
  AOI21_X1 U18516 ( .B1(n15194), .B2(n15198), .A(n15193), .ZN(n19226) );
  NAND2_X1 U18517 ( .A1(n19226), .A2(n15212), .ZN(n15196) );
  NAND2_X1 U18518 ( .A1(n9750), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15195) );
  OAI211_X1 U18519 ( .C1(n19063), .C2(n9750), .A(n15196), .B(n15195), .ZN(
        P2_U2871) );
  INV_X1 U18520 ( .A(n15197), .ZN(n15199) );
  OAI211_X1 U18521 ( .C1(n15143), .C2(n15199), .A(n15198), .B(n15212), .ZN(
        n15204) );
  OAI21_X1 U18522 ( .B1(n10515), .B2(n10514), .A(n15201), .ZN(n19070) );
  INV_X1 U18523 ( .A(n19070), .ZN(n15202) );
  NAND2_X1 U18524 ( .A1(n15202), .A2(n15205), .ZN(n15203) );
  OAI211_X1 U18525 ( .C1(n15205), .C2(n10920), .A(n15204), .B(n15203), .ZN(
        P2_U2872) );
  OR2_X1 U18526 ( .A1(n15207), .A2(n15206), .ZN(n15208) );
  AND2_X1 U18527 ( .A1(n15209), .A2(n15208), .ZN(n19080) );
  INV_X1 U18528 ( .A(n19080), .ZN(n15217) );
  INV_X1 U18529 ( .A(n14252), .ZN(n15214) );
  INV_X1 U18530 ( .A(n15210), .ZN(n15213) );
  OAI211_X1 U18531 ( .C1(n15214), .C2(n15213), .A(n15212), .B(n15211), .ZN(
        n15216) );
  NAND2_X1 U18532 ( .A1(n9750), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15215) );
  OAI211_X1 U18533 ( .C1(n15217), .C2(n9769), .A(n15216), .B(n15215), .ZN(
        P2_U2873) );
  AOI22_X1 U18534 ( .A1(n19222), .A2(BUF2_REG_28__SCAN_IN), .B1(n19221), .B2(
        n19233), .ZN(n15221) );
  INV_X1 U18535 ( .A(n16356), .ZN(n15218) );
  OAI22_X1 U18536 ( .A1(n15218), .A2(n15276), .B1(n19249), .B2(n13604), .ZN(
        n15219) );
  AOI21_X1 U18537 ( .B1(n19223), .B2(BUF1_REG_28__SCAN_IN), .A(n15219), .ZN(
        n15220) );
  OAI211_X1 U18538 ( .C1(n15222), .C2(n15282), .A(n15221), .B(n15220), .ZN(
        P2_U2891) );
  OAI22_X1 U18539 ( .A1(n15276), .A2(n15494), .B1(n19249), .B2(n15223), .ZN(
        n15228) );
  INV_X1 U18540 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15226) );
  OAI22_X1 U18541 ( .A1(n15278), .A2(n15226), .B1(n15225), .B2(n15224), .ZN(
        n15227) );
  AOI211_X1 U18542 ( .C1(n19223), .C2(BUF1_REG_27__SCAN_IN), .A(n15228), .B(
        n15227), .ZN(n15229) );
  OAI21_X1 U18543 ( .B1(n15230), .B2(n15282), .A(n15229), .ZN(P2_U2892) );
  AOI22_X1 U18544 ( .A1(n19222), .A2(BUF2_REG_26__SCAN_IN), .B1(n19221), .B2(
        n19236), .ZN(n15238) );
  INV_X1 U18545 ( .A(n15231), .ZN(n15235) );
  NAND2_X1 U18546 ( .A1(n15233), .A2(n15232), .ZN(n15234) );
  NAND2_X1 U18547 ( .A1(n15235), .A2(n15234), .ZN(n16364) );
  OAI22_X1 U18548 ( .A1(n15276), .A2(n16364), .B1(n19249), .B2(n13602), .ZN(
        n15236) );
  AOI21_X1 U18549 ( .B1(n19223), .B2(BUF1_REG_26__SCAN_IN), .A(n15236), .ZN(
        n15237) );
  OAI211_X1 U18550 ( .C1(n15239), .C2(n15282), .A(n15238), .B(n15237), .ZN(
        P2_U2893) );
  AOI22_X1 U18551 ( .A1(n19222), .A2(BUF2_REG_24__SCAN_IN), .B1(n19221), .B2(
        n19244), .ZN(n15246) );
  INV_X1 U18552 ( .A(n15240), .ZN(n15241) );
  AOI21_X1 U18553 ( .B1(n15242), .B2(n15050), .A(n15241), .ZN(n16386) );
  INV_X1 U18554 ( .A(n16386), .ZN(n15243) );
  OAI22_X1 U18555 ( .A1(n15276), .A2(n15243), .B1(n19249), .B2(n13608), .ZN(
        n15244) );
  AOI21_X1 U18556 ( .B1(n19223), .B2(BUF1_REG_24__SCAN_IN), .A(n15244), .ZN(
        n15245) );
  OAI211_X1 U18557 ( .C1(n15247), .C2(n15282), .A(n15246), .B(n15245), .ZN(
        P2_U2895) );
  NAND2_X1 U18558 ( .A1(n15248), .A2(n19225), .ZN(n15254) );
  INV_X1 U18559 ( .A(n15539), .ZN(n15249) );
  AOI22_X1 U18560 ( .A1(n19222), .A2(BUF2_REG_23__SCAN_IN), .B1(n13389), .B2(
        n15249), .ZN(n15253) );
  INV_X1 U18561 ( .A(n19370), .ZN(n15250) );
  AOI22_X1 U18562 ( .A1(n19221), .A2(n15250), .B1(n19239), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U18563 ( .A1(n19223), .A2(BUF1_REG_23__SCAN_IN), .ZN(n15251) );
  NAND4_X1 U18564 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        P2_U2896) );
  AOI22_X1 U18565 ( .A1(n19222), .A2(BUF2_REG_21__SCAN_IN), .B1(n13389), .B2(
        n15562), .ZN(n15258) );
  INV_X1 U18566 ( .A(n19359), .ZN(n15255) );
  AOI22_X1 U18567 ( .A1(n19221), .A2(n15255), .B1(n19239), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15257) );
  NAND2_X1 U18568 ( .A1(n19223), .A2(BUF1_REG_21__SCAN_IN), .ZN(n15256) );
  AND3_X1 U18569 ( .A1(n15258), .A2(n15257), .A3(n15256), .ZN(n15259) );
  OAI21_X1 U18570 ( .B1(n15260), .B2(n15282), .A(n15259), .ZN(P2_U2898) );
  NAND2_X1 U18571 ( .A1(n15261), .A2(n19225), .ZN(n15270) );
  NOR2_X1 U18572 ( .A1(n15264), .A2(n15263), .ZN(n15265) );
  AOI22_X1 U18573 ( .A1(n19222), .A2(BUF2_REG_19__SCAN_IN), .B1(n13389), .B2(
        n10207), .ZN(n15269) );
  AOI22_X1 U18574 ( .A1(n19221), .A2(n15266), .B1(n19239), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U18575 ( .A1(n19223), .A2(BUF1_REG_19__SCAN_IN), .ZN(n15267) );
  NAND4_X1 U18576 ( .A1(n15270), .A2(n15269), .A3(n15268), .A4(n15267), .ZN(
        P2_U2900) );
  NAND2_X1 U18577 ( .A1(n19221), .A2(n15271), .ZN(n15272) );
  OAI21_X1 U18578 ( .B1(n19249), .B2(n15273), .A(n15272), .ZN(n15280) );
  INV_X1 U18579 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n15277) );
  XNOR2_X1 U18580 ( .A(n15274), .B(n15275), .ZN(n19038) );
  OAI22_X1 U18581 ( .A1(n15278), .A2(n15277), .B1(n19038), .B2(n15276), .ZN(
        n15279) );
  AOI211_X1 U18582 ( .C1(n19223), .C2(BUF1_REG_18__SCAN_IN), .A(n15280), .B(
        n15279), .ZN(n15281) );
  OAI21_X1 U18583 ( .B1(n15283), .B2(n15282), .A(n15281), .ZN(P2_U2901) );
  NAND2_X1 U18584 ( .A1(n15284), .A2(n19225), .ZN(n15292) );
  INV_X1 U18585 ( .A(n15274), .ZN(n15286) );
  AOI21_X1 U18586 ( .B1(n15287), .B2(n15285), .A(n15286), .ZN(n19047) );
  AOI22_X1 U18587 ( .A1(n19222), .A2(BUF2_REG_17__SCAN_IN), .B1(n13389), .B2(
        n19047), .ZN(n15291) );
  AOI22_X1 U18588 ( .A1(n19221), .A2(n15288), .B1(n19239), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15290) );
  NAND2_X1 U18589 ( .A1(n19223), .A2(BUF1_REG_17__SCAN_IN), .ZN(n15289) );
  NAND4_X1 U18590 ( .A1(n15292), .A2(n15291), .A3(n15290), .A4(n15289), .ZN(
        P2_U2902) );
  NAND2_X1 U18591 ( .A1(n15294), .A2(n15293), .ZN(n15296) );
  XOR2_X1 U18592 ( .A(n15296), .B(n15295), .Z(n15489) );
  NAND2_X1 U18593 ( .A1(n15478), .A2(n19300), .ZN(n15303) );
  NAND2_X1 U18594 ( .A1(n15730), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15483) );
  OAI21_X1 U18595 ( .B1(n16462), .B2(n9972), .A(n15483), .ZN(n15301) );
  NOR2_X1 U18596 ( .A1(n16347), .A2(n19289), .ZN(n15300) );
  AOI211_X1 U18597 ( .C1(n16453), .C2(n16343), .A(n15301), .B(n15300), .ZN(
        n15302) );
  OAI211_X1 U18598 ( .C1(n15489), .C2(n19305), .A(n15303), .B(n15302), .ZN(
        P2_U2985) );
  XNOR2_X1 U18599 ( .A(n15304), .B(n15479), .ZN(n15500) );
  AOI21_X1 U18600 ( .B1(n15479), .B2(n15305), .A(n15306), .ZN(n15490) );
  NAND2_X1 U18601 ( .A1(n15730), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15493) );
  OAI21_X1 U18602 ( .B1(n16462), .B2(n15307), .A(n15493), .ZN(n15308) );
  AOI21_X1 U18603 ( .B1(n16453), .B2(n15309), .A(n15308), .ZN(n15310) );
  OAI21_X1 U18604 ( .B1(n15491), .B2(n19289), .A(n15310), .ZN(n15311) );
  AOI21_X1 U18605 ( .B1(n15490), .B2(n19300), .A(n15311), .ZN(n15312) );
  OAI21_X1 U18606 ( .B1(n15500), .B2(n19305), .A(n15312), .ZN(P2_U2987) );
  NOR2_X1 U18607 ( .A1(n15313), .A2(n15327), .ZN(n15326) );
  OAI21_X1 U18608 ( .B1(n15326), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15305), .ZN(n15512) );
  OAI21_X1 U18609 ( .B1(n9788), .B2(n15323), .A(n15322), .ZN(n15316) );
  XNOR2_X1 U18610 ( .A(n15316), .B(n15315), .ZN(n15510) );
  NOR2_X1 U18611 ( .A1(n16369), .A2(n19289), .ZN(n15320) );
  NAND2_X1 U18612 ( .A1(n15730), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15504) );
  NAND2_X1 U18613 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15317) );
  OAI211_X1 U18614 ( .C1(n19294), .C2(n15318), .A(n15504), .B(n15317), .ZN(
        n15319) );
  AOI211_X1 U18615 ( .C1(n15510), .C2(n19283), .A(n15320), .B(n15319), .ZN(
        n15321) );
  OAI21_X1 U18616 ( .B1(n15512), .B2(n16456), .A(n15321), .ZN(P2_U2988) );
  INV_X1 U18617 ( .A(n15322), .ZN(n15324) );
  NOR2_X1 U18618 ( .A1(n15324), .A2(n15323), .ZN(n15325) );
  XNOR2_X1 U18619 ( .A(n9788), .B(n15325), .ZN(n15524) );
  INV_X1 U18620 ( .A(n15326), .ZN(n15514) );
  NAND2_X1 U18621 ( .A1(n15313), .A2(n15327), .ZN(n15513) );
  NAND3_X1 U18622 ( .A1(n15514), .A2(n19300), .A3(n15513), .ZN(n15331) );
  NAND2_X1 U18623 ( .A1(n15730), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15516) );
  OAI21_X1 U18624 ( .B1(n16462), .B2(n16373), .A(n15516), .ZN(n15329) );
  NOR2_X1 U18625 ( .A1(n16380), .A2(n19289), .ZN(n15328) );
  AOI211_X1 U18626 ( .C1(n16453), .C2(n16372), .A(n15329), .B(n15328), .ZN(
        n15330) );
  OAI211_X1 U18627 ( .C1(n19305), .C2(n15524), .A(n15331), .B(n15330), .ZN(
        P2_U2989) );
  AND2_X1 U18628 ( .A1(n9804), .A2(n15332), .ZN(n15343) );
  OAI21_X1 U18629 ( .B1(n15343), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15313), .ZN(n15533) );
  XNOR2_X1 U18630 ( .A(n15334), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15335) );
  XNOR2_X1 U18631 ( .A(n15333), .B(n15335), .ZN(n15531) );
  INV_X1 U18632 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U18633 ( .A1(n19151), .A2(n15336), .ZN(n15527) );
  NOR2_X1 U18634 ( .A1(n19294), .A2(n15337), .ZN(n15338) );
  AOI211_X1 U18635 ( .C1(n19296), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15527), .B(n15338), .ZN(n15339) );
  OAI21_X1 U18636 ( .B1(n16390), .B2(n19289), .A(n15339), .ZN(n15340) );
  AOI21_X1 U18637 ( .B1(n15531), .B2(n19283), .A(n15340), .ZN(n15341) );
  OAI21_X1 U18638 ( .B1(n15533), .B2(n16456), .A(n15341), .ZN(P2_U2990) );
  NOR2_X1 U18639 ( .A1(n15392), .A2(n15342), .ZN(n15353) );
  INV_X1 U18640 ( .A(n15343), .ZN(n15344) );
  OAI21_X1 U18641 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15353), .A(
        n15344), .ZN(n15545) );
  XOR2_X1 U18642 ( .A(n15345), .B(n15346), .Z(n15542) );
  NAND2_X1 U18643 ( .A1(n15730), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15538) );
  OAI21_X1 U18644 ( .B1(n16462), .B2(n15347), .A(n15538), .ZN(n15348) );
  AOI21_X1 U18645 ( .B1(n16453), .B2(n15349), .A(n15348), .ZN(n15350) );
  OAI21_X1 U18646 ( .B1(n15534), .B2(n19289), .A(n15350), .ZN(n15351) );
  AOI21_X1 U18647 ( .B1(n15542), .B2(n19283), .A(n15351), .ZN(n15352) );
  OAI21_X1 U18648 ( .B1(n15545), .B2(n16456), .A(n15352), .ZN(P2_U2991) );
  NOR2_X1 U18649 ( .A1(n15392), .A2(n15564), .ZN(n15381) );
  INV_X1 U18650 ( .A(n15353), .ZN(n15354) );
  OAI21_X1 U18651 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15381), .A(
        n15354), .ZN(n15556) );
  INV_X1 U18652 ( .A(n15357), .ZN(n15359) );
  NOR2_X1 U18653 ( .A1(n15359), .A2(n15358), .ZN(n15360) );
  XNOR2_X1 U18654 ( .A(n15356), .B(n15360), .ZN(n15554) );
  NOR2_X1 U18655 ( .A1(n19151), .A2(n15361), .ZN(n15549) );
  NOR2_X1 U18656 ( .A1(n19294), .A2(n15362), .ZN(n15363) );
  AOI211_X1 U18657 ( .C1(n19296), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15549), .B(n15363), .ZN(n15364) );
  OAI21_X1 U18658 ( .B1(n15552), .B2(n19289), .A(n15364), .ZN(n15365) );
  AOI21_X1 U18659 ( .B1(n15554), .B2(n19283), .A(n15365), .ZN(n15366) );
  OAI21_X1 U18660 ( .B1(n15556), .B2(n16456), .A(n15366), .ZN(P2_U2992) );
  INV_X1 U18661 ( .A(n15646), .ZN(n15368) );
  INV_X1 U18662 ( .A(n15367), .ZN(n15645) );
  NAND2_X1 U18663 ( .A1(n15429), .A2(n15428), .ZN(n15427) );
  INV_X1 U18664 ( .A(n15370), .ZN(n15371) );
  NAND2_X1 U18665 ( .A1(n15371), .A2(n15372), .ZN(n15419) );
  INV_X1 U18666 ( .A(n15373), .ZN(n15374) );
  OAI211_X1 U18667 ( .C1(n15411), .C2(n15374), .A(n15410), .B(n15400), .ZN(
        n15390) );
  INV_X1 U18668 ( .A(n15389), .ZN(n15375) );
  INV_X1 U18669 ( .A(n15376), .ZN(n15377) );
  NOR2_X1 U18670 ( .A1(n15378), .A2(n15377), .ZN(n15379) );
  XNOR2_X1 U18671 ( .A(n15380), .B(n15379), .ZN(n15569) );
  AOI21_X1 U18672 ( .B1(n15564), .B2(n15392), .A(n15381), .ZN(n15567) );
  NAND2_X1 U18673 ( .A1(n15730), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15557) );
  OAI21_X1 U18674 ( .B1(n16462), .B2(n15382), .A(n15557), .ZN(n15383) );
  AOI21_X1 U18675 ( .B1(n16453), .B2(n15384), .A(n15383), .ZN(n15385) );
  OAI21_X1 U18676 ( .B1(n15559), .B2(n19289), .A(n15385), .ZN(n15386) );
  AOI21_X1 U18677 ( .B1(n15567), .B2(n19300), .A(n15386), .ZN(n15387) );
  OAI21_X1 U18678 ( .B1(n15569), .B2(n19305), .A(n15387), .ZN(P2_U2993) );
  NOR2_X1 U18679 ( .A1(n15389), .A2(n15388), .ZN(n15391) );
  XOR2_X1 U18680 ( .A(n15391), .B(n15390), .Z(n15583) );
  INV_X1 U18681 ( .A(n15392), .ZN(n15393) );
  AOI21_X1 U18682 ( .B1(n15575), .B2(n15405), .A(n15393), .ZN(n15581) );
  NOR2_X1 U18683 ( .A1(n19151), .A2(n19908), .ZN(n15577) );
  NOR2_X1 U18684 ( .A1(n19294), .A2(n19017), .ZN(n15394) );
  AOI211_X1 U18685 ( .C1(n19296), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15577), .B(n15394), .ZN(n15395) );
  OAI21_X1 U18686 ( .B1(n19010), .B2(n19289), .A(n15395), .ZN(n15396) );
  AOI21_X1 U18687 ( .B1(n15581), .B2(n19300), .A(n15396), .ZN(n15397) );
  OAI21_X1 U18688 ( .B1(n15583), .B2(n19305), .A(n15397), .ZN(P2_U2994) );
  INV_X1 U18689 ( .A(n15409), .ZN(n15398) );
  OAI21_X1 U18690 ( .B1(n9789), .B2(n15398), .A(n15410), .ZN(n15402) );
  NAND2_X1 U18691 ( .A1(n15400), .A2(n15399), .ZN(n15401) );
  XNOR2_X1 U18692 ( .A(n15402), .B(n15401), .ZN(n15593) );
  NAND2_X1 U18693 ( .A1(n16453), .A2(n19020), .ZN(n15403) );
  NAND2_X1 U18694 ( .A1(n15730), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15584) );
  OAI211_X1 U18695 ( .C1(n16462), .C2(n19021), .A(n15403), .B(n15584), .ZN(
        n15407) );
  NAND2_X1 U18696 ( .A1(n9794), .A2(n15574), .ZN(n15404) );
  NAND2_X1 U18697 ( .A1(n15405), .A2(n15404), .ZN(n15589) );
  NOR2_X1 U18698 ( .A1(n15589), .A2(n16456), .ZN(n15406) );
  OAI21_X1 U18699 ( .B1(n19305), .B2(n15593), .A(n15408), .ZN(P2_U2995) );
  INV_X1 U18700 ( .A(n15595), .ZN(n19035) );
  INV_X1 U18701 ( .A(n19032), .ZN(n15412) );
  NAND2_X1 U18702 ( .A1(n16453), .A2(n15412), .ZN(n15413) );
  NAND2_X1 U18703 ( .A1(n15730), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15599) );
  OAI211_X1 U18704 ( .C1(n16462), .C2(n15414), .A(n15413), .B(n15599), .ZN(
        n15417) );
  OAI21_X1 U18705 ( .B1(n15415), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n9794), .ZN(n15605) );
  NOR2_X1 U18706 ( .A1(n15605), .A2(n16456), .ZN(n15416) );
  AOI211_X1 U18707 ( .C1(n19302), .C2(n19035), .A(n15417), .B(n15416), .ZN(
        n15418) );
  OAI21_X1 U18708 ( .B1(n15594), .B2(n19305), .A(n15418), .ZN(P2_U2996) );
  XNOR2_X1 U18709 ( .A(n9786), .B(n15419), .ZN(n15620) );
  INV_X1 U18710 ( .A(n15608), .ZN(n19046) );
  NOR2_X1 U18711 ( .A1(n19151), .A2(n19902), .ZN(n15606) );
  AOI21_X1 U18712 ( .B1(n19296), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15606), .ZN(n15421) );
  OAI21_X1 U18713 ( .B1(n19294), .B2(n19050), .A(n15421), .ZN(n15425) );
  AOI211_X1 U18714 ( .C1(n15423), .C2(n15422), .A(n16456), .B(n15415), .ZN(
        n15424) );
  AOI211_X1 U18715 ( .C1(n19302), .C2(n19046), .A(n15425), .B(n15424), .ZN(
        n15426) );
  OAI21_X1 U18716 ( .B1(n15620), .B2(n19305), .A(n15426), .ZN(P2_U2997) );
  OAI21_X1 U18717 ( .B1(n9806), .B2(n15428), .A(n15427), .ZN(n15630) );
  INV_X1 U18718 ( .A(n19063), .ZN(n15626) );
  NAND2_X1 U18719 ( .A1(n15730), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15622) );
  NAND2_X1 U18720 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15430) );
  OAI211_X1 U18721 ( .C1(n19294), .C2(n19058), .A(n15622), .B(n15430), .ZN(
        n15431) );
  AOI21_X1 U18722 ( .B1(n19302), .B2(n15626), .A(n15431), .ZN(n15434) );
  INV_X1 U18723 ( .A(n15432), .ZN(n15610) );
  OAI211_X1 U18724 ( .C1(n15610), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n19300), .B(n15422), .ZN(n15433) );
  OAI211_X1 U18725 ( .C1(n15630), .C2(n19305), .A(n15434), .B(n15433), .ZN(
        P2_U2998) );
  OAI21_X1 U18726 ( .B1(n15436), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15432), .ZN(n15642) );
  INV_X1 U18727 ( .A(n15437), .ZN(n15438) );
  NOR2_X1 U18728 ( .A1(n15439), .A2(n15438), .ZN(n15440) );
  XNOR2_X1 U18729 ( .A(n15441), .B(n15440), .ZN(n15631) );
  NAND2_X1 U18730 ( .A1(n15631), .A2(n19283), .ZN(n15445) );
  NAND2_X1 U18731 ( .A1(n15730), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15636) );
  OAI21_X1 U18732 ( .B1(n16462), .B2(n10224), .A(n15636), .ZN(n15443) );
  NOR2_X1 U18733 ( .A1(n19070), .A2(n19289), .ZN(n15442) );
  AOI211_X1 U18734 ( .C1(n16453), .C2(n19065), .A(n15443), .B(n15442), .ZN(
        n15444) );
  OAI211_X1 U18735 ( .C1(n16456), .C2(n15642), .A(n15445), .B(n15444), .ZN(
        P2_U2999) );
  XNOR2_X1 U18736 ( .A(n16411), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15670) );
  INV_X1 U18737 ( .A(n15447), .ZN(n15448) );
  NOR2_X1 U18738 ( .A1(n15449), .A2(n15448), .ZN(n15450) );
  XNOR2_X1 U18739 ( .A(n9797), .B(n15450), .ZN(n15667) );
  NAND2_X1 U18740 ( .A1(n15730), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15663) );
  OAI21_X1 U18741 ( .B1(n16462), .B2(n15452), .A(n15663), .ZN(n15453) );
  AOI21_X1 U18742 ( .B1(n16453), .B2(n19093), .A(n15453), .ZN(n15454) );
  OAI21_X1 U18743 ( .B1(n19289), .B2(n15660), .A(n15454), .ZN(n15455) );
  AOI21_X1 U18744 ( .B1(n15667), .B2(n19283), .A(n15455), .ZN(n15456) );
  OAI21_X1 U18745 ( .B1(n15670), .B2(n16456), .A(n15456), .ZN(P2_U3001) );
  OAI21_X1 U18746 ( .B1(n15457), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15458), .ZN(n15715) );
  NAND2_X1 U18747 ( .A1(n15460), .A2(n15687), .ZN(n15461) );
  XNOR2_X1 U18748 ( .A(n15459), .B(n15461), .ZN(n15712) );
  INV_X1 U18749 ( .A(n19125), .ZN(n15462) );
  OAI22_X1 U18750 ( .A1(n16462), .A2(n15463), .B1(n19294), .B2(n15462), .ZN(
        n15466) );
  OAI22_X1 U18751 ( .A1(n19289), .A2(n15702), .B1(n19151), .B2(n15464), .ZN(
        n15465) );
  AOI211_X1 U18752 ( .C1(n15712), .C2(n19283), .A(n15466), .B(n15465), .ZN(
        n15467) );
  OAI21_X1 U18753 ( .B1(n15715), .B2(n16456), .A(n15467), .ZN(P2_U3005) );
  NAND2_X1 U18754 ( .A1(n16432), .A2(n16434), .ZN(n15469) );
  XOR2_X1 U18755 ( .A(n15469), .B(n15468), .Z(n15724) );
  OR2_X1 U18756 ( .A1(n15470), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15716) );
  NAND3_X1 U18757 ( .A1(n15716), .A2(n15472), .A3(n19300), .ZN(n15477) );
  OAI22_X1 U18758 ( .A1(n16462), .A2(n15473), .B1(n10477), .B2(n19151), .ZN(
        n15475) );
  NOR2_X1 U18759 ( .A1(n19289), .A2(n19145), .ZN(n15474) );
  AOI211_X1 U18760 ( .C1(n16453), .C2(n19141), .A(n15475), .B(n15474), .ZN(
        n15476) );
  OAI211_X1 U18761 ( .C1(n15724), .C2(n19305), .A(n15477), .B(n15476), .ZN(
        P2_U3007) );
  NAND2_X1 U18762 ( .A1(n15478), .A2(n19319), .ZN(n15488) );
  NOR2_X1 U18763 ( .A1(n16347), .A2(n19317), .ZN(n15485) );
  OAI21_X1 U18764 ( .B1(n15479), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15480) );
  OAI211_X1 U18765 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n15481), .B(n15480), .ZN(
        n15482) );
  OAI211_X1 U18766 ( .C1(n16340), .C2(n16466), .A(n15483), .B(n15482), .ZN(
        n15484) );
  AOI211_X1 U18767 ( .C1(n15486), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15485), .B(n15484), .ZN(n15487) );
  OAI211_X1 U18768 ( .C1(n15489), .C2(n15761), .A(n15488), .B(n15487), .ZN(
        P2_U3017) );
  NAND2_X1 U18769 ( .A1(n15490), .A2(n19319), .ZN(n15499) );
  NOR2_X1 U18770 ( .A1(n15491), .A2(n19317), .ZN(n15496) );
  OAI211_X1 U18771 ( .C1(n16466), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n15495) );
  AOI211_X1 U18772 ( .C1(n15497), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15496), .B(n15495), .ZN(n15498) );
  OAI211_X1 U18773 ( .C1(n15500), .C2(n15761), .A(n15499), .B(n15498), .ZN(
        P2_U3019) );
  INV_X1 U18774 ( .A(n16369), .ZN(n15506) );
  INV_X1 U18775 ( .A(n15517), .ZN(n15501) );
  OAI211_X1 U18776 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15502), .B(n15501), .ZN(
        n15503) );
  OAI211_X1 U18777 ( .C1(n16466), .C2(n16364), .A(n15504), .B(n15503), .ZN(
        n15505) );
  AOI21_X1 U18778 ( .B1(n15506), .B2(n16486), .A(n15505), .ZN(n15507) );
  OAI21_X1 U18779 ( .B1(n15515), .B2(n15508), .A(n15507), .ZN(n15509) );
  AOI21_X1 U18780 ( .B1(n15510), .B2(n19316), .A(n15509), .ZN(n15511) );
  OAI21_X1 U18781 ( .B1(n15512), .B2(n16496), .A(n15511), .ZN(P2_U3020) );
  NAND3_X1 U18782 ( .A1(n15514), .A2(n19319), .A3(n15513), .ZN(n15523) );
  INV_X1 U18783 ( .A(n15515), .ZN(n15521) );
  OAI21_X1 U18784 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15517), .A(
        n15516), .ZN(n15518) );
  AOI21_X1 U18785 ( .B1(n19326), .B2(n16376), .A(n15518), .ZN(n15519) );
  OAI21_X1 U18786 ( .B1(n16380), .B2(n19317), .A(n15519), .ZN(n15520) );
  AOI21_X1 U18787 ( .B1(n15521), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15520), .ZN(n15522) );
  OAI211_X1 U18788 ( .C1(n15524), .C2(n15761), .A(n15523), .B(n15522), .ZN(
        P2_U3021) );
  OAI21_X1 U18789 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15526), .A(
        n15525), .ZN(n15529) );
  AOI21_X1 U18790 ( .B1(n19326), .B2(n16386), .A(n15527), .ZN(n15528) );
  OAI211_X1 U18791 ( .C1(n19317), .C2(n16390), .A(n15529), .B(n15528), .ZN(
        n15530) );
  AOI21_X1 U18792 ( .B1(n15531), .B2(n19316), .A(n15530), .ZN(n15532) );
  OAI21_X1 U18793 ( .B1(n15533), .B2(n16496), .A(n15532), .ZN(P2_U3022) );
  NOR2_X1 U18794 ( .A1(n15534), .A2(n19317), .ZN(n15541) );
  INV_X1 U18795 ( .A(n15547), .ZN(n15536) );
  OAI211_X1 U18796 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15536), .B(n15535), .ZN(
        n15537) );
  OAI211_X1 U18797 ( .C1(n16466), .C2(n15539), .A(n15538), .B(n15537), .ZN(
        n15540) );
  AOI211_X1 U18798 ( .C1(n15546), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15541), .B(n15540), .ZN(n15544) );
  NAND2_X1 U18799 ( .A1(n15542), .A2(n19316), .ZN(n15543) );
  OAI211_X1 U18800 ( .C1(n15545), .C2(n16496), .A(n15544), .B(n15543), .ZN(
        P2_U3023) );
  NAND2_X1 U18801 ( .A1(n15546), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15551) );
  NOR2_X1 U18802 ( .A1(n15547), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15548) );
  AOI211_X1 U18803 ( .C1(n19326), .C2(n16392), .A(n15549), .B(n15548), .ZN(
        n15550) );
  OAI211_X1 U18804 ( .C1(n15552), .C2(n19317), .A(n15551), .B(n15550), .ZN(
        n15553) );
  AOI21_X1 U18805 ( .B1(n15554), .B2(n19316), .A(n15553), .ZN(n15555) );
  OAI21_X1 U18806 ( .B1(n15556), .B2(n16496), .A(n15555), .ZN(P2_U3024) );
  OAI21_X1 U18807 ( .B1(n15558), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15557), .ZN(n15561) );
  NOR2_X1 U18808 ( .A1(n15559), .A2(n19317), .ZN(n15560) );
  AOI211_X1 U18809 ( .C1(n19326), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15563) );
  OAI21_X1 U18810 ( .B1(n15565), .B2(n15564), .A(n15563), .ZN(n15566) );
  AOI21_X1 U18811 ( .B1(n15567), .B2(n19319), .A(n15566), .ZN(n15568) );
  OAI21_X1 U18812 ( .B1(n15569), .B2(n15761), .A(n15568), .ZN(P2_U3025) );
  NAND2_X1 U18813 ( .A1(n15602), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15579) );
  OAI21_X1 U18814 ( .B1(n15262), .B2(n15570), .A(n15080), .ZN(n15571) );
  INV_X1 U18815 ( .A(n15571), .ZN(n19009) );
  INV_X1 U18816 ( .A(n15572), .ZN(n15573) );
  AOI211_X1 U18817 ( .C1(n15575), .C2(n15574), .A(n15573), .B(n15585), .ZN(
        n15576) );
  AOI211_X1 U18818 ( .C1(n19326), .C2(n19009), .A(n15577), .B(n15576), .ZN(
        n15578) );
  OAI211_X1 U18819 ( .C1(n19010), .C2(n19317), .A(n15579), .B(n15578), .ZN(
        n15580) );
  AOI21_X1 U18820 ( .B1(n15581), .B2(n19319), .A(n15580), .ZN(n15582) );
  OAI21_X1 U18821 ( .B1(n15583), .B2(n15761), .A(n15582), .ZN(P2_U3026) );
  OAI21_X1 U18822 ( .B1(n15585), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15584), .ZN(n15586) );
  AOI21_X1 U18823 ( .B1(n19326), .B2(n10207), .A(n15586), .ZN(n15587) );
  OAI21_X1 U18824 ( .B1(n15588), .B2(n19317), .A(n15587), .ZN(n15591) );
  NOR2_X1 U18825 ( .A1(n15589), .A2(n16496), .ZN(n15590) );
  AOI211_X1 U18826 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15602), .A(
        n15591), .B(n15590), .ZN(n15592) );
  OAI21_X1 U18827 ( .B1(n15761), .B2(n15593), .A(n15592), .ZN(P2_U3027) );
  OR2_X1 U18828 ( .A1(n15594), .A2(n15761), .ZN(n15604) );
  NOR2_X1 U18829 ( .A1(n15595), .A2(n19317), .ZN(n15601) );
  NAND2_X1 U18830 ( .A1(n15597), .A2(n15596), .ZN(n15598) );
  OAI211_X1 U18831 ( .C1(n16466), .C2(n19038), .A(n15599), .B(n15598), .ZN(
        n15600) );
  AOI211_X1 U18832 ( .C1(n15602), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15601), .B(n15600), .ZN(n15603) );
  OAI211_X1 U18833 ( .C1(n15605), .C2(n16496), .A(n15604), .B(n15603), .ZN(
        P2_U3028) );
  INV_X1 U18834 ( .A(n15606), .ZN(n15607) );
  OAI21_X1 U18835 ( .B1(n15608), .B2(n19317), .A(n15607), .ZN(n15613) );
  INV_X1 U18836 ( .A(n15609), .ZN(n15634) );
  AOI22_X1 U18837 ( .A1(n15610), .A2(n19319), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15634), .ZN(n15623) );
  NOR3_X1 U18838 ( .A1(n15623), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15611), .ZN(n15612) );
  AOI211_X1 U18839 ( .C1(n19326), .C2(n19047), .A(n15613), .B(n15612), .ZN(
        n15619) );
  OAI21_X1 U18840 ( .B1(n19319), .B2(n19314), .A(n15422), .ZN(n15614) );
  OAI211_X1 U18841 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15615), .A(
        n15614), .B(n15632), .ZN(n15627) );
  NOR2_X1 U18842 ( .A1(n15616), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15617) );
  OAI21_X1 U18843 ( .B1(n15627), .B2(n15617), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15618) );
  OAI211_X1 U18844 ( .C1(n15620), .C2(n15761), .A(n15619), .B(n15618), .ZN(
        P2_U3029) );
  OAI21_X1 U18845 ( .B1(n14145), .B2(n15621), .A(n15285), .ZN(n19056) );
  OAI21_X1 U18846 ( .B1(n16466), .B2(n19056), .A(n15622), .ZN(n15625) );
  NOR2_X1 U18847 ( .A1(n15623), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15624) );
  AOI211_X1 U18848 ( .C1(n16486), .C2(n15626), .A(n15625), .B(n15624), .ZN(
        n15629) );
  NAND2_X1 U18849 ( .A1(n15627), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15628) );
  OAI211_X1 U18850 ( .C1(n15761), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        P2_U3030) );
  NAND2_X1 U18851 ( .A1(n15631), .A2(n19316), .ZN(n15641) );
  INV_X1 U18852 ( .A(n15632), .ZN(n15639) );
  NOR2_X1 U18853 ( .A1(n19070), .A2(n19317), .ZN(n15638) );
  NAND2_X1 U18854 ( .A1(n15634), .A2(n15633), .ZN(n15635) );
  OAI211_X1 U18855 ( .C1(n16466), .C2(n19069), .A(n15636), .B(n15635), .ZN(
        n15637) );
  AOI211_X1 U18856 ( .C1(n15639), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15638), .B(n15637), .ZN(n15640) );
  OAI211_X1 U18857 ( .C1(n15642), .C2(n16496), .A(n15641), .B(n15640), .ZN(
        P2_U3031) );
  AOI21_X1 U18858 ( .B1(n16411), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15643) );
  NOR2_X1 U18859 ( .A1(n15643), .A2(n15436), .ZN(n16403) );
  INV_X1 U18860 ( .A(n16403), .ZN(n15659) );
  OR2_X1 U18861 ( .A1(n15646), .A2(n15645), .ZN(n15647) );
  XNOR2_X1 U18862 ( .A(n9800), .B(n15647), .ZN(n16402) );
  INV_X1 U18863 ( .A(n16473), .ZN(n15648) );
  OAI21_X1 U18864 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15648), .A(
        n16467), .ZN(n15666) );
  AOI21_X1 U18865 ( .B1(n16473), .B2(n15661), .A(n15666), .ZN(n15656) );
  OAI21_X1 U18866 ( .B1(n13980), .B2(n15649), .A(n14143), .ZN(n15650) );
  INV_X1 U18867 ( .A(n15650), .ZN(n19231) );
  NAND2_X1 U18868 ( .A1(n19326), .A2(n19231), .ZN(n15652) );
  NAND4_X1 U18869 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16473), .A4(n15655), .ZN(
        n15651) );
  OAI211_X1 U18870 ( .C1(n10855), .C2(n19151), .A(n15652), .B(n15651), .ZN(
        n15653) );
  AOI21_X1 U18871 ( .B1(n16486), .B2(n19080), .A(n15653), .ZN(n15654) );
  OAI21_X1 U18872 ( .B1(n15656), .B2(n15655), .A(n15654), .ZN(n15657) );
  AOI21_X1 U18873 ( .B1(n16402), .B2(n19316), .A(n15657), .ZN(n15658) );
  OAI21_X1 U18874 ( .B1(n15659), .B2(n16496), .A(n15658), .ZN(P2_U3032) );
  NOR2_X1 U18875 ( .A1(n19317), .A2(n15660), .ZN(n15665) );
  NAND3_X1 U18876 ( .A1(n16473), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n15661), .ZN(n15662) );
  OAI211_X1 U18877 ( .C1(n16466), .C2(n19097), .A(n15663), .B(n15662), .ZN(
        n15664) );
  AOI211_X1 U18878 ( .C1(n15666), .C2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15665), .B(n15664), .ZN(n15669) );
  NAND2_X1 U18879 ( .A1(n15667), .A2(n19316), .ZN(n15668) );
  OAI211_X1 U18880 ( .C1(n15670), .C2(n16496), .A(n15669), .B(n15668), .ZN(
        P2_U3033) );
  INV_X1 U18881 ( .A(n15446), .ZN(n16423) );
  OAI21_X1 U18882 ( .B1(n16423), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16412), .ZN(n16417) );
  NAND2_X1 U18883 ( .A1(n15762), .A2(n15710), .ZN(n15671) );
  AND2_X1 U18884 ( .A1(n15704), .A2(n15671), .ZN(n15695) );
  INV_X1 U18885 ( .A(n15695), .ZN(n15679) );
  NAND2_X1 U18886 ( .A1(n16486), .A2(n16419), .ZN(n15676) );
  AOI211_X1 U18887 ( .C1(n15673), .C2(n15696), .A(n15672), .B(n15697), .ZN(
        n15674) );
  AOI21_X1 U18888 ( .B1(n15730), .B2(P2_REIP_REG_11__SCAN_IN), .A(n15674), 
        .ZN(n15675) );
  OAI211_X1 U18889 ( .C1(n16466), .C2(n15677), .A(n15676), .B(n15675), .ZN(
        n15678) );
  AOI21_X1 U18890 ( .B1(n15679), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15678), .ZN(n15686) );
  INV_X1 U18891 ( .A(n16407), .ZN(n15682) );
  NOR2_X1 U18892 ( .A1(n15683), .A2(n15682), .ZN(n15684) );
  XNOR2_X1 U18893 ( .A(n15681), .B(n15684), .ZN(n16416) );
  OR2_X1 U18894 ( .A1(n16416), .A2(n15761), .ZN(n15685) );
  OAI211_X1 U18895 ( .C1(n16417), .C2(n16496), .A(n15686), .B(n15685), .ZN(
        P2_U3035) );
  NAND2_X1 U18896 ( .A1(n15688), .A2(n15687), .ZN(n15691) );
  NOR2_X1 U18897 ( .A1(n15689), .A2(n10213), .ZN(n15690) );
  XNOR2_X1 U18898 ( .A(n15691), .B(n15690), .ZN(n16425) );
  INV_X1 U18899 ( .A(n15458), .ZN(n15692) );
  NOR2_X1 U18900 ( .A1(n15692), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16424) );
  OR3_X1 U18901 ( .A1(n16424), .A2(n16423), .A3(n16496), .ZN(n15701) );
  AOI21_X1 U18902 ( .B1(n15706), .B2(n15693), .A(n13444), .ZN(n19237) );
  NOR2_X1 U18903 ( .A1(n19317), .A2(n19119), .ZN(n15699) );
  NAND2_X1 U18904 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n15730), .ZN(n15694) );
  OAI221_X1 U18905 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15697), 
        .C1(n15696), .C2(n15695), .A(n15694), .ZN(n15698) );
  AOI211_X1 U18906 ( .C1(n19326), .C2(n19237), .A(n15699), .B(n15698), .ZN(
        n15700) );
  OAI211_X1 U18907 ( .C1(n16425), .C2(n15761), .A(n15701), .B(n15700), .ZN(
        P2_U3036) );
  INV_X1 U18908 ( .A(n15702), .ZN(n19127) );
  AOI22_X1 U18909 ( .A1(n16486), .A2(n19127), .B1(n15730), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n15703) );
  OAI21_X1 U18910 ( .B1(n15704), .B2(n15710), .A(n15703), .ZN(n15709) );
  OAI21_X1 U18911 ( .B1(n15705), .B2(n15707), .A(n15706), .ZN(n19242) );
  NOR2_X1 U18912 ( .A1(n19242), .A2(n16466), .ZN(n15708) );
  AOI211_X1 U18913 ( .C1(n15711), .C2(n15710), .A(n15709), .B(n15708), .ZN(
        n15714) );
  NAND2_X1 U18914 ( .A1(n15712), .A2(n19316), .ZN(n15713) );
  OAI211_X1 U18915 ( .C1(n15715), .C2(n16496), .A(n15714), .B(n15713), .ZN(
        P2_U3037) );
  NAND3_X1 U18916 ( .A1(n15716), .A2(n15472), .A3(n19319), .ZN(n15723) );
  INV_X1 U18917 ( .A(n16479), .ZN(n15721) );
  INV_X1 U18918 ( .A(n16490), .ZN(n15729) );
  NOR2_X1 U18919 ( .A1(n10477), .A2(n19151), .ZN(n15718) );
  NOR2_X1 U18920 ( .A1(n19317), .A2(n19145), .ZN(n15717) );
  AOI211_X1 U18921 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n15729), .A(
        n15718), .B(n15717), .ZN(n15719) );
  OAI21_X1 U18922 ( .B1(n19146), .B2(n16466), .A(n15719), .ZN(n15720) );
  AOI21_X1 U18923 ( .B1(n15721), .B2(n16481), .A(n15720), .ZN(n15722) );
  OAI211_X1 U18924 ( .C1(n15724), .C2(n15761), .A(n15723), .B(n15722), .ZN(
        P2_U3039) );
  XNOR2_X1 U18925 ( .A(n15726), .B(n15725), .ZN(n16449) );
  INV_X1 U18926 ( .A(n19163), .ZN(n15738) );
  NAND3_X1 U18927 ( .A1(n15749), .A2(n15728), .A3(n15727), .ZN(n15733) );
  AOI22_X1 U18928 ( .A1(n15730), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15729), .ZN(n15732) );
  NAND2_X1 U18929 ( .A1(n19159), .A2(n16486), .ZN(n15731) );
  NAND3_X1 U18930 ( .A1(n15733), .A2(n15732), .A3(n15731), .ZN(n15737) );
  OAI21_X1 U18931 ( .B1(n15734), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15735), .ZN(n16446) );
  NOR2_X1 U18932 ( .A1(n16446), .A2(n16496), .ZN(n15736) );
  AOI211_X1 U18933 ( .C1(n19326), .C2(n15738), .A(n15737), .B(n15736), .ZN(
        n15739) );
  OAI21_X1 U18934 ( .B1(n15761), .B2(n16449), .A(n15739), .ZN(P2_U3040) );
  XNOR2_X1 U18935 ( .A(n15740), .B(n15741), .ZN(n16457) );
  AND2_X1 U18936 ( .A1(n15743), .A2(n15742), .ZN(n15745) );
  OAI22_X1 U18937 ( .A1(n15747), .A2(n15746), .B1(n15745), .B2(n15744), .ZN(
        n16455) );
  INV_X1 U18938 ( .A(n16455), .ZN(n15759) );
  AOI211_X1 U18939 ( .C1(n15755), .C2(n15750), .A(n15749), .B(n15748), .ZN(
        n15758) );
  OAI22_X1 U18940 ( .A1(n16454), .A2(n19317), .B1(n19151), .B2(n15751), .ZN(
        n15752) );
  AOI21_X1 U18941 ( .B1(n15753), .B2(n19326), .A(n15752), .ZN(n15754) );
  OAI21_X1 U18942 ( .B1(n15756), .B2(n15755), .A(n15754), .ZN(n15757) );
  AOI211_X1 U18943 ( .C1(n15759), .C2(n19319), .A(n15758), .B(n15757), .ZN(
        n15760) );
  OAI21_X1 U18944 ( .B1(n15761), .B2(n16457), .A(n15760), .ZN(P2_U3041) );
  OAI211_X1 U18945 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15762), .B(n19322), .ZN(n15771) );
  AOI22_X1 U18946 ( .A1(n16486), .A2(n15764), .B1(n19319), .B2(n15763), .ZN(
        n15770) );
  AOI21_X1 U18947 ( .B1(n15766), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15765), .ZN(n15769) );
  AOI22_X1 U18948 ( .A1(n19316), .A2(n15767), .B1(n19326), .B2(n19966), .ZN(
        n15768) );
  NAND4_X1 U18949 ( .A1(n15771), .A2(n15770), .A3(n15769), .A4(n15768), .ZN(
        P2_U3045) );
  INV_X1 U18950 ( .A(n15772), .ZN(n15773) );
  OAI222_X1 U18951 ( .A1(n16508), .A2(n15775), .B1(n15787), .B2(n15774), .C1(
        n10456), .C2(n15773), .ZN(n15776) );
  MUX2_X1 U18952 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15776), .S(
        n15789), .Z(P2_U3601) );
  INV_X1 U18953 ( .A(n15777), .ZN(n15779) );
  AOI222_X1 U18954 ( .A1(n15781), .A2(n19941), .B1(n19963), .B2(n15780), .C1(
        n15779), .C2(n15778), .ZN(n15783) );
  NAND2_X1 U18955 ( .A1(n15784), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15782) );
  OAI21_X1 U18956 ( .B1(n15784), .B2(n15783), .A(n15782), .ZN(P2_U3600) );
  OAI22_X1 U18957 ( .A1(n19944), .A2(n16508), .B1(n15785), .B2(n15787), .ZN(
        n15786) );
  MUX2_X1 U18958 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15786), .S(
        n15789), .Z(P2_U3596) );
  NOR4_X1 U18959 ( .A1(n10983), .A2(n15788), .A3(n19990), .A4(n15787), .ZN(
        n15790) );
  MUX2_X1 U18960 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n15790), .S(
        n15789), .Z(P2_U3595) );
  INV_X1 U18961 ( .A(n15795), .ZN(n15792) );
  NAND2_X1 U18962 ( .A1(n19944), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19538) );
  INV_X1 U18963 ( .A(n19940), .ZN(n19669) );
  OAI21_X1 U18964 ( .B1(n19538), .B2(n19669), .A(n19942), .ZN(n15798) );
  NOR2_X1 U18965 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19401) );
  INV_X1 U18966 ( .A(n19401), .ZN(n19402) );
  NOR2_X1 U18967 ( .A1(n19968), .A2(n19402), .ZN(n15794) );
  NOR2_X1 U18968 ( .A1(n15798), .A2(n15794), .ZN(n15791) );
  AOI211_X1 U18969 ( .C1(n15792), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n15791), .ZN(n15793) );
  NOR2_X1 U18970 ( .A1(n19402), .A2(n19661), .ZN(n19445) );
  OAI21_X1 U18971 ( .B1(n15793), .B2(n19445), .A(n19738), .ZN(n19448) );
  INV_X1 U18972 ( .A(n19448), .ZN(n15803) );
  INV_X1 U18973 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15802) );
  INV_X1 U18974 ( .A(n15794), .ZN(n15797) );
  OAI21_X1 U18975 ( .B1(n15795), .B2(n19445), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15796) );
  OAI21_X1 U18976 ( .B1(n15798), .B2(n15797), .A(n15796), .ZN(n19447) );
  AOI22_X1 U18977 ( .A1(n19780), .A2(n19463), .B1(n19445), .B2(n19779), .ZN(
        n15799) );
  OAI21_X1 U18978 ( .B1(n19442), .B2(n19793), .A(n15799), .ZN(n15800) );
  AOI21_X1 U18979 ( .B1(n19790), .B2(n19447), .A(n15800), .ZN(n15801) );
  OAI21_X1 U18980 ( .B1(n15803), .B2(n15802), .A(n15801), .ZN(P2_U3072) );
  AOI22_X1 U18981 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15807) );
  AOI22_X1 U18982 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15806) );
  AOI22_X1 U18983 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15805) );
  AOI22_X1 U18984 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15804) );
  NAND4_X1 U18985 ( .A1(n15807), .A2(n15806), .A3(n15805), .A4(n15804), .ZN(
        n15814) );
  AOI22_X1 U18986 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U18987 ( .A1(n15869), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15811) );
  AOI22_X1 U18988 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15810) );
  AOI22_X1 U18989 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15809) );
  NAND4_X1 U18990 ( .A1(n15812), .A2(n15811), .A3(n15810), .A4(n15809), .ZN(
        n15813) );
  NOR2_X1 U18991 ( .A1(n15814), .A2(n15813), .ZN(n17071) );
  AOI22_X1 U18992 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15818) );
  AOI22_X1 U18993 ( .A1(n15826), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15817) );
  AOI22_X1 U18994 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15816) );
  AOI22_X1 U18995 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9773), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15815) );
  NAND4_X1 U18996 ( .A1(n15818), .A2(n15817), .A3(n15816), .A4(n15815), .ZN(
        n15825) );
  AOI22_X1 U18997 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15823) );
  AOI22_X1 U18998 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15822) );
  AOI22_X1 U18999 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15821) );
  AOI22_X1 U19000 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15820) );
  NAND4_X1 U19001 ( .A1(n15823), .A2(n15822), .A3(n15821), .A4(n15820), .ZN(
        n15824) );
  NOR2_X1 U19002 ( .A1(n15825), .A2(n15824), .ZN(n17080) );
  AOI22_X1 U19003 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15830) );
  AOI22_X1 U19004 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15829) );
  AOI22_X1 U19005 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15828) );
  AOI22_X1 U19006 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15827) );
  NAND4_X1 U19007 ( .A1(n15830), .A2(n15829), .A3(n15828), .A4(n15827), .ZN(
        n15836) );
  AOI22_X1 U19008 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15834) );
  AOI22_X1 U19009 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15833) );
  AOI22_X1 U19010 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15832) );
  AOI22_X1 U19011 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15831) );
  NAND4_X1 U19012 ( .A1(n15834), .A2(n15833), .A3(n15832), .A4(n15831), .ZN(
        n15835) );
  NOR2_X1 U19013 ( .A1(n15836), .A2(n15835), .ZN(n17089) );
  AOI22_X1 U19014 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17296), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17267), .ZN(n15840) );
  AOI22_X1 U19015 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17252), .ZN(n15839) );
  AOI22_X1 U19016 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17275), .ZN(n15838) );
  AOI22_X1 U19017 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n9773), .ZN(n15837) );
  NAND4_X1 U19018 ( .A1(n15840), .A2(n15839), .A3(n15838), .A4(n15837), .ZN(
        n15846) );
  AOI22_X1 U19019 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17268), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17270), .ZN(n15844) );
  AOI22_X1 U19020 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17288), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15843) );
  AOI22_X1 U19021 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17195), .B1(
        n17249), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15842) );
  AOI22_X1 U19022 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15841) );
  NAND4_X1 U19023 ( .A1(n15844), .A2(n15843), .A3(n15842), .A4(n15841), .ZN(
        n15845) );
  NOR2_X1 U19024 ( .A1(n15846), .A2(n15845), .ZN(n17090) );
  NOR2_X1 U19025 ( .A1(n17089), .A2(n17090), .ZN(n17088) );
  AOI22_X1 U19026 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15856) );
  AOI22_X1 U19027 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15855) );
  INV_X1 U19028 ( .A(n9822), .ZN(n15878) );
  AOI22_X1 U19029 ( .A1(n15826), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15847) );
  OAI21_X1 U19030 ( .B1(n10220), .B2(n18313), .A(n15847), .ZN(n15853) );
  AOI22_X1 U19031 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15851) );
  AOI22_X1 U19032 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15850) );
  AOI22_X1 U19033 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U19034 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15848) );
  NAND4_X1 U19035 ( .A1(n15851), .A2(n15850), .A3(n15849), .A4(n15848), .ZN(
        n15852) );
  AOI211_X1 U19036 ( .C1(n15878), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n15853), .B(n15852), .ZN(n15854) );
  NAND3_X1 U19037 ( .A1(n15856), .A2(n15855), .A3(n15854), .ZN(n17085) );
  NAND2_X1 U19038 ( .A1(n17088), .A2(n17085), .ZN(n17084) );
  NOR2_X1 U19039 ( .A1(n17080), .A2(n17084), .ZN(n17079) );
  AOI22_X1 U19040 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15867) );
  AOI22_X1 U19041 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15866) );
  INV_X1 U19042 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21082) );
  AOI22_X1 U19043 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15857) );
  OAI21_X1 U19044 ( .B1(n15858), .B2(n21082), .A(n15857), .ZN(n15864) );
  AOI22_X1 U19045 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15862) );
  AOI22_X1 U19046 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15861) );
  AOI22_X1 U19047 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15860) );
  AOI22_X1 U19048 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15859) );
  NAND4_X1 U19049 ( .A1(n15862), .A2(n15861), .A3(n15860), .A4(n15859), .ZN(
        n15863) );
  AOI211_X1 U19050 ( .C1(n17269), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n15864), .B(n15863), .ZN(n15865) );
  NAND3_X1 U19051 ( .A1(n15867), .A2(n15866), .A3(n15865), .ZN(n17076) );
  NAND2_X1 U19052 ( .A1(n17079), .A2(n17076), .ZN(n17075) );
  NOR2_X1 U19053 ( .A1(n17071), .A2(n17075), .ZN(n17070) );
  AOI22_X1 U19054 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17296), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15881) );
  AOI22_X1 U19055 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15880) );
  INV_X1 U19056 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15893) );
  AOI22_X1 U19057 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15870) );
  OAI21_X1 U19058 ( .B1(n16967), .B2(n15893), .A(n15870), .ZN(n15877) );
  AOI22_X1 U19059 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15875) );
  AOI22_X1 U19060 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15874) );
  AOI22_X1 U19061 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15873) );
  AOI22_X1 U19062 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15872) );
  NAND4_X1 U19063 ( .A1(n15875), .A2(n15874), .A3(n15873), .A4(n15872), .ZN(
        n15876) );
  AOI211_X1 U19064 ( .C1(n15878), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15877), .B(n15876), .ZN(n15879) );
  NAND3_X1 U19065 ( .A1(n15881), .A2(n15880), .A3(n15879), .ZN(n15882) );
  NAND2_X1 U19066 ( .A1(n17070), .A2(n15882), .ZN(n17064) );
  OAI21_X1 U19067 ( .B1(n17070), .B2(n15882), .A(n17064), .ZN(n17357) );
  NAND2_X1 U19068 ( .A1(n18343), .A2(n18326), .ZN(n15884) );
  NAND2_X1 U19069 ( .A1(n15883), .A2(n18749), .ZN(n15917) );
  OAI21_X1 U19070 ( .B1(n15885), .B2(n15884), .A(n15917), .ZN(n16009) );
  NAND4_X1 U19071 ( .A1(n18955), .A2(n15915), .A3(n17492), .A4(n16009), .ZN(
        n15888) );
  AND2_X1 U19072 ( .A1(n17337), .A2(n17459), .ZN(n17334) );
  INV_X2 U19073 ( .A(n17334), .ZN(n17329) );
  INV_X1 U19074 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17159) );
  INV_X1 U19075 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17188) );
  NAND2_X1 U19076 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17010) );
  INV_X1 U19077 ( .A(n17010), .ZN(n17326) );
  AND2_X1 U19078 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17326), .ZN(n17319) );
  NAND3_X1 U19079 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17319), .ZN(n17318) );
  NAND2_X1 U19080 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17309) );
  NAND2_X1 U19081 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n17244) );
  NAND2_X1 U19082 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .ZN(n17245) );
  NOR4_X1 U19083 ( .A1(n16883), .A2(n17309), .A3(n17244), .A4(n17245), .ZN(
        n15889) );
  INV_X1 U19084 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17216) );
  INV_X1 U19085 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n15890) );
  NOR3_X1 U19086 ( .A1(n17216), .A2(n17215), .A3(n15890), .ZN(n17202) );
  NAND3_X1 U19087 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n15889), .A3(n17202), 
        .ZN(n17187) );
  NOR3_X1 U19088 ( .A1(n17188), .A2(n17318), .A3(n17187), .ZN(n17172) );
  NAND3_X1 U19089 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17337), .A3(n17172), 
        .ZN(n17148) );
  NOR2_X1 U19090 ( .A1(n17159), .A2(n17148), .ZN(n17146) );
  NAND2_X1 U19091 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17146), .ZN(n17145) );
  NOR2_X1 U19092 ( .A1(n17459), .A2(n17145), .ZN(n17132) );
  NAND2_X1 U19093 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17132), .ZN(n17120) );
  NOR2_X1 U19094 ( .A1(n16767), .A2(n17120), .ZN(n17094) );
  NAND2_X1 U19095 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17083), .ZN(n17069) );
  INV_X1 U19096 ( .A(n17069), .ZN(n17078) );
  INV_X1 U19097 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n21212) );
  INV_X1 U19098 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17074) );
  NOR2_X1 U19099 ( .A1(n21212), .A2(n17074), .ZN(n17062) );
  NAND2_X1 U19100 ( .A1(n18343), .A2(n17337), .ZN(n17331) );
  OAI22_X1 U19101 ( .A1(n17334), .A2(n17078), .B1(n17062), .B2(n17331), .ZN(
        n17066) );
  NOR3_X1 U19102 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17074), .A3(n17069), .ZN(
        n15886) );
  AOI21_X1 U19103 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17066), .A(n15886), .ZN(
        n15887) );
  OAI21_X1 U19104 ( .B1(n17357), .B2(n17329), .A(n15887), .ZN(P3_U2675) );
  NOR2_X1 U19105 ( .A1(n15888), .A2(n17318), .ZN(n17315) );
  NAND2_X1 U19106 ( .A1(n15889), .A2(n17315), .ZN(n17246) );
  NOR3_X1 U19107 ( .A1(n17459), .A2(n15890), .A3(n17246), .ZN(n15905) );
  NOR2_X1 U19108 ( .A1(n17334), .A2(n15905), .ZN(n17231) );
  INV_X1 U19109 ( .A(n17231), .ZN(n15907) );
  AOI22_X1 U19110 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15904) );
  AOI22_X1 U19111 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15903) );
  AOI22_X1 U19112 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15892) );
  OAI21_X1 U19113 ( .B1(n9850), .B2(n15893), .A(n15892), .ZN(n15901) );
  AOI22_X1 U19114 ( .A1(n15894), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15899) );
  AOI22_X1 U19115 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15898) );
  AOI22_X1 U19116 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15895), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15897) );
  AOI22_X1 U19117 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15896) );
  NAND4_X1 U19118 ( .A1(n15899), .A2(n15898), .A3(n15897), .A4(n15896), .ZN(
        n15900) );
  AOI211_X1 U19119 ( .C1(n17269), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n15901), .B(n15900), .ZN(n15902) );
  NAND3_X1 U19120 ( .A1(n15904), .A2(n15903), .A3(n15902), .ZN(n17432) );
  AOI22_X1 U19121 ( .A1(n17334), .A2(n17432), .B1(n15905), .B2(n17215), .ZN(
        n15906) );
  OAI21_X1 U19122 ( .B1(n17215), .B2(n15907), .A(n15906), .ZN(P3_U2690) );
  NAND3_X1 U19123 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n18909)
         );
  NAND2_X1 U19124 ( .A1(n15922), .A2(n16966), .ZN(n15908) );
  NOR2_X1 U19125 ( .A1(n17296), .A2(n15908), .ZN(n18799) );
  INV_X1 U19126 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16655) );
  INV_X1 U19127 ( .A(n18661), .ZN(n18410) );
  OAI221_X1 U19128 ( .B1(n18909), .B2(n18799), .C1(n18909), .C2(n16655), .A(
        n18410), .ZN(n20995) );
  NAND2_X1 U19129 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n20991), .ZN(n20989) );
  NAND2_X1 U19130 ( .A1(n20995), .A2(n20989), .ZN(n15911) );
  INV_X1 U19131 ( .A(n15911), .ZN(n15910) );
  INV_X1 U19132 ( .A(n18601), .ZN(n18659) );
  INV_X1 U19133 ( .A(n17864), .ZN(n17923) );
  OAI22_X1 U19134 ( .A1(n20992), .A2(n17923), .B1(n20991), .B2(n18910), .ZN(
        n15913) );
  NAND3_X1 U19135 ( .A1(n18579), .A2(n20995), .A3(n15913), .ZN(n15909) );
  OAI221_X1 U19136 ( .B1(n18579), .B2(n15910), .C1(n18579), .C2(n18659), .A(
        n15909), .ZN(P3_U2864) );
  NAND2_X1 U19137 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18528) );
  NOR2_X1 U19138 ( .A1(n20992), .A2(n17923), .ZN(n15912) );
  AOI221_X1 U19139 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18528), .C1(n15912), 
        .C2(n18528), .A(n15911), .ZN(n18301) );
  OAI221_X1 U19140 ( .B1(n18601), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18601), .C2(n15913), .A(n20995), .ZN(n18299) );
  AOI22_X1 U19141 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18301), .B1(
        n18299), .B2(n18298), .ZN(P3_U2865) );
  INV_X1 U19142 ( .A(n9764), .ZN(n15914) );
  NAND2_X1 U19143 ( .A1(n18746), .A2(n18962), .ZN(n15919) );
  NOR2_X1 U19144 ( .A1(n15915), .A2(n15914), .ZN(n18798) );
  OAI21_X1 U19145 ( .B1(n15916), .B2(n18798), .A(n18822), .ZN(n17491) );
  OAI211_X1 U19146 ( .C1(n15919), .C2(n17491), .A(n15918), .B(n15917), .ZN(
        n15920) );
  NOR2_X1 U19147 ( .A1(n16011), .A2(n15920), .ZN(n18783) );
  INV_X1 U19148 ( .A(n18783), .ZN(n18782) );
  OAI22_X1 U19149 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18910), .B1(n18909), 
        .B2(n16655), .ZN(n15921) );
  AOI21_X1 U19150 ( .B1(n18955), .B2(n18782), .A(n15921), .ZN(n18941) );
  INV_X1 U19151 ( .A(n18941), .ZN(n18939) );
  AOI21_X1 U19152 ( .B1(n15922), .B2(n16966), .A(n18747), .ZN(n18756) );
  NAND3_X1 U19153 ( .A1(n18939), .A2(n18974), .A3(n18756), .ZN(n15923) );
  OAI21_X1 U19154 ( .B1(n18939), .B2(n16966), .A(n15923), .ZN(P3_U3284) );
  OAI22_X1 U19155 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17838), .B1(
        n15925), .B2(n15924), .ZN(n15926) );
  XNOR2_X1 U19156 ( .A(n16518), .B(n15926), .ZN(n16531) );
  AOI21_X1 U19157 ( .B1(n18181), .B2(n17622), .A(n15927), .ZN(n16549) );
  INV_X1 U19158 ( .A(n15928), .ZN(n18754) );
  NAND2_X1 U19159 ( .A1(n18754), .A2(n18288), .ZN(n18224) );
  NOR3_X1 U19160 ( .A1(n16517), .A2(n16534), .A3(n18224), .ZN(n15929) );
  AOI21_X1 U19161 ( .B1(n18292), .B2(n16528), .A(n15929), .ZN(n15984) );
  NAND2_X1 U19162 ( .A1(n18283), .A2(n16551), .ZN(n15930) );
  OAI211_X1 U19163 ( .C1(n9768), .C2(n16549), .A(n15984), .B(n15930), .ZN(
        n15935) );
  INV_X1 U19164 ( .A(n16527), .ZN(n15933) );
  INV_X1 U19165 ( .A(n18204), .ZN(n18106) );
  OAI21_X1 U19166 ( .B1(n18106), .B2(n17974), .A(n15931), .ZN(n15932) );
  AOI22_X1 U19167 ( .A1(n17976), .A2(n18292), .B1(n18288), .B2(n15932), .ZN(
        n15991) );
  OAI21_X1 U19168 ( .B1(n15933), .B2(n15991), .A(n16518), .ZN(n15934) );
  OAI21_X1 U19169 ( .B1(n16518), .B2(n15935), .A(n15934), .ZN(n15936) );
  NAND2_X1 U19170 ( .A1(n9768), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16521) );
  OAI211_X1 U19171 ( .C1(n18200), .C2(n16531), .A(n15936), .B(n16521), .ZN(
        P3_U2833) );
  OR2_X1 U19172 ( .A1(n15938), .A2(n15937), .ZN(n15944) );
  AOI21_X1 U19173 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15940), .A(
        n15939), .ZN(n15941) );
  AOI22_X1 U19174 ( .A1(n15944), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n15941), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15942) );
  INV_X1 U19175 ( .A(n15942), .ZN(n15943) );
  OAI21_X1 U19176 ( .B1(n15944), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15943), .ZN(n15946) );
  OAI22_X1 U19177 ( .A1(n15946), .A2(n20611), .B1(n15947), .B2(n20652), .ZN(
        n15950) );
  AOI21_X1 U19178 ( .B1(n15946), .B2(n20611), .A(n15945), .ZN(n15949) );
  INV_X1 U19179 ( .A(n15947), .ZN(n15948) );
  OAI22_X1 U19180 ( .A1(n15950), .A2(n15949), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15948), .ZN(n15959) );
  INV_X1 U19181 ( .A(n15951), .ZN(n15955) );
  OAI21_X1 U19182 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15952), .ZN(n15953) );
  NAND4_X1 U19183 ( .A1(n15956), .A2(n15955), .A3(n15954), .A4(n15953), .ZN(
        n15957) );
  AOI211_X1 U19184 ( .C1(n15959), .C2(n20250), .A(n15958), .B(n15957), .ZN(
        n15975) );
  INV_X1 U19185 ( .A(n15975), .ZN(n15966) );
  NAND2_X1 U19186 ( .A1(n15961), .A2(n15960), .ZN(n15964) );
  NOR3_X1 U19187 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20888), .A3(n20978), 
        .ZN(n15962) );
  OAI22_X1 U19188 ( .A1(n15965), .A2(n15964), .B1(n15963), .B2(n15962), .ZN(
        n16323) );
  AOI221_X1 U19189 ( .B1(n20885), .B2(n20884), .C1(n15966), .C2(n20884), .A(
        n16323), .ZN(n16325) );
  INV_X1 U19190 ( .A(n20983), .ZN(n16321) );
  NOR2_X1 U19191 ( .A1(n16321), .A2(n15967), .ZN(n15968) );
  NOR2_X1 U19192 ( .A1(n16325), .A2(n15968), .ZN(n15973) );
  INV_X1 U19193 ( .A(n16320), .ZN(n15969) );
  AOI211_X1 U19194 ( .C1(n20890), .C2(n20888), .A(n15970), .B(n15969), .ZN(
        n15971) );
  NAND2_X1 U19195 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15971), .ZN(n15972) );
  OAI22_X1 U19196 ( .A1(n15973), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n16325), 
        .B2(n15972), .ZN(n15974) );
  OAI21_X1 U19197 ( .B1(n15975), .B2(n20012), .A(n15974), .ZN(P1_U3161) );
  AOI22_X1 U19198 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16191), .B1(
        n20236), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15982) );
  NOR3_X1 U19199 ( .A1(n15976), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16134), .ZN(n15977) );
  AOI21_X1 U19200 ( .B1(n15978), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15977), .ZN(n15979) );
  XNOR2_X1 U19201 ( .A(n15979), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16098) );
  AOI22_X1 U19202 ( .A1(n16098), .A2(n20243), .B1(n16195), .B2(n15980), .ZN(
        n15981) );
  OAI211_X1 U19203 ( .C1(n20230), .C2(n16039), .A(n15982), .B(n15981), .ZN(
        P1_U3010) );
  AOI21_X1 U19204 ( .B1(n15985), .B2(n15984), .A(n15983), .ZN(n15986) );
  AOI21_X1 U19205 ( .B1(n9895), .B2(n15987), .A(n15986), .ZN(n15989) );
  OAI211_X1 U19206 ( .C1(n15991), .C2(n15990), .A(n15989), .B(n15988), .ZN(
        P3_U2832) );
  INV_X1 U19207 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20894) );
  INV_X1 U19208 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20898) );
  NOR2_X1 U19209 ( .A1(n20897), .A2(n20898), .ZN(n15992) );
  INV_X1 U19210 ( .A(HOLD), .ZN(n20902) );
  INV_X1 U19211 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20905) );
  OAI222_X1 U19212 ( .A1(n15992), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n15992), 
        .B2(HOLD), .C1(n20902), .C2(n20905), .ZN(n15994) );
  OAI211_X1 U19213 ( .C1(n20978), .C2(n20894), .A(n15994), .B(n15993), .ZN(
        P1_U3195) );
  INV_X1 U19214 ( .A(n15995), .ZN(n15998) );
  INV_X1 U19215 ( .A(n15996), .ZN(n16199) );
  AOI221_X1 U19216 ( .B1(n15999), .B2(n15998), .C1(n15997), .C2(n15998), .A(
        n16199), .ZN(n16005) );
  AOI21_X1 U19217 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16200), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16004) );
  AOI22_X1 U19218 ( .A1(n16001), .A2(n20243), .B1(n20238), .B2(n16000), .ZN(
        n16003) );
  OAI211_X1 U19219 ( .C1(n16005), .C2(n16004), .A(n16003), .B(n16002), .ZN(
        P1_U3011) );
  NOR3_X1 U19220 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16007) );
  NOR2_X1 U19221 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16006) );
  AND2_X1 U19222 ( .A1(n19996), .A2(n18982), .ZN(n16505) );
  NOR4_X1 U19223 ( .A1(n16007), .A2(n16006), .A3(n16505), .A4(n16507), .ZN(
        P2_U3178) );
  INV_X1 U19224 ( .A(n19977), .ZN(n19974) );
  NOR2_X1 U19225 ( .A1(n16008), .A2(n19974), .ZN(P2_U3047) );
  OAI221_X1 U19226 ( .B1(n16011), .B2(n16010), .C1(n16011), .C2(n16009), .A(
        n18955), .ZN(n16012) );
  INV_X1 U19227 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17561) );
  INV_X1 U19228 ( .A(n16012), .ZN(n17340) );
  NAND2_X1 U19229 ( .A1(n18343), .A2(n17340), .ZN(n17385) );
  NAND2_X1 U19230 ( .A1(n16013), .A2(n17340), .ZN(n17483) );
  INV_X1 U19231 ( .A(n17483), .ZN(n17485) );
  NAND2_X1 U19232 ( .A1(n16014), .A2(n17340), .ZN(n17480) );
  AOI22_X1 U19233 ( .A1(n17485), .A2(BUF2_REG_0__SCAN_IN), .B1(n17484), .B2(
        n17959), .ZN(n16015) );
  OAI221_X1 U19234 ( .B1(n17488), .B2(n17561), .C1(n17488), .C2(n17385), .A(
        n16015), .ZN(P3_U2735) );
  AOI22_X1 U19235 ( .A1(n20071), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20051), .ZN(n16025) );
  OAI22_X1 U19236 ( .A1(n16183), .A2(n20061), .B1(n16088), .B2(n20107), .ZN(
        n16017) );
  AOI21_X1 U19237 ( .B1(n16085), .B2(n20066), .A(n16017), .ZN(n16024) );
  OAI21_X1 U19238 ( .B1(n16019), .B2(n16018), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n16023) );
  INV_X1 U19239 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21204) );
  NAND3_X1 U19240 ( .A1(n16021), .A2(n21204), .A3(n16020), .ZN(n16022) );
  NAND4_X1 U19241 ( .A1(n16025), .A2(n16024), .A3(n16023), .A4(n16022), .ZN(
        P1_U2815) );
  AOI21_X1 U19242 ( .B1(n16027), .B2(n16026), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n16031) );
  AOI22_X1 U19243 ( .A1(n20071), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20051), .ZN(n16030) );
  OAI22_X1 U19244 ( .A1(n16190), .A2(n20061), .B1(n20107), .B2(n16096), .ZN(
        n16028) );
  AOI21_X1 U19245 ( .B1(n16093), .B2(n20066), .A(n16028), .ZN(n16029) );
  OAI211_X1 U19246 ( .C1(n16032), .C2(n16031), .A(n16030), .B(n16029), .ZN(
        P1_U2817) );
  INV_X1 U19247 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16043) );
  NOR3_X1 U19248 ( .A1(n20101), .A2(n16033), .A3(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n16036) );
  INV_X1 U19249 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20937) );
  NOR2_X1 U19250 ( .A1(n16034), .A2(n20937), .ZN(n16035) );
  AOI211_X1 U19251 ( .C1(n20071), .C2(P1_EBX_REG_21__SCAN_IN), .A(n16036), .B(
        n16035), .ZN(n16042) );
  INV_X1 U19252 ( .A(n16101), .ZN(n16037) );
  NAND2_X1 U19253 ( .A1(n20039), .A2(n16037), .ZN(n16038) );
  OAI21_X1 U19254 ( .B1(n16039), .B2(n20061), .A(n16038), .ZN(n16040) );
  AOI21_X1 U19255 ( .B1(n16097), .B2(n20066), .A(n16040), .ZN(n16041) );
  OAI211_X1 U19256 ( .C1(n16043), .C2(n20093), .A(n16042), .B(n16041), .ZN(
        P1_U2819) );
  OAI22_X1 U19257 ( .A1(n20094), .A2(n16045), .B1(n16044), .B2(n20093), .ZN(
        n16046) );
  AOI211_X1 U19258 ( .C1(n20039), .C2(n16114), .A(n20050), .B(n16046), .ZN(
        n16051) );
  INV_X1 U19259 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20929) );
  OAI21_X1 U19260 ( .B1(n16047), .B2(n16054), .A(n20929), .ZN(n16049) );
  AOI22_X1 U19261 ( .A1(n16115), .A2(n20066), .B1(n16049), .B2(n16048), .ZN(
        n16050) );
  OAI211_X1 U19262 ( .C1(n20061), .C2(n16217), .A(n16051), .B(n16050), .ZN(
        P1_U2823) );
  INV_X1 U19263 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16052) );
  OAI21_X1 U19264 ( .B1(n20093), .B2(n16052), .A(n20091), .ZN(n16056) );
  OAI22_X1 U19265 ( .A1(n16054), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n16053), 
        .B2(n20094), .ZN(n16055) );
  AOI211_X1 U19266 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16057), .A(n16056), 
        .B(n16055), .ZN(n16059) );
  AOI22_X1 U19267 ( .A1(n16125), .A2(n20066), .B1(n20039), .B2(n16124), .ZN(
        n16058) );
  OAI211_X1 U19268 ( .C1(n20061), .C2(n16231), .A(n16059), .B(n16058), .ZN(
        P1_U2825) );
  NOR2_X1 U19269 ( .A1(n20101), .A2(n16060), .ZN(n16067) );
  AOI21_X1 U19270 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16067), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16065) );
  OAI22_X1 U19271 ( .A1(n20094), .A2(n16077), .B1(n16061), .B2(n20093), .ZN(
        n16062) );
  AOI211_X1 U19272 ( .C1(n16075), .C2(n20099), .A(n20050), .B(n16062), .ZN(
        n16064) );
  AOI22_X1 U19273 ( .A1(n16129), .A2(n20039), .B1(n20066), .B2(n16128), .ZN(
        n16063) );
  OAI211_X1 U19274 ( .C1(n16066), .C2(n16065), .A(n16064), .B(n16063), .ZN(
        P1_U2828) );
  INV_X1 U19275 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21111) );
  AOI22_X1 U19276 ( .A1(n16067), .A2(n21111), .B1(n20071), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16074) );
  XOR2_X1 U19277 ( .A(n16069), .B(n16068), .Z(n16255) );
  AOI22_X1 U19278 ( .A1(n20099), .A2(n16255), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n16070), .ZN(n16071) );
  OAI211_X1 U19279 ( .C1(n20093), .C2(n12162), .A(n16071), .B(n20091), .ZN(
        n16072) );
  AOI21_X1 U19280 ( .B1(n20066), .B2(n16139), .A(n16072), .ZN(n16073) );
  OAI211_X1 U19281 ( .C1(n16142), .C2(n20107), .A(n16074), .B(n16073), .ZN(
        P1_U2829) );
  AOI22_X1 U19282 ( .A1(n16128), .A2(n20113), .B1(n20112), .B2(n16075), .ZN(
        n16076) );
  OAI21_X1 U19283 ( .B1(n20115), .B2(n16077), .A(n16076), .ZN(P1_U2860) );
  AOI22_X1 U19284 ( .A1(n16139), .A2(n20113), .B1(n20112), .B2(n16255), .ZN(
        n16078) );
  OAI21_X1 U19285 ( .B1(n20115), .B2(n16079), .A(n16078), .ZN(P1_U2861) );
  AOI22_X1 U19286 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n16087) );
  MUX2_X1 U19287 ( .A(n12813), .B(n16080), .S(n16121), .Z(n16081) );
  AOI21_X1 U19288 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16082), .A(
        n16081), .ZN(n16084) );
  XNOR2_X1 U19289 ( .A(n16084), .B(n16083), .ZN(n16180) );
  AOI22_X1 U19290 ( .A1(n16180), .A2(n20186), .B1(n20194), .B2(n16085), .ZN(
        n16086) );
  OAI211_X1 U19291 ( .C1(n20179), .C2(n16088), .A(n16087), .B(n16086), .ZN(
        P1_U2974) );
  AOI22_X1 U19292 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16095) );
  MUX2_X1 U19293 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n16089), .S(
        n16121), .Z(n16091) );
  NAND2_X1 U19294 ( .A1(n16134), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16090) );
  MUX2_X1 U19295 ( .A(n16091), .B(n16090), .S(n14884), .Z(n16092) );
  OAI21_X1 U19296 ( .B1(n16080), .B2(n16134), .A(n16092), .ZN(n16188) );
  AOI22_X1 U19297 ( .A1(n16188), .A2(n20186), .B1(n20194), .B2(n16093), .ZN(
        n16094) );
  OAI211_X1 U19298 ( .C1(n20179), .C2(n16096), .A(n16095), .B(n16094), .ZN(
        P1_U2976) );
  AOI22_X1 U19299 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16100) );
  AOI22_X1 U19300 ( .A1(n16098), .A2(n20186), .B1(n20194), .B2(n16097), .ZN(
        n16099) );
  OAI211_X1 U19301 ( .C1(n20179), .C2(n16101), .A(n16100), .B(n16099), .ZN(
        P1_U2978) );
  AOI22_X1 U19302 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16107) );
  MUX2_X1 U19303 ( .A(n16102), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n16121), .Z(n16103) );
  XNOR2_X1 U19304 ( .A(n16104), .B(n16103), .ZN(n16201) );
  AOI22_X1 U19305 ( .A1(n16201), .A2(n20186), .B1(n20194), .B2(n16105), .ZN(
        n16106) );
  OAI211_X1 U19306 ( .C1(n20179), .C2(n16108), .A(n16107), .B(n16106), .ZN(
        P1_U2980) );
  NOR2_X1 U19307 ( .A1(n16134), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16112) );
  AOI21_X1 U19308 ( .B1(n16110), .B2(n16133), .A(n16109), .ZN(n16111) );
  MUX2_X1 U19309 ( .A(n16112), .B(n16134), .S(n16111), .Z(n16113) );
  XNOR2_X1 U19310 ( .A(n16113), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16218) );
  AOI22_X1 U19311 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16117) );
  AOI22_X1 U19312 ( .A1(n16115), .A2(n20194), .B1(n16114), .B2(n20185), .ZN(
        n16116) );
  OAI211_X1 U19313 ( .C1(n16218), .C2(n20198), .A(n16117), .B(n16116), .ZN(
        P1_U2982) );
  NAND2_X1 U19314 ( .A1(n16119), .A2(n16118), .ZN(n16123) );
  AOI21_X1 U19315 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16121), .A(
        n16120), .ZN(n16122) );
  XNOR2_X1 U19316 ( .A(n16123), .B(n16122), .ZN(n16232) );
  AOI22_X1 U19317 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16127) );
  AOI22_X1 U19318 ( .A1(n16125), .A2(n20194), .B1(n20185), .B2(n16124), .ZN(
        n16126) );
  OAI211_X1 U19319 ( .C1(n16232), .C2(n20198), .A(n16127), .B(n16126), .ZN(
        P1_U2984) );
  AOI22_X1 U19320 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16131) );
  AOI22_X1 U19321 ( .A1(n20185), .A2(n16129), .B1(n20194), .B2(n16128), .ZN(
        n16130) );
  OAI211_X1 U19322 ( .C1(n16132), .C2(n20198), .A(n16131), .B(n16130), .ZN(
        P1_U2987) );
  AOI22_X1 U19323 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16141) );
  NOR2_X1 U19324 ( .A1(n14967), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16136) );
  NOR2_X1 U19325 ( .A1(n16133), .A2(n12778), .ZN(n16135) );
  MUX2_X1 U19326 ( .A(n16136), .B(n16135), .S(n16134), .Z(n16138) );
  XNOR2_X1 U19327 ( .A(n16138), .B(n16137), .ZN(n16257) );
  AOI22_X1 U19328 ( .A1(n20186), .A2(n16257), .B1(n20194), .B2(n16139), .ZN(
        n16140) );
  OAI211_X1 U19329 ( .C1(n20179), .C2(n16142), .A(n16141), .B(n16140), .ZN(
        P1_U2988) );
  NAND2_X1 U19330 ( .A1(n16144), .A2(n16145), .ZN(n16146) );
  NAND2_X1 U19331 ( .A1(n16143), .A2(n16146), .ZN(n16289) );
  OAI22_X1 U19332 ( .A1(n20052), .A2(n20258), .B1(n20059), .B2(n20179), .ZN(
        n16147) );
  AOI21_X1 U19333 ( .B1(n16289), .B2(n20186), .A(n16147), .ZN(n16148) );
  NAND2_X1 U19334 ( .A1(n20236), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n16295) );
  OAI211_X1 U19335 ( .C1(n16149), .C2(n20190), .A(n16148), .B(n16295), .ZN(
        P1_U2992) );
  AOI22_X1 U19336 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16155) );
  XNOR2_X1 U19337 ( .A(n16151), .B(n16150), .ZN(n16152) );
  XNOR2_X1 U19338 ( .A(n16153), .B(n16152), .ZN(n16303) );
  AOI22_X1 U19339 ( .A1(n16303), .A2(n20186), .B1(n20194), .B2(n20109), .ZN(
        n16154) );
  OAI211_X1 U19340 ( .C1(n20179), .C2(n20070), .A(n16155), .B(n16154), .ZN(
        P1_U2993) );
  AOI22_X1 U19341 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16161) );
  OAI21_X1 U19342 ( .B1(n16158), .B2(n16157), .A(n16156), .ZN(n16159) );
  INV_X1 U19343 ( .A(n16159), .ZN(n16308) );
  AOI22_X1 U19344 ( .A1(n16308), .A2(n20186), .B1(n20194), .B2(n20082), .ZN(
        n16160) );
  OAI211_X1 U19345 ( .C1(n20179), .C2(n20084), .A(n16161), .B(n16160), .ZN(
        P1_U2994) );
  NAND2_X1 U19346 ( .A1(n20236), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16165) );
  NAND2_X1 U19347 ( .A1(n16163), .A2(n9809), .ZN(n16164) );
  OAI211_X1 U19348 ( .C1(n16166), .C2(n9809), .A(n16165), .B(n16164), .ZN(
        n16167) );
  AOI21_X1 U19349 ( .B1(n9808), .B2(n20243), .A(n16167), .ZN(n16168) );
  OAI21_X1 U19350 ( .B1(n20230), .B2(n16169), .A(n16168), .ZN(P1_U3004) );
  AOI22_X1 U19351 ( .A1(n16171), .A2(n20243), .B1(n20238), .B2(n16170), .ZN(
        n16177) );
  NOR3_X1 U19352 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n16172), .A3(
        n16186), .ZN(n16178) );
  INV_X1 U19353 ( .A(n16173), .ZN(n16174) );
  OAI22_X1 U19354 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16175), .B1(
        n16178), .B2(n16174), .ZN(n16176) );
  OAI211_X1 U19355 ( .C1(n20944), .C2(n16230), .A(n16177), .B(n16176), .ZN(
        P1_U3005) );
  AOI21_X1 U19356 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n20236), .A(n16178), 
        .ZN(n16182) );
  AOI22_X1 U19357 ( .A1(n16180), .A2(n20243), .B1(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16179), .ZN(n16181) );
  OAI211_X1 U19358 ( .C1(n20230), .C2(n16183), .A(n16182), .B(n16181), .ZN(
        P1_U3006) );
  NAND2_X1 U19359 ( .A1(n20236), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n16184) );
  OAI221_X1 U19360 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16186), 
        .C1(n16089), .C2(n16185), .A(n16184), .ZN(n16187) );
  AOI21_X1 U19361 ( .B1(n16188), .B2(n20243), .A(n16187), .ZN(n16189) );
  OAI21_X1 U19362 ( .B1(n20230), .B2(n16190), .A(n16189), .ZN(P1_U3008) );
  AOI22_X1 U19363 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16191), .B1(
        n20236), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16198) );
  AOI22_X1 U19364 ( .A1(n16193), .A2(n20243), .B1(n20238), .B2(n16192), .ZN(
        n16197) );
  OAI211_X1 U19365 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16195), .B(n16194), .ZN(
        n16196) );
  NAND3_X1 U19366 ( .A1(n16198), .A2(n16197), .A3(n16196), .ZN(P1_U3009) );
  AOI22_X1 U19367 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16199), .B1(
        n20236), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16203) );
  AOI22_X1 U19368 ( .A1(n16201), .A2(n20243), .B1(n16102), .B2(n16200), .ZN(
        n16202) );
  OAI211_X1 U19369 ( .C1(n20230), .C2(n16204), .A(n16203), .B(n16202), .ZN(
        P1_U3012) );
  NAND2_X1 U19370 ( .A1(n16223), .A2(n16208), .ZN(n16214) );
  OAI21_X1 U19371 ( .B1(n12903), .B2(n16239), .A(n20219), .ZN(n16205) );
  OAI211_X1 U19372 ( .C1(n16207), .C2(n20205), .A(n16206), .B(n16205), .ZN(
        n16241) );
  AOI21_X1 U19373 ( .B1(n16263), .B2(n16215), .A(n16241), .ZN(n16222) );
  OAI22_X1 U19374 ( .A1(n16209), .A2(n16291), .B1(n16222), .B2(n16208), .ZN(
        n16210) );
  AOI21_X1 U19375 ( .B1(n20238), .B2(n16211), .A(n16210), .ZN(n16213) );
  NAND2_X1 U19376 ( .A1(n20236), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16212) );
  OAI211_X1 U19377 ( .C1(n16215), .C2(n16214), .A(n16213), .B(n16212), .ZN(
        P1_U3013) );
  NOR3_X1 U19378 ( .A1(n14945), .A2(n16224), .A3(n12775), .ZN(n16216) );
  AOI21_X1 U19379 ( .B1(n16216), .B2(n16223), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16221) );
  OAI22_X1 U19380 ( .A1(n16218), .A2(n16291), .B1(n20230), .B2(n16217), .ZN(
        n16219) );
  AOI21_X1 U19381 ( .B1(n20236), .B2(P1_REIP_REG_17__SCAN_IN), .A(n16219), 
        .ZN(n16220) );
  OAI21_X1 U19382 ( .B1(n16222), .B2(n16221), .A(n16220), .ZN(P1_U3014) );
  NAND2_X1 U19383 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16223), .ZN(
        n16237) );
  AOI22_X1 U19384 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n12775), .B1(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16224), .ZN(n16229) );
  INV_X1 U19385 ( .A(n16241), .ZN(n16249) );
  OAI21_X1 U19386 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n20239), .A(
        n16249), .ZN(n16235) );
  AOI22_X1 U19387 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16235), .B1(
        n20236), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16228) );
  AOI22_X1 U19388 ( .A1(n16226), .A2(n20243), .B1(n20238), .B2(n16225), .ZN(
        n16227) );
  OAI211_X1 U19389 ( .C1(n16237), .C2(n16229), .A(n16228), .B(n16227), .ZN(
        P1_U3015) );
  INV_X1 U19390 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20927) );
  NOR2_X1 U19391 ( .A1(n16230), .A2(n20927), .ZN(n16234) );
  OAI22_X1 U19392 ( .A1(n16232), .A2(n16291), .B1(n20230), .B2(n16231), .ZN(
        n16233) );
  AOI211_X1 U19393 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16235), .A(
        n16234), .B(n16233), .ZN(n16236) );
  OAI21_X1 U19394 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16237), .A(
        n16236), .ZN(P1_U3016) );
  NAND2_X1 U19395 ( .A1(n16238), .A2(n16302), .ZN(n16260) );
  NOR2_X1 U19396 ( .A1(n12903), .A2(n16239), .ZN(n16240) );
  NAND2_X1 U19397 ( .A1(n16240), .A2(n14945), .ZN(n16247) );
  AOI22_X1 U19398 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16241), .B1(
        n20236), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16246) );
  INV_X1 U19399 ( .A(n16242), .ZN(n16244) );
  AOI22_X1 U19400 ( .A1(n16244), .A2(n20243), .B1(n20238), .B2(n16243), .ZN(
        n16245) );
  OAI211_X1 U19401 ( .C1(n16260), .C2(n16247), .A(n16246), .B(n16245), .ZN(
        P1_U3017) );
  NAND2_X1 U19402 ( .A1(n20236), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16248) );
  OAI221_X1 U19403 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16250), 
        .C1(n12903), .C2(n16249), .A(n16248), .ZN(n16251) );
  AOI21_X1 U19404 ( .B1(n16252), .B2(n20243), .A(n16251), .ZN(n16253) );
  OAI21_X1 U19405 ( .B1(n20230), .B2(n16254), .A(n16253), .ZN(P1_U3018) );
  AOI22_X1 U19406 ( .A1(n20236), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20238), 
        .B2(n16255), .ZN(n16259) );
  AOI22_X1 U19407 ( .A1(n16257), .A2(n20243), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16256), .ZN(n16258) );
  OAI211_X1 U19408 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16260), .A(
        n16259), .B(n16258), .ZN(P1_U3020) );
  AOI21_X1 U19409 ( .B1(n16283), .B2(n16281), .A(n16261), .ZN(n16264) );
  AOI221_X1 U19410 ( .B1(n16264), .B2(n16263), .C1(n16262), .C2(n16263), .A(
        n20218), .ZN(n16274) );
  AOI22_X1 U19411 ( .A1(n20236), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n20238), 
        .B2(n16265), .ZN(n16270) );
  INV_X1 U19412 ( .A(n16266), .ZN(n16268) );
  NAND4_X1 U19413 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16302), .ZN(n16276) );
  AOI221_X1 U19414 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12778), .C2(n16275), .A(
        n16276), .ZN(n16267) );
  AOI21_X1 U19415 ( .B1(n16268), .B2(n20243), .A(n16267), .ZN(n16269) );
  OAI211_X1 U19416 ( .C1(n12778), .C2(n16274), .A(n16270), .B(n16269), .ZN(
        P1_U3021) );
  AOI222_X1 U19417 ( .A1(n16272), .A2(n20243), .B1(n20238), .B2(n16271), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(n20236), .ZN(n16273) );
  OAI221_X1 U19418 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16276), .C1(
        n16275), .C2(n16274), .A(n16273), .ZN(P1_U3022) );
  NAND2_X1 U19419 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16302), .ZN(
        n16290) );
  NAND2_X1 U19420 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16277) );
  OAI21_X1 U19421 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16277), .ZN(n16288) );
  AOI22_X1 U19422 ( .A1(n20236), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n20238), 
        .B2(n16278), .ZN(n16287) );
  NAND2_X1 U19423 ( .A1(n16279), .A2(n20199), .ZN(n16311) );
  INV_X1 U19424 ( .A(n16311), .ZN(n16284) );
  AOI21_X1 U19425 ( .B1(n20219), .B2(n16280), .A(n20218), .ZN(n20204) );
  OR2_X1 U19426 ( .A1(n20205), .A2(n16281), .ZN(n16282) );
  OAI211_X1 U19427 ( .C1(n16283), .C2(n20199), .A(n20204), .B(n16282), .ZN(
        n16307) );
  AOI21_X1 U19428 ( .B1(n20217), .B2(n16284), .A(n16307), .ZN(n16306) );
  OAI21_X1 U19429 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n20239), .A(
        n16306), .ZN(n16294) );
  AOI22_X1 U19430 ( .A1(n16285), .A2(n20243), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16294), .ZN(n16286) );
  OAI211_X1 U19431 ( .C1(n16290), .C2(n16288), .A(n16287), .B(n16286), .ZN(
        P1_U3023) );
  INV_X1 U19432 ( .A(n16289), .ZN(n16292) );
  OAI22_X1 U19433 ( .A1(n16292), .A2(n16291), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16290), .ZN(n16293) );
  AOI21_X1 U19434 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16294), .A(
        n16293), .ZN(n16296) );
  OAI211_X1 U19435 ( .C1(n20230), .C2(n20048), .A(n16296), .B(n16295), .ZN(
        P1_U3024) );
  INV_X1 U19436 ( .A(n13990), .ZN(n16299) );
  AOI21_X1 U19437 ( .B1(n16299), .B2(n16298), .A(n16297), .ZN(n16301) );
  OR2_X1 U19438 ( .A1(n16301), .A2(n16300), .ZN(n20060) );
  INV_X1 U19439 ( .A(n20060), .ZN(n20108) );
  AOI22_X1 U19440 ( .A1(n20236), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20238), 
        .B2(n20108), .ZN(n16305) );
  AOI22_X1 U19441 ( .A1(n16303), .A2(n20243), .B1(n16150), .B2(n16302), .ZN(
        n16304) );
  OAI211_X1 U19442 ( .C1(n16306), .C2(n16150), .A(n16305), .B(n16304), .ZN(
        P1_U3025) );
  AOI22_X1 U19443 ( .A1(n20236), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20238), 
        .B2(n20079), .ZN(n16310) );
  AOI22_X1 U19444 ( .A1(n16308), .A2(n20243), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16307), .ZN(n16309) );
  OAI211_X1 U19445 ( .C1(n20216), .C2(n16311), .A(n16310), .B(n16309), .ZN(
        P1_U3026) );
  OR4_X1 U19446 ( .A1(n20096), .A2(n16313), .A3(n16312), .A4(n13617), .ZN(
        n16314) );
  OAI21_X1 U19447 ( .B1(n16316), .B2(n16315), .A(n16314), .ZN(P1_U3468) );
  NAND4_X1 U19448 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20888), .A4(n20978), .ZN(n16317) );
  OAI21_X1 U19449 ( .B1(n16318), .B2(n20789), .A(n16317), .ZN(n20886) );
  OAI21_X1 U19450 ( .B1(n16325), .B2(n20885), .A(n20884), .ZN(n16319) );
  OAI211_X1 U19451 ( .C1(n16321), .C2(n20978), .A(n16320), .B(n16319), .ZN(
        n16322) );
  AOI221_X1 U19452 ( .B1(n16324), .B2(n16323), .C1(n20886), .C2(n16323), .A(
        n16322), .ZN(P1_U3162) );
  NOR2_X1 U19453 ( .A1(n16325), .A2(n20885), .ZN(n16327) );
  OAI22_X1 U19454 ( .A1(n20701), .A2(n16327), .B1(n16326), .B2(n20885), .ZN(
        P1_U3466) );
  INV_X1 U19455 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n16332) );
  INV_X1 U19456 ( .A(n16328), .ZN(n16331) );
  OAI222_X1 U19457 ( .A1(n19204), .A2(n16332), .B1(n19201), .B2(n16331), .C1(
        n16330), .C2(n16329), .ZN(n16333) );
  AOI21_X1 U19458 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19213), .A(
        n16333), .ZN(n16335) );
  AOI22_X1 U19459 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19167), .ZN(n16339) );
  AOI22_X1 U19460 ( .A1(n16337), .A2(n19185), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19207), .ZN(n16338) );
  OAI211_X1 U19461 ( .C1(n16340), .C2(n19203), .A(n16339), .B(n16338), .ZN(
        n16345) );
  AOI211_X1 U19462 ( .C1(n16343), .C2(n16342), .A(n16341), .B(n19216), .ZN(
        n16344) );
  NOR2_X1 U19463 ( .A1(n16345), .A2(n16344), .ZN(n16346) );
  OAI21_X1 U19464 ( .B1(n16347), .B2(n19209), .A(n16346), .ZN(P2_U2826) );
  AOI211_X1 U19465 ( .C1(n10206), .C2(n16349), .A(n16348), .B(n19216), .ZN(
        n16355) );
  INV_X1 U19466 ( .A(n16350), .ZN(n16353) );
  NAND2_X1 U19467 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19207), .ZN(n16352) );
  AOI22_X1 U19468 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19167), .ZN(n16351) );
  OAI211_X1 U19469 ( .C1(n16353), .C2(n19201), .A(n16352), .B(n16351), .ZN(
        n16354) );
  AOI211_X1 U19470 ( .C1(n19182), .C2(n16356), .A(n16355), .B(n16354), .ZN(
        n16357) );
  OAI21_X1 U19471 ( .B1(n16358), .B2(n19209), .A(n16357), .ZN(P2_U2827) );
  AOI211_X1 U19472 ( .C1(n16361), .C2(n16360), .A(n16359), .B(n19216), .ZN(
        n16363) );
  OAI22_X1 U19473 ( .A1(n10545), .A2(n19178), .B1(n19918), .B2(n19204), .ZN(
        n16362) );
  AOI211_X1 U19474 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n19207), .A(n16363), .B(
        n16362), .ZN(n16368) );
  OAI22_X1 U19475 ( .A1(n16365), .A2(n19201), .B1(n16364), .B2(n19203), .ZN(
        n16366) );
  INV_X1 U19476 ( .A(n16366), .ZN(n16367) );
  OAI211_X1 U19477 ( .C1(n16369), .C2(n19209), .A(n16368), .B(n16367), .ZN(
        P2_U2829) );
  AOI211_X1 U19478 ( .C1(n16372), .C2(n16371), .A(n16370), .B(n19216), .ZN(
        n16375) );
  OAI22_X1 U19479 ( .A1(n16373), .A2(n19178), .B1(n19916), .B2(n19204), .ZN(
        n16374) );
  AOI211_X1 U19480 ( .C1(P2_EBX_REG_25__SCAN_IN), .C2(n19207), .A(n16375), .B(
        n16374), .ZN(n16379) );
  AOI22_X1 U19481 ( .A1(n16377), .A2(n19185), .B1(n19182), .B2(n16376), .ZN(
        n16378) );
  OAI211_X1 U19482 ( .C1(n16380), .C2(n19209), .A(n16379), .B(n16378), .ZN(
        P2_U2830) );
  AOI211_X1 U19483 ( .C1(n16383), .C2(n16382), .A(n16381), .B(n19216), .ZN(
        n16385) );
  OAI22_X1 U19484 ( .A1(n19188), .A2(n15136), .B1(n15336), .B2(n19204), .ZN(
        n16384) );
  AOI211_X1 U19485 ( .C1(n19213), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16385), .B(n16384), .ZN(n16389) );
  AOI22_X1 U19486 ( .A1(n16387), .A2(n19185), .B1(n16386), .B2(n19182), .ZN(
        n16388) );
  OAI211_X1 U19487 ( .C1(n16390), .C2(n19209), .A(n16389), .B(n16388), .ZN(
        P2_U2831) );
  INV_X1 U19488 ( .A(n19362), .ZN(n16391) );
  AOI22_X1 U19489 ( .A1(n19221), .A2(n16391), .B1(n19239), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16396) );
  AOI22_X1 U19490 ( .A1(n19223), .A2(BUF1_REG_22__SCAN_IN), .B1(n19222), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16395) );
  AOI22_X1 U19491 ( .A1(n16393), .A2(n19225), .B1(n13389), .B2(n16392), .ZN(
        n16394) );
  NAND3_X1 U19492 ( .A1(n16396), .A2(n16395), .A3(n16394), .ZN(P2_U2897) );
  AOI22_X1 U19493 ( .A1(n19221), .A2(n16397), .B1(n19239), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16401) );
  AOI22_X1 U19494 ( .A1(n19223), .A2(BUF1_REG_20__SCAN_IN), .B1(n19222), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16400) );
  AOI22_X1 U19495 ( .A1(n16398), .A2(n19225), .B1(n13389), .B2(n19009), .ZN(
        n16399) );
  NAND3_X1 U19496 ( .A1(n16401), .A2(n16400), .A3(n16399), .ZN(P2_U2899) );
  AOI22_X1 U19497 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n11352), .ZN(n16405) );
  AOI222_X1 U19498 ( .A1(n16403), .A2(n19300), .B1(n19283), .B2(n16402), .C1(
        n19302), .C2(n19080), .ZN(n16404) );
  OAI211_X1 U19499 ( .C1(n19294), .C2(n19075), .A(n16405), .B(n16404), .ZN(
        P2_U3000) );
  AOI22_X1 U19500 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n11352), .ZN(n16414) );
  NAND2_X1 U19501 ( .A1(n16406), .A2(n16407), .ZN(n16410) );
  NAND2_X1 U19502 ( .A1(n16410), .A2(n16409), .ZN(n16408) );
  OAI21_X1 U19503 ( .B1(n16410), .B2(n16409), .A(n16408), .ZN(n16471) );
  AOI21_X1 U19504 ( .B1(n16472), .B2(n16412), .A(n16411), .ZN(n16469) );
  AOI222_X1 U19505 ( .A1(n16471), .A2(n19283), .B1(n19302), .B2(n16470), .C1(
        n19300), .C2(n16469), .ZN(n16413) );
  OAI211_X1 U19506 ( .C1(n19294), .C2(n19103), .A(n16414), .B(n16413), .ZN(
        P2_U3002) );
  AOI22_X1 U19507 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n11352), .B1(n16453), 
        .B2(n16415), .ZN(n16421) );
  OAI22_X1 U19508 ( .A1(n16417), .A2(n16456), .B1(n16416), .B2(n19305), .ZN(
        n16418) );
  AOI21_X1 U19509 ( .B1(n19302), .B2(n16419), .A(n16418), .ZN(n16420) );
  OAI211_X1 U19510 ( .C1(n16462), .C2(n16422), .A(n16421), .B(n16420), .ZN(
        P2_U3003) );
  AOI22_X1 U19511 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n11352), .ZN(n16429) );
  NOR3_X1 U19512 ( .A1(n16424), .A2(n16423), .A3(n16456), .ZN(n16427) );
  OAI22_X1 U19513 ( .A1(n16425), .A2(n19305), .B1(n19289), .B2(n19119), .ZN(
        n16426) );
  NOR2_X1 U19514 ( .A1(n16427), .A2(n16426), .ZN(n16428) );
  OAI211_X1 U19515 ( .C1(n19294), .C2(n19114), .A(n16429), .B(n16428), .ZN(
        P2_U3004) );
  AOI22_X1 U19516 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n11352), .ZN(n16445) );
  NAND2_X1 U19517 ( .A1(n16431), .A2(n16430), .ZN(n16436) );
  INV_X1 U19518 ( .A(n16432), .ZN(n16433) );
  AOI21_X1 U19519 ( .B1(n15468), .B2(n16434), .A(n16433), .ZN(n16435) );
  XOR2_X1 U19520 ( .A(n16436), .B(n16435), .Z(n16487) );
  INV_X1 U19521 ( .A(n19139), .ZN(n16485) );
  NAND2_X1 U19522 ( .A1(n15472), .A2(n16437), .ZN(n16442) );
  AND2_X1 U19523 ( .A1(n16439), .A2(n16438), .ZN(n16441) );
  NAND2_X1 U19524 ( .A1(n16442), .A2(n16441), .ZN(n16440) );
  OAI21_X1 U19525 ( .B1(n16442), .B2(n16441), .A(n16440), .ZN(n16443) );
  INV_X1 U19526 ( .A(n16443), .ZN(n16484) );
  AOI222_X1 U19527 ( .A1(n16487), .A2(n19283), .B1(n19302), .B2(n16485), .C1(
        n19300), .C2(n16484), .ZN(n16444) );
  OAI211_X1 U19528 ( .C1(n19294), .C2(n19134), .A(n16445), .B(n16444), .ZN(
        P2_U3006) );
  AOI22_X1 U19529 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n11352), .ZN(n16452) );
  OR2_X1 U19530 ( .A1(n16446), .A2(n16456), .ZN(n16448) );
  NAND2_X1 U19531 ( .A1(n19159), .A2(n19302), .ZN(n16447) );
  OAI211_X1 U19532 ( .C1(n16449), .C2(n19305), .A(n16448), .B(n16447), .ZN(
        n16450) );
  INV_X1 U19533 ( .A(n16450), .ZN(n16451) );
  OAI211_X1 U19534 ( .C1(n19294), .C2(n19157), .A(n16452), .B(n16451), .ZN(
        P2_U3008) );
  AOI22_X1 U19535 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n11352), .B1(n16453), 
        .B2(n19170), .ZN(n16460) );
  INV_X1 U19536 ( .A(n16454), .ZN(n19171) );
  OAI22_X1 U19537 ( .A1(n16457), .A2(n19305), .B1(n16456), .B2(n16455), .ZN(
        n16458) );
  AOI21_X1 U19538 ( .B1(n19302), .B2(n19171), .A(n16458), .ZN(n16459) );
  OAI211_X1 U19539 ( .C1(n16462), .C2(n16461), .A(n16460), .B(n16459), .ZN(
        P2_U3009) );
  NAND2_X1 U19540 ( .A1(n16463), .A2(n13445), .ZN(n16464) );
  AND2_X1 U19541 ( .A1(n16464), .A2(n9866), .ZN(n19234) );
  INV_X1 U19542 ( .A(n19234), .ZN(n16465) );
  OAI22_X1 U19543 ( .A1(n16467), .A2(n16472), .B1(n16466), .B2(n16465), .ZN(
        n16468) );
  INV_X1 U19544 ( .A(n16468), .ZN(n16477) );
  AOI222_X1 U19545 ( .A1(n16471), .A2(n19316), .B1(n16486), .B2(n16470), .C1(
        n19319), .C2(n16469), .ZN(n16476) );
  NAND2_X1 U19546 ( .A1(n16473), .A2(n16472), .ZN(n16475) );
  NAND2_X1 U19547 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n15730), .ZN(n16474) );
  NAND4_X1 U19548 ( .A1(n16477), .A2(n16476), .A3(n16475), .A4(n16474), .ZN(
        P2_U3034) );
  AOI21_X1 U19549 ( .B1(n16478), .B2(n13690), .A(n15705), .ZN(n19246) );
  AOI211_X1 U19550 ( .C1(n16481), .C2(n16491), .A(n16480), .B(n16479), .ZN(
        n16483) );
  NOR2_X1 U19551 ( .A1(n19151), .A2(n10481), .ZN(n16482) );
  AOI211_X1 U19552 ( .C1(n19326), .C2(n19246), .A(n16483), .B(n16482), .ZN(
        n16489) );
  AOI222_X1 U19553 ( .A1(n16487), .A2(n19316), .B1(n16486), .B2(n16485), .C1(
        n19319), .C2(n16484), .ZN(n16488) );
  OAI211_X1 U19554 ( .C1(n16491), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        P2_U3038) );
  INV_X1 U19555 ( .A(n16492), .ZN(n16502) );
  OAI21_X1 U19556 ( .B1(n19317), .B2(n13727), .A(n16493), .ZN(n16494) );
  AOI21_X1 U19557 ( .B1(n19948), .B2(n19326), .A(n16494), .ZN(n16495) );
  OAI21_X1 U19558 ( .B1(n16497), .B2(n16496), .A(n16495), .ZN(n16498) );
  AOI21_X1 U19559 ( .B1(n16499), .B2(n19316), .A(n16498), .ZN(n16500) );
  OAI221_X1 U19560 ( .B1(n16502), .B2(n10459), .C1(n16502), .C2(n16501), .A(
        n16500), .ZN(P2_U3043) );
  INV_X1 U19561 ( .A(n16503), .ZN(n18985) );
  INV_X1 U19562 ( .A(n19983), .ZN(n16506) );
  AOI211_X1 U19563 ( .C1(n16507), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        n16514) );
  MUX2_X1 U19564 ( .A(n16508), .B(n16510), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16512) );
  NAND3_X1 U19565 ( .A1(n16510), .A2(n19996), .A3(n16509), .ZN(n16511) );
  OAI21_X1 U19566 ( .B1(n16512), .B2(n19993), .A(n16511), .ZN(n16513) );
  OAI211_X1 U19567 ( .C1(n16515), .C2(n18985), .A(n16514), .B(n16513), .ZN(
        P2_U3176) );
  OAI21_X1 U19568 ( .B1(n18411), .B2(n16516), .A(n20999), .ZN(n16525) );
  INV_X1 U19569 ( .A(n17974), .ZN(n17596) );
  NAND2_X1 U19570 ( .A1(n17596), .A2(n16527), .ZN(n16543) );
  AOI211_X1 U19571 ( .C1(n16518), .C2(n16543), .A(n16517), .B(n17878), .ZN(
        n16524) );
  AOI21_X1 U19572 ( .B1(n20999), .B2(n16673), .A(n16519), .ZN(n16696) );
  OAI21_X1 U19573 ( .B1(n16520), .B2(n17812), .A(n16696), .ZN(n16522) );
  NAND2_X1 U19574 ( .A1(n16522), .A2(n16521), .ZN(n16523) );
  AOI211_X1 U19575 ( .C1(n16526), .C2(n16525), .A(n16524), .B(n16523), .ZN(
        n16530) );
  AND2_X1 U19576 ( .A1(n16527), .A2(n17976), .ZN(n16545) );
  OAI211_X1 U19577 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16545), .A(
        n17950), .B(n16528), .ZN(n16529) );
  OAI211_X1 U19578 ( .C1(n16531), .C2(n17853), .A(n16530), .B(n16529), .ZN(
        P3_U2801) );
  INV_X1 U19579 ( .A(n16532), .ZN(n16533) );
  AOI22_X1 U19580 ( .A1(n17873), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n16551), .B2(n17838), .ZN(n17608) );
  NOR2_X1 U19581 ( .A1(n18217), .A2(n16542), .ZN(n16540) );
  INV_X1 U19582 ( .A(n16535), .ZN(n18031) );
  INV_X1 U19583 ( .A(n18750), .ZN(n18028) );
  INV_X1 U19584 ( .A(n17827), .ZN(n18168) );
  AOI22_X1 U19585 ( .A1(n18028), .A2(n18168), .B1(n16536), .B2(n18204), .ZN(
        n18073) );
  OAI21_X1 U19586 ( .B1(n18073), .B2(n16538), .A(n16537), .ZN(n18017) );
  NAND2_X1 U19587 ( .A1(n18288), .A2(n18017), .ZN(n18042) );
  NOR2_X1 U19588 ( .A1(n18031), .A2(n18042), .ZN(n18034) );
  AOI22_X1 U19589 ( .A1(n16541), .A2(n16540), .B1(n16539), .B2(n18034), .ZN(
        n16556) );
  INV_X1 U19590 ( .A(n16542), .ZN(n16548) );
  INV_X1 U19591 ( .A(n15924), .ZN(n16547) );
  NAND2_X1 U19592 ( .A1(n16543), .A2(n18204), .ZN(n16544) );
  OAI21_X1 U19593 ( .B1(n16545), .B2(n18750), .A(n16544), .ZN(n16546) );
  NOR2_X1 U19594 ( .A1(n9768), .A2(n16551), .ZN(n16553) );
  NAND2_X1 U19595 ( .A1(n9768), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17601) );
  OAI21_X1 U19596 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n16556), .A(
        n16555), .ZN(P3_U2834) );
  NOR3_X1 U19597 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16558) );
  NOR4_X1 U19598 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16557) );
  NAND4_X1 U19599 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16558), .A3(n16557), .A4(
        U215), .ZN(U213) );
  INV_X1 U19600 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16642) );
  NOR2_X1 U19601 ( .A1(n16606), .A2(n16559), .ZN(n16604) );
  INV_X1 U19602 ( .A(n16604), .ZN(n16608) );
  INV_X1 U19603 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16641) );
  OAI222_X1 U19604 ( .A1(U212), .A2(n16642), .B1(n16608), .B2(n16560), .C1(
        U214), .C2(n16641), .ZN(U216) );
  INV_X1 U19605 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16562) );
  AOI22_X1 U19606 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16606), .ZN(n16561) );
  OAI21_X1 U19607 ( .B1(n16562), .B2(n16608), .A(n16561), .ZN(U217) );
  AOI22_X1 U19608 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16606), .ZN(n16563) );
  OAI21_X1 U19609 ( .B1(n16564), .B2(n16608), .A(n16563), .ZN(U218) );
  INV_X1 U19610 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20290) );
  AOI22_X1 U19611 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16606), .ZN(n16565) );
  OAI21_X1 U19612 ( .B1(n20290), .B2(n16608), .A(n16565), .ZN(U219) );
  INV_X1 U19613 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16567) );
  AOI22_X1 U19614 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16606), .ZN(n16566) );
  OAI21_X1 U19615 ( .B1(n16567), .B2(n16608), .A(n16566), .ZN(U220) );
  INV_X1 U19616 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U19617 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16606), .ZN(n16568) );
  OAI21_X1 U19618 ( .B1(n16569), .B2(n16608), .A(n16568), .ZN(U221) );
  INV_X1 U19619 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16571) );
  AOI22_X1 U19620 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16606), .ZN(n16570) );
  OAI21_X1 U19621 ( .B1(n16571), .B2(n16608), .A(n16570), .ZN(U222) );
  AOI222_X1 U19622 ( .A1(n16606), .A2(P1_DATAO_REG_24__SCAN_IN), .B1(n16604), 
        .B2(BUF1_REG_24__SCAN_IN), .C1(n16602), .C2(P2_DATAO_REG_24__SCAN_IN), 
        .ZN(n16572) );
  INV_X1 U19623 ( .A(n16572), .ZN(U223) );
  AOI222_X1 U19624 ( .A1(n16606), .A2(P1_DATAO_REG_23__SCAN_IN), .B1(n16604), 
        .B2(BUF1_REG_23__SCAN_IN), .C1(n16602), .C2(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n16573) );
  INV_X1 U19625 ( .A(n16573), .ZN(U224) );
  INV_X1 U19626 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16575) );
  AOI22_X1 U19627 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16606), .ZN(n16574) );
  OAI21_X1 U19628 ( .B1(n16575), .B2(n16608), .A(n16574), .ZN(U225) );
  INV_X1 U19629 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20301) );
  AOI22_X1 U19630 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16606), .ZN(n16576) );
  OAI21_X1 U19631 ( .B1(n20301), .B2(n16608), .A(n16576), .ZN(U226) );
  INV_X1 U19632 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16578) );
  AOI22_X1 U19633 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16606), .ZN(n16577) );
  OAI21_X1 U19634 ( .B1(n16578), .B2(n16608), .A(n16577), .ZN(U227) );
  AOI222_X1 U19635 ( .A1(n16606), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n16604), 
        .B2(BUF1_REG_19__SCAN_IN), .C1(n16602), .C2(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n16579) );
  INV_X1 U19636 ( .A(n16579), .ZN(U228) );
  INV_X1 U19637 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U19638 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16606), .ZN(n16580) );
  OAI21_X1 U19639 ( .B1(n16581), .B2(n16608), .A(n16580), .ZN(U229) );
  INV_X1 U19640 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20275) );
  AOI22_X1 U19641 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16606), .ZN(n16582) );
  OAI21_X1 U19642 ( .B1(n20275), .B2(n16608), .A(n16582), .ZN(U230) );
  INV_X1 U19643 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16584) );
  AOI22_X1 U19644 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16606), .ZN(n16583) );
  OAI21_X1 U19645 ( .B1(n16584), .B2(n16608), .A(n16583), .ZN(U231) );
  AOI22_X1 U19646 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16606), .ZN(n16585) );
  OAI21_X1 U19647 ( .B1(n13697), .B2(n16608), .A(n16585), .ZN(U232) );
  AOI22_X1 U19648 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16606), .ZN(n16586) );
  OAI21_X1 U19649 ( .B1(n14771), .B2(n16608), .A(n16586), .ZN(U233) );
  INV_X1 U19650 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n21125) );
  AOI22_X1 U19651 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16604), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16606), .ZN(n16587) );
  OAI21_X1 U19652 ( .B1(n21125), .B2(U212), .A(n16587), .ZN(U234) );
  AOI22_X1 U19653 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16606), .ZN(n16588) );
  OAI21_X1 U19654 ( .B1(n16589), .B2(n16608), .A(n16588), .ZN(U235) );
  INV_X1 U19655 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16619) );
  AOI22_X1 U19656 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16604), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16606), .ZN(n16590) );
  OAI21_X1 U19657 ( .B1(n16619), .B2(U212), .A(n16590), .ZN(U236) );
  AOI22_X1 U19658 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16606), .ZN(n16591) );
  OAI21_X1 U19659 ( .B1(n13693), .B2(n16608), .A(n16591), .ZN(U237) );
  INV_X1 U19660 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n21161) );
  INV_X1 U19661 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16617) );
  OAI222_X1 U19662 ( .A1(U214), .A2(n21161), .B1(n16608), .B2(n16592), .C1(
        U212), .C2(n16617), .ZN(U238) );
  AOI22_X1 U19663 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16606), .ZN(n16593) );
  OAI21_X1 U19664 ( .B1(n14230), .B2(n16608), .A(n16593), .ZN(U239) );
  AOI22_X1 U19665 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16606), .ZN(n16594) );
  OAI21_X1 U19666 ( .B1(n16595), .B2(n16608), .A(n16594), .ZN(U240) );
  INV_X1 U19667 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16597) );
  AOI22_X1 U19668 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16606), .ZN(n16596) );
  OAI21_X1 U19669 ( .B1(n16597), .B2(n16608), .A(n16596), .ZN(U241) );
  INV_X1 U19670 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16613) );
  AOI22_X1 U19671 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16604), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16606), .ZN(n16598) );
  OAI21_X1 U19672 ( .B1(n16613), .B2(U212), .A(n16598), .ZN(U242) );
  INV_X1 U19673 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16600) );
  AOI22_X1 U19674 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16606), .ZN(n16599) );
  OAI21_X1 U19675 ( .B1(n16600), .B2(n16608), .A(n16599), .ZN(U243) );
  INV_X1 U19676 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n21238) );
  AOI22_X1 U19677 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16604), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16606), .ZN(n16601) );
  OAI21_X1 U19678 ( .B1(n21238), .B2(U212), .A(n16601), .ZN(U244) );
  INV_X1 U19679 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n21195) );
  AOI22_X1 U19680 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16606), .ZN(n16603) );
  OAI21_X1 U19681 ( .B1(n21195), .B2(n16608), .A(n16603), .ZN(U245) );
  INV_X1 U19682 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n21062) );
  AOI22_X1 U19683 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16604), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16606), .ZN(n16605) );
  OAI21_X1 U19684 ( .B1(n21062), .B2(U212), .A(n16605), .ZN(U246) );
  AOI22_X1 U19685 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16602), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16606), .ZN(n16607) );
  OAI21_X1 U19686 ( .B1(n16609), .B2(n16608), .A(n16607), .ZN(U247) );
  INV_X1 U19687 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16610) );
  AOI22_X1 U19688 ( .A1(n16634), .A2(n16610), .B1(n18304), .B2(U215), .ZN(U251) );
  INV_X1 U19689 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n21207) );
  AOI22_X1 U19690 ( .A1(n16634), .A2(n21062), .B1(n21207), .B2(U215), .ZN(U252) );
  INV_X1 U19691 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16611) );
  INV_X1 U19692 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18314) );
  AOI22_X1 U19693 ( .A1(n16634), .A2(n16611), .B1(n18314), .B2(U215), .ZN(U253) );
  INV_X1 U19694 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18320) );
  AOI22_X1 U19695 ( .A1(n16634), .A2(n21238), .B1(n18320), .B2(U215), .ZN(U254) );
  INV_X1 U19696 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16612) );
  INV_X1 U19697 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18325) );
  AOI22_X1 U19698 ( .A1(n16634), .A2(n16612), .B1(n18325), .B2(U215), .ZN(U255) );
  INV_X1 U19699 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U19700 ( .A1(n16634), .A2(n16613), .B1(n18330), .B2(U215), .ZN(U256) );
  INV_X1 U19701 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16614) );
  INV_X1 U19702 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18335) );
  AOI22_X1 U19703 ( .A1(n16638), .A2(n16614), .B1(n18335), .B2(U215), .ZN(U257) );
  INV_X1 U19704 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16615) );
  INV_X1 U19705 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18340) );
  AOI22_X1 U19706 ( .A1(n16638), .A2(n16615), .B1(n18340), .B2(U215), .ZN(U258) );
  OAI22_X1 U19707 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16634), .ZN(n16616) );
  INV_X1 U19708 ( .A(n16616), .ZN(U259) );
  INV_X1 U19709 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U19710 ( .A1(n16638), .A2(n16617), .B1(n17453), .B2(U215), .ZN(U260) );
  OAI22_X1 U19711 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16634), .ZN(n16618) );
  INV_X1 U19712 ( .A(n16618), .ZN(U261) );
  INV_X1 U19713 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21224) );
  AOI22_X1 U19714 ( .A1(n16634), .A2(n16619), .B1(n21224), .B2(U215), .ZN(U262) );
  INV_X1 U19715 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16620) );
  INV_X1 U19716 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U19717 ( .A1(n16634), .A2(n16620), .B1(n17441), .B2(U215), .ZN(U263) );
  INV_X1 U19718 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n16621) );
  AOI22_X1 U19719 ( .A1(n16638), .A2(n21125), .B1(n16621), .B2(U215), .ZN(U264) );
  INV_X1 U19720 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16622) );
  INV_X1 U19721 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U19722 ( .A1(n16634), .A2(n16622), .B1(n17430), .B2(U215), .ZN(U265) );
  OAI22_X1 U19723 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16634), .ZN(n16623) );
  INV_X1 U19724 ( .A(n16623), .ZN(U266) );
  OAI22_X1 U19725 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16634), .ZN(n16624) );
  INV_X1 U19726 ( .A(n16624), .ZN(U267) );
  OAI22_X1 U19727 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16634), .ZN(n16625) );
  INV_X1 U19728 ( .A(n16625), .ZN(U268) );
  OAI22_X1 U19729 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16634), .ZN(n16626) );
  INV_X1 U19730 ( .A(n16626), .ZN(U269) );
  INV_X1 U19731 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n21148) );
  INV_X1 U19732 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18319) );
  AOI22_X1 U19733 ( .A1(n16634), .A2(n21148), .B1(n18319), .B2(U215), .ZN(U270) );
  OAI22_X1 U19734 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16634), .ZN(n16627) );
  INV_X1 U19735 ( .A(n16627), .ZN(U271) );
  OAI22_X1 U19736 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16634), .ZN(n16628) );
  INV_X1 U19737 ( .A(n16628), .ZN(U272) );
  OAI22_X1 U19738 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16634), .ZN(n16629) );
  INV_X1 U19739 ( .A(n16629), .ZN(U273) );
  INV_X1 U19740 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n21049) );
  INV_X1 U19741 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U19742 ( .A1(n16634), .A2(n21049), .B1(n18339), .B2(U215), .ZN(U274) );
  OAI22_X1 U19743 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16634), .ZN(n16630) );
  INV_X1 U19744 ( .A(n16630), .ZN(U275) );
  OAI22_X1 U19745 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16638), .ZN(n16631) );
  INV_X1 U19746 ( .A(n16631), .ZN(U276) );
  OAI22_X1 U19747 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16638), .ZN(n16632) );
  INV_X1 U19748 ( .A(n16632), .ZN(U277) );
  INV_X1 U19749 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16633) );
  AOI22_X1 U19750 ( .A1(n16634), .A2(n16633), .B1(n15226), .B2(U215), .ZN(U278) );
  OAI22_X1 U19751 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16638), .ZN(n16635) );
  INV_X1 U19752 ( .A(n16635), .ZN(U279) );
  OAI22_X1 U19753 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16638), .ZN(n16636) );
  INV_X1 U19754 ( .A(n16636), .ZN(U280) );
  OAI22_X1 U19755 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16638), .ZN(n16637) );
  INV_X1 U19756 ( .A(n16637), .ZN(U281) );
  OAI22_X1 U19757 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16638), .ZN(n16639) );
  INV_X1 U19758 ( .A(n16639), .ZN(U282) );
  INV_X1 U19759 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16640) );
  AOI222_X1 U19760 ( .A1(n16642), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16641), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16640), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16643) );
  INV_X1 U19761 ( .A(n16645), .ZN(n16644) );
  INV_X1 U19762 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18852) );
  INV_X1 U19763 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U19764 ( .A1(n16644), .A2(n18852), .B1(n19894), .B2(n16645), .ZN(
        U347) );
  INV_X1 U19765 ( .A(n16645), .ZN(n16646) );
  INV_X1 U19766 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18850) );
  INV_X1 U19767 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U19768 ( .A1(n16646), .A2(n18850), .B1(n19893), .B2(n16645), .ZN(
        U348) );
  INV_X1 U19769 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18847) );
  INV_X1 U19770 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U19771 ( .A1(n16644), .A2(n18847), .B1(n19892), .B2(n16645), .ZN(
        U349) );
  INV_X1 U19772 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18846) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19774 ( .A1(n16644), .A2(n18846), .B1(n19891), .B2(n16645), .ZN(
        U350) );
  INV_X1 U19775 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18844) );
  INV_X1 U19776 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U19777 ( .A1(n16644), .A2(n18844), .B1(n19890), .B2(n16645), .ZN(
        U351) );
  INV_X1 U19778 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18842) );
  INV_X1 U19779 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U19780 ( .A1(n16644), .A2(n18842), .B1(n19889), .B2(n16645), .ZN(
        U352) );
  INV_X1 U19781 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18840) );
  AOI22_X1 U19782 ( .A1(n16646), .A2(n18840), .B1(n19888), .B2(n16645), .ZN(
        U353) );
  INV_X1 U19783 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18838) );
  INV_X1 U19784 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U19785 ( .A1(n16644), .A2(n18838), .B1(n19887), .B2(n16645), .ZN(
        U354) );
  INV_X1 U19786 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18893) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19925) );
  AOI22_X1 U19788 ( .A1(n16644), .A2(n18893), .B1(n19925), .B2(n16645), .ZN(
        U355) );
  INV_X1 U19789 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18890) );
  INV_X1 U19790 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19922) );
  AOI22_X1 U19791 ( .A1(n16644), .A2(n18890), .B1(n19922), .B2(n16645), .ZN(
        U356) );
  INV_X1 U19792 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18887) );
  INV_X1 U19793 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19920) );
  AOI22_X1 U19794 ( .A1(n16644), .A2(n18887), .B1(n19920), .B2(n16645), .ZN(
        U357) );
  INV_X1 U19795 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18885) );
  INV_X1 U19796 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21236) );
  AOI22_X1 U19797 ( .A1(n16644), .A2(n18885), .B1(n21236), .B2(n16645), .ZN(
        U358) );
  INV_X1 U19798 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18883) );
  INV_X1 U19799 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n21027) );
  AOI22_X1 U19800 ( .A1(n16644), .A2(n18883), .B1(n21027), .B2(n16645), .ZN(
        U359) );
  INV_X1 U19801 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18881) );
  INV_X1 U19802 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19917) );
  AOI22_X1 U19803 ( .A1(n16644), .A2(n18881), .B1(n19917), .B2(n16645), .ZN(
        U360) );
  INV_X1 U19804 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18879) );
  INV_X1 U19805 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U19806 ( .A1(n16644), .A2(n18879), .B1(n19915), .B2(n16645), .ZN(
        U361) );
  INV_X1 U19807 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18877) );
  INV_X1 U19808 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U19809 ( .A1(n16644), .A2(n18877), .B1(n19914), .B2(n16645), .ZN(
        U362) );
  INV_X1 U19810 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18875) );
  INV_X1 U19811 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19912) );
  AOI22_X1 U19812 ( .A1(n16644), .A2(n18875), .B1(n19912), .B2(n16645), .ZN(
        U363) );
  INV_X1 U19813 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18873) );
  INV_X1 U19814 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19911) );
  AOI22_X1 U19815 ( .A1(n16644), .A2(n18873), .B1(n19911), .B2(n16645), .ZN(
        U364) );
  INV_X1 U19816 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18836) );
  INV_X1 U19817 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19886) );
  AOI22_X1 U19818 ( .A1(n16644), .A2(n18836), .B1(n19886), .B2(n16645), .ZN(
        U365) );
  INV_X1 U19819 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18870) );
  INV_X1 U19820 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U19821 ( .A1(n16644), .A2(n18870), .B1(n19909), .B2(n16645), .ZN(
        U366) );
  INV_X1 U19822 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18869) );
  INV_X1 U19823 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U19824 ( .A1(n16644), .A2(n18869), .B1(n19907), .B2(n16645), .ZN(
        U367) );
  INV_X1 U19825 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18867) );
  INV_X1 U19826 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19827 ( .A1(n16644), .A2(n18867), .B1(n19905), .B2(n16645), .ZN(
        U368) );
  INV_X1 U19828 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18864) );
  INV_X1 U19829 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U19830 ( .A1(n16644), .A2(n18864), .B1(n19903), .B2(n16645), .ZN(
        U369) );
  INV_X1 U19831 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18863) );
  INV_X1 U19832 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U19833 ( .A1(n16644), .A2(n18863), .B1(n19901), .B2(n16645), .ZN(
        U370) );
  INV_X1 U19834 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18861) );
  INV_X1 U19835 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19900) );
  AOI22_X1 U19836 ( .A1(n16646), .A2(n18861), .B1(n19900), .B2(n16645), .ZN(
        U371) );
  INV_X1 U19837 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18858) );
  INV_X1 U19838 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19898) );
  AOI22_X1 U19839 ( .A1(n16646), .A2(n18858), .B1(n19898), .B2(n16645), .ZN(
        U372) );
  INV_X1 U19840 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18857) );
  INV_X1 U19841 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19842 ( .A1(n16646), .A2(n18857), .B1(n19897), .B2(n16645), .ZN(
        U373) );
  INV_X1 U19843 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18856) );
  INV_X1 U19844 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U19845 ( .A1(n16646), .A2(n18856), .B1(n19896), .B2(n16645), .ZN(
        U374) );
  INV_X1 U19846 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18854) );
  INV_X1 U19847 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19895) );
  AOI22_X1 U19848 ( .A1(n16646), .A2(n18854), .B1(n19895), .B2(n16645), .ZN(
        U375) );
  INV_X1 U19849 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18834) );
  INV_X1 U19850 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n21094) );
  AOI22_X1 U19851 ( .A1(n16646), .A2(n18834), .B1(n21094), .B2(n16645), .ZN(
        U376) );
  INV_X1 U19852 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16647) );
  INV_X1 U19853 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18818) );
  NOR2_X1 U19854 ( .A1(n18818), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18820) );
  OAI22_X1 U19855 ( .A1(n18830), .A2(n18820), .B1(n18818), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18904) );
  OAI21_X1 U19856 ( .B1(n18830), .B2(n16647), .A(n18904), .ZN(P3_U2633) );
  NOR2_X1 U19857 ( .A1(n9764), .A2(n16653), .ZN(n16648) );
  OAI21_X1 U19858 ( .B1(n16648), .B2(n17530), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16649) );
  OAI21_X1 U19859 ( .B1(n16650), .B2(n18805), .A(n16649), .ZN(P3_U2634) );
  AOI21_X1 U19860 ( .B1(n18830), .B2(n18833), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16651) );
  AOI22_X1 U19861 ( .A1(n18972), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16651), 
        .B2(n18970), .ZN(P3_U2635) );
  INV_X1 U19862 ( .A(n18904), .ZN(n18907) );
  OAI21_X1 U19863 ( .B1(n18816), .B2(BS16), .A(n18907), .ZN(n18905) );
  OAI21_X1 U19864 ( .B1(n18907), .B2(n18960), .A(n18905), .ZN(P3_U2636) );
  OAI211_X1 U19865 ( .C1(n9764), .C2(n16653), .A(n18746), .B(n16652), .ZN(
        n18791) );
  NAND2_X1 U19866 ( .A1(n18791), .A2(n18955), .ZN(n18954) );
  INV_X1 U19867 ( .A(n18954), .ZN(n16656) );
  OAI21_X1 U19868 ( .B1(n16656), .B2(n16655), .A(n16654), .ZN(P3_U2637) );
  NOR4_X1 U19869 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16660) );
  NOR4_X1 U19870 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16659) );
  NOR4_X1 U19871 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16658) );
  NOR4_X1 U19872 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16657) );
  NAND4_X1 U19873 ( .A1(n16660), .A2(n16659), .A3(n16658), .A4(n16657), .ZN(
        n16666) );
  NOR4_X1 U19874 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16664) );
  AOI211_X1 U19875 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_13__SCAN_IN), .B(
        P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(n16663) );
  NOR4_X1 U19876 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n16662) );
  NOR4_X1 U19877 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16661) );
  NAND4_X1 U19878 ( .A1(n16664), .A2(n16663), .A3(n16662), .A4(n16661), .ZN(
        n16665) );
  NOR2_X1 U19879 ( .A1(n16666), .A2(n16665), .ZN(n18946) );
  INV_X1 U19880 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18900) );
  NOR3_X1 U19881 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16668) );
  OAI21_X1 U19882 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16668), .A(n18946), .ZN(
        n16667) );
  OAI21_X1 U19883 ( .B1(n18946), .B2(n18900), .A(n16667), .ZN(P3_U2638) );
  INV_X1 U19884 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18942) );
  INV_X1 U19885 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18906) );
  AOI21_X1 U19886 ( .B1(n18942), .B2(n18906), .A(n16668), .ZN(n16669) );
  INV_X1 U19887 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18897) );
  INV_X1 U19888 ( .A(n18946), .ZN(n18949) );
  AOI22_X1 U19889 ( .A1(n18946), .A2(n16669), .B1(n18897), .B2(n18949), .ZN(
        P3_U2639) );
  INV_X1 U19890 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17618) );
  INV_X1 U19891 ( .A(n16670), .ZN(n16671) );
  NOR2_X1 U19892 ( .A1(n17618), .A2(n16671), .ZN(n16674) );
  AOI21_X1 U19893 ( .B1(n17618), .B2(n16671), .A(n16674), .ZN(n17614) );
  NOR2_X1 U19894 ( .A1(n16672), .A2(n9920), .ZN(n16714) );
  OAI21_X1 U19896 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16674), .A(
        n16673), .ZN(n17603) );
  INV_X1 U19897 ( .A(n17603), .ZN(n16706) );
  NOR2_X1 U19898 ( .A1(n16704), .A2(n9920), .ZN(n16695) );
  NAND2_X1 U19900 ( .A1(n9921), .A2(n16987), .ZN(n17014) );
  NOR3_X1 U19901 ( .A1(n16684), .A2(n16683), .A3(n17014), .ZN(n16678) );
  NOR2_X1 U19902 ( .A1(n17015), .A2(n16675), .ZN(n16702) );
  NAND4_X1 U19903 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16702), .ZN(n16685) );
  INV_X1 U19904 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18894) );
  AOI22_X1 U19905 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18894), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n18892), .ZN(n16676) );
  OAI22_X1 U19906 ( .A1(n9910), .A2(n17013), .B1(n16685), .B2(n16676), .ZN(
        n16677) );
  AOI211_X1 U19907 ( .C1(n17006), .C2(P3_EBX_REG_31__SCAN_IN), .A(n16678), .B(
        n16677), .ZN(n16681) );
  INV_X1 U19908 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18889) );
  NAND2_X1 U19909 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16690) );
  NOR2_X1 U19910 ( .A1(n18889), .A2(n16690), .ZN(n16679) );
  OAI21_X1 U19911 ( .B1(n16679), .B2(n17015), .A(n16722), .ZN(n16699) );
  NAND2_X1 U19912 ( .A1(n16719), .A2(n17074), .ZN(n16718) );
  NOR2_X1 U19913 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16718), .ZN(n16703) );
  INV_X1 U19914 ( .A(n16703), .ZN(n16693) );
  OR2_X1 U19915 ( .A1(n16693), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n16682) );
  NOR2_X1 U19916 ( .A1(n17022), .A2(n16682), .ZN(n16687) );
  INV_X1 U19917 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U19918 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n16699), .B1(n16687), 
        .B2(n17037), .ZN(n16680) );
  NAND2_X1 U19919 ( .A1(n16681), .A2(n16680), .ZN(P3_U2640) );
  NAND2_X1 U19920 ( .A1(n16977), .A2(n16682), .ZN(n16692) );
  OAI22_X1 U19921 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16685), .B1(n9912), 
        .B2(n17013), .ZN(n16686) );
  OAI21_X1 U19922 ( .B1(n17006), .B2(n16687), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16688) );
  OAI211_X1 U19923 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16692), .A(n16689), .B(
        n16688), .ZN(P3_U2641) );
  NOR2_X1 U19924 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16690), .ZN(n16691) );
  AOI22_X1 U19925 ( .A1(n17006), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16702), 
        .B2(n16691), .ZN(n16701) );
  AOI21_X1 U19926 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16693), .A(n16692), .ZN(
        n16698) );
  AOI211_X1 U19927 ( .C1(n16696), .C2(n16695), .A(n16694), .B(n18811), .ZN(
        n16697) );
  AOI211_X1 U19928 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16699), .A(n16698), 
        .B(n16697), .ZN(n16700) );
  OAI211_X1 U19929 ( .C1(n20999), .C2(n17013), .A(n16701), .B(n16700), .ZN(
        P3_U2642) );
  NAND2_X1 U19930 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16702), .ZN(n16712) );
  AOI22_X1 U19931 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16903), .B1(
        n17006), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16711) );
  INV_X1 U19932 ( .A(n16702), .ZN(n16715) );
  OAI21_X1 U19933 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16715), .A(n16722), 
        .ZN(n16709) );
  AOI211_X1 U19934 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16718), .A(n16703), .B(
        n17022), .ZN(n16708) );
  AOI211_X1 U19935 ( .C1(n16706), .C2(n16705), .A(n16704), .B(n18811), .ZN(
        n16707) );
  AOI211_X1 U19936 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16709), .A(n16708), 
        .B(n16707), .ZN(n16710) );
  OAI211_X1 U19937 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16712), .A(n16711), 
        .B(n16710), .ZN(P3_U2643) );
  INV_X1 U19938 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18884) );
  AOI211_X1 U19939 ( .C1(n17614), .C2(n16714), .A(n16713), .B(n18811), .ZN(
        n16717) );
  OAI22_X1 U19940 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16715), .B1(n17618), 
        .B2(n17013), .ZN(n16716) );
  AOI211_X1 U19941 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17006), .A(n16717), .B(
        n16716), .ZN(n16721) );
  OAI211_X1 U19942 ( .C1(n16719), .C2(n17074), .A(n16977), .B(n16718), .ZN(
        n16720) );
  OAI211_X1 U19943 ( .C1(n16722), .C2(n18884), .A(n16721), .B(n16720), .ZN(
        P3_U2644) );
  OR2_X1 U19944 ( .A1(n17022), .A2(n16723), .ZN(n16732) );
  AOI21_X1 U19945 ( .B1(n16977), .B2(n16723), .A(n17006), .ZN(n16731) );
  AOI21_X1 U19946 ( .B1(n17001), .B2(n16741), .A(n17012), .ZN(n16744) );
  OAI21_X1 U19947 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17015), .A(n16744), 
        .ZN(n16729) );
  AOI211_X1 U19948 ( .C1(n16725), .C2(n16724), .A(n9826), .B(n18811), .ZN(
        n16728) );
  INV_X1 U19949 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17641) );
  OAI22_X1 U19950 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16726), .B1(n17641), 
        .B2(n17013), .ZN(n16727) );
  AOI211_X1 U19951 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16729), .A(n16728), 
        .B(n16727), .ZN(n16730) );
  OAI221_X1 U19952 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16732), .C1(n17031), 
        .C2(n16731), .A(n16730), .ZN(P3_U2646) );
  NAND2_X1 U19953 ( .A1(n17001), .A2(n18878), .ZN(n16740) );
  AOI22_X1 U19954 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16903), .B1(
        n17006), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16739) );
  INV_X1 U19955 ( .A(n16744), .ZN(n16737) );
  AOI21_X1 U19956 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16747), .A(n16732), .ZN(
        n16736) );
  AOI211_X1 U19957 ( .C1(n17660), .C2(n16734), .A(n16733), .B(n18811), .ZN(
        n16735) );
  AOI211_X1 U19958 ( .C1(n16737), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16736), 
        .B(n16735), .ZN(n16738) );
  OAI211_X1 U19959 ( .C1(n16741), .C2(n16740), .A(n16739), .B(n16738), .ZN(
        P3_U2647) );
  INV_X1 U19960 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18876) );
  NAND2_X1 U19961 ( .A1(n16752), .A2(n18876), .ZN(n16751) );
  NAND2_X1 U19962 ( .A1(n17001), .A2(n16823), .ZN(n16824) );
  INV_X1 U19963 ( .A(n16824), .ZN(n16808) );
  NAND2_X1 U19964 ( .A1(n16754), .A2(n16808), .ZN(n16761) );
  AOI211_X1 U19965 ( .C1(n17669), .C2(n16743), .A(n16742), .B(n18811), .ZN(
        n16746) );
  OAI22_X1 U19966 ( .A1(n17023), .A2(n16748), .B1(n18876), .B2(n16744), .ZN(
        n16745) );
  AOI211_X1 U19967 ( .C1(n16903), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16746), .B(n16745), .ZN(n16750) );
  OAI211_X1 U19968 ( .C1(n16755), .C2(n16748), .A(n16977), .B(n16747), .ZN(
        n16749) );
  OAI211_X1 U19969 ( .C1(n16751), .C2(n16761), .A(n16750), .B(n16749), .ZN(
        P3_U2648) );
  AOI211_X1 U19970 ( .C1(n18874), .C2(n18872), .A(n16752), .B(n16761), .ZN(
        n16753) );
  AOI21_X1 U19971 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17006), .A(n16753), .ZN(
        n16760) );
  AND2_X1 U19972 ( .A1(n17025), .A2(n16823), .ZN(n16839) );
  NOR2_X1 U19973 ( .A1(n17012), .A2(n17001), .ZN(n17028) );
  AOI21_X1 U19974 ( .B1(n16754), .B2(n16839), .A(n17028), .ZN(n16771) );
  AOI211_X1 U19975 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16766), .A(n16755), .B(
        n17022), .ZN(n16758) );
  AOI211_X1 U19976 ( .C1(n17685), .C2(n16756), .A(n9872), .B(n18811), .ZN(
        n16757) );
  AOI211_X1 U19977 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16771), .A(n16758), 
        .B(n16757), .ZN(n16759) );
  OAI211_X1 U19978 ( .C1(n17694), .C2(n17013), .A(n16760), .B(n16759), .ZN(
        P3_U2649) );
  AOI22_X1 U19979 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16903), .B1(
        n17006), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16770) );
  INV_X1 U19980 ( .A(n16761), .ZN(n16765) );
  AOI211_X1 U19981 ( .C1(n17699), .C2(n16763), .A(n16762), .B(n18811), .ZN(
        n16764) );
  AOI221_X1 U19982 ( .B1(n16765), .B2(n18872), .C1(n16771), .C2(
        P3_REIP_REG_21__SCAN_IN), .A(n16764), .ZN(n16769) );
  OAI211_X1 U19983 ( .C1(n16775), .C2(n16767), .A(n16977), .B(n16766), .ZN(
        n16768) );
  NAND3_X1 U19984 ( .A1(n16770), .A2(n16769), .A3(n16768), .ZN(P3_U2650) );
  INV_X1 U19985 ( .A(n16771), .ZN(n16780) );
  NOR2_X1 U19986 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16772), .ZN(n16773) );
  AOI22_X1 U19987 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16903), .B1(
        n16808), .B2(n16773), .ZN(n16779) );
  AOI211_X1 U19988 ( .C1(n17713), .C2(n16781), .A(n16774), .B(n18811), .ZN(
        n16777) );
  AOI211_X1 U19989 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16786), .A(n16775), .B(
        n17022), .ZN(n16776) );
  AOI211_X1 U19990 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17006), .A(n16777), .B(
        n16776), .ZN(n16778) );
  OAI211_X1 U19991 ( .C1(n16780), .C2(n18871), .A(n16779), .B(n16778), .ZN(
        P3_U2651) );
  AOI21_X1 U19992 ( .B1(n16791), .B2(n16839), .A(n17028), .ZN(n16815) );
  INV_X1 U19993 ( .A(n16815), .ZN(n16794) );
  INV_X1 U19994 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18868) );
  INV_X1 U19995 ( .A(n16781), .ZN(n16785) );
  INV_X1 U19996 ( .A(n17723), .ZN(n16797) );
  NOR2_X1 U19997 ( .A1(n17726), .A2(n16797), .ZN(n16782) );
  OAI21_X1 U19998 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16782), .A(
        n17679), .ZN(n17727) );
  NAND2_X1 U19999 ( .A1(n16987), .A2(n9920), .ZN(n17009) );
  OAI21_X1 U20000 ( .B1(n16783), .B2(n17727), .A(n16987), .ZN(n16784) );
  AOI22_X1 U20001 ( .A1(n16785), .A2(n17727), .B1(n17009), .B2(n16784), .ZN(
        n16790) );
  OAI211_X1 U20002 ( .C1(n16795), .C2(n16788), .A(n16977), .B(n16786), .ZN(
        n16787) );
  OAI211_X1 U20003 ( .C1(n17023), .C2(n16788), .A(n18289), .B(n16787), .ZN(
        n16789) );
  AOI211_X1 U20004 ( .C1(n16903), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16790), .B(n16789), .ZN(n16793) );
  INV_X1 U20005 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18866) );
  AND2_X1 U20006 ( .A1(n16791), .A2(n16808), .ZN(n16802) );
  OAI221_X1 U20007 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n18868), .C2(n18866), .A(n16802), .ZN(n16792) );
  OAI211_X1 U20008 ( .C1(n16794), .C2(n18868), .A(n16793), .B(n16792), .ZN(
        P3_U2652) );
  AOI211_X1 U20009 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16809), .A(n16795), .B(
        n17022), .ZN(n16796) );
  AOI211_X1 U20010 ( .C1(n17006), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9768), .B(
        n16796), .ZN(n16804) );
  AOI22_X1 U20011 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16797), .B1(
        n17723), .B2(n17726), .ZN(n17738) );
  NAND2_X1 U20012 ( .A1(n9921), .A2(n16798), .ZN(n16800) );
  OAI21_X1 U20013 ( .B1(n17738), .B2(n16800), .A(n16987), .ZN(n16799) );
  AOI21_X1 U20014 ( .B1(n17738), .B2(n16800), .A(n16799), .ZN(n16801) );
  AOI221_X1 U20015 ( .B1(n16815), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16802), 
        .C2(n18866), .A(n16801), .ZN(n16803) );
  OAI211_X1 U20016 ( .C1(n17726), .C2(n17013), .A(n16804), .B(n16803), .ZN(
        P3_U2653) );
  INV_X1 U20017 ( .A(n16828), .ZN(n16805) );
  NAND2_X1 U20018 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16805), .ZN(
        n16806) );
  OAI21_X1 U20019 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16805), .A(
        n16806), .ZN(n17766) );
  AOI21_X1 U20020 ( .B1(n16818), .B2(n17766), .A(n9920), .ZN(n16807) );
  AOI21_X1 U20021 ( .B1(n17750), .B2(n16806), .A(n17723), .ZN(n17752) );
  XNOR2_X1 U20022 ( .A(n16807), .B(n17752), .ZN(n16817) );
  OAI22_X1 U20023 ( .A1(n17750), .A2(n17013), .B1(n17023), .B2(n21210), .ZN(
        n16814) );
  NAND2_X1 U20024 ( .A1(n16808), .A2(n18865), .ZN(n16811) );
  OAI211_X1 U20025 ( .C1(n16819), .C2(n21210), .A(n16977), .B(n16809), .ZN(
        n16810) );
  OAI211_X1 U20026 ( .C1(n16812), .C2(n16811), .A(n18289), .B(n16810), .ZN(
        n16813) );
  AOI211_X1 U20027 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n16815), .A(n16814), 
        .B(n16813), .ZN(n16816) );
  OAI21_X1 U20028 ( .B1(n18811), .B2(n16817), .A(n16816), .ZN(P3_U2654) );
  NOR2_X1 U20029 ( .A1(n16818), .A2(n9920), .ZN(n16832) );
  XOR2_X1 U20030 ( .A(n16832), .B(n17766), .Z(n16827) );
  AOI211_X1 U20031 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16833), .A(n16819), .B(
        n17022), .ZN(n16822) );
  INV_X1 U20032 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18860) );
  NOR3_X1 U20033 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18860), .A3(n16824), 
        .ZN(n16821) );
  INV_X1 U20034 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17761) );
  OAI22_X1 U20035 ( .A1(n17761), .A2(n17013), .B1(n17023), .B2(n17188), .ZN(
        n16820) );
  NOR4_X1 U20036 ( .A1(n9768), .A2(n16822), .A3(n16821), .A4(n16820), .ZN(
        n16826) );
  OAI21_X1 U20037 ( .B1(n16823), .B2(n17015), .A(n17025), .ZN(n16841) );
  NOR2_X1 U20038 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16824), .ZN(n16830) );
  OAI21_X1 U20039 ( .B1(n16841), .B2(n16830), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16825) );
  OAI211_X1 U20040 ( .C1(n18811), .C2(n16827), .A(n16826), .B(n16825), .ZN(
        P3_U2655) );
  AOI22_X1 U20041 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16903), .B1(
        P3_REIP_REG_15__SCAN_IN), .B2(n16841), .ZN(n16838) );
  AOI21_X1 U20042 ( .B1(n9921), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18811), .ZN(n17019) );
  OAI21_X1 U20043 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17764), .A(
        n16828), .ZN(n17772) );
  AOI21_X1 U20044 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17009), .A(
        n17772), .ZN(n16831) );
  OAI21_X1 U20045 ( .B1(n17023), .B2(n16834), .A(n18289), .ZN(n16829) );
  AOI211_X1 U20046 ( .C1(n17019), .C2(n16831), .A(n16830), .B(n16829), .ZN(
        n16837) );
  NAND3_X1 U20047 ( .A1(n16987), .A2(n16832), .A3(n17772), .ZN(n16836) );
  OAI211_X1 U20048 ( .C1(n16840), .C2(n16834), .A(n16977), .B(n16833), .ZN(
        n16835) );
  NAND4_X1 U20049 ( .A1(n16838), .A2(n16837), .A3(n16836), .A4(n16835), .ZN(
        P3_U2656) );
  AOI21_X1 U20050 ( .B1(n17787), .B2(n16850), .A(n17764), .ZN(n17789) );
  INV_X1 U20051 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21127) );
  NAND2_X1 U20052 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n21127), .ZN(
        n16999) );
  INV_X1 U20053 ( .A(n17014), .ZN(n16976) );
  OAI21_X1 U20054 ( .B1(n17786), .B2(n16999), .A(n16976), .ZN(n16862) );
  NOR4_X1 U20055 ( .A1(n16839), .A2(n21048), .A3(n17015), .A4(n16852), .ZN(
        n16846) );
  AOI211_X1 U20056 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16854), .A(n16840), .B(
        n17022), .ZN(n16845) );
  OAI21_X1 U20057 ( .B1(n17023), .B2(n17216), .A(n18289), .ZN(n16844) );
  AOI22_X1 U20058 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16903), .B1(
        P3_REIP_REG_14__SCAN_IN), .B2(n16841), .ZN(n16842) );
  INV_X1 U20059 ( .A(n16842), .ZN(n16843) );
  NOR4_X1 U20060 ( .A1(n16846), .A2(n16845), .A3(n16844), .A4(n16843), .ZN(
        n16849) );
  NOR2_X1 U20061 ( .A1(n17786), .A2(n16999), .ZN(n16847) );
  OAI211_X1 U20062 ( .C1(n16847), .C2(n9920), .A(n16987), .B(n17789), .ZN(
        n16848) );
  OAI211_X1 U20063 ( .C1(n17789), .C2(n16862), .A(n16849), .B(n16848), .ZN(
        P3_U2657) );
  INV_X1 U20064 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16865) );
  INV_X1 U20065 ( .A(n17801), .ZN(n16876) );
  NOR2_X1 U20066 ( .A1(n16865), .A2(n16876), .ZN(n16864) );
  OAI21_X1 U20067 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16864), .A(
        n16850), .ZN(n17803) );
  INV_X1 U20068 ( .A(n17803), .ZN(n16863) );
  INV_X1 U20069 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16851) );
  OAI21_X1 U20070 ( .B1(n16851), .B2(n9920), .A(n17019), .ZN(n16861) );
  NOR2_X1 U20071 ( .A1(n17015), .A2(n16852), .ZN(n16859) );
  INV_X1 U20072 ( .A(n16869), .ZN(n16853) );
  AOI21_X1 U20073 ( .B1(n17001), .B2(n16853), .A(n17012), .ZN(n16880) );
  OAI21_X1 U20074 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17015), .A(n16880), 
        .ZN(n16858) );
  AOI21_X1 U20075 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16903), .A(
        n9768), .ZN(n16856) );
  OAI211_X1 U20076 ( .C1(n16867), .C2(n17215), .A(n16977), .B(n16854), .ZN(
        n16855) );
  OAI211_X1 U20077 ( .C1(n17215), .C2(n17023), .A(n16856), .B(n16855), .ZN(
        n16857) );
  AOI221_X1 U20078 ( .B1(n16859), .B2(n21048), .C1(n16858), .C2(
        P3_REIP_REG_13__SCAN_IN), .A(n16857), .ZN(n16860) );
  OAI221_X1 U20079 ( .B1(n16863), .B2(n16862), .C1(n17803), .C2(n16861), .A(
        n16860), .ZN(P3_U2658) );
  OAI21_X1 U20080 ( .B1(n17799), .B2(n16999), .A(n9921), .ZN(n16866) );
  AOI21_X1 U20081 ( .B1(n16865), .B2(n16876), .A(n16864), .ZN(n17811) );
  XOR2_X1 U20082 ( .A(n16866), .B(n17811), .Z(n16874) );
  AOI211_X1 U20083 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16882), .A(n16867), .B(
        n17022), .ZN(n16872) );
  INV_X1 U20084 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18855) );
  NOR2_X1 U20085 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17015), .ZN(n16868) );
  AOI22_X1 U20086 ( .A1(n17006), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16869), 
        .B2(n16868), .ZN(n16870) );
  OAI211_X1 U20087 ( .C1(n16880), .C2(n18855), .A(n16870), .B(n18289), .ZN(
        n16871) );
  AOI211_X1 U20088 ( .C1(n16903), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16872), .B(n16871), .ZN(n16873) );
  OAI21_X1 U20089 ( .B1(n16874), .B2(n18811), .A(n16873), .ZN(P3_U2659) );
  INV_X1 U20090 ( .A(n16888), .ZN(n16875) );
  NOR2_X1 U20091 ( .A1(n17015), .A2(n16886), .ZN(n16899) );
  AOI21_X1 U20092 ( .B1(n16875), .B2(n16899), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16879) );
  NOR2_X1 U20093 ( .A1(n17018), .A2(n17822), .ZN(n16894) );
  OAI21_X1 U20094 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16894), .A(
        n16876), .ZN(n17823) );
  OAI21_X1 U20095 ( .B1(n17822), .B2(n16999), .A(n9921), .ZN(n16877) );
  XNOR2_X1 U20096 ( .A(n17823), .B(n16877), .ZN(n16878) );
  OAI22_X1 U20097 ( .A1(n16880), .A2(n16879), .B1(n18811), .B2(n16878), .ZN(
        n16881) );
  AOI211_X1 U20098 ( .C1(n17006), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9768), .B(
        n16881), .ZN(n16885) );
  OAI211_X1 U20099 ( .C1(n16887), .C2(n16883), .A(n16977), .B(n16882), .ZN(
        n16884) );
  OAI211_X1 U20100 ( .C1(n17013), .C2(n17825), .A(n16885), .B(n16884), .ZN(
        P3_U2660) );
  AOI21_X1 U20101 ( .B1(n17001), .B2(n16886), .A(n17012), .ZN(n16923) );
  INV_X1 U20102 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18851) );
  AOI211_X1 U20103 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16900), .A(n16887), .B(
        n17022), .ZN(n16892) );
  INV_X1 U20104 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16890) );
  OAI211_X1 U20105 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16899), .B(n16888), .ZN(n16889) );
  OAI211_X1 U20106 ( .C1(n17023), .C2(n16890), .A(n18289), .B(n16889), .ZN(
        n16891) );
  AOI211_X1 U20107 ( .C1(n16903), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16892), .B(n16891), .ZN(n16898) );
  INV_X1 U20108 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16905) );
  NAND2_X1 U20109 ( .A1(n17863), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17862) );
  NOR2_X1 U20110 ( .A1(n17018), .A2(n17862), .ZN(n16924) );
  NAND2_X1 U20111 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16924), .ZN(
        n16918) );
  NOR2_X1 U20112 ( .A1(n16905), .A2(n16918), .ZN(n16904) );
  INV_X1 U20113 ( .A(n16904), .ZN(n16893) );
  OAI21_X1 U20114 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16893), .A(
        n9921), .ZN(n16906) );
  INV_X1 U20115 ( .A(n16894), .ZN(n16895) );
  OAI21_X1 U20116 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16904), .A(
        n16895), .ZN(n17842) );
  AOI21_X1 U20117 ( .B1(n16906), .B2(n17842), .A(n18811), .ZN(n16896) );
  OAI21_X1 U20118 ( .B1(n16906), .B2(n17842), .A(n16896), .ZN(n16897) );
  OAI211_X1 U20119 ( .C1(n16923), .C2(n18851), .A(n16898), .B(n16897), .ZN(
        P3_U2661) );
  INV_X1 U20120 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18849) );
  AOI22_X1 U20121 ( .A1(n17006), .A2(P3_EBX_REG_9__SCAN_IN), .B1(n16899), .B2(
        n18849), .ZN(n16912) );
  OAI211_X1 U20122 ( .C1(n16913), .C2(n17263), .A(n16977), .B(n16900), .ZN(
        n16901) );
  OAI21_X1 U20123 ( .B1(n16923), .B2(n18849), .A(n16901), .ZN(n16902) );
  AOI21_X1 U20124 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16903), .A(
        n16902), .ZN(n16911) );
  INV_X1 U20125 ( .A(n17861), .ZN(n16907) );
  AOI21_X1 U20126 ( .B1(n16905), .B2(n16918), .A(n16904), .ZN(n17849) );
  INV_X1 U20127 ( .A(n16999), .ZN(n16964) );
  NAND2_X1 U20128 ( .A1(n17863), .A2(n16964), .ZN(n16932) );
  AOI221_X1 U20129 ( .B1(n16907), .B2(n17849), .C1(n16932), .C2(n17849), .A(
        n16906), .ZN(n16909) );
  INV_X1 U20130 ( .A(n17009), .ZN(n16908) );
  AOI22_X1 U20131 ( .A1(n16987), .A2(n16909), .B1(n17849), .B2(n16908), .ZN(
        n16910) );
  NAND4_X1 U20132 ( .A1(n16912), .A2(n16911), .A3(n16910), .A4(n18289), .ZN(
        P3_U2662) );
  INV_X1 U20133 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18848) );
  AOI211_X1 U20134 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16928), .A(n16913), .B(
        n17022), .ZN(n16917) );
  NAND3_X1 U20135 ( .A1(n17001), .A2(n16914), .A3(n18848), .ZN(n16915) );
  OAI211_X1 U20136 ( .C1(n17865), .C2(n17013), .A(n18289), .B(n16915), .ZN(
        n16916) );
  AOI211_X1 U20137 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17006), .A(n16917), .B(
        n16916), .ZN(n16922) );
  OAI21_X1 U20138 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16924), .A(
        n16918), .ZN(n17867) );
  OAI21_X1 U20139 ( .B1(n17862), .B2(n16999), .A(n9921), .ZN(n16920) );
  AOI21_X1 U20140 ( .B1(n17867), .B2(n16920), .A(n18811), .ZN(n16919) );
  OAI21_X1 U20141 ( .B1(n17867), .B2(n16920), .A(n16919), .ZN(n16921) );
  OAI211_X1 U20142 ( .C1(n16923), .C2(n18848), .A(n16922), .B(n16921), .ZN(
        P3_U2663) );
  NOR2_X1 U20143 ( .A1(n17018), .A2(n17832), .ZN(n16950) );
  NAND2_X1 U20144 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16950), .ZN(
        n16936) );
  AOI21_X1 U20145 ( .B1(n17883), .B2(n16936), .A(n16924), .ZN(n17887) );
  NAND2_X1 U20146 ( .A1(n16976), .A2(n16932), .ZN(n16945) );
  INV_X1 U20147 ( .A(n16925), .ZN(n16947) );
  NOR3_X1 U20148 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17015), .A3(n16947), .ZN(
        n16941) );
  OAI21_X1 U20149 ( .B1(n16925), .B2(n17015), .A(n17025), .ZN(n16939) );
  NOR3_X1 U20150 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17015), .A3(n16926), .ZN(
        n16927) );
  AOI211_X1 U20151 ( .C1(n17006), .C2(P3_EBX_REG_7__SCAN_IN), .A(n9768), .B(
        n16927), .ZN(n16930) );
  OAI211_X1 U20152 ( .C1(n16937), .C2(n17306), .A(n16977), .B(n16928), .ZN(
        n16929) );
  OAI211_X1 U20153 ( .C1(n17013), .C2(n17883), .A(n16930), .B(n16929), .ZN(
        n16931) );
  AOI221_X1 U20154 ( .B1(n16941), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n16939), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n16931), .ZN(n16935) );
  INV_X1 U20155 ( .A(n16932), .ZN(n16933) );
  OAI211_X1 U20156 ( .C1(n16933), .C2(n9920), .A(n16987), .B(n17887), .ZN(
        n16934) );
  OAI211_X1 U20157 ( .C1(n17887), .C2(n16945), .A(n16935), .B(n16934), .ZN(
        P3_U2664) );
  OAI21_X1 U20158 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16950), .A(
        n16936), .ZN(n17897) );
  INV_X1 U20159 ( .A(n17897), .ZN(n16946) );
  AOI211_X1 U20160 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16956), .A(n16937), .B(
        n17022), .ZN(n16938) );
  AOI211_X1 U20161 ( .C1(n17006), .C2(P3_EBX_REG_6__SCAN_IN), .A(n9768), .B(
        n16938), .ZN(n16944) );
  AOI21_X1 U20162 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9921), .A(
        n17897), .ZN(n16942) );
  INV_X1 U20163 ( .A(n16939), .ZN(n16953) );
  INV_X1 U20164 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18843) );
  OAI22_X1 U20165 ( .A1(n16953), .A2(n18843), .B1(n17896), .B2(n17013), .ZN(
        n16940) );
  AOI211_X1 U20166 ( .C1(n17019), .C2(n16942), .A(n16941), .B(n16940), .ZN(
        n16943) );
  OAI211_X1 U20167 ( .C1(n16946), .C2(n16945), .A(n16944), .B(n16943), .ZN(
        P3_U2665) );
  INV_X1 U20168 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16959) );
  NAND2_X1 U20169 ( .A1(n17001), .A2(n16947), .ZN(n16948) );
  OAI22_X1 U20170 ( .A1(n17023), .A2(n17312), .B1(n16949), .B2(n16948), .ZN(
        n16955) );
  NAND2_X1 U20171 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17901), .ZN(
        n16960) );
  AOI21_X1 U20172 ( .B1(n16959), .B2(n16960), .A(n16950), .ZN(n17909) );
  INV_X1 U20173 ( .A(n16960), .ZN(n16951) );
  AOI21_X1 U20174 ( .B1(n21127), .B2(n16951), .A(n9920), .ZN(n16963) );
  XNOR2_X1 U20175 ( .A(n17909), .B(n16963), .ZN(n16952) );
  OAI22_X1 U20176 ( .A1(n16953), .A2(n18841), .B1(n18811), .B2(n16952), .ZN(
        n16954) );
  NOR3_X1 U20177 ( .A1(n9768), .A2(n16955), .A3(n16954), .ZN(n16958) );
  OAI211_X1 U20178 ( .C1(n16965), .C2(n17312), .A(n16977), .B(n16956), .ZN(
        n16957) );
  OAI211_X1 U20179 ( .C1(n17013), .C2(n16959), .A(n16958), .B(n16957), .ZN(
        P3_U2666) );
  NOR2_X1 U20180 ( .A1(n17018), .A2(n17922), .ZN(n16975) );
  OAI21_X1 U20181 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16975), .A(
        n16960), .ZN(n17925) );
  OAI21_X1 U20182 ( .B1(n16961), .B2(n17015), .A(n17025), .ZN(n16986) );
  NAND2_X1 U20183 ( .A1(n17001), .A2(n16961), .ZN(n16962) );
  OAI22_X1 U20184 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16962), .B1(n17924), 
        .B2(n17013), .ZN(n16973) );
  NOR2_X1 U20185 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17922), .ZN(
        n17918) );
  AOI22_X1 U20186 ( .A1(n16964), .A2(n17918), .B1(n16963), .B2(n17925), .ZN(
        n16971) );
  AOI211_X1 U20187 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16978), .A(n16965), .B(
        n17022), .ZN(n16969) );
  NAND2_X1 U20188 ( .A1(n18307), .A2(n18976), .ZN(n16992) );
  AOI21_X1 U20189 ( .B1(n16967), .B2(n16966), .A(n16992), .ZN(n16968) );
  AOI211_X1 U20190 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17006), .A(n16969), .B(
        n16968), .ZN(n16970) );
  OAI211_X1 U20191 ( .C1(n16971), .C2(n18811), .A(n16970), .B(n18289), .ZN(
        n16972) );
  AOI211_X1 U20192 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16986), .A(n16973), .B(
        n16972), .ZN(n16974) );
  OAI21_X1 U20193 ( .B1(n17925), .B2(n17009), .A(n16974), .ZN(P3_U2667) );
  INV_X1 U20194 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16982) );
  NAND2_X1 U20195 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16991) );
  AOI21_X1 U20196 ( .B1(n16982), .B2(n16991), .A(n16975), .ZN(n17935) );
  INV_X1 U20197 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17948) );
  OAI21_X1 U20198 ( .B1(n17948), .B2(n16999), .A(n16976), .ZN(n16998) );
  OAI21_X1 U20199 ( .B1(n17015), .B2(n17002), .A(n18837), .ZN(n16985) );
  OAI21_X1 U20200 ( .B1(n16994), .B2(n17320), .A(n16977), .ZN(n16980) );
  INV_X1 U20201 ( .A(n16978), .ZN(n16979) );
  AOI221_X1 U20202 ( .B1(n17320), .B2(n16980), .C1(n17023), .C2(n16980), .A(
        n16979), .ZN(n16984) );
  NAND2_X1 U20203 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18775) );
  NOR2_X1 U20204 ( .A1(n16981), .A2(n18775), .ZN(n16993) );
  INV_X1 U20205 ( .A(n16993), .ZN(n18760) );
  AOI21_X1 U20206 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18760), .A(
        n15871), .ZN(n18912) );
  OAI22_X1 U20207 ( .A1(n18912), .A2(n16992), .B1(n16982), .B2(n17013), .ZN(
        n16983) );
  AOI211_X1 U20208 ( .C1(n16986), .C2(n16985), .A(n16984), .B(n16983), .ZN(
        n16990) );
  NOR2_X1 U20209 ( .A1(n17948), .A2(n16999), .ZN(n16988) );
  OAI211_X1 U20210 ( .C1(n16988), .C2(n9920), .A(n16987), .B(n17935), .ZN(
        n16989) );
  OAI211_X1 U20211 ( .C1(n17935), .C2(n16998), .A(n16990), .B(n16989), .ZN(
        P3_U2668) );
  OAI21_X1 U20212 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16991), .ZN(n17945) );
  INV_X1 U20213 ( .A(n16992), .ZN(n18978) );
  AOI21_X1 U20214 ( .B1(n11534), .B2(n18778), .A(n16993), .ZN(n18924) );
  INV_X1 U20215 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17336) );
  INV_X1 U20216 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17330) );
  NAND2_X1 U20217 ( .A1(n17336), .A2(n17330), .ZN(n16995) );
  AOI211_X1 U20218 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16995), .A(n16994), .B(
        n17022), .ZN(n16997) );
  INV_X1 U20219 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18835) );
  OAI22_X1 U20220 ( .A1(n17948), .A2(n17013), .B1(n17025), .B2(n18835), .ZN(
        n16996) );
  AOI211_X1 U20221 ( .C1(n18978), .C2(n18924), .A(n16997), .B(n16996), .ZN(
        n17008) );
  INV_X1 U20222 ( .A(n17945), .ZN(n17000) );
  AOI21_X1 U20223 ( .B1(n17000), .B2(n16999), .A(n16998), .ZN(n17005) );
  OAI211_X1 U20224 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17002), .B(n17001), .ZN(n17003) );
  INV_X1 U20225 ( .A(n17003), .ZN(n17004) );
  AOI211_X1 U20226 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17006), .A(n17005), .B(
        n17004), .ZN(n17007) );
  OAI211_X1 U20227 ( .C1(n17945), .C2(n17009), .A(n17008), .B(n17007), .ZN(
        P3_U2669) );
  OAI21_X1 U20228 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17010), .ZN(n17332) );
  AND2_X1 U20229 ( .A1(n18778), .A2(n17011), .ZN(n18931) );
  AOI22_X1 U20230 ( .A1(n17012), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18931), 
        .B2(n18978), .ZN(n17021) );
  OAI21_X1 U20231 ( .B1(n21127), .B2(n17014), .A(n17013), .ZN(n17017) );
  OAI22_X1 U20232 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17015), .B1(n17023), 
        .B2(n17330), .ZN(n17016) );
  AOI221_X1 U20233 ( .B1(n17019), .B2(n17018), .C1(n17017), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17016), .ZN(n17020) );
  OAI211_X1 U20234 ( .C1(n17022), .C2(n17332), .A(n17021), .B(n17020), .ZN(
        P3_U2670) );
  INV_X1 U20235 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18948) );
  NAND2_X1 U20236 ( .A1(n17023), .A2(n17022), .ZN(n17024) );
  AOI22_X1 U20237 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17024), .B1(n18978), .B2(
        n16981), .ZN(n17027) );
  NAND3_X1 U20238 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18913), .A3(
        n17025), .ZN(n17026) );
  OAI211_X1 U20239 ( .C1(n17028), .C2(n18948), .A(n17027), .B(n17026), .ZN(
        P3_U2671) );
  INV_X1 U20240 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17029) );
  NOR2_X1 U20241 ( .A1(n17029), .A2(n17145), .ZN(n17108) );
  NAND4_X1 U20242 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17062), .A4(n17108), .ZN(n17030) );
  NOR3_X1 U20243 ( .A1(n17032), .A2(n17031), .A3(n17030), .ZN(n17033) );
  NAND4_X1 U20244 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(n17033), .ZN(n17036) );
  NOR2_X1 U20245 ( .A1(n17037), .A2(n17036), .ZN(n17061) );
  NAND2_X1 U20246 ( .A1(n17329), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17035) );
  NAND2_X1 U20247 ( .A1(n17061), .A2(n18343), .ZN(n17034) );
  OAI22_X1 U20248 ( .A1(n17061), .A2(n17035), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17034), .ZN(P3_U2672) );
  NAND2_X1 U20249 ( .A1(n17037), .A2(n17036), .ZN(n17038) );
  NAND2_X1 U20250 ( .A1(n17038), .A2(n17329), .ZN(n17060) );
  AOI22_X1 U20251 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20252 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20253 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20254 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17039) );
  NAND4_X1 U20255 ( .A1(n17042), .A2(n17041), .A3(n17040), .A4(n17039), .ZN(
        n17048) );
  AOI22_X1 U20256 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20257 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20258 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20259 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17043) );
  NAND4_X1 U20260 ( .A1(n17046), .A2(n17045), .A3(n17044), .A4(n17043), .ZN(
        n17047) );
  NOR2_X1 U20261 ( .A1(n17048), .A2(n17047), .ZN(n17065) );
  NOR2_X1 U20262 ( .A1(n17065), .A2(n17064), .ZN(n17063) );
  AOI22_X1 U20263 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17270), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17268), .ZN(n17052) );
  AOI22_X1 U20264 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U20265 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17296), .ZN(n17050) );
  AOI22_X1 U20266 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17252), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17049) );
  NAND4_X1 U20267 ( .A1(n17052), .A2(n17051), .A3(n17050), .A4(n17049), .ZN(
        n17058) );
  AOI22_X1 U20268 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20269 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n15869), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17267), .ZN(n17055) );
  AOI22_X1 U20270 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17288), .ZN(n17054) );
  AOI22_X1 U20271 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11477), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17053) );
  NAND4_X1 U20272 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        n17057) );
  NOR2_X1 U20273 ( .A1(n17058), .A2(n17057), .ZN(n17059) );
  XOR2_X1 U20274 ( .A(n17063), .B(n17059), .Z(n17347) );
  OAI22_X1 U20275 ( .A1(n17061), .A2(n17060), .B1(n17347), .B2(n17329), .ZN(
        P3_U2673) );
  NAND2_X1 U20276 ( .A1(n17078), .A2(n17062), .ZN(n17068) );
  AOI21_X1 U20277 ( .B1(n17065), .B2(n17064), .A(n17063), .ZN(n17351) );
  AOI22_X1 U20278 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17066), .B1(n17351), 
        .B2(n17334), .ZN(n17067) );
  OAI21_X1 U20279 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17068), .A(n17067), .ZN(
        P3_U2674) );
  NAND2_X1 U20280 ( .A1(n17329), .A2(n17069), .ZN(n17073) );
  AOI21_X1 U20281 ( .B1(n17071), .B2(n17075), .A(n17070), .ZN(n17358) );
  AOI22_X1 U20282 ( .A1(n17334), .A2(n17358), .B1(n17078), .B2(n17074), .ZN(
        n17072) );
  OAI21_X1 U20283 ( .B1(n17074), .B2(n17073), .A(n17072), .ZN(P3_U2676) );
  AOI21_X1 U20284 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17329), .A(n17083), .ZN(
        n17077) );
  OAI21_X1 U20285 ( .B1(n17079), .B2(n17076), .A(n17075), .ZN(n17366) );
  OAI22_X1 U20286 ( .A1(n17078), .A2(n17077), .B1(n17366), .B2(n17329), .ZN(
        P3_U2677) );
  AOI21_X1 U20287 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17329), .A(n17087), .ZN(
        n17082) );
  AOI21_X1 U20288 ( .B1(n17080), .B2(n17084), .A(n17079), .ZN(n17367) );
  INV_X1 U20289 ( .A(n17367), .ZN(n17081) );
  OAI22_X1 U20290 ( .A1(n17083), .A2(n17082), .B1(n17081), .B2(n17329), .ZN(
        P3_U2678) );
  AOI21_X1 U20291 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17329), .A(n17093), .ZN(
        n17086) );
  OAI21_X1 U20292 ( .B1(n17088), .B2(n17085), .A(n17084), .ZN(n17376) );
  OAI22_X1 U20293 ( .A1(n17087), .A2(n17086), .B1(n17376), .B2(n17329), .ZN(
        P3_U2679) );
  AOI22_X1 U20294 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17329), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n17094), .ZN(n17092) );
  AOI21_X1 U20295 ( .B1(n17090), .B2(n17089), .A(n17088), .ZN(n17377) );
  INV_X1 U20296 ( .A(n17377), .ZN(n17091) );
  OAI22_X1 U20297 ( .A1(n17093), .A2(n17092), .B1(n17091), .B2(n17329), .ZN(
        P3_U2680) );
  INV_X1 U20298 ( .A(n17094), .ZN(n17107) );
  AOI22_X1 U20299 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20300 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17103) );
  INV_X1 U20301 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U20302 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17095) );
  OAI21_X1 U20303 ( .B1(n9849), .B2(n21018), .A(n17095), .ZN(n17101) );
  AOI22_X1 U20304 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20305 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20306 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20307 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17096) );
  NAND4_X1 U20308 ( .A1(n17099), .A2(n17098), .A3(n17097), .A4(n17096), .ZN(
        n17100) );
  AOI211_X1 U20309 ( .C1(n15871), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17101), .B(n17100), .ZN(n17102) );
  NAND3_X1 U20310 ( .A1(n17104), .A2(n17103), .A3(n17102), .ZN(n17383) );
  INV_X1 U20311 ( .A(n17383), .ZN(n17106) );
  NAND3_X1 U20312 ( .A1(n17107), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17329), 
        .ZN(n17105) );
  OAI221_X1 U20313 ( .B1(n17107), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17329), 
        .C2(n17106), .A(n17105), .ZN(P3_U2681) );
  NOR2_X1 U20314 ( .A1(n17334), .A2(n17108), .ZN(n17131) );
  AOI22_X1 U20315 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20316 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20317 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20318 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17109) );
  NAND4_X1 U20319 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        n17118) );
  AOI22_X1 U20320 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20321 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20322 ( .A1(n15808), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20323 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17113) );
  NAND4_X1 U20324 ( .A1(n17116), .A2(n17115), .A3(n17114), .A4(n17113), .ZN(
        n17117) );
  OR2_X1 U20325 ( .A1(n17118), .A2(n17117), .ZN(n17391) );
  AOI22_X1 U20326 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17131), .B1(n17334), 
        .B2(n17391), .ZN(n17119) );
  OAI21_X1 U20327 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17120), .A(n17119), .ZN(
        P3_U2682) );
  AOI22_X1 U20328 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20329 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17129) );
  AOI22_X1 U20330 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17121) );
  OAI21_X1 U20331 ( .B1(n9849), .B2(n18329), .A(n17121), .ZN(n17127) );
  AOI22_X1 U20332 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20333 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20334 ( .A1(n17275), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20335 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17122) );
  NAND4_X1 U20336 ( .A1(n17125), .A2(n17124), .A3(n17123), .A4(n17122), .ZN(
        n17126) );
  AOI211_X1 U20337 ( .C1(n15871), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17127), .B(n17126), .ZN(n17128) );
  NAND3_X1 U20338 ( .A1(n17130), .A2(n17129), .A3(n17128), .ZN(n17396) );
  INV_X1 U20339 ( .A(n17396), .ZN(n17134) );
  OAI21_X1 U20340 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17132), .A(n17131), .ZN(
        n17133) );
  OAI21_X1 U20341 ( .B1(n17134), .B2(n17329), .A(n17133), .ZN(P3_U2683) );
  AOI22_X1 U20342 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20343 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20344 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20345 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17135) );
  NAND4_X1 U20346 ( .A1(n17138), .A2(n17137), .A3(n17136), .A4(n17135), .ZN(
        n17144) );
  AOI22_X1 U20347 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20348 ( .A1(n17275), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15819), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20349 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20350 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17139) );
  NAND4_X1 U20351 ( .A1(n17142), .A2(n17141), .A3(n17140), .A4(n17139), .ZN(
        n17143) );
  NOR2_X1 U20352 ( .A1(n17144), .A2(n17143), .ZN(n17405) );
  OAI21_X1 U20353 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17146), .A(n17145), .ZN(
        n17147) );
  AOI22_X1 U20354 ( .A1(n17334), .A2(n17405), .B1(n17147), .B2(n17329), .ZN(
        P3_U2684) );
  NAND2_X1 U20355 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17148), .ZN(n17161) );
  AOI22_X1 U20356 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20357 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20358 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20359 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9773), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17149) );
  NAND4_X1 U20360 ( .A1(n17152), .A2(n17151), .A3(n17150), .A4(n17149), .ZN(
        n17158) );
  AOI22_X1 U20361 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20362 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20363 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20364 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17153) );
  NAND4_X1 U20365 ( .A1(n17156), .A2(n17155), .A3(n17154), .A4(n17153), .ZN(
        n17157) );
  NOR2_X1 U20366 ( .A1(n17158), .A2(n17157), .ZN(n17409) );
  INV_X1 U20367 ( .A(n17331), .ZN(n17333) );
  NAND4_X1 U20368 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17172), .A3(n17333), 
        .A4(n17159), .ZN(n17160) );
  OAI221_X1 U20369 ( .B1(n17334), .B2(n17161), .C1(n17329), .C2(n17409), .A(
        n17160), .ZN(P3_U2685) );
  AOI22_X1 U20370 ( .A1(n15869), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20371 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20372 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20373 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15819), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17162) );
  NAND4_X1 U20374 ( .A1(n17165), .A2(n17164), .A3(n17163), .A4(n17162), .ZN(
        n17171) );
  AOI22_X1 U20375 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20376 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20377 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15891), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17167) );
  AOI22_X1 U20378 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17166) );
  NAND4_X1 U20379 ( .A1(n17169), .A2(n17168), .A3(n17167), .A4(n17166), .ZN(
        n17170) );
  NOR2_X1 U20380 ( .A1(n17171), .A2(n17170), .ZN(n17415) );
  AND2_X1 U20381 ( .A1(n17172), .A2(n17333), .ZN(n17174) );
  NOR2_X1 U20382 ( .A1(n17172), .A2(n17459), .ZN(n17176) );
  NAND2_X1 U20383 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17337), .ZN(n17173) );
  OAI22_X1 U20384 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17174), .B1(n17176), 
        .B2(n17173), .ZN(n17175) );
  OAI21_X1 U20385 ( .B1(n17415), .B2(n17329), .A(n17175), .ZN(P3_U2686) );
  INV_X1 U20386 ( .A(n17176), .ZN(n17190) );
  INV_X1 U20387 ( .A(n17315), .ZN(n17305) );
  OR2_X1 U20388 ( .A1(n17187), .A2(n17305), .ZN(n17189) );
  AOI22_X1 U20389 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20390 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20391 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20392 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17177) );
  NAND4_X1 U20393 ( .A1(n17180), .A2(n17179), .A3(n17178), .A4(n17177), .ZN(
        n17186) );
  AOI22_X1 U20394 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20395 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20396 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U20397 ( .A1(n15869), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17181) );
  NAND4_X1 U20398 ( .A1(n17184), .A2(n17183), .A3(n17182), .A4(n17181), .ZN(
        n17185) );
  NOR2_X1 U20399 ( .A1(n17186), .A2(n17185), .ZN(n17421) );
  OAI21_X1 U20400 ( .B1(n17187), .B2(n17305), .A(n17329), .ZN(n17203) );
  OAI222_X1 U20401 ( .A1(n17190), .A2(n17189), .B1(n17329), .B2(n17421), .C1(
        n17188), .C2(n17203), .ZN(P3_U2687) );
  AOI22_X1 U20402 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17275), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20403 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17288), .B1(
        n17249), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20404 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17268), .ZN(n17192) );
  AOI22_X1 U20405 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9773), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17191) );
  NAND4_X1 U20406 ( .A1(n17194), .A2(n17193), .A3(n17192), .A4(n17191), .ZN(
        n17201) );
  AOI22_X1 U20407 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17270), .ZN(n17199) );
  AOI22_X1 U20408 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17252), .ZN(n17198) );
  AOI22_X1 U20409 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9775), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20410 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17196) );
  NAND4_X1 U20411 ( .A1(n17199), .A2(n17198), .A3(n17197), .A4(n17196), .ZN(
        n17200) );
  NOR2_X1 U20412 ( .A1(n17201), .A2(n17200), .ZN(n17424) );
  INV_X1 U20413 ( .A(n17246), .ZN(n17232) );
  AOI21_X1 U20414 ( .B1(n17202), .B2(n17232), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n17204) );
  OAI22_X1 U20415 ( .A1(n17424), .A2(n17329), .B1(n17204), .B2(n17203), .ZN(
        P3_U2688) );
  AOI22_X1 U20416 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15819), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20417 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U20418 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20419 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17205) );
  NAND4_X1 U20420 ( .A1(n17208), .A2(n17207), .A3(n17206), .A4(n17205), .ZN(
        n17214) );
  AOI22_X1 U20421 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20422 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20423 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20424 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17209) );
  NAND4_X1 U20425 ( .A1(n17212), .A2(n17211), .A3(n17210), .A4(n17209), .ZN(
        n17213) );
  NOR2_X1 U20426 ( .A1(n17214), .A2(n17213), .ZN(n17427) );
  OAI221_X1 U20427 ( .B1(n17231), .B2(n17333), .C1(n17231), .C2(n17215), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n17219) );
  NOR2_X1 U20428 ( .A1(n17459), .A2(n17246), .ZN(n17217) );
  NAND4_X1 U20429 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17217), .A4(n17216), .ZN(n17218) );
  OAI211_X1 U20430 ( .C1(n17427), .C2(n17329), .A(n17219), .B(n17218), .ZN(
        P3_U2689) );
  AOI22_X1 U20431 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20432 ( .A1(n15871), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20433 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20434 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9773), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17220) );
  NAND4_X1 U20435 ( .A1(n17223), .A2(n17222), .A3(n17221), .A4(n17220), .ZN(
        n17230) );
  AOI22_X1 U20436 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20437 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20438 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20439 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17225) );
  NAND4_X1 U20440 ( .A1(n17228), .A2(n17227), .A3(n17226), .A4(n17225), .ZN(
        n17229) );
  NOR2_X1 U20441 ( .A1(n17230), .A2(n17229), .ZN(n17438) );
  OAI21_X1 U20442 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17232), .A(n17231), .ZN(
        n17233) );
  OAI21_X1 U20443 ( .B1(n17438), .B2(n17329), .A(n17233), .ZN(P3_U2691) );
  AOI22_X1 U20444 ( .A1(n15869), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20445 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20446 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17234) );
  OAI21_X1 U20447 ( .B1(n10200), .B2(n21082), .A(n17234), .ZN(n17240) );
  AOI22_X1 U20448 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20449 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20450 ( .A1(n15808), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20451 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17235) );
  NAND4_X1 U20452 ( .A1(n17238), .A2(n17237), .A3(n17236), .A4(n17235), .ZN(
        n17239) );
  AOI211_X1 U20453 ( .C1(n17276), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n17240), .B(n17239), .ZN(n17241) );
  NAND3_X1 U20454 ( .A1(n17243), .A2(n17242), .A3(n17241), .ZN(n17442) );
  INV_X1 U20455 ( .A(n17442), .ZN(n17248) );
  NOR3_X1 U20456 ( .A1(n17309), .A2(n17244), .A3(n17305), .ZN(n17283) );
  INV_X1 U20457 ( .A(n17283), .ZN(n17307) );
  NOR2_X1 U20458 ( .A1(n17245), .A2(n17307), .ZN(n17265) );
  OAI21_X1 U20459 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17265), .A(n17246), .ZN(
        n17247) );
  AOI22_X1 U20460 ( .A1(n17334), .A2(n17248), .B1(n17247), .B2(n17329), .ZN(
        P3_U2692) );
  AOI22_X1 U20461 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17249), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17262) );
  AOI22_X1 U20462 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U20463 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U20464 ( .B1(n9850), .B2(n21233), .A(n17251), .ZN(n17258) );
  AOI22_X1 U20465 ( .A1(n9775), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20466 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20467 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20468 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17253) );
  NAND4_X1 U20469 ( .A1(n17256), .A2(n17255), .A3(n17254), .A4(n17253), .ZN(
        n17257) );
  AOI211_X1 U20470 ( .C1(n17259), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n17258), .B(n17257), .ZN(n17260) );
  NAND3_X1 U20471 ( .A1(n17262), .A2(n17261), .A3(n17260), .ZN(n17445) );
  INV_X1 U20472 ( .A(n17445), .ZN(n17266) );
  NOR2_X1 U20473 ( .A1(n17263), .A2(n17307), .ZN(n17285) );
  OAI21_X1 U20474 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17285), .A(n17329), .ZN(
        n17264) );
  OAI22_X1 U20475 ( .A1(n17266), .A2(n17329), .B1(n17265), .B2(n17264), .ZN(
        P3_U2693) );
  AOI22_X1 U20476 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15869), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20477 ( .A1(n15808), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15868), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U20478 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U20479 ( .A1(n9773), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17271) );
  NAND4_X1 U20480 ( .A1(n17274), .A2(n17273), .A3(n17272), .A4(n17271), .ZN(
        n17282) );
  AOI22_X1 U20481 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20482 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17279) );
  AOI22_X1 U20483 ( .A1(n15878), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U20484 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17277) );
  NAND4_X1 U20485 ( .A1(n17280), .A2(n17279), .A3(n17278), .A4(n17277), .ZN(
        n17281) );
  NOR2_X1 U20486 ( .A1(n17282), .A2(n17281), .ZN(n17450) );
  OAI21_X1 U20487 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17283), .A(n17329), .ZN(
        n17284) );
  OAI22_X1 U20488 ( .A1(n17450), .A2(n17329), .B1(n17285), .B2(n17284), .ZN(
        P3_U2694) );
  AOI22_X1 U20489 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9775), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U20490 ( .A1(n17249), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20491 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9773), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20492 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11477), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17290) );
  NAND4_X1 U20493 ( .A1(n17293), .A2(n17292), .A3(n17291), .A4(n17290), .ZN(
        n17304) );
  AOI22_X1 U20494 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20495 ( .A1(n17259), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20496 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15819), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20497 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17299) );
  NAND4_X1 U20498 ( .A1(n17302), .A2(n17301), .A3(n17300), .A4(n17299), .ZN(
        n17303) );
  NOR2_X1 U20499 ( .A1(n17304), .A2(n17303), .ZN(n17458) );
  NOR3_X1 U20500 ( .A1(n17306), .A2(n17309), .A3(n17305), .ZN(n17311) );
  OAI21_X1 U20501 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17311), .A(n17307), .ZN(
        n17308) );
  AOI22_X1 U20502 ( .A1(n17334), .A2(n17458), .B1(n17308), .B2(n17329), .ZN(
        P3_U2695) );
  NOR3_X1 U20503 ( .A1(n17318), .A2(n17309), .A3(n17331), .ZN(n17314) );
  OAI21_X1 U20504 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17314), .A(n17329), .ZN(
        n17310) );
  INV_X1 U20505 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18347) );
  OAI22_X1 U20506 ( .A1(n17311), .A2(n17310), .B1(n18347), .B2(n17329), .ZN(
        P3_U2696) );
  NOR3_X1 U20507 ( .A1(n17312), .A2(n17318), .A3(n17331), .ZN(n17317) );
  AOI21_X1 U20508 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17329), .A(n17317), .ZN(
        n17313) );
  OAI22_X1 U20509 ( .A1(n17314), .A2(n17313), .B1(n21018), .B2(n17329), .ZN(
        P3_U2697) );
  OAI21_X1 U20510 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17315), .A(n17329), .ZN(
        n17316) );
  INV_X1 U20511 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18334) );
  OAI22_X1 U20512 ( .A1(n17317), .A2(n17316), .B1(n18334), .B2(n17329), .ZN(
        P3_U2698) );
  NOR2_X1 U20513 ( .A1(n17318), .A2(n17331), .ZN(n17322) );
  NAND2_X1 U20514 ( .A1(n17319), .A2(n17333), .ZN(n17323) );
  NOR2_X1 U20515 ( .A1(n17320), .A2(n17323), .ZN(n17325) );
  AOI21_X1 U20516 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17329), .A(n17325), .ZN(
        n17321) );
  OAI22_X1 U20517 ( .A1(n17322), .A2(n17321), .B1(n18329), .B2(n17329), .ZN(
        P3_U2699) );
  INV_X1 U20518 ( .A(n17323), .ZN(n17327) );
  AOI21_X1 U20519 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17329), .A(n17327), .ZN(
        n17324) );
  INV_X1 U20520 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18324) );
  OAI22_X1 U20521 ( .A1(n17325), .A2(n17324), .B1(n18324), .B2(n17329), .ZN(
        P3_U2700) );
  INV_X1 U20522 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18318) );
  AOI221_X1 U20523 ( .B1(n17326), .B2(n17337), .C1(n17459), .C2(n17337), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17328) );
  AOI211_X1 U20524 ( .C1(n17334), .C2(n18318), .A(n17328), .B(n17327), .ZN(
        P3_U2701) );
  OAI222_X1 U20525 ( .A1(n17332), .A2(n17331), .B1(n17330), .B2(n17337), .C1(
        n18313), .C2(n17329), .ZN(P3_U2702) );
  AOI22_X1 U20526 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17334), .B1(
        n17333), .B2(n17336), .ZN(n17335) );
  OAI21_X1 U20527 ( .B1(n17337), .B2(n17336), .A(n17335), .ZN(P3_U2703) );
  INV_X1 U20528 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17558) );
  INV_X1 U20529 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17552) );
  INV_X1 U20530 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17595) );
  INV_X1 U20531 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17565) );
  INV_X1 U20532 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17569) );
  INV_X1 U20533 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17567) );
  NOR2_X1 U20534 ( .A1(n17569), .A2(n17567), .ZN(n17338) );
  NAND4_X1 U20535 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(n17338), .ZN(n17460) );
  NAND4_X1 U20536 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .A4(P3_EAX_REG_12__SCAN_IN), .ZN(n17339)
         );
  INV_X1 U20537 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17579) );
  INV_X1 U20538 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17541) );
  INV_X1 U20539 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17539) );
  INV_X1 U20540 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17537) );
  NOR3_X1 U20541 ( .A1(n17541), .A2(n17539), .A3(n17537), .ZN(n17384) );
  NAND3_X1 U20542 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(n17384), .ZN(n17390) );
  INV_X1 U20543 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17545) );
  NAND2_X1 U20544 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17379), .ZN(n17378) );
  NAND2_X1 U20545 ( .A1(n17348), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17344) );
  NOR2_X2 U20546 ( .A1(n18336), .A2(n17487), .ZN(n17416) );
  OAI22_X1 U20547 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17385), .B1(n17434), 
        .B2(n17348), .ZN(n17341) );
  AOI22_X1 U20548 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17416), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17341), .ZN(n17342) );
  OAI21_X1 U20549 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17344), .A(n17342), .ZN(
        P3_U2704) );
  NOR2_X2 U20550 ( .A1(n17343), .A2(n17487), .ZN(n17417) );
  AOI22_X1 U20551 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17416), .ZN(n17346) );
  OAI211_X1 U20552 ( .C1(n17348), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17487), .B(
        n17344), .ZN(n17345) );
  OAI211_X1 U20553 ( .C1(n17347), .C2(n17480), .A(n17346), .B(n17345), .ZN(
        P3_U2705) );
  INV_X1 U20554 ( .A(n17348), .ZN(n17350) );
  OAI21_X1 U20555 ( .B1(n17434), .B2(n17558), .A(n9845), .ZN(n17349) );
  AOI22_X1 U20556 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17416), .B1(n17350), .B2(
        n17349), .ZN(n17353) );
  AOI22_X1 U20557 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17417), .B1(n17484), .B2(
        n17351), .ZN(n17352) );
  NAND2_X1 U20558 ( .A1(n17353), .A2(n17352), .ZN(P3_U2706) );
  AOI22_X1 U20559 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17416), .ZN(n17356) );
  OAI211_X1 U20560 ( .C1(n17354), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17487), .B(
        n9845), .ZN(n17355) );
  OAI211_X1 U20561 ( .C1(n17357), .C2(n17480), .A(n17356), .B(n17355), .ZN(
        P3_U2707) );
  INV_X1 U20562 ( .A(n17416), .ZN(n17382) );
  AOI22_X1 U20563 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17417), .B1(n17484), .B2(
        n17358), .ZN(n17361) );
  OAI211_X1 U20564 ( .C1(n17362), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17487), .B(
        n17359), .ZN(n17360) );
  OAI211_X1 U20565 ( .C1(n17382), .C2(n15226), .A(n17361), .B(n17360), .ZN(
        P3_U2708) );
  AOI22_X1 U20566 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17416), .ZN(n17365) );
  AOI211_X1 U20567 ( .C1(n17552), .C2(n17368), .A(n17362), .B(n17434), .ZN(
        n17363) );
  INV_X1 U20568 ( .A(n17363), .ZN(n17364) );
  OAI211_X1 U20569 ( .C1(n17366), .C2(n17480), .A(n17365), .B(n17364), .ZN(
        P3_U2709) );
  INV_X1 U20570 ( .A(n17417), .ZN(n17393) );
  AOI22_X1 U20571 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n17416), .B1(n17484), .B2(
        n17367), .ZN(n17371) );
  OAI211_X1 U20572 ( .C1(n17369), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17487), .B(
        n17368), .ZN(n17370) );
  OAI211_X1 U20573 ( .C1(n17393), .C2(n17453), .A(n17371), .B(n17370), .ZN(
        P3_U2710) );
  AOI22_X1 U20574 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17416), .ZN(n17375) );
  OAI211_X1 U20575 ( .C1(n17373), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17487), .B(
        n17372), .ZN(n17374) );
  OAI211_X1 U20576 ( .C1(n17376), .C2(n17480), .A(n17375), .B(n17374), .ZN(
        P3_U2711) );
  AOI22_X1 U20577 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17417), .B1(n17484), .B2(
        n17377), .ZN(n17381) );
  OAI211_X1 U20578 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17379), .A(n17487), .B(
        n17378), .ZN(n17380) );
  OAI211_X1 U20579 ( .C1(n17382), .C2(n18339), .A(n17381), .B(n17380), .ZN(
        P3_U2712) );
  NOR2_X1 U20580 ( .A1(n17459), .A2(n17418), .ZN(n17412) );
  NAND2_X1 U20581 ( .A1(n17412), .A2(n17545), .ZN(n17389) );
  AOI22_X1 U20582 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17416), .B1(n17484), .B2(
        n17383), .ZN(n17388) );
  INV_X1 U20583 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17535) );
  NAND2_X1 U20584 ( .A1(n17384), .A2(n17410), .ZN(n17397) );
  NAND2_X1 U20585 ( .A1(n17487), .A2(n17397), .ZN(n17400) );
  OAI21_X1 U20586 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17385), .A(n17400), .ZN(
        n17386) );
  AOI22_X1 U20587 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17417), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17386), .ZN(n17387) );
  OAI211_X1 U20588 ( .C1(n17390), .C2(n17389), .A(n17388), .B(n17387), .ZN(
        P3_U2713) );
  INV_X1 U20589 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U20590 ( .A1(n17391), .A2(n17484), .B1(BUF2_REG_21__SCAN_IN), .B2(
        n17416), .ZN(n17392) );
  OAI21_X1 U20591 ( .B1(n18330), .B2(n17393), .A(n17392), .ZN(n17394) );
  INV_X1 U20592 ( .A(n17394), .ZN(n17395) );
  OAI221_X1 U20593 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17397), .C1(n17543), 
        .C2(n17400), .A(n17395), .ZN(P3_U2714) );
  AOI22_X1 U20594 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17416), .B1(n17484), .B2(
        n17396), .ZN(n17399) );
  NAND2_X1 U20595 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17410), .ZN(n17406) );
  NOR2_X1 U20596 ( .A1(n17539), .A2(n17406), .ZN(n17401) );
  AOI22_X1 U20597 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17417), .B1(n17401), .B2(
        n17397), .ZN(n17398) );
  OAI211_X1 U20598 ( .C1(n17541), .C2(n17400), .A(n17399), .B(n17398), .ZN(
        P3_U2715) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17416), .ZN(n17404) );
  AOI211_X1 U20600 ( .C1(n17539), .C2(n17406), .A(n17401), .B(n17434), .ZN(
        n17402) );
  INV_X1 U20601 ( .A(n17402), .ZN(n17403) );
  OAI211_X1 U20602 ( .C1(n17405), .C2(n17480), .A(n17404), .B(n17403), .ZN(
        P3_U2716) );
  AOI22_X1 U20603 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17416), .ZN(n17408) );
  OAI211_X1 U20604 ( .C1(n17410), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17487), .B(
        n17406), .ZN(n17407) );
  OAI211_X1 U20605 ( .C1(n17409), .C2(n17480), .A(n17408), .B(n17407), .ZN(
        P3_U2717) );
  AOI22_X1 U20606 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17416), .ZN(n17414) );
  INV_X1 U20607 ( .A(n17410), .ZN(n17411) );
  OAI211_X1 U20608 ( .C1(n17412), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17487), .B(
        n17411), .ZN(n17413) );
  OAI211_X1 U20609 ( .C1(n17415), .C2(n17480), .A(n17414), .B(n17413), .ZN(
        P3_U2718) );
  AOI22_X1 U20610 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17417), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17416), .ZN(n17420) );
  OAI211_X1 U20611 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n9865), .A(n17487), .B(
        n17418), .ZN(n17419) );
  OAI211_X1 U20612 ( .C1(n17421), .C2(n17480), .A(n17420), .B(n17419), .ZN(
        P3_U2719) );
  AOI211_X1 U20613 ( .C1(n17595), .C2(n17425), .A(n17434), .B(n9865), .ZN(
        n17422) );
  AOI21_X1 U20614 ( .B1(n17485), .B2(BUF2_REG_15__SCAN_IN), .A(n17422), .ZN(
        n17423) );
  OAI21_X1 U20615 ( .B1(n17424), .B2(n17480), .A(n17423), .ZN(P3_U2720) );
  INV_X1 U20616 ( .A(n17425), .ZN(n17429) );
  AOI22_X1 U20617 ( .A1(n18343), .A2(n17426), .B1(P3_EAX_REG_14__SCAN_IN), 
        .B2(n17487), .ZN(n17428) );
  OAI222_X1 U20618 ( .A1(n17483), .A2(n17430), .B1(n17429), .B2(n17428), .C1(
        n17480), .C2(n17427), .ZN(P3_U2721) );
  NAND2_X1 U20619 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n17431) );
  NOR2_X1 U20620 ( .A1(n17459), .A2(n17454), .ZN(n17449) );
  NAND2_X1 U20621 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17449), .ZN(n17447) );
  NOR2_X1 U20622 ( .A1(n17431), .A2(n17447), .ZN(n17437) );
  NAND2_X1 U20623 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17437), .ZN(n17436) );
  NAND2_X1 U20624 ( .A1(n17436), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20625 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17485), .B1(n17484), .B2(
        n17432), .ZN(n17433) );
  OAI221_X1 U20626 ( .B1(n17436), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17435), 
        .C2(n17434), .A(n17433), .ZN(P3_U2722) );
  INV_X1 U20627 ( .A(n17436), .ZN(n17440) );
  AOI21_X1 U20628 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17487), .A(n17437), .ZN(
        n17439) );
  OAI222_X1 U20629 ( .A1(n17483), .A2(n17441), .B1(n17440), .B2(n17439), .C1(
        n17480), .C2(n17438), .ZN(P3_U2723) );
  INV_X1 U20630 ( .A(n17447), .ZN(n17452) );
  NAND2_X1 U20631 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17452), .ZN(n17444) );
  INV_X1 U20632 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17583) );
  INV_X1 U20633 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17581) );
  OAI21_X1 U20634 ( .B1(n17581), .B2(n17447), .A(n17487), .ZN(n17448) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17485), .B1(n17484), .B2(
        n17442), .ZN(n17443) );
  OAI221_X1 U20636 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17444), .C1(n17583), 
        .C2(n17448), .A(n17443), .ZN(P3_U2724) );
  AOI22_X1 U20637 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17485), .B1(n17484), .B2(
        n17445), .ZN(n17446) );
  OAI221_X1 U20638 ( .B1(n17448), .B2(n17581), .C1(n17448), .C2(n17447), .A(
        n17446), .ZN(P3_U2725) );
  AOI21_X1 U20639 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17487), .A(n17449), .ZN(
        n17451) );
  OAI222_X1 U20640 ( .A1(n17483), .A2(n17453), .B1(n17452), .B2(n17451), .C1(
        n17480), .C2(n17450), .ZN(P3_U2726) );
  NAND2_X1 U20641 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17485), .ZN(n17457) );
  OAI211_X1 U20642 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17455), .A(n17487), .B(
        n17454), .ZN(n17456) );
  OAI211_X1 U20643 ( .C1(n17458), .C2(n17480), .A(n17457), .B(n17456), .ZN(
        P3_U2727) );
  NOR2_X1 U20644 ( .A1(n17459), .A2(n17486), .ZN(n17478) );
  NAND2_X1 U20645 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17478), .ZN(n17474) );
  NOR2_X1 U20646 ( .A1(n17460), .A2(n17474), .ZN(n17463) );
  INV_X1 U20647 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17573) );
  NOR2_X1 U20648 ( .A1(n17567), .A2(n17474), .ZN(n17477) );
  AND2_X1 U20649 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17477), .ZN(n17473) );
  NAND2_X1 U20650 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17473), .ZN(n17464) );
  NOR2_X1 U20651 ( .A1(n17573), .A2(n17464), .ZN(n17467) );
  AOI21_X1 U20652 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17487), .A(n17467), .ZN(
        n17462) );
  OAI222_X1 U20653 ( .A1(n17483), .A2(n18340), .B1(n17463), .B2(n17462), .C1(
        n17480), .C2(n17461), .ZN(P3_U2728) );
  INV_X1 U20654 ( .A(n17464), .ZN(n17470) );
  AOI21_X1 U20655 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17487), .A(n17470), .ZN(
        n17466) );
  OAI222_X1 U20656 ( .A1(n18335), .A2(n17483), .B1(n17467), .B2(n17466), .C1(
        n17480), .C2(n17465), .ZN(P3_U2729) );
  AOI21_X1 U20657 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17487), .A(n17473), .ZN(
        n17469) );
  OAI222_X1 U20658 ( .A1(n18330), .A2(n17483), .B1(n17470), .B2(n17469), .C1(
        n17480), .C2(n17468), .ZN(P3_U2730) );
  AOI21_X1 U20659 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17487), .A(n17477), .ZN(
        n17472) );
  OAI222_X1 U20660 ( .A1(n18325), .A2(n17483), .B1(n17473), .B2(n17472), .C1(
        n17480), .C2(n17471), .ZN(P3_U2731) );
  INV_X1 U20661 ( .A(n17474), .ZN(n17482) );
  AOI21_X1 U20662 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17487), .A(n17482), .ZN(
        n17476) );
  OAI222_X1 U20663 ( .A1(n18320), .A2(n17483), .B1(n17477), .B2(n17476), .C1(
        n17480), .C2(n17475), .ZN(P3_U2732) );
  AOI21_X1 U20664 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17487), .A(n17478), .ZN(
        n17481) );
  OAI222_X1 U20665 ( .A1(n18314), .A2(n17483), .B1(n17482), .B2(n17481), .C1(
        n17480), .C2(n17479), .ZN(P3_U2733) );
  OAI211_X1 U20666 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17488), .A(n17487), .B(
        n17486), .ZN(n17489) );
  NAND2_X1 U20667 ( .A1(n17490), .A2(n17489), .ZN(P3_U2734) );
  NAND2_X1 U20668 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17680), .ZN(n18956) );
  NOR2_X1 U20669 ( .A1(n17530), .A2(n17491), .ZN(n17509) );
  AND2_X1 U20670 ( .A1(n17519), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20671 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n21041) );
  NAND2_X1 U20672 ( .A1(n17509), .A2(n17492), .ZN(n17508) );
  AOI22_X1 U20673 ( .A1(n17527), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17493) );
  OAI21_X1 U20674 ( .B1(n21041), .B2(n17508), .A(n17493), .ZN(P3_U2737) );
  AOI22_X1 U20675 ( .A1(n17527), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17494) );
  OAI21_X1 U20676 ( .B1(n17558), .B2(n17508), .A(n17494), .ZN(P3_U2738) );
  INV_X1 U20677 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U20678 ( .A1(n17527), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17495) );
  OAI21_X1 U20679 ( .B1(n17556), .B2(n17508), .A(n17495), .ZN(P3_U2739) );
  INV_X1 U20680 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20681 ( .A1(n17527), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17496) );
  OAI21_X1 U20682 ( .B1(n17554), .B2(n17508), .A(n17496), .ZN(P3_U2740) );
  AOI22_X1 U20683 ( .A1(n17527), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17497) );
  OAI21_X1 U20684 ( .B1(n17552), .B2(n17508), .A(n17497), .ZN(P3_U2741) );
  INV_X1 U20685 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U20686 ( .A1(n17527), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17498) );
  OAI21_X1 U20687 ( .B1(n17550), .B2(n17508), .A(n17498), .ZN(P3_U2742) );
  INV_X1 U20688 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n21145) );
  AOI22_X1 U20689 ( .A1(n17527), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17499) );
  OAI21_X1 U20690 ( .B1(n21145), .B2(n17508), .A(n17499), .ZN(P3_U2743) );
  INV_X1 U20691 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17547) );
  AOI22_X1 U20692 ( .A1(n17527), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17500) );
  OAI21_X1 U20693 ( .B1(n17547), .B2(n17508), .A(n17500), .ZN(P3_U2744) );
  AOI22_X1 U20694 ( .A1(n17527), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17501) );
  OAI21_X1 U20695 ( .B1(n17545), .B2(n17508), .A(n17501), .ZN(P3_U2745) );
  AOI22_X1 U20696 ( .A1(n17527), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17502) );
  OAI21_X1 U20697 ( .B1(n17543), .B2(n17508), .A(n17502), .ZN(P3_U2746) );
  AOI22_X1 U20698 ( .A1(n17527), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17503) );
  OAI21_X1 U20699 ( .B1(n17541), .B2(n17508), .A(n17503), .ZN(P3_U2747) );
  AOI22_X1 U20700 ( .A1(n17527), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17504) );
  OAI21_X1 U20701 ( .B1(n17539), .B2(n17508), .A(n17504), .ZN(P3_U2748) );
  AOI22_X1 U20702 ( .A1(n17527), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U20703 ( .B1(n17537), .B2(n17508), .A(n17505), .ZN(P3_U2749) );
  AOI22_X1 U20704 ( .A1(n17527), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U20705 ( .B1(n17535), .B2(n17508), .A(n17506), .ZN(P3_U2750) );
  AOI22_X1 U20706 ( .A1(n17527), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17507) );
  OAI21_X1 U20707 ( .B1(n9991), .B2(n17508), .A(n17507), .ZN(P3_U2751) );
  INV_X1 U20708 ( .A(n17509), .ZN(n17529) );
  AOI22_X1 U20709 ( .A1(n17527), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17510) );
  OAI21_X1 U20710 ( .B1(n17595), .B2(n17529), .A(n17510), .ZN(P3_U2752) );
  AOI22_X1 U20711 ( .A1(n17527), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17511) );
  OAI21_X1 U20712 ( .B1(n9990), .B2(n17529), .A(n17511), .ZN(P3_U2753) );
  INV_X1 U20713 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U20714 ( .A1(n17527), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17512) );
  OAI21_X1 U20715 ( .B1(n17588), .B2(n17529), .A(n17512), .ZN(P3_U2754) );
  INV_X1 U20716 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17586) );
  AOI22_X1 U20717 ( .A1(n17527), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17513) );
  OAI21_X1 U20718 ( .B1(n17586), .B2(n17529), .A(n17513), .ZN(P3_U2755) );
  AOI22_X1 U20719 ( .A1(n17527), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17514) );
  OAI21_X1 U20720 ( .B1(n17583), .B2(n17529), .A(n17514), .ZN(P3_U2756) );
  AOI22_X1 U20721 ( .A1(n17527), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17515) );
  OAI21_X1 U20722 ( .B1(n17581), .B2(n17529), .A(n17515), .ZN(P3_U2757) );
  AOI22_X1 U20723 ( .A1(n17527), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17516) );
  OAI21_X1 U20724 ( .B1(n17579), .B2(n17529), .A(n17516), .ZN(P3_U2758) );
  INV_X1 U20725 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17577) );
  AOI22_X1 U20726 ( .A1(n17527), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U20727 ( .B1(n17577), .B2(n17529), .A(n17517), .ZN(P3_U2759) );
  INV_X1 U20728 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17575) );
  AOI22_X1 U20729 ( .A1(n17527), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17518) );
  OAI21_X1 U20730 ( .B1(n17575), .B2(n17529), .A(n17518), .ZN(P3_U2760) );
  AOI22_X1 U20731 ( .A1(n17527), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17519), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17520) );
  OAI21_X1 U20732 ( .B1(n17573), .B2(n17529), .A(n17520), .ZN(P3_U2761) );
  INV_X1 U20733 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17571) );
  AOI22_X1 U20734 ( .A1(n17527), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U20735 ( .B1(n17571), .B2(n17529), .A(n17521), .ZN(P3_U2762) );
  AOI22_X1 U20736 ( .A1(n17527), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17522) );
  OAI21_X1 U20737 ( .B1(n17569), .B2(n17529), .A(n17522), .ZN(P3_U2763) );
  AOI22_X1 U20738 ( .A1(n17527), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U20739 ( .B1(n17567), .B2(n17529), .A(n17523), .ZN(P3_U2764) );
  AOI22_X1 U20740 ( .A1(n17527), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U20741 ( .B1(n17565), .B2(n17529), .A(n17524), .ZN(P3_U2765) );
  INV_X1 U20742 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U20743 ( .A1(n17527), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U20744 ( .B1(n17563), .B2(n17529), .A(n17525), .ZN(P3_U2766) );
  AOI22_X1 U20745 ( .A1(n17527), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17526), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U20746 ( .B1(n17561), .B2(n17529), .A(n17528), .ZN(P3_U2767) );
  INV_X1 U20747 ( .A(n17530), .ZN(n17531) );
  OAI211_X1 U20748 ( .C1(n18961), .C2(n18962), .A(n9764), .B(n17531), .ZN(
        n17584) );
  AOI22_X1 U20749 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17589), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17591), .ZN(n17533) );
  OAI21_X1 U20750 ( .B1(n9991), .B2(n17594), .A(n17533), .ZN(P3_U2768) );
  AOI22_X1 U20751 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17589), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17591), .ZN(n17534) );
  OAI21_X1 U20752 ( .B1(n17535), .B2(n17594), .A(n17534), .ZN(P3_U2769) );
  AOI22_X1 U20753 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17589), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17591), .ZN(n17536) );
  OAI21_X1 U20754 ( .B1(n17537), .B2(n17594), .A(n17536), .ZN(P3_U2770) );
  AOI22_X1 U20755 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17589), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17591), .ZN(n17538) );
  OAI21_X1 U20756 ( .B1(n17539), .B2(n17594), .A(n17538), .ZN(P3_U2771) );
  AOI22_X1 U20757 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17591), .ZN(n17540) );
  OAI21_X1 U20758 ( .B1(n17541), .B2(n17594), .A(n17540), .ZN(P3_U2772) );
  AOI22_X1 U20759 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17591), .ZN(n17542) );
  OAI21_X1 U20760 ( .B1(n17543), .B2(n17594), .A(n17542), .ZN(P3_U2773) );
  AOI22_X1 U20761 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17591), .ZN(n17544) );
  OAI21_X1 U20762 ( .B1(n17545), .B2(n17594), .A(n17544), .ZN(P3_U2774) );
  AOI22_X1 U20763 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17591), .ZN(n17546) );
  OAI21_X1 U20764 ( .B1(n17547), .B2(n17594), .A(n17546), .ZN(P3_U2775) );
  AOI22_X1 U20765 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17591), .ZN(n17548) );
  OAI21_X1 U20766 ( .B1(n21145), .B2(n17594), .A(n17548), .ZN(P3_U2776) );
  AOI22_X1 U20767 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17591), .ZN(n17549) );
  OAI21_X1 U20768 ( .B1(n17550), .B2(n17594), .A(n17549), .ZN(P3_U2777) );
  AOI22_X1 U20769 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17591), .ZN(n17551) );
  OAI21_X1 U20770 ( .B1(n17552), .B2(n17594), .A(n17551), .ZN(P3_U2778) );
  AOI22_X1 U20771 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17592), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17591), .ZN(n17553) );
  OAI21_X1 U20772 ( .B1(n17554), .B2(n17594), .A(n17553), .ZN(P3_U2779) );
  AOI22_X1 U20773 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17589), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17591), .ZN(n17555) );
  OAI21_X1 U20774 ( .B1(n17556), .B2(n17594), .A(n17555), .ZN(P3_U2780) );
  AOI22_X1 U20775 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17589), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17591), .ZN(n17557) );
  OAI21_X1 U20776 ( .B1(n17558), .B2(n17594), .A(n17557), .ZN(P3_U2781) );
  AOI22_X1 U20777 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17589), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17591), .ZN(n17559) );
  OAI21_X1 U20778 ( .B1(n21041), .B2(n17594), .A(n17559), .ZN(P3_U2782) );
  AOI22_X1 U20779 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17591), .ZN(n17560) );
  OAI21_X1 U20780 ( .B1(n17561), .B2(n17594), .A(n17560), .ZN(P3_U2783) );
  AOI22_X1 U20781 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17591), .ZN(n17562) );
  OAI21_X1 U20782 ( .B1(n17563), .B2(n17594), .A(n17562), .ZN(P3_U2784) );
  AOI22_X1 U20783 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17591), .ZN(n17564) );
  OAI21_X1 U20784 ( .B1(n17565), .B2(n17594), .A(n17564), .ZN(P3_U2785) );
  AOI22_X1 U20785 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17584), .ZN(n17566) );
  OAI21_X1 U20786 ( .B1(n17567), .B2(n17594), .A(n17566), .ZN(P3_U2786) );
  AOI22_X1 U20787 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17584), .ZN(n17568) );
  OAI21_X1 U20788 ( .B1(n17569), .B2(n17594), .A(n17568), .ZN(P3_U2787) );
  AOI22_X1 U20789 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17584), .ZN(n17570) );
  OAI21_X1 U20790 ( .B1(n17571), .B2(n17594), .A(n17570), .ZN(P3_U2788) );
  AOI22_X1 U20791 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17584), .ZN(n17572) );
  OAI21_X1 U20792 ( .B1(n17573), .B2(n17594), .A(n17572), .ZN(P3_U2789) );
  AOI22_X1 U20793 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17584), .ZN(n17574) );
  OAI21_X1 U20794 ( .B1(n17575), .B2(n17594), .A(n17574), .ZN(P3_U2790) );
  AOI22_X1 U20795 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17584), .ZN(n17576) );
  OAI21_X1 U20796 ( .B1(n17577), .B2(n17594), .A(n17576), .ZN(P3_U2791) );
  AOI22_X1 U20797 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17584), .ZN(n17578) );
  OAI21_X1 U20798 ( .B1(n17579), .B2(n17594), .A(n17578), .ZN(P3_U2792) );
  AOI22_X1 U20799 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17592), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17584), .ZN(n17580) );
  OAI21_X1 U20800 ( .B1(n17581), .B2(n17594), .A(n17580), .ZN(P3_U2793) );
  AOI22_X1 U20801 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17584), .ZN(n17582) );
  OAI21_X1 U20802 ( .B1(n17583), .B2(n17594), .A(n17582), .ZN(P3_U2794) );
  AOI22_X1 U20803 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17584), .ZN(n17585) );
  OAI21_X1 U20804 ( .B1(n17586), .B2(n17594), .A(n17585), .ZN(P3_U2795) );
  AOI22_X1 U20805 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17592), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17591), .ZN(n17587) );
  OAI21_X1 U20806 ( .B1(n17588), .B2(n17594), .A(n17587), .ZN(P3_U2796) );
  AOI22_X1 U20807 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17589), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17591), .ZN(n17590) );
  OAI21_X1 U20808 ( .B1(n9990), .B2(n17594), .A(n17590), .ZN(P3_U2797) );
  AOI22_X1 U20809 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17592), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17591), .ZN(n17593) );
  OAI21_X1 U20810 ( .B1(n17595), .B2(n17594), .A(n17593), .ZN(P3_U2798) );
  OAI22_X1 U20811 ( .A1(n17596), .A2(n17878), .B1(n17976), .B2(n17965), .ZN(
        n17632) );
  NOR2_X1 U20812 ( .A1(n17622), .A2(n17632), .ZN(n17623) );
  NAND2_X1 U20813 ( .A1(n17878), .A2(n17965), .ZN(n17709) );
  NAND2_X1 U20814 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17709), .ZN(
        n17611) );
  OAI21_X1 U20815 ( .B1(n17599), .B2(n17864), .A(n17960), .ZN(n17597) );
  AOI21_X1 U20816 ( .B1(n17680), .B2(n17598), .A(n17597), .ZN(n17626) );
  OAI21_X1 U20817 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17678), .A(
        n17626), .ZN(n17615) );
  NOR3_X1 U20818 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17622), .A3(
        n17621), .ZN(n17605) );
  AND2_X1 U20819 ( .A1(n17809), .A2(n17599), .ZN(n17619) );
  OAI211_X1 U20820 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17619), .B(n17600), .ZN(n17602) );
  OAI211_X1 U20821 ( .C1(n17802), .C2(n17603), .A(n17602), .B(n17601), .ZN(
        n17604) );
  AOI211_X1 U20822 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17615), .A(
        n17605), .B(n17604), .ZN(n17610) );
  OAI211_X1 U20823 ( .C1(n17608), .C2(n17607), .A(n17874), .B(n17606), .ZN(
        n17609) );
  OAI211_X1 U20824 ( .C1(n17623), .C2(n17611), .A(n17610), .B(n17609), .ZN(
        P3_U2802) );
  NAND2_X1 U20825 ( .A1(n16532), .A2(n17612), .ZN(n17613) );
  XNOR2_X1 U20826 ( .A(n17613), .B(n17873), .ZN(n17983) );
  AOI22_X1 U20827 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17615), .B1(
        n17812), .B2(n17614), .ZN(n17616) );
  NAND2_X1 U20828 ( .A1(n9768), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17981) );
  OAI211_X1 U20829 ( .C1(n17983), .C2(n17853), .A(n17616), .B(n17981), .ZN(
        n17617) );
  AOI21_X1 U20830 ( .B1(n17619), .B2(n17618), .A(n17617), .ZN(n17620) );
  OAI221_X1 U20831 ( .B1(n17623), .B2(n17622), .C1(n17623), .C2(n17621), .A(
        n17620), .ZN(P3_U2803) );
  AOI21_X1 U20832 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17625), .A(
        n17624), .ZN(n17991) );
  NAND2_X1 U20833 ( .A1(n17802), .A2(n17678), .ZN(n17934) );
  NOR2_X1 U20834 ( .A1(n18289), .A2(n18882), .ZN(n17989) );
  AOI221_X1 U20835 ( .B1(n18411), .B2(n17628), .C1(n17627), .C2(n17628), .A(
        n17626), .ZN(n17629) );
  AOI211_X1 U20836 ( .C1(n17630), .C2(n17934), .A(n17989), .B(n17629), .ZN(
        n17634) );
  AOI22_X1 U20837 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17632), .B1(
        n17631), .B2(n17985), .ZN(n17633) );
  OAI211_X1 U20838 ( .C1(n17991), .C2(n17853), .A(n17634), .B(n17633), .ZN(
        P3_U2804) );
  OAI21_X1 U20839 ( .B1(n17838), .B2(n17636), .A(n17635), .ZN(n17637) );
  XNOR2_X1 U20840 ( .A(n17637), .B(n17996), .ZN(n18002) );
  NOR2_X1 U20841 ( .A1(n17640), .A2(n18411), .ZN(n17662) );
  AOI211_X1 U20842 ( .C1(n17680), .C2(n17639), .A(n17921), .B(n17662), .ZN(
        n17667) );
  OAI21_X1 U20843 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17678), .A(
        n17667), .ZN(n17651) );
  NAND2_X1 U20844 ( .A1(n17640), .A2(n17809), .ZN(n17654) );
  AOI221_X1 U20845 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C1(n17653), .C2(n17641), .A(
        n17654), .ZN(n17644) );
  OAI22_X1 U20846 ( .A1(n18289), .A2(n18880), .B1(n17802), .B2(n17642), .ZN(
        n17643) );
  AOI211_X1 U20847 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17651), .A(
        n17644), .B(n17643), .ZN(n17649) );
  INV_X1 U20848 ( .A(n17878), .ZN(n17828) );
  AOI21_X1 U20849 ( .B1(n17996), .B2(n17646), .A(n17645), .ZN(n17994) );
  NOR2_X1 U20850 ( .A1(n17996), .A2(n17968), .ZN(n17966) );
  AOI22_X1 U20851 ( .A1(n17966), .A2(n18026), .B1(n17996), .B2(n17647), .ZN(
        n17998) );
  AOI22_X1 U20852 ( .A1(n17828), .A2(n17994), .B1(n17950), .B2(n17998), .ZN(
        n17648) );
  OAI211_X1 U20853 ( .C1(n17853), .C2(n18002), .A(n17649), .B(n17648), .ZN(
        P3_U2805) );
  NAND2_X1 U20854 ( .A1(n17650), .A2(n18010), .ZN(n18016) );
  INV_X1 U20855 ( .A(n17651), .ZN(n17652) );
  NAND2_X1 U20856 ( .A1(n9768), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18014) );
  OAI221_X1 U20857 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17654), .C1(
        n17653), .C2(n17652), .A(n18014), .ZN(n17659) );
  AOI22_X1 U20858 ( .A1(n17828), .A2(n17655), .B1(n17950), .B2(n18007), .ZN(
        n17677) );
  AOI21_X1 U20859 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17657), .A(
        n17656), .ZN(n18003) );
  OAI22_X1 U20860 ( .A1(n17677), .A2(n18010), .B1(n18003), .B2(n17853), .ZN(
        n17658) );
  AOI211_X1 U20861 ( .C1(n17812), .C2(n17660), .A(n17659), .B(n17658), .ZN(
        n17661) );
  OAI21_X1 U20862 ( .B1(n17771), .B2(n18016), .A(n17661), .ZN(P3_U2806) );
  NOR2_X1 U20863 ( .A1(n18289), .A2(n18876), .ZN(n18019) );
  NOR2_X1 U20864 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17678), .ZN(
        n17663) );
  AOI21_X1 U20865 ( .B1(n17663), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n17662), .ZN(n17665) );
  OAI22_X1 U20866 ( .A1(n17667), .A2(n17666), .B1(n17665), .B2(n17664), .ZN(
        n17668) );
  AOI211_X1 U20867 ( .C1(n17669), .C2(n17812), .A(n18019), .B(n17668), .ZN(
        n17676) );
  NOR2_X1 U20868 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17771), .ZN(
        n17674) );
  AOI22_X1 U20869 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17838), .B1(
        n17671), .B2(n17687), .ZN(n17672) );
  NAND2_X1 U20870 ( .A1(n17670), .A2(n17672), .ZN(n17673) );
  XNOR2_X1 U20871 ( .A(n17673), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18020) );
  AOI22_X1 U20872 ( .A1(n18018), .A2(n17674), .B1(n17874), .B2(n18020), .ZN(
        n17675) );
  OAI211_X1 U20873 ( .C1(n17677), .C2(n18023), .A(n17676), .B(n17675), .ZN(
        P3_U2807) );
  INV_X1 U20874 ( .A(n17678), .ZN(n17712) );
  AOI21_X1 U20875 ( .B1(n17680), .B2(n17679), .A(n17921), .ZN(n17681) );
  OAI21_X1 U20876 ( .B1(n17682), .B2(n17864), .A(n17681), .ZN(n17717) );
  AOI21_X1 U20877 ( .B1(n17712), .B2(n17710), .A(n17717), .ZN(n17695) );
  NOR2_X1 U20878 ( .A1(n18289), .A2(n18874), .ZN(n18038) );
  NAND2_X1 U20879 ( .A1(n17682), .A2(n17809), .ZN(n17697) );
  AOI211_X1 U20880 ( .C1(n17696), .C2(n17694), .A(n17683), .B(n17697), .ZN(
        n17684) );
  AOI211_X1 U20881 ( .C1(n17685), .C2(n17812), .A(n18038), .B(n17684), .ZN(
        n17693) );
  INV_X1 U20882 ( .A(n17670), .ZN(n17686) );
  AOI221_X1 U20883 ( .B1(n17759), .B2(n17687), .C1(n18031), .C2(n17687), .A(
        n17686), .ZN(n17688) );
  XNOR2_X1 U20884 ( .A(n17688), .B(n18041), .ZN(n18039) );
  NOR2_X1 U20885 ( .A1(n18031), .A2(n17771), .ZN(n17690) );
  NAND2_X1 U20886 ( .A1(n17828), .A2(n18027), .ZN(n17783) );
  OAI21_X1 U20887 ( .B1(n18026), .B2(n17965), .A(n17783), .ZN(n17742) );
  AOI21_X1 U20888 ( .B1(n18031), .B2(n17709), .A(n17742), .ZN(n17708) );
  INV_X1 U20889 ( .A(n17708), .ZN(n17689) );
  MUX2_X1 U20890 ( .A(n17690), .B(n17689), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17691) );
  AOI21_X1 U20891 ( .B1(n17874), .B2(n18039), .A(n17691), .ZN(n17692) );
  OAI211_X1 U20892 ( .C1(n17695), .C2(n17694), .A(n17693), .B(n17692), .ZN(
        P3_U2808) );
  NAND2_X1 U20893 ( .A1(n9768), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18051) );
  OAI221_X1 U20894 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17697), .C1(
        n17696), .C2(n17695), .A(n18051), .ZN(n17698) );
  AOI21_X1 U20895 ( .B1(n17812), .B2(n17699), .A(n17698), .ZN(n17706) );
  INV_X1 U20896 ( .A(n17704), .ZN(n18048) );
  NOR3_X1 U20897 ( .A1(n17838), .A2(n17737), .A3(n17700), .ZN(n17730) );
  INV_X1 U20898 ( .A(n17701), .ZN(n17731) );
  AOI22_X1 U20899 ( .A1(n18048), .A2(n17730), .B1(n17731), .B2(n17702), .ZN(
        n17703) );
  XNOR2_X1 U20900 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17703), .ZN(
        n18045) );
  NOR2_X1 U20901 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17704), .ZN(
        n18044) );
  NOR2_X1 U20902 ( .A1(n18043), .A2(n17771), .ZN(n17733) );
  AOI22_X1 U20903 ( .A1(n17874), .A2(n18045), .B1(n18044), .B2(n17733), .ZN(
        n17705) );
  OAI211_X1 U20904 ( .C1(n17708), .C2(n17707), .A(n17706), .B(n17705), .ZN(
        P3_U2809) );
  INV_X1 U20905 ( .A(n18043), .ZN(n18046) );
  NAND2_X1 U20906 ( .A1(n18046), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18053) );
  AOI21_X1 U20907 ( .B1(n17709), .B2(n18053), .A(n17742), .ZN(n17736) );
  INV_X1 U20908 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18058) );
  OAI21_X1 U20909 ( .B1(n17711), .B2(n18411), .A(n17710), .ZN(n17716) );
  INV_X1 U20910 ( .A(n17713), .ZN(n17714) );
  AOI21_X1 U20911 ( .B1(n17802), .B2(n17678), .A(n17714), .ZN(n17715) );
  NOR2_X1 U20912 ( .A1(n18289), .A2(n18871), .ZN(n18061) );
  AOI211_X1 U20913 ( .C1(n17717), .C2(n17716), .A(n17715), .B(n18061), .ZN(
        n17721) );
  OAI221_X1 U20914 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17744), 
        .C1(n18070), .C2(n17730), .A(n17670), .ZN(n17718) );
  XOR2_X1 U20915 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17718), .Z(
        n18064) );
  INV_X1 U20916 ( .A(n18064), .ZN(n17719) );
  NOR2_X1 U20917 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18070), .ZN(
        n18062) );
  AOI22_X1 U20918 ( .A1(n17874), .A2(n17719), .B1(n17733), .B2(n18062), .ZN(
        n17720) );
  OAI211_X1 U20919 ( .C1(n17736), .C2(n18058), .A(n17721), .B(n17720), .ZN(
        P3_U2810) );
  OAI21_X1 U20920 ( .B1(n17921), .B2(n17722), .A(n17954), .ZN(n17748) );
  OAI21_X1 U20921 ( .B1(n17723), .B2(n17961), .A(n17748), .ZN(n17741) );
  INV_X1 U20922 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17725) );
  NAND2_X1 U20923 ( .A1(n17724), .A2(n17809), .ZN(n17739) );
  AOI221_X1 U20924 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n17726), .C2(n17725), .A(
        n17739), .ZN(n17729) );
  OAI22_X1 U20925 ( .A1(n18289), .A2(n18868), .B1(n17802), .B2(n17727), .ZN(
        n17728) );
  AOI211_X1 U20926 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17741), .A(
        n17729), .B(n17728), .ZN(n17735) );
  AOI21_X1 U20927 ( .B1(n17744), .B2(n17731), .A(n17730), .ZN(n17732) );
  XNOR2_X1 U20928 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17732), .ZN(
        n18066) );
  AOI22_X1 U20929 ( .A1(n17874), .A2(n18066), .B1(n17733), .B2(n18070), .ZN(
        n17734) );
  OAI211_X1 U20930 ( .C1(n17736), .C2(n18070), .A(n17735), .B(n17734), .ZN(
        P3_U2811) );
  NAND2_X1 U20931 ( .A1(n17743), .A2(n17737), .ZN(n18088) );
  NOR2_X1 U20932 ( .A1(n18289), .A2(n18866), .ZN(n18085) );
  OAI22_X1 U20933 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17739), .B1(
        n17738), .B2(n17802), .ZN(n17740) );
  AOI211_X1 U20934 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17741), .A(
        n18085), .B(n17740), .ZN(n17747) );
  INV_X1 U20935 ( .A(n17742), .ZN(n17770) );
  OAI21_X1 U20936 ( .B1(n17743), .B2(n17771), .A(n17770), .ZN(n17755) );
  AOI21_X1 U20937 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17873), .A(
        n17744), .ZN(n17745) );
  XNOR2_X1 U20938 ( .A(n17745), .B(n17701), .ZN(n18083) );
  AOI22_X1 U20939 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17755), .B1(
        n17874), .B2(n18083), .ZN(n17746) );
  OAI211_X1 U20940 ( .C1(n17771), .C2(n18088), .A(n17747), .B(n17746), .ZN(
        P3_U2812) );
  NAND2_X1 U20941 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18089), .ZN(
        n18095) );
  NOR2_X1 U20942 ( .A1(n18289), .A2(n18865), .ZN(n18092) );
  AOI221_X1 U20943 ( .B1(n18411), .B2(n17750), .C1(n17749), .C2(n17750), .A(
        n17748), .ZN(n17751) );
  AOI211_X1 U20944 ( .C1(n17752), .C2(n17934), .A(n18092), .B(n17751), .ZN(
        n17757) );
  OAI21_X1 U20945 ( .B1(n17754), .B2(n18089), .A(n17753), .ZN(n18093) );
  AOI22_X1 U20946 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17755), .B1(
        n17874), .B2(n18093), .ZN(n17756) );
  OAI211_X1 U20947 ( .C1(n17771), .C2(n18095), .A(n17757), .B(n17756), .ZN(
        P3_U2813) );
  AOI21_X1 U20948 ( .B1(n17873), .B2(n17759), .A(n17758), .ZN(n17760) );
  XNOR2_X1 U20949 ( .A(n17760), .B(n21097), .ZN(n18102) );
  INV_X1 U20950 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17762) );
  NAND2_X1 U20951 ( .A1(n17763), .A2(n17809), .ZN(n17773) );
  AOI221_X1 U20952 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n17762), .C2(n17761), .A(
        n17773), .ZN(n17768) );
  AOI21_X1 U20953 ( .B1(n17923), .B2(n9915), .A(n17921), .ZN(n17785) );
  OAI21_X1 U20954 ( .B1(n17764), .B2(n17961), .A(n17785), .ZN(n17775) );
  AOI22_X1 U20955 ( .A1(n9768), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17775), .ZN(n17765) );
  OAI21_X1 U20956 ( .B1(n17802), .B2(n17766), .A(n17765), .ZN(n17767) );
  AOI211_X1 U20957 ( .C1(n18102), .C2(n17874), .A(n17768), .B(n17767), .ZN(
        n17769) );
  OAI221_X1 U20958 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17771), 
        .C1(n21097), .C2(n17770), .A(n17769), .ZN(P3_U2814) );
  NOR2_X1 U20959 ( .A1(n18170), .A2(n18126), .ZN(n17790) );
  NOR2_X1 U20960 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17790), .ZN(
        n18108) );
  NOR2_X1 U20961 ( .A1(n18289), .A2(n18860), .ZN(n18117) );
  OAI22_X1 U20962 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17773), .B1(
        n17772), .B2(n17802), .ZN(n17774) );
  AOI211_X1 U20963 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17775), .A(
        n18117), .B(n17774), .ZN(n17782) );
  INV_X1 U20964 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18128) );
  OAI21_X1 U20965 ( .B1(n17777), .B2(n17837), .A(n17776), .ZN(n17778) );
  OAI221_X1 U20966 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18128), 
        .C1(n18160), .C2(n17873), .A(n17778), .ZN(n17779) );
  XNOR2_X1 U20967 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17779), .ZN(
        n18118) );
  NOR2_X1 U20968 ( .A1(n18026), .A2(n17965), .ZN(n17780) );
  NAND2_X1 U20969 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18141), .ZN(
        n18154) );
  NOR2_X1 U20970 ( .A1(n17827), .A2(n18154), .ZN(n18145) );
  NAND3_X1 U20971 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n18145), .ZN(n17784) );
  NAND2_X1 U20972 ( .A1(n18115), .A2(n17784), .ZN(n18119) );
  AOI22_X1 U20973 ( .A1(n17874), .A2(n18118), .B1(n17780), .B2(n18119), .ZN(
        n17781) );
  OAI211_X1 U20974 ( .C1(n18108), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        P3_U2815) );
  OAI221_X1 U20975 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18145), .A(n17784), .ZN(
        n18134) );
  AOI221_X1 U20976 ( .B1(n18411), .B2(n17787), .C1(n17786), .C2(n17787), .A(
        n17785), .ZN(n17788) );
  NOR2_X1 U20977 ( .A1(n18289), .A2(n18859), .ZN(n18133) );
  AOI211_X1 U20978 ( .C1(n17789), .C2(n17934), .A(n17788), .B(n18133), .ZN(
        n17795) );
  NOR2_X1 U20979 ( .A1(n18146), .A2(n18154), .ZN(n17792) );
  INV_X1 U20980 ( .A(n17792), .ZN(n18109) );
  AOI221_X1 U20981 ( .B1(n18170), .B2(n18128), .C1(n18109), .C2(n18128), .A(
        n17790), .ZN(n18132) );
  NOR2_X1 U20982 ( .A1(n17838), .A2(n18170), .ZN(n17835) );
  AOI21_X1 U20983 ( .B1(n17792), .B2(n17835), .A(n17791), .ZN(n17793) );
  XNOR2_X1 U20984 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17793), .ZN(
        n18135) );
  AOI22_X1 U20985 ( .A1(n17828), .A2(n18132), .B1(n17874), .B2(n18135), .ZN(
        n17794) );
  OAI211_X1 U20986 ( .C1(n17965), .C2(n18134), .A(n17795), .B(n17794), .ZN(
        P3_U2816) );
  OAI22_X1 U20987 ( .A1(n17873), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18154), .B2(n17837), .ZN(n17797) );
  OAI21_X1 U20988 ( .B1(n17873), .B2(n17796), .A(n17797), .ZN(n17798) );
  XNOR2_X1 U20989 ( .A(n17798), .B(n18146), .ZN(n18153) );
  AOI21_X1 U20990 ( .B1(n17923), .B2(n17799), .A(n17921), .ZN(n17800) );
  OAI21_X1 U20991 ( .B1(n17801), .B2(n17961), .A(n17800), .ZN(n17813) );
  NOR2_X1 U20992 ( .A1(n18289), .A2(n21048), .ZN(n18150) );
  OAI211_X1 U20993 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17810), .B(n17809), .ZN(n17804) );
  OAI22_X1 U20994 ( .A1(n10217), .A2(n17804), .B1(n17803), .B2(n17802), .ZN(
        n17805) );
  AOI211_X1 U20995 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17813), .A(
        n18150), .B(n17805), .ZN(n17807) );
  NOR2_X1 U20996 ( .A1(n18170), .A2(n18154), .ZN(n18140) );
  OAI22_X1 U20997 ( .A1(n18140), .A2(n17878), .B1(n18145), .B2(n17965), .ZN(
        n17817) );
  NOR2_X1 U20998 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18154), .ZN(
        n18151) );
  AOI22_X1 U20999 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17817), .B1(
        n18151), .B2(n17856), .ZN(n17806) );
  OAI211_X1 U21000 ( .C1(n17853), .C2(n18153), .A(n17807), .B(n17806), .ZN(
        P3_U2817) );
  AOI21_X1 U21001 ( .B1(n17835), .B2(n18141), .A(n17796), .ZN(n17808) );
  XOR2_X1 U21002 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17808), .Z(
        n18165) );
  NAND2_X1 U21003 ( .A1(n17810), .A2(n17809), .ZN(n17815) );
  AOI22_X1 U21004 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17813), .B1(
        n17812), .B2(n17811), .ZN(n17814) );
  NAND2_X1 U21005 ( .A1(n9768), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18163) );
  OAI211_X1 U21006 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17815), .A(
        n17814), .B(n18163), .ZN(n17816) );
  AOI21_X1 U21007 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17817), .A(
        n17816), .ZN(n17819) );
  NAND3_X1 U21008 ( .A1(n18141), .A2(n18160), .A3(n17856), .ZN(n17818) );
  OAI211_X1 U21009 ( .C1(n18165), .C2(n17853), .A(n17819), .B(n17818), .ZN(
        P3_U2818) );
  NAND2_X1 U21010 ( .A1(n18174), .A2(n17835), .ZN(n17840) );
  NAND2_X1 U21011 ( .A1(n17840), .A2(n17820), .ZN(n17821) );
  XNOR2_X1 U21012 ( .A(n17821), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18180) );
  NOR2_X1 U21013 ( .A1(n18411), .A2(n17822), .ZN(n17848) );
  NOR2_X1 U21014 ( .A1(n17825), .A2(n17848), .ZN(n17826) );
  OAI22_X1 U21015 ( .A1(n17958), .A2(n17823), .B1(n18289), .B2(n18853), .ZN(
        n17824) );
  AOI221_X1 U21016 ( .B1(n17954), .B2(n17826), .C1(n17825), .C2(n17848), .A(
        n17824), .ZN(n17831) );
  INV_X1 U21017 ( .A(n17856), .ZN(n17833) );
  AOI22_X1 U21018 ( .A1(n17828), .A2(n18170), .B1(n17950), .B2(n17827), .ZN(
        n17854) );
  OAI21_X1 U21019 ( .B1(n18174), .B2(n17833), .A(n17854), .ZN(n17845) );
  INV_X1 U21020 ( .A(n18174), .ZN(n17829) );
  NOR2_X1 U21021 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17829), .ZN(
        n18166) );
  AOI22_X1 U21022 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17845), .B1(
        n18166), .B2(n17856), .ZN(n17830) );
  OAI211_X1 U21023 ( .C1(n18180), .C2(n17853), .A(n17831), .B(n17830), .ZN(
        P3_U2819) );
  NOR2_X1 U21024 ( .A1(n18411), .A2(n17832), .ZN(n17892) );
  INV_X1 U21025 ( .A(n17892), .ZN(n17895) );
  NOR2_X1 U21026 ( .A1(n17896), .A2(n17895), .ZN(n17884) );
  AND3_X1 U21027 ( .A1(n17861), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17884), .ZN(n17860) );
  AOI21_X1 U21028 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17954), .A(
        n17860), .ZN(n17847) );
  OAI21_X1 U21029 ( .B1(n17833), .B2(n18189), .A(n17836), .ZN(n17844) );
  INV_X1 U21030 ( .A(n17834), .ZN(n17850) );
  INV_X1 U21031 ( .A(n17835), .ZN(n17851) );
  OAI221_X1 U21032 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17850), .C1(
        n18189), .C2(n17851), .A(n17836), .ZN(n17841) );
  NAND4_X1 U21033 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17838), .A3(
        n18189), .A4(n17837), .ZN(n17839) );
  NAND3_X1 U21034 ( .A1(n17841), .A2(n17840), .A3(n17839), .ZN(n18188) );
  OAI22_X1 U21035 ( .A1(n17958), .A2(n17842), .B1(n17853), .B2(n18188), .ZN(
        n17843) );
  AOI21_X1 U21036 ( .B1(n17845), .B2(n17844), .A(n17843), .ZN(n17846) );
  NAND2_X1 U21037 ( .A1(n9768), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18186) );
  OAI211_X1 U21038 ( .C1(n17848), .C2(n17847), .A(n17846), .B(n18186), .ZN(
        P3_U2820) );
  AOI22_X1 U21039 ( .A1(n17861), .A2(n17884), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17954), .ZN(n17859) );
  AOI22_X1 U21040 ( .A1(n9768), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17849), .B2(
        n17934), .ZN(n17858) );
  NAND2_X1 U21041 ( .A1(n17851), .A2(n17850), .ZN(n17852) );
  XNOR2_X1 U21042 ( .A(n17852), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18201) );
  OAI22_X1 U21043 ( .A1(n17854), .A2(n18189), .B1(n18201), .B2(n17853), .ZN(
        n17855) );
  AOI21_X1 U21044 ( .B1(n18189), .B2(n17856), .A(n17855), .ZN(n17857) );
  OAI211_X1 U21045 ( .C1(n17860), .C2(n17859), .A(n17858), .B(n17857), .ZN(
        P3_U2821) );
  AOI211_X1 U21046 ( .C1(n17865), .C2(n17862), .A(n17861), .B(n18411), .ZN(
        n17869) );
  OAI21_X1 U21047 ( .B1(n17864), .B2(n17863), .A(n17960), .ZN(n17882) );
  INV_X1 U21048 ( .A(n17882), .ZN(n17866) );
  OAI22_X1 U21049 ( .A1(n17958), .A2(n17867), .B1(n17866), .B2(n17865), .ZN(
        n17868) );
  AOI211_X1 U21050 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n9768), .A(n17869), .B(
        n17868), .ZN(n17876) );
  AOI21_X1 U21051 ( .B1(n17871), .B2(n18193), .A(n17870), .ZN(n18214) );
  OAI21_X1 U21052 ( .B1(n17873), .B2(n18205), .A(n17872), .ZN(n18212) );
  AOI22_X1 U21053 ( .A1(n17950), .A2(n18214), .B1(n17874), .B2(n18212), .ZN(
        n17875) );
  OAI211_X1 U21054 ( .C1(n17878), .C2(n17877), .A(n17876), .B(n17875), .ZN(
        P3_U2822) );
  NAND2_X1 U21055 ( .A1(n17880), .A2(n17879), .ZN(n17881) );
  XNOR2_X1 U21056 ( .A(n17881), .B(n18222), .ZN(n18229) );
  NOR2_X1 U21057 ( .A1(n18289), .A2(n18845), .ZN(n18219) );
  AOI221_X1 U21058 ( .B1(n17884), .B2(n17883), .C1(n17882), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18219), .ZN(n17889) );
  AOI21_X1 U21059 ( .B1(n17886), .B2(n18222), .A(n17885), .ZN(n18225) );
  AOI22_X1 U21060 ( .A1(n17955), .A2(n18225), .B1(n17887), .B2(n17934), .ZN(
        n17888) );
  OAI211_X1 U21061 ( .C1(n17965), .C2(n18229), .A(n17889), .B(n17888), .ZN(
        P3_U2823) );
  AOI21_X1 U21062 ( .B1(n17891), .B2(n17890), .A(n9890), .ZN(n18234) );
  AOI22_X1 U21063 ( .A1(n17955), .A2(n18234), .B1(n17892), .B2(n17896), .ZN(
        n17900) );
  AOI21_X1 U21064 ( .B1(n18238), .B2(n17894), .A(n17893), .ZN(n18235) );
  NAND2_X1 U21065 ( .A1(n17954), .A2(n17895), .ZN(n17912) );
  OAI22_X1 U21066 ( .A1(n17958), .A2(n17897), .B1(n17896), .B2(n17912), .ZN(
        n17898) );
  AOI21_X1 U21067 ( .B1(n17950), .B2(n18235), .A(n17898), .ZN(n17899) );
  OAI211_X1 U21068 ( .C1(n18289), .C2(n18843), .A(n17900), .B(n17899), .ZN(
        P3_U2824) );
  AOI21_X1 U21069 ( .B1(n17901), .B2(n17960), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17913) );
  OAI21_X1 U21070 ( .B1(n17904), .B2(n17903), .A(n17902), .ZN(n17905) );
  XNOR2_X1 U21071 ( .A(n17905), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18241) );
  AOI22_X1 U21072 ( .A1(n17955), .A2(n18241), .B1(n9768), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17911) );
  AOI21_X1 U21073 ( .B1(n17908), .B2(n17907), .A(n17906), .ZN(n18239) );
  AOI22_X1 U21074 ( .A1(n17950), .A2(n18239), .B1(n17909), .B2(n17934), .ZN(
        n17910) );
  OAI211_X1 U21075 ( .C1(n17913), .C2(n17912), .A(n17911), .B(n17910), .ZN(
        P3_U2825) );
  OAI21_X1 U21076 ( .B1(n17916), .B2(n17915), .A(n17914), .ZN(n17917) );
  XNOR2_X1 U21077 ( .A(n17917), .B(n21099), .ZN(n18247) );
  AOI22_X1 U21078 ( .A1(n9768), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18692), .B2(
        n17918), .ZN(n17928) );
  AOI21_X1 U21079 ( .B1(n9894), .B2(n17920), .A(n17919), .ZN(n18250) );
  AOI21_X1 U21080 ( .B1(n17923), .B2(n17922), .A(n17921), .ZN(n17938) );
  OAI22_X1 U21081 ( .A1(n17958), .A2(n17925), .B1(n17924), .B2(n17938), .ZN(
        n17926) );
  AOI21_X1 U21082 ( .B1(n17955), .B2(n18250), .A(n17926), .ZN(n17927) );
  OAI211_X1 U21083 ( .C1(n17965), .C2(n18247), .A(n17928), .B(n17927), .ZN(
        P3_U2826) );
  AOI21_X1 U21084 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17960), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17939) );
  AOI21_X1 U21085 ( .B1(n18246), .B2(n17930), .A(n17929), .ZN(n18255) );
  AOI22_X1 U21086 ( .A1(n17955), .A2(n18255), .B1(n9768), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17937) );
  AOI21_X1 U21087 ( .B1(n17933), .B2(n17932), .A(n17931), .ZN(n18256) );
  AOI22_X1 U21088 ( .A1(n17950), .A2(n18256), .B1(n17935), .B2(n17934), .ZN(
        n17936) );
  OAI211_X1 U21089 ( .C1(n17939), .C2(n17938), .A(n17937), .B(n17936), .ZN(
        P3_U2827) );
  AOI21_X1 U21090 ( .B1(n17942), .B2(n17941), .A(n17940), .ZN(n18273) );
  NOR2_X1 U21091 ( .A1(n18289), .A2(n18835), .ZN(n18275) );
  XNOR2_X1 U21092 ( .A(n17944), .B(n17943), .ZN(n18272) );
  OAI22_X1 U21093 ( .A1(n17958), .A2(n17945), .B1(n17965), .B2(n18272), .ZN(
        n17946) );
  AOI211_X1 U21094 ( .C1(n17955), .C2(n18273), .A(n18275), .B(n17946), .ZN(
        n17947) );
  OAI221_X1 U21095 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18411), .C1(
        n17948), .C2(n17960), .A(n17947), .ZN(P3_U2828) );
  NOR2_X1 U21096 ( .A1(n17959), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17949) );
  XNOR2_X1 U21097 ( .A(n17953), .B(n17949), .ZN(n18282) );
  AOI22_X1 U21098 ( .A1(n17950), .A2(n18282), .B1(n9768), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17957) );
  AOI21_X1 U21099 ( .B1(n17951), .B2(n17953), .A(n17952), .ZN(n18281) );
  AOI22_X1 U21100 ( .A1(n17955), .A2(n18281), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17954), .ZN(n17956) );
  OAI211_X1 U21101 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17958), .A(
        n17957), .B(n17956), .ZN(P3_U2829) );
  OAI21_X1 U21102 ( .B1(n17959), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17951), .ZN(n18291) );
  INV_X1 U21103 ( .A(n18291), .ZN(n18293) );
  NAND3_X1 U21104 ( .A1(n18921), .A2(n17961), .A3(n17960), .ZN(n17962) );
  AOI22_X1 U21105 ( .A1(n9768), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17962), .ZN(n17963) );
  OAI221_X1 U21106 ( .B1(n18293), .B2(n17965), .C1(n18291), .C2(n17964), .A(
        n17963), .ZN(P3_U2830) );
  NAND2_X1 U21107 ( .A1(n17966), .A2(n18017), .ZN(n17986) );
  NOR2_X1 U21108 ( .A1(n17985), .A2(n17986), .ZN(n17979) );
  NOR2_X1 U21109 ( .A1(n18771), .A2(n18192), .ZN(n18082) );
  INV_X1 U21110 ( .A(n18082), .ZN(n18262) );
  NOR2_X1 U21111 ( .A1(n18769), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18263) );
  AOI21_X1 U21112 ( .B1(n18262), .B2(n17967), .A(n18263), .ZN(n18004) );
  OAI21_X1 U21113 ( .B1(n17969), .B2(n17968), .A(n18268), .ZN(n17970) );
  OAI211_X1 U21114 ( .C1(n18082), .C2(n17971), .A(n18004), .B(n17970), .ZN(
        n17992) );
  NOR2_X1 U21115 ( .A1(n18268), .A2(n18192), .ZN(n18124) );
  OAI22_X1 U21116 ( .A1(n18763), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n17972), .B2(n18124), .ZN(n17973) );
  AOI211_X1 U21117 ( .C1(n18204), .C2(n17974), .A(n17992), .B(n17973), .ZN(
        n17975) );
  OAI21_X1 U21118 ( .B1(n17976), .B2(n18750), .A(n17975), .ZN(n17984) );
  AOI21_X1 U21119 ( .B1(n18771), .B2(n17985), .A(n17984), .ZN(n17977) );
  INV_X1 U21120 ( .A(n17977), .ZN(n17978) );
  MUX2_X1 U21121 ( .A(n17979), .B(n17978), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17980) );
  AOI22_X1 U21122 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18254), .B1(
        n18288), .B2(n17980), .ZN(n17982) );
  OAI211_X1 U21123 ( .C1(n17983), .C2(n18200), .A(n17982), .B(n17981), .ZN(
        P3_U2835) );
  INV_X1 U21124 ( .A(n17984), .ZN(n17987) );
  AOI221_X1 U21125 ( .B1(n17987), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n17986), .C2(n17985), .A(n18217), .ZN(n17988) );
  AOI211_X1 U21126 ( .C1(n18254), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17989), .B(n17988), .ZN(n17990) );
  OAI21_X1 U21127 ( .B1(n17991), .B2(n18200), .A(n17990), .ZN(P3_U2836) );
  AOI22_X1 U21128 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18254), .B1(
        n9768), .B2(P3_REIP_REG_25__SCAN_IN), .ZN(n18001) );
  INV_X1 U21129 ( .A(n17992), .ZN(n17997) );
  AOI22_X1 U21130 ( .A1(n17994), .A2(n18204), .B1(n17993), .B2(n17996), .ZN(
        n17995) );
  OAI21_X1 U21131 ( .B1(n17997), .B2(n17996), .A(n17995), .ZN(n17999) );
  AOI22_X1 U21132 ( .A1(n18288), .A2(n17999), .B1(n18292), .B2(n17998), .ZN(
        n18000) );
  OAI211_X1 U21133 ( .C1(n18200), .C2(n18002), .A(n18001), .B(n18000), .ZN(
        P3_U2837) );
  INV_X1 U21134 ( .A(n18003), .ZN(n18013) );
  OAI21_X1 U21135 ( .B1(n18005), .B2(n18106), .A(n18004), .ZN(n18006) );
  AOI211_X1 U21136 ( .C1(n18028), .C2(n18007), .A(n18254), .B(n18006), .ZN(
        n18011) );
  NAND2_X1 U21137 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18011), .ZN(
        n18008) );
  OAI21_X1 U21138 ( .B1(n18009), .B2(n18008), .A(n18289), .ZN(n18024) );
  AOI211_X1 U21139 ( .C1(n18230), .C2(n18011), .A(n18010), .B(n18024), .ZN(
        n18012) );
  AOI21_X1 U21140 ( .B1(n9895), .B2(n18013), .A(n18012), .ZN(n18015) );
  OAI211_X1 U21141 ( .C1(n18016), .C2(n18042), .A(n18015), .B(n18014), .ZN(
        P3_U2838) );
  INV_X1 U21142 ( .A(n18254), .ZN(n18280) );
  NAND3_X1 U21143 ( .A1(n18018), .A2(n18280), .A3(n18017), .ZN(n18022) );
  AOI21_X1 U21144 ( .B1(n18020), .B2(n9895), .A(n18019), .ZN(n18021) );
  OAI221_X1 U21145 ( .B1(n18024), .B2(n18023), .C1(n18024), .C2(n18022), .A(
        n18021), .ZN(P3_U2839) );
  NAND2_X1 U21146 ( .A1(n18750), .A2(n18106), .ZN(n18080) );
  INV_X1 U21147 ( .A(n18025), .ZN(n18076) );
  INV_X1 U21148 ( .A(n18026), .ZN(n18120) );
  AOI22_X1 U21149 ( .A1(n18028), .A2(n18120), .B1(n18204), .B2(n18027), .ZN(
        n18096) );
  OAI221_X1 U21150 ( .B1(n18781), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n18781), .C2(n18075), .A(n18096), .ZN(n18029) );
  AOI221_X1 U21151 ( .B1(n18076), .B2(n18771), .C1(n18053), .C2(n18771), .A(
        n18029), .ZN(n18054) );
  OAI21_X1 U21152 ( .B1(n18763), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n18054), .ZN(n18030) );
  AOI21_X1 U21153 ( .B1(n18031), .B2(n18080), .A(n18030), .ZN(n18047) );
  AOI211_X1 U21154 ( .C1(n18181), .C2(n18033), .A(n18032), .B(n18041), .ZN(
        n18036) );
  AOI21_X1 U21155 ( .B1(n18288), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n18034), .ZN(n18035) );
  AOI21_X1 U21156 ( .B1(n18047), .B2(n18036), .A(n18035), .ZN(n18037) );
  AOI211_X1 U21157 ( .C1(n18039), .C2(n9895), .A(n18038), .B(n18037), .ZN(
        n18040) );
  OAI21_X1 U21158 ( .B1(n18041), .B2(n18280), .A(n18040), .ZN(P3_U2840) );
  NOR2_X1 U21159 ( .A1(n18043), .A2(n18042), .ZN(n18065) );
  AOI22_X1 U21160 ( .A1(n9895), .A2(n18045), .B1(n18044), .B2(n18065), .ZN(
        n18052) );
  OAI221_X1 U21161 ( .B1(n18769), .B2(n18046), .C1(n18769), .C2(n18100), .A(
        n18288), .ZN(n18057) );
  OAI21_X1 U21162 ( .B1(n18048), .B2(n18124), .A(n18047), .ZN(n18049) );
  OAI211_X1 U21163 ( .C1(n18057), .C2(n18049), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18289), .ZN(n18050) );
  NAND3_X1 U21164 ( .A1(n18052), .A2(n18051), .A3(n18050), .ZN(P3_U2841) );
  INV_X1 U21165 ( .A(n18053), .ZN(n18055) );
  INV_X1 U21166 ( .A(n18080), .ZN(n18173) );
  OAI21_X1 U21167 ( .B1(n18055), .B2(n18173), .A(n18054), .ZN(n18056) );
  OAI21_X1 U21168 ( .B1(n18057), .B2(n18056), .A(n18289), .ZN(n18069) );
  INV_X1 U21169 ( .A(n18124), .ZN(n18279) );
  NAND3_X1 U21170 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18070), .A3(n18279), 
        .ZN(n18059) );
  AOI21_X1 U21171 ( .B1(n18069), .B2(n18059), .A(n18058), .ZN(n18060) );
  AOI211_X1 U21172 ( .C1(n18062), .C2(n18065), .A(n18061), .B(n18060), .ZN(
        n18063) );
  OAI21_X1 U21173 ( .B1(n18200), .B2(n18064), .A(n18063), .ZN(P3_U2842) );
  AOI22_X1 U21174 ( .A1(n9895), .A2(n18066), .B1(n18065), .B2(n18070), .ZN(
        n18068) );
  NAND2_X1 U21175 ( .A1(n9768), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18067) );
  OAI211_X1 U21176 ( .C1(n18070), .C2(n18069), .A(n18068), .B(n18067), .ZN(
        P3_U2843) );
  INV_X1 U21177 ( .A(n18208), .ZN(n18267) );
  INV_X1 U21178 ( .A(n18269), .ZN(n18071) );
  OAI22_X1 U21179 ( .A1(n18267), .A2(n18781), .B1(n18071), .B2(n18206), .ZN(
        n18258) );
  NAND2_X1 U21180 ( .A1(n18072), .A2(n18258), .ZN(n18110) );
  AND2_X1 U21181 ( .A1(n18073), .A2(n18110), .ZN(n18161) );
  NAND2_X1 U21182 ( .A1(n18074), .A2(n18190), .ZN(n18105) );
  NOR2_X1 U21183 ( .A1(n18075), .A2(n18781), .ZN(n18079) );
  NOR3_X1 U21184 ( .A1(n18263), .A2(n18076), .A3(n21097), .ZN(n18077) );
  OAI211_X1 U21185 ( .C1(n18082), .C2(n18077), .A(n18288), .B(n18096), .ZN(
        n18078) );
  AOI211_X1 U21186 ( .C1(n18081), .C2(n18080), .A(n18079), .B(n18078), .ZN(
        n18090) );
  AOI221_X1 U21187 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18090), 
        .C1(n18082), .C2(n18090), .A(n9768), .ZN(n18084) );
  AOI22_X1 U21188 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18084), .B1(
        n9895), .B2(n18083), .ZN(n18087) );
  INV_X1 U21189 ( .A(n18085), .ZN(n18086) );
  OAI211_X1 U21190 ( .C1(n18088), .C2(n18105), .A(n18087), .B(n18086), .ZN(
        P3_U2844) );
  NOR3_X1 U21191 ( .A1(n9768), .A2(n18090), .A3(n18089), .ZN(n18091) );
  AOI211_X1 U21192 ( .C1(n9895), .C2(n18093), .A(n18092), .B(n18091), .ZN(
        n18094) );
  OAI21_X1 U21193 ( .B1(n18105), .B2(n18095), .A(n18094), .ZN(P3_U2845) );
  NAND2_X1 U21194 ( .A1(n18288), .A2(n18096), .ZN(n18101) );
  NAND2_X1 U21195 ( .A1(n18268), .A2(n18097), .ZN(n18167) );
  OAI21_X1 U21196 ( .B1(n18763), .B2(n18098), .A(n18167), .ZN(n18142) );
  AOI21_X1 U21197 ( .B1(n18181), .B2(n18126), .A(n18142), .ZN(n18099) );
  OAI211_X1 U21198 ( .C1(n18100), .C2(n18769), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18099), .ZN(n18112) );
  OAI221_X1 U21199 ( .B1(n18101), .B2(n18209), .C1(n18101), .C2(n18112), .A(
        n18289), .ZN(n18104) );
  AOI22_X1 U21200 ( .A1(n9768), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n9895), .B2(
        n18102), .ZN(n18103) );
  OAI221_X1 U21201 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18105), 
        .C1(n21097), .C2(n18104), .A(n18103), .ZN(P3_U2846) );
  NOR2_X1 U21202 ( .A1(n18107), .A2(n18106), .ZN(n18114) );
  INV_X1 U21203 ( .A(n18108), .ZN(n18113) );
  OR2_X1 U21204 ( .A1(n18110), .A2(n18109), .ZN(n18127) );
  OAI21_X1 U21205 ( .B1(n18128), .B2(n18127), .A(n18115), .ZN(n18111) );
  AOI22_X1 U21206 ( .A1(n18114), .A2(n18113), .B1(n18112), .B2(n18111), .ZN(
        n18123) );
  NOR2_X1 U21207 ( .A1(n18115), .A2(n18280), .ZN(n18116) );
  AOI211_X1 U21208 ( .C1(n18118), .C2(n9895), .A(n18117), .B(n18116), .ZN(
        n18122) );
  NAND3_X1 U21209 ( .A1(n18292), .A2(n18120), .A3(n18119), .ZN(n18121) );
  OAI211_X1 U21210 ( .C1(n18123), .C2(n18217), .A(n18122), .B(n18121), .ZN(
        P3_U2847) );
  OAI21_X1 U21211 ( .B1(n18191), .B2(n18154), .A(n18192), .ZN(n18147) );
  AOI21_X1 U21212 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18147), .A(
        n18124), .ZN(n18125) );
  AOI211_X1 U21213 ( .C1(n18268), .C2(n18154), .A(n18125), .B(n18142), .ZN(
        n18130) );
  OAI21_X1 U21214 ( .B1(n18128), .B2(n18771), .A(n18126), .ZN(n18129) );
  AOI22_X1 U21215 ( .A1(n18130), .A2(n18129), .B1(n18128), .B2(n18127), .ZN(
        n18131) );
  AOI21_X1 U21216 ( .B1(n18132), .B2(n18204), .A(n18131), .ZN(n18139) );
  AOI21_X1 U21217 ( .B1(n18254), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18133), .ZN(n18138) );
  INV_X1 U21218 ( .A(n18134), .ZN(n18136) );
  AOI22_X1 U21219 ( .A1(n18292), .A2(n18136), .B1(n9895), .B2(n18135), .ZN(
        n18137) );
  OAI211_X1 U21220 ( .C1(n18139), .C2(n18217), .A(n18138), .B(n18137), .ZN(
        P3_U2848) );
  OAI21_X1 U21221 ( .B1(n18763), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18155) );
  INV_X1 U21222 ( .A(n18140), .ZN(n18143) );
  OAI22_X1 U21223 ( .A1(n18763), .A2(n18174), .B1(n18141), .B2(n18781), .ZN(
        n18177) );
  AOI211_X1 U21224 ( .C1(n18204), .C2(n18143), .A(n18142), .B(n18177), .ZN(
        n18144) );
  OAI21_X1 U21225 ( .B1(n18145), .B2(n18750), .A(n18144), .ZN(n18156) );
  AOI211_X1 U21226 ( .C1(n18181), .C2(n18155), .A(n18217), .B(n18156), .ZN(
        n18148) );
  AOI211_X1 U21227 ( .C1(n18148), .C2(n18147), .A(n9768), .B(n18146), .ZN(
        n18149) );
  AOI211_X1 U21228 ( .C1(n18151), .C2(n18190), .A(n18150), .B(n18149), .ZN(
        n18152) );
  OAI21_X1 U21229 ( .B1(n18200), .B2(n18153), .A(n18152), .ZN(P3_U2849) );
  OR2_X1 U21230 ( .A1(n18191), .A2(n18154), .ZN(n18157) );
  AOI211_X1 U21231 ( .C1(n18157), .C2(n18192), .A(n18156), .B(n18155), .ZN(
        n18158) );
  AOI221_X1 U21232 ( .B1(n18161), .B2(n18160), .C1(n18159), .C2(n18160), .A(
        n18158), .ZN(n18162) );
  AOI22_X1 U21233 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18254), .B1(
        n18288), .B2(n18162), .ZN(n18164) );
  OAI211_X1 U21234 ( .C1(n18165), .C2(n18200), .A(n18164), .B(n18163), .ZN(
        P3_U2850) );
  AOI22_X1 U21235 ( .A1(n9768), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18190), 
        .B2(n18166), .ZN(n18179) );
  OAI211_X1 U21236 ( .C1(n18168), .C2(n18750), .A(n18288), .B(n18167), .ZN(
        n18169) );
  AOI21_X1 U21237 ( .B1(n18204), .B2(n18170), .A(n18169), .ZN(n18195) );
  NAND2_X1 U21238 ( .A1(n18771), .A2(n18171), .ZN(n18172) );
  OAI211_X1 U21239 ( .C1(n18174), .C2(n18173), .A(n18195), .B(n18172), .ZN(
        n18175) );
  AOI221_X1 U21240 ( .B1(n18189), .B2(n18192), .C1(n18191), .C2(n18192), .A(
        n18175), .ZN(n18182) );
  OAI21_X1 U21241 ( .B1(n18769), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18182), .ZN(n18176) );
  OAI211_X1 U21242 ( .C1(n18177), .C2(n18176), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18289), .ZN(n18178) );
  OAI211_X1 U21243 ( .C1(n18180), .C2(n18200), .A(n18179), .B(n18178), .ZN(
        P3_U2851) );
  INV_X1 U21244 ( .A(n18181), .ZN(n18183) );
  AOI221_X1 U21245 ( .B1(n18183), .B2(n18182), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18182), .A(n9768), .ZN(n18185) );
  NOR2_X1 U21246 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18189), .ZN(
        n18184) );
  AOI22_X1 U21247 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18185), .B1(
        n18190), .B2(n18184), .ZN(n18187) );
  OAI211_X1 U21248 ( .C1(n18200), .C2(n18188), .A(n18187), .B(n18186), .ZN(
        P3_U2852) );
  AOI22_X1 U21249 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n9768), .B1(n18190), .B2(
        n18189), .ZN(n18199) );
  OAI211_X1 U21250 ( .C1(n18193), .C2(n18192), .A(n18262), .B(n18191), .ZN(
        n18194) );
  OAI211_X1 U21251 ( .C1(n18763), .C2(n18196), .A(n18195), .B(n18194), .ZN(
        n18197) );
  NAND3_X1 U21252 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18289), .A3(
        n18197), .ZN(n18198) );
  OAI211_X1 U21253 ( .C1(n18201), .C2(n18200), .A(n18199), .B(n18198), .ZN(
        P3_U2853) );
  NOR2_X1 U21254 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18202), .ZN(
        n18203) );
  AOI22_X1 U21255 ( .A1(n18205), .A2(n18204), .B1(n18203), .B2(n18258), .ZN(
        n18218) );
  OAI21_X1 U21256 ( .B1(n18263), .B2(n18206), .A(n18262), .ZN(n18207) );
  OAI21_X1 U21257 ( .B1(n18208), .B2(n18781), .A(n18207), .ZN(n18245) );
  AOI211_X1 U21258 ( .C1(n18209), .C2(n18221), .A(n18222), .B(n18245), .ZN(
        n18220) );
  OAI21_X1 U21259 ( .B1(n18220), .B2(n18210), .A(n18280), .ZN(n18211) );
  AOI22_X1 U21260 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18211), .B1(
        n9768), .B2(P3_REIP_REG_8__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U21261 ( .A1(n18292), .A2(n18214), .B1(n9895), .B2(n18212), .ZN(
        n18215) );
  OAI211_X1 U21262 ( .C1(n18218), .C2(n18217), .A(n18216), .B(n18215), .ZN(
        P3_U2854) );
  INV_X1 U21263 ( .A(n18292), .ZN(n18248) );
  AOI21_X1 U21264 ( .B1(n18254), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18219), .ZN(n18228) );
  INV_X1 U21265 ( .A(n18258), .ZN(n18223) );
  AOI221_X1 U21266 ( .B1(n18223), .B2(n18222), .C1(n18221), .C2(n18222), .A(
        n18220), .ZN(n18226) );
  AOI22_X1 U21267 ( .A1(n18288), .A2(n18226), .B1(n18294), .B2(n18225), .ZN(
        n18227) );
  OAI211_X1 U21268 ( .C1(n18248), .C2(n18229), .A(n18228), .B(n18227), .ZN(
        P3_U2855) );
  OAI21_X1 U21269 ( .B1(n18230), .B2(n18232), .A(n18288), .ZN(n18231) );
  OAI21_X1 U21270 ( .B1(n18245), .B2(n18231), .A(n18289), .ZN(n18244) );
  AND4_X1 U21271 ( .A1(n18238), .A2(n18258), .A3(n18288), .A4(n18232), .ZN(
        n18233) );
  AOI21_X1 U21272 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n9768), .A(n18233), .ZN(
        n18237) );
  AOI22_X1 U21273 ( .A1(n18292), .A2(n18235), .B1(n18294), .B2(n18234), .ZN(
        n18236) );
  OAI211_X1 U21274 ( .C1(n18238), .C2(n18244), .A(n18237), .B(n18236), .ZN(
        P3_U2856) );
  AOI22_X1 U21275 ( .A1(n9768), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18292), .B2(
        n18239), .ZN(n18243) );
  NAND3_X1 U21276 ( .A1(n18288), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18258), .ZN(n18253) );
  NOR3_X1 U21277 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21099), .A3(
        n18253), .ZN(n18240) );
  AOI21_X1 U21278 ( .B1(n18241), .B2(n18294), .A(n18240), .ZN(n18242) );
  OAI211_X1 U21279 ( .C1(n10115), .C2(n18244), .A(n18243), .B(n18242), .ZN(
        P3_U2857) );
  OR2_X1 U21280 ( .A1(n18246), .A2(n18245), .ZN(n18257) );
  AOI21_X1 U21281 ( .B1(n18283), .B2(n18257), .A(n18254), .ZN(n18252) );
  INV_X1 U21282 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18839) );
  OAI22_X1 U21283 ( .A1(n18289), .A2(n18839), .B1(n18248), .B2(n18247), .ZN(
        n18249) );
  AOI21_X1 U21284 ( .B1(n18294), .B2(n18250), .A(n18249), .ZN(n18251) );
  OAI221_X1 U21285 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18253), .C1(
        n21099), .C2(n18252), .A(n18251), .ZN(P3_U2858) );
  AOI22_X1 U21286 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18254), .B1(
        n9768), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U21287 ( .A1(n18292), .A2(n18256), .B1(n18294), .B2(n18255), .ZN(
        n18260) );
  OAI211_X1 U21288 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18258), .A(
        n18288), .B(n18257), .ZN(n18259) );
  NAND3_X1 U21289 ( .A1(n18261), .A2(n18260), .A3(n18259), .ZN(P3_U2859) );
  NAND2_X1 U21290 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18265) );
  OAI21_X1 U21291 ( .B1(n18263), .B2(n18923), .A(n18262), .ZN(n18264) );
  OAI21_X1 U21292 ( .B1(n18265), .B2(n18781), .A(n18264), .ZN(n18266) );
  AOI22_X1 U21293 ( .A1(n18268), .A2(n18267), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18266), .ZN(n18271) );
  NAND3_X1 U21294 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18269), .A3(
        n18278), .ZN(n18270) );
  OAI211_X1 U21295 ( .C1(n18272), .C2(n18750), .A(n18271), .B(n18270), .ZN(
        n18274) );
  AOI22_X1 U21296 ( .A1(n18288), .A2(n18274), .B1(n18294), .B2(n18273), .ZN(
        n18277) );
  INV_X1 U21297 ( .A(n18275), .ZN(n18276) );
  OAI211_X1 U21298 ( .C1(n18280), .C2(n18278), .A(n18277), .B(n18276), .ZN(
        P3_U2860) );
  NAND3_X1 U21299 ( .A1(n18288), .A2(n18938), .A3(n18279), .ZN(n18296) );
  NAND2_X1 U21300 ( .A1(n18280), .A2(n18296), .ZN(n18287) );
  AOI22_X1 U21301 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18287), .B1(
        n9768), .B2(P3_REIP_REG_1__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U21302 ( .A1(n18292), .A2(n18282), .B1(n18294), .B2(n18281), .ZN(
        n18285) );
  OAI211_X1 U21303 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18771), .A(
        n18283), .B(n18923), .ZN(n18284) );
  NAND3_X1 U21304 ( .A1(n18286), .A2(n18285), .A3(n18284), .ZN(P3_U2861) );
  AOI21_X1 U21305 ( .B1(n18288), .B2(n18771), .A(n18287), .ZN(n18297) );
  NOR2_X1 U21306 ( .A1(n18289), .A2(n18948), .ZN(n18290) );
  AOI221_X1 U21307 ( .B1(n18294), .B2(n18293), .C1(n18292), .C2(n18291), .A(
        n18290), .ZN(n18295) );
  OAI211_X1 U21308 ( .C1(n18297), .C2(n18938), .A(n18296), .B(n18295), .ZN(
        P3_U2862) );
  INV_X1 U21309 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18787) );
  NOR2_X1 U21310 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18787), .ZN(
        n18600) );
  NOR2_X1 U21311 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18298), .ZN(
        n18479) );
  NOR2_X1 U21312 ( .A1(n18600), .A2(n18479), .ZN(n18300) );
  OAI22_X1 U21313 ( .A1(n18301), .A2(n18787), .B1(n18300), .B2(n18299), .ZN(
        P3_U2866) );
  NOR2_X1 U21314 ( .A1(n21096), .A2(n20995), .ZN(P3_U2867) );
  NAND2_X1 U21315 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18305) );
  NAND2_X1 U21316 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20991), .ZN(
        n18553) );
  NAND2_X1 U21317 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18579), .ZN(
        n18532) );
  AND2_X1 U21318 ( .A1(n18553), .A2(n18532), .ZN(n18603) );
  OR2_X1 U21319 ( .A1(n18305), .A2(n18603), .ZN(n18657) );
  NOR2_X1 U21320 ( .A1(n18579), .A2(n20991), .ZN(n18772) );
  INV_X1 U21321 ( .A(n18772), .ZN(n18481) );
  NOR2_X2 U21322 ( .A1(n18481), .A2(n18305), .ZN(n18739) );
  NOR2_X1 U21323 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18773) );
  NOR2_X1 U21324 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18389) );
  NAND2_X1 U21325 ( .A1(n18773), .A2(n18389), .ZN(n18409) );
  INV_X1 U21326 ( .A(n18409), .ZN(n18402) );
  NOR2_X1 U21327 ( .A1(n18739), .A2(n18402), .ZN(n18367) );
  INV_X1 U21328 ( .A(n18367), .ZN(n18302) );
  OAI211_X1 U21329 ( .C1(n18910), .C2(n20991), .A(n18661), .B(n18302), .ZN(
        n18303) );
  OAI21_X1 U21330 ( .B1(n18657), .B2(n18411), .A(n18303), .ZN(n18346) );
  NAND2_X1 U21331 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18692), .ZN(n18696) );
  INV_X1 U21332 ( .A(n18696), .ZN(n18632) );
  NOR2_X1 U21333 ( .A1(n18305), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18691) );
  NAND2_X1 U21334 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18691), .ZN(
        n18734) );
  INV_X1 U21335 ( .A(n18734), .ZN(n18738) );
  NOR2_X2 U21336 ( .A1(n18410), .A2(n18304), .ZN(n18687) );
  INV_X1 U21337 ( .A(n18806), .ZN(n18658) );
  NOR2_X1 U21338 ( .A1(n18658), .A2(n18367), .ZN(n18341) );
  AOI22_X1 U21339 ( .A1(n18632), .A2(n18738), .B1(n18687), .B2(n18341), .ZN(
        n18309) );
  NOR2_X1 U21340 ( .A1(n18305), .A2(n18553), .ZN(n18673) );
  NAND2_X1 U21341 ( .A1(n18692), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18636) );
  INV_X1 U21342 ( .A(n18636), .ZN(n18688) );
  OR3_X1 U21343 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18306), .A3(n18910), 
        .ZN(n18342) );
  NOR2_X2 U21344 ( .A1(n18307), .A2(n18342), .ZN(n18693) );
  AOI22_X1 U21345 ( .A1(n18673), .A2(n18688), .B1(n18693), .B2(n18402), .ZN(
        n18308) );
  OAI211_X1 U21346 ( .C1(n18310), .C2(n18346), .A(n18309), .B(n18308), .ZN(
        P3_U2868) );
  CLKBUF_X1 U21347 ( .A(n18673), .Z(n18682) );
  NAND2_X1 U21348 ( .A1(n18692), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18702) );
  INV_X1 U21349 ( .A(n18702), .ZN(n18637) );
  NOR2_X2 U21350 ( .A1(n18410), .A2(n21207), .ZN(n18697) );
  AOI22_X1 U21351 ( .A1(n18682), .A2(n18637), .B1(n18697), .B2(n18341), .ZN(
        n18312) );
  NAND2_X1 U21352 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18692), .ZN(n18640) );
  INV_X1 U21353 ( .A(n18640), .ZN(n18698) );
  NOR2_X2 U21354 ( .A1(n18961), .A2(n18342), .ZN(n18699) );
  AOI22_X1 U21355 ( .A1(n18738), .A2(n18698), .B1(n18699), .B2(n18402), .ZN(
        n18311) );
  OAI211_X1 U21356 ( .C1(n18313), .C2(n18346), .A(n18312), .B(n18311), .ZN(
        P3_U2869) );
  NAND2_X1 U21357 ( .A1(n18692), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18708) );
  INV_X1 U21358 ( .A(n18708), .ZN(n18667) );
  NOR2_X2 U21359 ( .A1(n18410), .A2(n18314), .ZN(n18703) );
  AOI22_X1 U21360 ( .A1(n18682), .A2(n18667), .B1(n18703), .B2(n18341), .ZN(
        n18317) );
  NAND2_X1 U21361 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18692), .ZN(n18670) );
  INV_X1 U21362 ( .A(n18670), .ZN(n18704) );
  NOR2_X2 U21363 ( .A1(n18315), .A2(n18342), .ZN(n18705) );
  AOI22_X1 U21364 ( .A1(n18738), .A2(n18704), .B1(n18705), .B2(n18402), .ZN(
        n18316) );
  OAI211_X1 U21365 ( .C1(n18318), .C2(n18346), .A(n18317), .B(n18316), .ZN(
        P3_U2870) );
  NOR2_X2 U21366 ( .A1(n18410), .A2(n18320), .ZN(n18709) );
  AOI22_X1 U21367 ( .A1(n18673), .A2(n18710), .B1(n18709), .B2(n18341), .ZN(
        n18323) );
  NAND2_X1 U21368 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18692), .ZN(n18714) );
  INV_X1 U21369 ( .A(n18714), .ZN(n18511) );
  NOR2_X2 U21370 ( .A1(n18321), .A2(n18342), .ZN(n18711) );
  AOI22_X1 U21371 ( .A1(n18738), .A2(n18511), .B1(n18711), .B2(n18402), .ZN(
        n18322) );
  OAI211_X1 U21372 ( .C1(n18324), .C2(n18346), .A(n18323), .B(n18322), .ZN(
        P3_U2871) );
  NAND2_X1 U21373 ( .A1(n18692), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18720) );
  INV_X1 U21374 ( .A(n18720), .ZN(n18613) );
  NOR2_X2 U21375 ( .A1(n18410), .A2(n18325), .ZN(n18715) );
  AOI22_X1 U21376 ( .A1(n18673), .A2(n18613), .B1(n18715), .B2(n18341), .ZN(
        n18328) );
  NAND2_X1 U21377 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18692), .ZN(n18616) );
  INV_X1 U21378 ( .A(n18616), .ZN(n18716) );
  NOR2_X2 U21379 ( .A1(n18326), .A2(n18342), .ZN(n18717) );
  AOI22_X1 U21380 ( .A1(n18738), .A2(n18716), .B1(n18717), .B2(n18402), .ZN(
        n18327) );
  OAI211_X1 U21381 ( .C1(n18329), .C2(n18346), .A(n18328), .B(n18327), .ZN(
        P3_U2872) );
  NAND2_X1 U21382 ( .A1(n18692), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18726) );
  INV_X1 U21383 ( .A(n18726), .ZN(n18566) );
  NOR2_X2 U21384 ( .A1(n18410), .A2(n18330), .ZN(n18721) );
  AOI22_X1 U21385 ( .A1(n18682), .A2(n18566), .B1(n18721), .B2(n18341), .ZN(
        n18333) );
  NAND2_X1 U21386 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18692), .ZN(n18570) );
  INV_X1 U21387 ( .A(n18570), .ZN(n18722) );
  NOR2_X2 U21388 ( .A1(n18331), .A2(n18342), .ZN(n18723) );
  AOI22_X1 U21389 ( .A1(n18738), .A2(n18722), .B1(n18723), .B2(n18402), .ZN(
        n18332) );
  OAI211_X1 U21390 ( .C1(n18334), .C2(n18346), .A(n18333), .B(n18332), .ZN(
        P3_U2873) );
  NAND2_X1 U21391 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18692), .ZN(n18623) );
  INV_X1 U21392 ( .A(n18623), .ZN(n18728) );
  NOR2_X2 U21393 ( .A1(n18410), .A2(n18335), .ZN(n18727) );
  AOI22_X1 U21394 ( .A1(n18738), .A2(n18728), .B1(n18727), .B2(n18341), .ZN(
        n18338) );
  NAND2_X1 U21395 ( .A1(n18692), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18733) );
  INV_X1 U21396 ( .A(n18733), .ZN(n18619) );
  NOR2_X2 U21397 ( .A1(n18336), .A2(n18342), .ZN(n18730) );
  AOI22_X1 U21398 ( .A1(n18682), .A2(n18619), .B1(n18730), .B2(n18402), .ZN(
        n18337) );
  OAI211_X1 U21399 ( .C1(n21018), .C2(n18346), .A(n18338), .B(n18337), .ZN(
        P3_U2874) );
  NOR2_X1 U21400 ( .A1(n18339), .A2(n18411), .ZN(n18737) );
  NOR2_X2 U21401 ( .A1(n18340), .A2(n18410), .ZN(n18736) );
  AOI22_X1 U21402 ( .A1(n18673), .A2(n18737), .B1(n18736), .B2(n18341), .ZN(
        n18345) );
  NAND2_X1 U21403 ( .A1(n18692), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18744) );
  INV_X1 U21404 ( .A(n18744), .ZN(n18626) );
  NOR2_X2 U21405 ( .A1(n18343), .A2(n18342), .ZN(n18740) );
  AOI22_X1 U21406 ( .A1(n18738), .A2(n18626), .B1(n18740), .B2(n18402), .ZN(
        n18344) );
  OAI211_X1 U21407 ( .C1(n18347), .C2(n18346), .A(n18345), .B(n18344), .ZN(
        P3_U2875) );
  INV_X1 U21408 ( .A(n18673), .ZN(n18360) );
  INV_X1 U21409 ( .A(n18389), .ZN(n18388) );
  NAND2_X1 U21410 ( .A1(n18579), .A2(n18806), .ZN(n18527) );
  NOR2_X1 U21411 ( .A1(n18388), .A2(n18527), .ZN(n18363) );
  AOI22_X1 U21412 ( .A1(n18688), .A2(n18739), .B1(n18687), .B2(n18363), .ZN(
        n18349) );
  NOR2_X1 U21413 ( .A1(n18787), .A2(n18528), .ZN(n18689) );
  NAND2_X1 U21414 ( .A1(n18661), .A2(n20989), .ZN(n18529) );
  NOR2_X1 U21415 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18529), .ZN(
        n18434) );
  AOI22_X1 U21416 ( .A1(n18692), .A2(n18689), .B1(n18389), .B2(n18434), .ZN(
        n18364) );
  NOR2_X2 U21417 ( .A1(n18532), .A2(n18388), .ZN(n18430) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18364), .B1(
        n18693), .B2(n18430), .ZN(n18348) );
  OAI211_X1 U21419 ( .C1(n18696), .C2(n18360), .A(n18349), .B(n18348), .ZN(
        P3_U2876) );
  INV_X1 U21420 ( .A(n18739), .ZN(n18381) );
  AOI22_X1 U21421 ( .A1(n18673), .A2(n18698), .B1(n18697), .B2(n18363), .ZN(
        n18351) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18364), .B1(
        n18699), .B2(n18430), .ZN(n18350) );
  OAI211_X1 U21423 ( .C1(n18702), .C2(n18381), .A(n18351), .B(n18350), .ZN(
        P3_U2877) );
  AOI22_X1 U21424 ( .A1(n18703), .A2(n18363), .B1(n18667), .B2(n18739), .ZN(
        n18353) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18364), .B1(
        n18705), .B2(n18430), .ZN(n18352) );
  OAI211_X1 U21426 ( .C1(n18360), .C2(n18670), .A(n18353), .B(n18352), .ZN(
        P3_U2878) );
  INV_X1 U21427 ( .A(n18710), .ZN(n18514) );
  AOI22_X1 U21428 ( .A1(n18682), .A2(n18511), .B1(n18709), .B2(n18363), .ZN(
        n18355) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18364), .B1(
        n18711), .B2(n18430), .ZN(n18354) );
  OAI211_X1 U21430 ( .C1(n18514), .C2(n18381), .A(n18355), .B(n18354), .ZN(
        P3_U2879) );
  AOI22_X1 U21431 ( .A1(n18613), .A2(n18739), .B1(n18715), .B2(n18363), .ZN(
        n18357) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18364), .B1(
        n18717), .B2(n18430), .ZN(n18356) );
  OAI211_X1 U21433 ( .C1(n18360), .C2(n18616), .A(n18357), .B(n18356), .ZN(
        P3_U2880) );
  AOI22_X1 U21434 ( .A1(n18566), .A2(n18739), .B1(n18721), .B2(n18363), .ZN(
        n18359) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18364), .B1(
        n18723), .B2(n18430), .ZN(n18358) );
  OAI211_X1 U21436 ( .C1(n18360), .C2(n18570), .A(n18359), .B(n18358), .ZN(
        P3_U2881) );
  AOI22_X1 U21437 ( .A1(n18682), .A2(n18728), .B1(n18727), .B2(n18363), .ZN(
        n18362) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18364), .B1(
        n18730), .B2(n18430), .ZN(n18361) );
  OAI211_X1 U21439 ( .C1(n18733), .C2(n18381), .A(n18362), .B(n18361), .ZN(
        P3_U2882) );
  INV_X1 U21440 ( .A(n18737), .ZN(n18630) );
  AOI22_X1 U21441 ( .A1(n18673), .A2(n18626), .B1(n18736), .B2(n18363), .ZN(
        n18366) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18364), .B1(
        n18740), .B2(n18430), .ZN(n18365) );
  OAI211_X1 U21443 ( .C1(n18630), .C2(n18381), .A(n18366), .B(n18365), .ZN(
        P3_U2883) );
  INV_X1 U21444 ( .A(n18430), .ZN(n18428) );
  NOR2_X2 U21445 ( .A1(n18553), .A2(n18388), .ZN(n18452) );
  INV_X1 U21446 ( .A(n18452), .ZN(n18450) );
  AOI21_X1 U21447 ( .B1(n18428), .B2(n18450), .A(n18658), .ZN(n18384) );
  AOI22_X1 U21448 ( .A1(n18632), .A2(n18739), .B1(n18687), .B2(n18384), .ZN(
        n18370) );
  AOI221_X1 U21449 ( .B1(n18367), .B2(n18428), .C1(n18659), .C2(n18428), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18368) );
  OAI21_X1 U21450 ( .B1(n18452), .B2(n18368), .A(n18661), .ZN(n18385) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18385), .B1(
        n18693), .B2(n18452), .ZN(n18369) );
  OAI211_X1 U21452 ( .C1(n18636), .C2(n18409), .A(n18370), .B(n18369), .ZN(
        P3_U2884) );
  AOI22_X1 U21453 ( .A1(n18697), .A2(n18384), .B1(n18698), .B2(n18739), .ZN(
        n18372) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18385), .B1(
        n18699), .B2(n18452), .ZN(n18371) );
  OAI211_X1 U21455 ( .C1(n18702), .C2(n18409), .A(n18372), .B(n18371), .ZN(
        P3_U2885) );
  AOI22_X1 U21456 ( .A1(n18704), .A2(n18739), .B1(n18703), .B2(n18384), .ZN(
        n18374) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18385), .B1(
        n18705), .B2(n18452), .ZN(n18373) );
  OAI211_X1 U21458 ( .C1(n18708), .C2(n18409), .A(n18374), .B(n18373), .ZN(
        P3_U2886) );
  AOI22_X1 U21459 ( .A1(n18709), .A2(n18384), .B1(n18710), .B2(n18402), .ZN(
        n18376) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18385), .B1(
        n18711), .B2(n18452), .ZN(n18375) );
  OAI211_X1 U21461 ( .C1(n18714), .C2(n18381), .A(n18376), .B(n18375), .ZN(
        P3_U2887) );
  AOI22_X1 U21462 ( .A1(n18715), .A2(n18384), .B1(n18716), .B2(n18739), .ZN(
        n18378) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18385), .B1(
        n18717), .B2(n18452), .ZN(n18377) );
  OAI211_X1 U21464 ( .C1(n18720), .C2(n18409), .A(n18378), .B(n18377), .ZN(
        P3_U2888) );
  AOI22_X1 U21465 ( .A1(n18566), .A2(n18402), .B1(n18721), .B2(n18384), .ZN(
        n18380) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18385), .B1(
        n18723), .B2(n18452), .ZN(n18379) );
  OAI211_X1 U21467 ( .C1(n18570), .C2(n18381), .A(n18380), .B(n18379), .ZN(
        P3_U2889) );
  AOI22_X1 U21468 ( .A1(n18727), .A2(n18384), .B1(n18728), .B2(n18739), .ZN(
        n18383) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18385), .B1(
        n18730), .B2(n18452), .ZN(n18382) );
  OAI211_X1 U21470 ( .C1(n18733), .C2(n18409), .A(n18383), .B(n18382), .ZN(
        P3_U2890) );
  AOI22_X1 U21471 ( .A1(n18626), .A2(n18739), .B1(n18736), .B2(n18384), .ZN(
        n18387) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18385), .B1(
        n18740), .B2(n18452), .ZN(n18386) );
  OAI211_X1 U21473 ( .C1(n18630), .C2(n18409), .A(n18387), .B(n18386), .ZN(
        P3_U2891) );
  NOR2_X1 U21474 ( .A1(n18579), .A2(n18388), .ZN(n18435) );
  AND2_X1 U21475 ( .A1(n18806), .A2(n18435), .ZN(n18405) );
  AOI22_X1 U21476 ( .A1(n18632), .A2(n18402), .B1(n18687), .B2(n18405), .ZN(
        n18391) );
  AOI21_X1 U21477 ( .B1(n18579), .B2(n18659), .A(n18529), .ZN(n18478) );
  NAND2_X1 U21478 ( .A1(n18389), .A2(n18478), .ZN(n18406) );
  NAND2_X1 U21479 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18435), .ZN(
        n18477) );
  INV_X1 U21480 ( .A(n18477), .ZN(n18470) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18406), .B1(
        n18693), .B2(n18470), .ZN(n18390) );
  OAI211_X1 U21482 ( .C1(n18636), .C2(n18428), .A(n18391), .B(n18390), .ZN(
        P3_U2892) );
  AOI22_X1 U21483 ( .A1(n18637), .A2(n18430), .B1(n18697), .B2(n18405), .ZN(
        n18393) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18406), .B1(
        n18699), .B2(n18470), .ZN(n18392) );
  OAI211_X1 U21485 ( .C1(n18640), .C2(n18409), .A(n18393), .B(n18392), .ZN(
        P3_U2893) );
  AOI22_X1 U21486 ( .A1(n18703), .A2(n18405), .B1(n18667), .B2(n18430), .ZN(
        n18395) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18406), .B1(
        n18705), .B2(n18470), .ZN(n18394) );
  OAI211_X1 U21488 ( .C1(n18670), .C2(n18409), .A(n18395), .B(n18394), .ZN(
        P3_U2894) );
  AOI22_X1 U21489 ( .A1(n18709), .A2(n18405), .B1(n18710), .B2(n18430), .ZN(
        n18397) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18406), .B1(
        n18711), .B2(n18470), .ZN(n18396) );
  OAI211_X1 U21491 ( .C1(n18714), .C2(n18409), .A(n18397), .B(n18396), .ZN(
        P3_U2895) );
  AOI22_X1 U21492 ( .A1(n18613), .A2(n18430), .B1(n18715), .B2(n18405), .ZN(
        n18399) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18406), .B1(
        n18717), .B2(n18470), .ZN(n18398) );
  OAI211_X1 U21494 ( .C1(n18616), .C2(n18409), .A(n18399), .B(n18398), .ZN(
        P3_U2896) );
  AOI22_X1 U21495 ( .A1(n18566), .A2(n18430), .B1(n18721), .B2(n18405), .ZN(
        n18401) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18406), .B1(
        n18723), .B2(n18470), .ZN(n18400) );
  OAI211_X1 U21497 ( .C1(n18570), .C2(n18409), .A(n18401), .B(n18400), .ZN(
        P3_U2897) );
  AOI22_X1 U21498 ( .A1(n18727), .A2(n18405), .B1(n18728), .B2(n18402), .ZN(
        n18404) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18406), .B1(
        n18730), .B2(n18470), .ZN(n18403) );
  OAI211_X1 U21500 ( .C1(n18733), .C2(n18428), .A(n18404), .B(n18403), .ZN(
        P3_U2898) );
  AOI22_X1 U21501 ( .A1(n18737), .A2(n18430), .B1(n18736), .B2(n18405), .ZN(
        n18408) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18406), .B1(
        n18740), .B2(n18470), .ZN(n18407) );
  OAI211_X1 U21503 ( .C1(n18744), .C2(n18409), .A(n18408), .B(n18407), .ZN(
        P3_U2899) );
  INV_X1 U21504 ( .A(n18773), .ZN(n18502) );
  INV_X1 U21505 ( .A(n18479), .ZN(n18480) );
  NOR2_X2 U21506 ( .A1(n18502), .A2(n18480), .ZN(n18492) );
  NOR2_X1 U21507 ( .A1(n18470), .A2(n18492), .ZN(n18456) );
  NOR2_X1 U21508 ( .A1(n18658), .A2(n18456), .ZN(n18429) );
  AOI22_X1 U21509 ( .A1(n18632), .A2(n18430), .B1(n18687), .B2(n18429), .ZN(
        n18415) );
  NOR2_X1 U21510 ( .A1(n18430), .A2(n18452), .ZN(n18412) );
  OAI22_X1 U21511 ( .A1(n18412), .A2(n18411), .B1(n18456), .B2(n18410), .ZN(
        n18413) );
  OAI21_X1 U21512 ( .B1(n18492), .B2(n18910), .A(n18413), .ZN(n18431) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18431), .B1(
        n18693), .B2(n18492), .ZN(n18414) );
  OAI211_X1 U21514 ( .C1(n18636), .C2(n18450), .A(n18415), .B(n18414), .ZN(
        P3_U2900) );
  AOI22_X1 U21515 ( .A1(n18697), .A2(n18429), .B1(n18698), .B2(n18430), .ZN(
        n18417) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18431), .B1(
        n18699), .B2(n18492), .ZN(n18416) );
  OAI211_X1 U21517 ( .C1(n18702), .C2(n18450), .A(n18417), .B(n18416), .ZN(
        P3_U2901) );
  AOI22_X1 U21518 ( .A1(n18703), .A2(n18429), .B1(n18667), .B2(n18452), .ZN(
        n18419) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18431), .B1(
        n18705), .B2(n18492), .ZN(n18418) );
  OAI211_X1 U21520 ( .C1(n18670), .C2(n18428), .A(n18419), .B(n18418), .ZN(
        P3_U2902) );
  AOI22_X1 U21521 ( .A1(n18511), .A2(n18430), .B1(n18709), .B2(n18429), .ZN(
        n18421) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18431), .B1(
        n18711), .B2(n18492), .ZN(n18420) );
  OAI211_X1 U21523 ( .C1(n18514), .C2(n18450), .A(n18421), .B(n18420), .ZN(
        P3_U2903) );
  AOI22_X1 U21524 ( .A1(n18613), .A2(n18452), .B1(n18715), .B2(n18429), .ZN(
        n18423) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18431), .B1(
        n18717), .B2(n18492), .ZN(n18422) );
  OAI211_X1 U21526 ( .C1(n18616), .C2(n18428), .A(n18423), .B(n18422), .ZN(
        P3_U2904) );
  AOI22_X1 U21527 ( .A1(n18566), .A2(n18452), .B1(n18721), .B2(n18429), .ZN(
        n18425) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18431), .B1(
        n18723), .B2(n18492), .ZN(n18424) );
  OAI211_X1 U21529 ( .C1(n18570), .C2(n18428), .A(n18425), .B(n18424), .ZN(
        P3_U2905) );
  AOI22_X1 U21530 ( .A1(n18619), .A2(n18452), .B1(n18727), .B2(n18429), .ZN(
        n18427) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18431), .B1(
        n18730), .B2(n18492), .ZN(n18426) );
  OAI211_X1 U21532 ( .C1(n18623), .C2(n18428), .A(n18427), .B(n18426), .ZN(
        P3_U2906) );
  AOI22_X1 U21533 ( .A1(n18626), .A2(n18430), .B1(n18736), .B2(n18429), .ZN(
        n18433) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18431), .B1(
        n18740), .B2(n18492), .ZN(n18432) );
  OAI211_X1 U21535 ( .C1(n18630), .C2(n18450), .A(n18433), .B(n18432), .ZN(
        P3_U2907) );
  NOR2_X1 U21536 ( .A1(n18480), .A2(n18527), .ZN(n18451) );
  AOI22_X1 U21537 ( .A1(n18688), .A2(n18470), .B1(n18687), .B2(n18451), .ZN(
        n18437) );
  AOI22_X1 U21538 ( .A1(n18692), .A2(n18435), .B1(n18479), .B2(n18434), .ZN(
        n18453) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18453), .B1(
        n18693), .B2(n9747), .ZN(n18436) );
  OAI211_X1 U21540 ( .C1(n18696), .C2(n18450), .A(n18437), .B(n18436), .ZN(
        P3_U2908) );
  AOI22_X1 U21541 ( .A1(n18637), .A2(n18470), .B1(n18697), .B2(n18451), .ZN(
        n18439) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18453), .B1(
        n18699), .B2(n9747), .ZN(n18438) );
  OAI211_X1 U21543 ( .C1(n18640), .C2(n18450), .A(n18439), .B(n18438), .ZN(
        P3_U2909) );
  AOI22_X1 U21544 ( .A1(n18703), .A2(n18451), .B1(n18667), .B2(n18470), .ZN(
        n18441) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18453), .B1(
        n18705), .B2(n9747), .ZN(n18440) );
  OAI211_X1 U21546 ( .C1(n18670), .C2(n18450), .A(n18441), .B(n18440), .ZN(
        P3_U2910) );
  AOI22_X1 U21547 ( .A1(n18709), .A2(n18451), .B1(n18710), .B2(n18470), .ZN(
        n18443) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18453), .B1(
        n18711), .B2(n9747), .ZN(n18442) );
  OAI211_X1 U21549 ( .C1(n18714), .C2(n18450), .A(n18443), .B(n18442), .ZN(
        P3_U2911) );
  AOI22_X1 U21550 ( .A1(n18715), .A2(n18451), .B1(n18716), .B2(n18452), .ZN(
        n18445) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18453), .B1(
        n18717), .B2(n9747), .ZN(n18444) );
  OAI211_X1 U21552 ( .C1(n18720), .C2(n18477), .A(n18445), .B(n18444), .ZN(
        P3_U2912) );
  AOI22_X1 U21553 ( .A1(n18721), .A2(n18451), .B1(n18722), .B2(n18452), .ZN(
        n18447) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18453), .B1(
        n18723), .B2(n9747), .ZN(n18446) );
  OAI211_X1 U21555 ( .C1(n18726), .C2(n18477), .A(n18447), .B(n18446), .ZN(
        P3_U2913) );
  AOI22_X1 U21556 ( .A1(n18619), .A2(n18470), .B1(n18727), .B2(n18451), .ZN(
        n18449) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18453), .B1(
        n18730), .B2(n9747), .ZN(n18448) );
  OAI211_X1 U21558 ( .C1(n18623), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        P3_U2914) );
  AOI22_X1 U21559 ( .A1(n18626), .A2(n18452), .B1(n18736), .B2(n18451), .ZN(
        n18455) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18453), .B1(
        n18740), .B2(n9747), .ZN(n18454) );
  OAI211_X1 U21561 ( .C1(n18630), .C2(n18477), .A(n18455), .B(n18454), .ZN(
        P3_U2915) );
  NOR2_X2 U21562 ( .A1(n18553), .A2(n18480), .ZN(n18549) );
  NOR2_X1 U21563 ( .A1(n9747), .A2(n18549), .ZN(n18503) );
  NOR2_X1 U21564 ( .A1(n18658), .A2(n18503), .ZN(n18473) );
  AOI22_X1 U21565 ( .A1(n18688), .A2(n18492), .B1(n18687), .B2(n18473), .ZN(
        n18459) );
  OAI21_X1 U21566 ( .B1(n18456), .B2(n18659), .A(n18503), .ZN(n18457) );
  OAI211_X1 U21567 ( .C1(n18549), .C2(n18910), .A(n18661), .B(n18457), .ZN(
        n18474) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18474), .B1(
        n18693), .B2(n18549), .ZN(n18458) );
  OAI211_X1 U21569 ( .C1(n18696), .C2(n18477), .A(n18459), .B(n18458), .ZN(
        P3_U2916) );
  INV_X1 U21570 ( .A(n18492), .ZN(n18501) );
  AOI22_X1 U21571 ( .A1(n18697), .A2(n18473), .B1(n18698), .B2(n18470), .ZN(
        n18461) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18474), .B1(
        n18699), .B2(n18549), .ZN(n18460) );
  OAI211_X1 U21573 ( .C1(n18702), .C2(n18501), .A(n18461), .B(n18460), .ZN(
        P3_U2917) );
  AOI22_X1 U21574 ( .A1(n18703), .A2(n18473), .B1(n18667), .B2(n18492), .ZN(
        n18463) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18474), .B1(
        n18705), .B2(n18549), .ZN(n18462) );
  OAI211_X1 U21576 ( .C1(n18670), .C2(n18477), .A(n18463), .B(n18462), .ZN(
        P3_U2918) );
  AOI22_X1 U21577 ( .A1(n18511), .A2(n18470), .B1(n18709), .B2(n18473), .ZN(
        n18465) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18474), .B1(
        n18711), .B2(n18549), .ZN(n18464) );
  OAI211_X1 U21579 ( .C1(n18514), .C2(n18501), .A(n18465), .B(n18464), .ZN(
        P3_U2919) );
  AOI22_X1 U21580 ( .A1(n18613), .A2(n18492), .B1(n18715), .B2(n18473), .ZN(
        n18467) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18474), .B1(
        n18717), .B2(n18549), .ZN(n18466) );
  OAI211_X1 U21582 ( .C1(n18616), .C2(n18477), .A(n18467), .B(n18466), .ZN(
        P3_U2920) );
  AOI22_X1 U21583 ( .A1(n18721), .A2(n18473), .B1(n18722), .B2(n18470), .ZN(
        n18469) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18474), .B1(
        n18723), .B2(n18549), .ZN(n18468) );
  OAI211_X1 U21585 ( .C1(n18726), .C2(n18501), .A(n18469), .B(n18468), .ZN(
        P3_U2921) );
  AOI22_X1 U21586 ( .A1(n18727), .A2(n18473), .B1(n18728), .B2(n18470), .ZN(
        n18472) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18474), .B1(
        n18730), .B2(n18549), .ZN(n18471) );
  OAI211_X1 U21588 ( .C1(n18733), .C2(n18501), .A(n18472), .B(n18471), .ZN(
        P3_U2922) );
  AOI22_X1 U21589 ( .A1(n18737), .A2(n18492), .B1(n18736), .B2(n18473), .ZN(
        n18476) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18474), .B1(
        n18740), .B2(n18549), .ZN(n18475) );
  OAI211_X1 U21591 ( .C1(n18744), .C2(n18477), .A(n18476), .B(n18475), .ZN(
        P3_U2923) );
  AOI22_X1 U21592 ( .A1(n18688), .A2(n9747), .B1(n18687), .B2(n18497), .ZN(
        n18483) );
  NAND2_X1 U21593 ( .A1(n18479), .A2(n18478), .ZN(n18498) );
  NOR2_X2 U21594 ( .A1(n18481), .A2(n18480), .ZN(n18574) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18498), .B1(
        n18693), .B2(n18574), .ZN(n18482) );
  OAI211_X1 U21596 ( .C1(n18696), .C2(n18501), .A(n18483), .B(n18482), .ZN(
        P3_U2924) );
  AOI22_X1 U21597 ( .A1(n18637), .A2(n9747), .B1(n18697), .B2(n18497), .ZN(
        n18485) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18498), .B1(
        n18699), .B2(n18574), .ZN(n18484) );
  OAI211_X1 U21599 ( .C1(n18640), .C2(n18501), .A(n18485), .B(n18484), .ZN(
        P3_U2925) );
  INV_X1 U21600 ( .A(n9747), .ZN(n18519) );
  AOI22_X1 U21601 ( .A1(n18704), .A2(n18492), .B1(n18703), .B2(n18497), .ZN(
        n18487) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18498), .B1(
        n18705), .B2(n18574), .ZN(n18486) );
  OAI211_X1 U21603 ( .C1(n18708), .C2(n18519), .A(n18487), .B(n18486), .ZN(
        P3_U2926) );
  AOI22_X1 U21604 ( .A1(n18709), .A2(n18497), .B1(n18710), .B2(n9747), .ZN(
        n18489) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18498), .B1(
        n18711), .B2(n18574), .ZN(n18488) );
  OAI211_X1 U21606 ( .C1(n18714), .C2(n18501), .A(n18489), .B(n18488), .ZN(
        P3_U2927) );
  AOI22_X1 U21607 ( .A1(n18613), .A2(n9747), .B1(n18715), .B2(n18497), .ZN(
        n18491) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18498), .B1(
        n18717), .B2(n18574), .ZN(n18490) );
  OAI211_X1 U21609 ( .C1(n18616), .C2(n18501), .A(n18491), .B(n18490), .ZN(
        P3_U2928) );
  AOI22_X1 U21610 ( .A1(n18721), .A2(n18497), .B1(n18722), .B2(n18492), .ZN(
        n18494) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18498), .B1(
        n18723), .B2(n18574), .ZN(n18493) );
  OAI211_X1 U21612 ( .C1(n18726), .C2(n18519), .A(n18494), .B(n18493), .ZN(
        P3_U2929) );
  AOI22_X1 U21613 ( .A1(n18619), .A2(n9747), .B1(n18727), .B2(n18497), .ZN(
        n18496) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18498), .B1(
        n18730), .B2(n18574), .ZN(n18495) );
  OAI211_X1 U21615 ( .C1(n18623), .C2(n18501), .A(n18496), .B(n18495), .ZN(
        P3_U2930) );
  AOI22_X1 U21616 ( .A1(n18737), .A2(n9747), .B1(n18736), .B2(n18497), .ZN(
        n18500) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18498), .B1(
        n18740), .B2(n18574), .ZN(n18499) );
  OAI211_X1 U21618 ( .C1(n18744), .C2(n18501), .A(n18500), .B(n18499), .ZN(
        P3_U2931) );
  INV_X1 U21619 ( .A(n18600), .ZN(n18578) );
  NOR2_X2 U21620 ( .A1(n18502), .A2(n18578), .ZN(n18590) );
  NOR2_X1 U21621 ( .A1(n18574), .A2(n18590), .ZN(n18554) );
  OAI21_X1 U21622 ( .B1(n18503), .B2(n18659), .A(n18554), .ZN(n18504) );
  OAI211_X1 U21623 ( .C1(n18590), .C2(n18910), .A(n18661), .B(n18504), .ZN(
        n18524) );
  NOR2_X1 U21624 ( .A1(n18658), .A2(n18554), .ZN(n18522) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18524), .B1(
        n18687), .B2(n18522), .ZN(n18506) );
  AOI22_X1 U21626 ( .A1(n18693), .A2(n18590), .B1(n18688), .B2(n18549), .ZN(
        n18505) );
  OAI211_X1 U21627 ( .C1(n18696), .C2(n18519), .A(n18506), .B(n18505), .ZN(
        P3_U2932) );
  INV_X1 U21628 ( .A(n18549), .ZN(n18547) );
  AOI22_X1 U21629 ( .A1(n18697), .A2(n18522), .B1(n18698), .B2(n9747), .ZN(
        n18508) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18524), .B1(
        n18699), .B2(n18590), .ZN(n18507) );
  OAI211_X1 U21631 ( .C1(n18702), .C2(n18547), .A(n18508), .B(n18507), .ZN(
        P3_U2933) );
  AOI22_X1 U21632 ( .A1(n18704), .A2(n9747), .B1(n18703), .B2(n18522), .ZN(
        n18510) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18524), .B1(
        n18705), .B2(n18590), .ZN(n18509) );
  OAI211_X1 U21634 ( .C1(n18708), .C2(n18547), .A(n18510), .B(n18509), .ZN(
        P3_U2934) );
  AOI22_X1 U21635 ( .A1(n18511), .A2(n9747), .B1(n18709), .B2(n18522), .ZN(
        n18513) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18524), .B1(
        n18711), .B2(n18590), .ZN(n18512) );
  OAI211_X1 U21637 ( .C1(n18514), .C2(n18547), .A(n18513), .B(n18512), .ZN(
        P3_U2935) );
  AOI22_X1 U21638 ( .A1(n18715), .A2(n18522), .B1(n18716), .B2(n9747), .ZN(
        n18516) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18524), .B1(
        n18717), .B2(n18590), .ZN(n18515) );
  OAI211_X1 U21640 ( .C1(n18720), .C2(n18547), .A(n18516), .B(n18515), .ZN(
        P3_U2936) );
  AOI22_X1 U21641 ( .A1(n18566), .A2(n18549), .B1(n18721), .B2(n18522), .ZN(
        n18518) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18524), .B1(
        n18723), .B2(n18590), .ZN(n18517) );
  OAI211_X1 U21643 ( .C1(n18570), .C2(n18519), .A(n18518), .B(n18517), .ZN(
        P3_U2937) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18524), .B1(
        n18727), .B2(n18522), .ZN(n18521) );
  AOI22_X1 U21645 ( .A1(n18730), .A2(n18590), .B1(n18728), .B2(n9747), .ZN(
        n18520) );
  OAI211_X1 U21646 ( .C1(n18733), .C2(n18547), .A(n18521), .B(n18520), .ZN(
        P3_U2938) );
  AOI22_X1 U21647 ( .A1(n18626), .A2(n9747), .B1(n18736), .B2(n18522), .ZN(
        n18526) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18524), .B1(
        n18740), .B2(n18590), .ZN(n18525) );
  OAI211_X1 U21649 ( .C1(n18630), .C2(n18547), .A(n18526), .B(n18525), .ZN(
        P3_U2939) );
  NOR2_X1 U21650 ( .A1(n18578), .A2(n18527), .ZN(n18548) );
  AOI22_X1 U21651 ( .A1(n18688), .A2(n18574), .B1(n18687), .B2(n18548), .ZN(
        n18534) );
  NOR2_X1 U21652 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18528), .ZN(
        n18531) );
  INV_X1 U21653 ( .A(n18529), .ZN(n18690) );
  NOR2_X1 U21654 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18578), .ZN(
        n18530) );
  AOI22_X1 U21655 ( .A1(n18692), .A2(n18531), .B1(n18690), .B2(n18530), .ZN(
        n18550) );
  NOR2_X2 U21656 ( .A1(n18578), .A2(n18532), .ZN(n18625) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18550), .B1(
        n18693), .B2(n18625), .ZN(n18533) );
  OAI211_X1 U21658 ( .C1(n18696), .C2(n18547), .A(n18534), .B(n18533), .ZN(
        P3_U2940) );
  INV_X1 U21659 ( .A(n18574), .ZN(n18569) );
  AOI22_X1 U21660 ( .A1(n18697), .A2(n18548), .B1(n18698), .B2(n18549), .ZN(
        n18536) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18550), .B1(
        n18699), .B2(n18625), .ZN(n18535) );
  OAI211_X1 U21662 ( .C1(n18702), .C2(n18569), .A(n18536), .B(n18535), .ZN(
        P3_U2941) );
  AOI22_X1 U21663 ( .A1(n18704), .A2(n18549), .B1(n18703), .B2(n18548), .ZN(
        n18538) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18550), .B1(
        n18705), .B2(n18625), .ZN(n18537) );
  OAI211_X1 U21665 ( .C1(n18708), .C2(n18569), .A(n18538), .B(n18537), .ZN(
        P3_U2942) );
  AOI22_X1 U21666 ( .A1(n18709), .A2(n18548), .B1(n18710), .B2(n18574), .ZN(
        n18540) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18550), .B1(
        n18711), .B2(n18625), .ZN(n18539) );
  OAI211_X1 U21668 ( .C1(n18714), .C2(n18547), .A(n18540), .B(n18539), .ZN(
        P3_U2943) );
  AOI22_X1 U21669 ( .A1(n18715), .A2(n18548), .B1(n18716), .B2(n18549), .ZN(
        n18542) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18550), .B1(
        n18717), .B2(n18625), .ZN(n18541) );
  OAI211_X1 U21671 ( .C1(n18720), .C2(n18569), .A(n18542), .B(n18541), .ZN(
        P3_U2944) );
  AOI22_X1 U21672 ( .A1(n18566), .A2(n18574), .B1(n18721), .B2(n18548), .ZN(
        n18544) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18550), .B1(
        n18723), .B2(n18625), .ZN(n18543) );
  OAI211_X1 U21674 ( .C1(n18570), .C2(n18547), .A(n18544), .B(n18543), .ZN(
        P3_U2945) );
  AOI22_X1 U21675 ( .A1(n18619), .A2(n18574), .B1(n18727), .B2(n18548), .ZN(
        n18546) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18550), .B1(
        n18730), .B2(n18625), .ZN(n18545) );
  OAI211_X1 U21677 ( .C1(n18623), .C2(n18547), .A(n18546), .B(n18545), .ZN(
        P3_U2946) );
  AOI22_X1 U21678 ( .A1(n18626), .A2(n18549), .B1(n18736), .B2(n18548), .ZN(
        n18552) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18550), .B1(
        n18740), .B2(n18625), .ZN(n18551) );
  OAI211_X1 U21680 ( .C1(n18630), .C2(n18569), .A(n18552), .B(n18551), .ZN(
        P3_U2947) );
  AOI22_X1 U21681 ( .A1(n18688), .A2(n18590), .B1(n18687), .B2(n18573), .ZN(
        n18557) );
  NOR2_X2 U21682 ( .A1(n18578), .A2(n18553), .ZN(n18649) );
  INV_X1 U21683 ( .A(n18625), .ZN(n18622) );
  AOI221_X1 U21684 ( .B1(n18554), .B2(n18622), .C1(n18659), .C2(n18622), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18555) );
  OAI21_X1 U21685 ( .B1(n18649), .B2(n18555), .A(n18661), .ZN(n18575) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18575), .B1(
        n18693), .B2(n18649), .ZN(n18556) );
  OAI211_X1 U21687 ( .C1(n18696), .C2(n18569), .A(n18557), .B(n18556), .ZN(
        P3_U2948) );
  AOI22_X1 U21688 ( .A1(n18637), .A2(n18590), .B1(n18697), .B2(n18573), .ZN(
        n18559) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18575), .B1(
        n18699), .B2(n18649), .ZN(n18558) );
  OAI211_X1 U21690 ( .C1(n18640), .C2(n18569), .A(n18559), .B(n18558), .ZN(
        P3_U2949) );
  AOI22_X1 U21691 ( .A1(n18703), .A2(n18573), .B1(n18667), .B2(n18590), .ZN(
        n18561) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18575), .B1(
        n18705), .B2(n18649), .ZN(n18560) );
  OAI211_X1 U21693 ( .C1(n18670), .C2(n18569), .A(n18561), .B(n18560), .ZN(
        P3_U2950) );
  AOI22_X1 U21694 ( .A1(n18709), .A2(n18573), .B1(n18710), .B2(n18590), .ZN(
        n18563) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18575), .B1(
        n18711), .B2(n18649), .ZN(n18562) );
  OAI211_X1 U21696 ( .C1(n18714), .C2(n18569), .A(n18563), .B(n18562), .ZN(
        P3_U2951) );
  INV_X1 U21697 ( .A(n18590), .ZN(n18599) );
  AOI22_X1 U21698 ( .A1(n18715), .A2(n18573), .B1(n18716), .B2(n18574), .ZN(
        n18565) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18575), .B1(
        n18717), .B2(n18649), .ZN(n18564) );
  OAI211_X1 U21700 ( .C1(n18720), .C2(n18599), .A(n18565), .B(n18564), .ZN(
        P3_U2952) );
  AOI22_X1 U21701 ( .A1(n18566), .A2(n18590), .B1(n18721), .B2(n18573), .ZN(
        n18568) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18575), .B1(
        n18723), .B2(n18649), .ZN(n18567) );
  OAI211_X1 U21703 ( .C1(n18570), .C2(n18569), .A(n18568), .B(n18567), .ZN(
        P3_U2953) );
  AOI22_X1 U21704 ( .A1(n18727), .A2(n18573), .B1(n18728), .B2(n18574), .ZN(
        n18572) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18575), .B1(
        n18730), .B2(n18649), .ZN(n18571) );
  OAI211_X1 U21706 ( .C1(n18733), .C2(n18599), .A(n18572), .B(n18571), .ZN(
        P3_U2954) );
  AOI22_X1 U21707 ( .A1(n18626), .A2(n18574), .B1(n18736), .B2(n18573), .ZN(
        n18577) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18575), .B1(
        n18740), .B2(n18649), .ZN(n18576) );
  OAI211_X1 U21709 ( .C1(n18630), .C2(n18599), .A(n18577), .B(n18576), .ZN(
        P3_U2955) );
  NOR2_X1 U21710 ( .A1(n18579), .A2(n18578), .ZN(n18633) );
  AND2_X1 U21711 ( .A1(n18806), .A2(n18633), .ZN(n18595) );
  AOI22_X1 U21712 ( .A1(n18688), .A2(n18625), .B1(n18687), .B2(n18595), .ZN(
        n18581) );
  OAI211_X1 U21713 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18692), .A(
        n18690), .B(n18600), .ZN(n18596) );
  NAND2_X1 U21714 ( .A1(n18772), .A2(n18600), .ZN(n18686) );
  INV_X1 U21715 ( .A(n18686), .ZN(n18678) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18693), .ZN(n18580) );
  OAI211_X1 U21717 ( .C1(n18696), .C2(n18599), .A(n18581), .B(n18580), .ZN(
        P3_U2956) );
  AOI22_X1 U21718 ( .A1(n18697), .A2(n18595), .B1(n18698), .B2(n18590), .ZN(
        n18583) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18699), .ZN(n18582) );
  OAI211_X1 U21720 ( .C1(n18702), .C2(n18622), .A(n18583), .B(n18582), .ZN(
        P3_U2957) );
  AOI22_X1 U21721 ( .A1(n18703), .A2(n18595), .B1(n18667), .B2(n18625), .ZN(
        n18585) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18705), .ZN(n18584) );
  OAI211_X1 U21723 ( .C1(n18670), .C2(n18599), .A(n18585), .B(n18584), .ZN(
        P3_U2958) );
  AOI22_X1 U21724 ( .A1(n18709), .A2(n18595), .B1(n18710), .B2(n18625), .ZN(
        n18587) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18711), .ZN(n18586) );
  OAI211_X1 U21726 ( .C1(n18714), .C2(n18599), .A(n18587), .B(n18586), .ZN(
        P3_U2959) );
  AOI22_X1 U21727 ( .A1(n18613), .A2(n18625), .B1(n18715), .B2(n18595), .ZN(
        n18589) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18717), .ZN(n18588) );
  OAI211_X1 U21729 ( .C1(n18616), .C2(n18599), .A(n18589), .B(n18588), .ZN(
        P3_U2960) );
  AOI22_X1 U21730 ( .A1(n18721), .A2(n18595), .B1(n18722), .B2(n18590), .ZN(
        n18592) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18723), .ZN(n18591) );
  OAI211_X1 U21732 ( .C1(n18726), .C2(n18622), .A(n18592), .B(n18591), .ZN(
        P3_U2961) );
  AOI22_X1 U21733 ( .A1(n18619), .A2(n18625), .B1(n18727), .B2(n18595), .ZN(
        n18594) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18730), .ZN(n18593) );
  OAI211_X1 U21735 ( .C1(n18623), .C2(n18599), .A(n18594), .B(n18593), .ZN(
        P3_U2962) );
  AOI22_X1 U21736 ( .A1(n18737), .A2(n18625), .B1(n18736), .B2(n18595), .ZN(
        n18598) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18596), .B1(
        n18678), .B2(n18740), .ZN(n18597) );
  OAI211_X1 U21738 ( .C1(n18744), .C2(n18599), .A(n18598), .B(n18597), .ZN(
        P3_U2963) );
  INV_X1 U21739 ( .A(n18691), .ZN(n18631) );
  NOR2_X2 U21740 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18631), .ZN(
        n18729) );
  NOR2_X1 U21741 ( .A1(n18678), .A2(n18729), .ZN(n18660) );
  NOR2_X1 U21742 ( .A1(n18658), .A2(n18660), .ZN(n18624) );
  AOI22_X1 U21743 ( .A1(n18688), .A2(n18649), .B1(n18687), .B2(n18624), .ZN(
        n18606) );
  NAND2_X1 U21744 ( .A1(n18601), .A2(n18600), .ZN(n18602) );
  OAI21_X1 U21745 ( .B1(n18603), .B2(n18602), .A(n18660), .ZN(n18604) );
  OAI211_X1 U21746 ( .C1(n18729), .C2(n18910), .A(n18661), .B(n18604), .ZN(
        n18627) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18627), .B1(
        n18729), .B2(n18693), .ZN(n18605) );
  OAI211_X1 U21748 ( .C1(n18696), .C2(n18622), .A(n18606), .B(n18605), .ZN(
        P3_U2964) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18627), .B1(
        n18697), .B2(n18624), .ZN(n18608) );
  AOI22_X1 U21750 ( .A1(n18729), .A2(n18699), .B1(n18637), .B2(n18649), .ZN(
        n18607) );
  OAI211_X1 U21751 ( .C1(n18640), .C2(n18622), .A(n18608), .B(n18607), .ZN(
        P3_U2965) );
  AOI22_X1 U21752 ( .A1(n18703), .A2(n18624), .B1(n18667), .B2(n18649), .ZN(
        n18610) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18627), .B1(
        n18729), .B2(n18705), .ZN(n18609) );
  OAI211_X1 U21754 ( .C1(n18670), .C2(n18622), .A(n18610), .B(n18609), .ZN(
        P3_U2966) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18627), .B1(
        n18709), .B2(n18624), .ZN(n18612) );
  AOI22_X1 U21756 ( .A1(n18729), .A2(n18711), .B1(n18710), .B2(n18649), .ZN(
        n18611) );
  OAI211_X1 U21757 ( .C1(n18714), .C2(n18622), .A(n18612), .B(n18611), .ZN(
        P3_U2967) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18627), .B1(
        n18715), .B2(n18624), .ZN(n18615) );
  AOI22_X1 U21759 ( .A1(n18729), .A2(n18717), .B1(n18613), .B2(n18649), .ZN(
        n18614) );
  OAI211_X1 U21760 ( .C1(n18616), .C2(n18622), .A(n18615), .B(n18614), .ZN(
        P3_U2968) );
  INV_X1 U21761 ( .A(n18649), .ZN(n18656) );
  AOI22_X1 U21762 ( .A1(n18721), .A2(n18624), .B1(n18722), .B2(n18625), .ZN(
        n18618) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18627), .B1(
        n18729), .B2(n18723), .ZN(n18617) );
  OAI211_X1 U21764 ( .C1(n18726), .C2(n18656), .A(n18618), .B(n18617), .ZN(
        P3_U2969) );
  AOI22_X1 U21765 ( .A1(n18619), .A2(n18649), .B1(n18727), .B2(n18624), .ZN(
        n18621) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18627), .B1(
        n18729), .B2(n18730), .ZN(n18620) );
  OAI211_X1 U21767 ( .C1(n18623), .C2(n18622), .A(n18621), .B(n18620), .ZN(
        P3_U2970) );
  AOI22_X1 U21768 ( .A1(n18626), .A2(n18625), .B1(n18736), .B2(n18624), .ZN(
        n18629) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18627), .B1(
        n18729), .B2(n18740), .ZN(n18628) );
  OAI211_X1 U21770 ( .C1(n18630), .C2(n18656), .A(n18629), .B(n18628), .ZN(
        P3_U2971) );
  NOR2_X1 U21771 ( .A1(n18658), .A2(n18631), .ZN(n18652) );
  AOI22_X1 U21772 ( .A1(n18632), .A2(n18649), .B1(n18687), .B2(n18652), .ZN(
        n18635) );
  AOI22_X1 U21773 ( .A1(n18692), .A2(n18633), .B1(n18691), .B2(n18690), .ZN(
        n18653) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18693), .ZN(n18634) );
  OAI211_X1 U21775 ( .C1(n18686), .C2(n18636), .A(n18635), .B(n18634), .ZN(
        P3_U2972) );
  AOI22_X1 U21776 ( .A1(n18678), .A2(n18637), .B1(n18697), .B2(n18652), .ZN(
        n18639) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18699), .ZN(n18638) );
  OAI211_X1 U21778 ( .C1(n18640), .C2(n18656), .A(n18639), .B(n18638), .ZN(
        P3_U2973) );
  AOI22_X1 U21779 ( .A1(n18704), .A2(n18649), .B1(n18703), .B2(n18652), .ZN(
        n18642) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18705), .ZN(n18641) );
  OAI211_X1 U21781 ( .C1(n18686), .C2(n18708), .A(n18642), .B(n18641), .ZN(
        P3_U2974) );
  AOI22_X1 U21782 ( .A1(n18678), .A2(n18710), .B1(n18709), .B2(n18652), .ZN(
        n18644) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18711), .ZN(n18643) );
  OAI211_X1 U21784 ( .C1(n18714), .C2(n18656), .A(n18644), .B(n18643), .ZN(
        P3_U2975) );
  AOI22_X1 U21785 ( .A1(n18715), .A2(n18652), .B1(n18716), .B2(n18649), .ZN(
        n18646) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18717), .ZN(n18645) );
  OAI211_X1 U21787 ( .C1(n18686), .C2(n18720), .A(n18646), .B(n18645), .ZN(
        P3_U2976) );
  AOI22_X1 U21788 ( .A1(n18721), .A2(n18652), .B1(n18722), .B2(n18649), .ZN(
        n18648) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18723), .ZN(n18647) );
  OAI211_X1 U21790 ( .C1(n18686), .C2(n18726), .A(n18648), .B(n18647), .ZN(
        P3_U2977) );
  AOI22_X1 U21791 ( .A1(n18727), .A2(n18652), .B1(n18728), .B2(n18649), .ZN(
        n18651) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18730), .ZN(n18650) );
  OAI211_X1 U21793 ( .C1(n18686), .C2(n18733), .A(n18651), .B(n18650), .ZN(
        P3_U2978) );
  AOI22_X1 U21794 ( .A1(n18678), .A2(n18737), .B1(n18736), .B2(n18652), .ZN(
        n18655) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18653), .B1(
        n18738), .B2(n18740), .ZN(n18654) );
  OAI211_X1 U21796 ( .C1(n18744), .C2(n18656), .A(n18655), .B(n18654), .ZN(
        P3_U2979) );
  NOR2_X1 U21797 ( .A1(n18658), .A2(n18657), .ZN(n18681) );
  AOI22_X1 U21798 ( .A1(n18729), .A2(n18688), .B1(n18687), .B2(n18681), .ZN(
        n18664) );
  AOI221_X1 U21799 ( .B1(n18660), .B2(n18734), .C1(n18659), .C2(n18734), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18662) );
  OAI21_X1 U21800 ( .B1(n18682), .B2(n18662), .A(n18661), .ZN(n18683) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18683), .B1(
        n18673), .B2(n18693), .ZN(n18663) );
  OAI211_X1 U21802 ( .C1(n18696), .C2(n18686), .A(n18664), .B(n18663), .ZN(
        P3_U2980) );
  INV_X1 U21803 ( .A(n18729), .ZN(n18745) );
  AOI22_X1 U21804 ( .A1(n18678), .A2(n18698), .B1(n18681), .B2(n18697), .ZN(
        n18666) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18683), .B1(
        n18673), .B2(n18699), .ZN(n18665) );
  OAI211_X1 U21806 ( .C1(n18745), .C2(n18702), .A(n18666), .B(n18665), .ZN(
        P3_U2981) );
  AOI22_X1 U21807 ( .A1(n18729), .A2(n18667), .B1(n18681), .B2(n18703), .ZN(
        n18669) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18683), .B1(
        n18682), .B2(n18705), .ZN(n18668) );
  OAI211_X1 U21809 ( .C1(n18686), .C2(n18670), .A(n18669), .B(n18668), .ZN(
        P3_U2982) );
  AOI22_X1 U21810 ( .A1(n18729), .A2(n18710), .B1(n18681), .B2(n18709), .ZN(
        n18672) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18683), .B1(
        n18682), .B2(n18711), .ZN(n18671) );
  OAI211_X1 U21812 ( .C1(n18686), .C2(n18714), .A(n18672), .B(n18671), .ZN(
        P3_U2983) );
  AOI22_X1 U21813 ( .A1(n18678), .A2(n18716), .B1(n18681), .B2(n18715), .ZN(
        n18675) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18683), .B1(
        n18673), .B2(n18717), .ZN(n18674) );
  OAI211_X1 U21815 ( .C1(n18745), .C2(n18720), .A(n18675), .B(n18674), .ZN(
        P3_U2984) );
  AOI22_X1 U21816 ( .A1(n18678), .A2(n18722), .B1(n18681), .B2(n18721), .ZN(
        n18677) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18683), .B1(
        n18682), .B2(n18723), .ZN(n18676) );
  OAI211_X1 U21818 ( .C1(n18745), .C2(n18726), .A(n18677), .B(n18676), .ZN(
        P3_U2985) );
  AOI22_X1 U21819 ( .A1(n18678), .A2(n18728), .B1(n18681), .B2(n18727), .ZN(
        n18680) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18683), .B1(
        n18682), .B2(n18730), .ZN(n18679) );
  OAI211_X1 U21821 ( .C1(n18745), .C2(n18733), .A(n18680), .B(n18679), .ZN(
        P3_U2986) );
  AOI22_X1 U21822 ( .A1(n18729), .A2(n18737), .B1(n18681), .B2(n18736), .ZN(
        n18685) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18683), .B1(
        n18682), .B2(n18740), .ZN(n18684) );
  OAI211_X1 U21824 ( .C1(n18686), .C2(n18744), .A(n18685), .B(n18684), .ZN(
        P3_U2987) );
  AND2_X1 U21825 ( .A1(n18806), .A2(n18689), .ZN(n18735) );
  AOI22_X1 U21826 ( .A1(n18738), .A2(n18688), .B1(n18687), .B2(n18735), .ZN(
        n18695) );
  AOI22_X1 U21827 ( .A1(n18692), .A2(n18691), .B1(n18690), .B2(n18689), .ZN(
        n18741) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18741), .B1(
        n18693), .B2(n18739), .ZN(n18694) );
  OAI211_X1 U21829 ( .C1(n18696), .C2(n18745), .A(n18695), .B(n18694), .ZN(
        P3_U2988) );
  AOI22_X1 U21830 ( .A1(n18729), .A2(n18698), .B1(n18697), .B2(n18735), .ZN(
        n18701) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18741), .B1(
        n18699), .B2(n18739), .ZN(n18700) );
  OAI211_X1 U21832 ( .C1(n18734), .C2(n18702), .A(n18701), .B(n18700), .ZN(
        P3_U2989) );
  AOI22_X1 U21833 ( .A1(n18729), .A2(n18704), .B1(n18703), .B2(n18735), .ZN(
        n18707) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18741), .B1(
        n18705), .B2(n18739), .ZN(n18706) );
  OAI211_X1 U21835 ( .C1(n18734), .C2(n18708), .A(n18707), .B(n18706), .ZN(
        P3_U2990) );
  AOI22_X1 U21836 ( .A1(n18738), .A2(n18710), .B1(n18709), .B2(n18735), .ZN(
        n18713) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18741), .B1(
        n18711), .B2(n18739), .ZN(n18712) );
  OAI211_X1 U21838 ( .C1(n18745), .C2(n18714), .A(n18713), .B(n18712), .ZN(
        P3_U2991) );
  AOI22_X1 U21839 ( .A1(n18729), .A2(n18716), .B1(n18715), .B2(n18735), .ZN(
        n18719) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18741), .B1(
        n18717), .B2(n18739), .ZN(n18718) );
  OAI211_X1 U21841 ( .C1(n18734), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P3_U2992) );
  AOI22_X1 U21842 ( .A1(n18729), .A2(n18722), .B1(n18721), .B2(n18735), .ZN(
        n18725) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18741), .B1(
        n18723), .B2(n18739), .ZN(n18724) );
  OAI211_X1 U21844 ( .C1(n18734), .C2(n18726), .A(n18725), .B(n18724), .ZN(
        P3_U2993) );
  AOI22_X1 U21845 ( .A1(n18729), .A2(n18728), .B1(n18727), .B2(n18735), .ZN(
        n18732) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18741), .B1(
        n18730), .B2(n18739), .ZN(n18731) );
  OAI211_X1 U21847 ( .C1(n18734), .C2(n18733), .A(n18732), .B(n18731), .ZN(
        P3_U2994) );
  AOI22_X1 U21848 ( .A1(n18738), .A2(n18737), .B1(n18736), .B2(n18735), .ZN(
        n18743) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18741), .B1(
        n18740), .B2(n18739), .ZN(n18742) );
  OAI211_X1 U21850 ( .C1(n18745), .C2(n18744), .A(n18743), .B(n18742), .ZN(
        P3_U2995) );
  INV_X1 U21851 ( .A(n18962), .ZN(n18957) );
  INV_X1 U21852 ( .A(n18955), .ZN(n18796) );
  AOI21_X1 U21853 ( .B1(n18748), .B2(n18747), .A(n18746), .ZN(n18752) );
  AOI21_X1 U21854 ( .B1(n18781), .B2(n18750), .A(n18749), .ZN(n18751) );
  AOI211_X1 U21855 ( .C1(n18754), .C2(n18753), .A(n18752), .B(n18751), .ZN(
        n18953) );
  AOI211_X1 U21856 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18783), .A(
        n18756), .B(n18755), .ZN(n18795) );
  OAI21_X1 U21857 ( .B1(n18759), .B2(n18758), .A(n18757), .ZN(n18777) );
  AOI22_X1 U21858 ( .A1(n18771), .A2(n18775), .B1(n18760), .B2(n18777), .ZN(
        n18761) );
  NAND2_X1 U21859 ( .A1(n11534), .A2(n18778), .ZN(n18762) );
  NAND2_X1 U21860 ( .A1(n18761), .A2(n18762), .ZN(n18917) );
  NOR2_X1 U21861 ( .A1(n18783), .A2(n18917), .ZN(n18767) );
  INV_X1 U21862 ( .A(n18762), .ZN(n18765) );
  OAI21_X1 U21863 ( .B1(n16981), .B2(n18769), .A(n18763), .ZN(n18776) );
  INV_X1 U21864 ( .A(n18776), .ZN(n18764) );
  OAI22_X1 U21865 ( .A1(n18765), .A2(n18781), .B1(n18764), .B2(n18775), .ZN(
        n18914) );
  NAND2_X1 U21866 ( .A1(n18918), .A2(n18914), .ZN(n18766) );
  OAI22_X1 U21867 ( .A1(n18767), .A2(n18918), .B1(n18783), .B2(n18766), .ZN(
        n18790) );
  NAND2_X1 U21868 ( .A1(n18769), .A2(n18768), .ZN(n18770) );
  AOI22_X1 U21869 ( .A1(n18931), .A2(n18770), .B1(n18776), .B2(n18934), .ZN(
        n18927) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18771), .B1(
        n18770), .B2(n16981), .ZN(n18935) );
  AOI222_X1 U21871 ( .A1(n18927), .A2(n18935), .B1(n18927), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18935), .C2(n18772), .ZN(
        n18774) );
  AOI21_X1 U21872 ( .B1(n18774), .B2(n18782), .A(n18773), .ZN(n18785) );
  OAI211_X1 U21873 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18776), .B(n18775), .ZN(
        n18780) );
  NAND3_X1 U21874 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18778), .A3(
        n18777), .ZN(n18779) );
  OAI211_X1 U21875 ( .C1(n18924), .C2(n18781), .A(n18780), .B(n18779), .ZN(
        n18925) );
  AOI22_X1 U21876 ( .A1(n18783), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18925), .B2(n18782), .ZN(n18786) );
  OR2_X1 U21877 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18786), .ZN(
        n18784) );
  AOI221_X1 U21878 ( .B1(n18785), .B2(n18784), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18786), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18789) );
  OAI21_X1 U21879 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18786), .ZN(n18788) );
  AOI222_X1 U21880 ( .A1(n18790), .A2(n18789), .B1(n18790), .B2(n18788), .C1(
        n18789), .C2(n18787), .ZN(n18794) );
  INV_X1 U21881 ( .A(n18791), .ZN(n18792) );
  OAI21_X1 U21882 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n18792), .ZN(n18793) );
  NAND4_X1 U21883 ( .A1(n18953), .A2(n18795), .A3(n18794), .A4(n18793), .ZN(
        n18802) );
  AOI211_X1 U21884 ( .C1(n18798), .C2(n18797), .A(n18796), .B(n18802), .ZN(
        n18908) );
  AOI21_X1 U21885 ( .B1(n18957), .B2(n18973), .A(n18908), .ZN(n18807) );
  OAI211_X1 U21886 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18799), .A(
        P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .ZN(n20990)
         );
  NOR2_X1 U21887 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18965) );
  NOR2_X1 U21888 ( .A1(n18962), .A2(n18956), .ZN(n18804) );
  AOI211_X1 U21889 ( .C1(n18936), .C2(n18965), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18804), .ZN(n18800) );
  AOI211_X1 U21890 ( .C1(n18955), .C2(n18802), .A(n18801), .B(n18800), .ZN(
        n18803) );
  OAI221_X1 U21891 ( .B1(n20997), .B2(n18807), .C1(n20997), .C2(n20990), .A(
        n18803), .ZN(P3_U2996) );
  INV_X1 U21892 ( .A(n18804), .ZN(n18810) );
  NAND4_X1 U21893 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18957), .A4(n18973), .ZN(n18812) );
  INV_X1 U21894 ( .A(n18805), .ZN(n18808) );
  NAND3_X1 U21895 ( .A1(n18808), .A2(n18807), .A3(n18806), .ZN(n18809) );
  NAND4_X1 U21896 ( .A1(n18811), .A2(n18810), .A3(n18812), .A4(n18809), .ZN(
        P3_U2997) );
  INV_X1 U21897 ( .A(n18965), .ZN(n18814) );
  AND4_X1 U21898 ( .A1(n18814), .A2(n18813), .A3(n18812), .A4(n18909), .ZN(
        P3_U2998) );
  AND2_X1 U21899 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18904), .ZN(
        P3_U2999) );
  INV_X1 U21900 ( .A(n18907), .ZN(n18815) );
  AND2_X1 U21901 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18815), .ZN(
        P3_U3000) );
  AND2_X1 U21902 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18815), .ZN(
        P3_U3001) );
  AND2_X1 U21903 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18815), .ZN(
        P3_U3002) );
  INV_X1 U21904 ( .A(P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21228) );
  NOR2_X1 U21905 ( .A1(n21228), .A2(n18907), .ZN(P3_U3003) );
  AND2_X1 U21906 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18815), .ZN(
        P3_U3004) );
  AND2_X1 U21907 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18815), .ZN(
        P3_U3005) );
  AND2_X1 U21908 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18815), .ZN(
        P3_U3006) );
  AND2_X1 U21909 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18815), .ZN(
        P3_U3007) );
  AND2_X1 U21910 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18815), .ZN(
        P3_U3008) );
  AND2_X1 U21911 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18815), .ZN(
        P3_U3009) );
  AND2_X1 U21912 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18815), .ZN(
        P3_U3010) );
  AND2_X1 U21913 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18815), .ZN(
        P3_U3011) );
  AND2_X1 U21914 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18815), .ZN(
        P3_U3012) );
  AND2_X1 U21915 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18815), .ZN(
        P3_U3013) );
  AND2_X1 U21916 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18815), .ZN(
        P3_U3014) );
  AND2_X1 U21917 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18815), .ZN(
        P3_U3015) );
  AND2_X1 U21918 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18815), .ZN(
        P3_U3016) );
  AND2_X1 U21919 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18815), .ZN(
        P3_U3017) );
  AND2_X1 U21920 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18815), .ZN(
        P3_U3018) );
  AND2_X1 U21921 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18815), .ZN(
        P3_U3019) );
  AND2_X1 U21922 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18815), .ZN(
        P3_U3020) );
  AND2_X1 U21923 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18815), .ZN(P3_U3021) );
  AND2_X1 U21924 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18815), .ZN(P3_U3022) );
  AND2_X1 U21925 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18815), .ZN(P3_U3023) );
  AND2_X1 U21926 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18904), .ZN(P3_U3024) );
  AND2_X1 U21927 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18904), .ZN(P3_U3025) );
  AND2_X1 U21928 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18904), .ZN(P3_U3026) );
  AND2_X1 U21929 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18904), .ZN(P3_U3027) );
  AND2_X1 U21930 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18904), .ZN(P3_U3028) );
  NOR2_X1 U21931 ( .A1(n18962), .A2(n18818), .ZN(n18824) );
  OAI21_X1 U21932 ( .B1(n18816), .B2(n20902), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18817) );
  AOI22_X1 U21933 ( .A1(n18824), .A2(n18833), .B1(n18970), .B2(n18817), .ZN(
        n18819) );
  NAND3_X1 U21934 ( .A1(NA), .A2(n18830), .A3(n18818), .ZN(n18825) );
  OAI211_X1 U21935 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18819), .B(n18825), .ZN(P3_U3029) );
  NOR2_X1 U21936 ( .A1(n18833), .A2(n20902), .ZN(n18828) );
  INV_X1 U21937 ( .A(n18828), .ZN(n18821) );
  AOI22_X1 U21938 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18821), .B1(HOLD), 
        .B2(n18820), .ZN(n18823) );
  INV_X1 U21939 ( .A(n18824), .ZN(n18826) );
  INV_X1 U21940 ( .A(n18822), .ZN(n18959) );
  OAI211_X1 U21941 ( .C1(n18823), .C2(n18830), .A(n18826), .B(n18959), .ZN(
        P3_U3030) );
  AOI21_X1 U21942 ( .B1(n18830), .B2(n18825), .A(n18824), .ZN(n18831) );
  OAI22_X1 U21943 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18826), .ZN(n18827) );
  OAI22_X1 U21944 ( .A1(n18828), .A2(n18827), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18829) );
  OAI22_X1 U21945 ( .A1(n18831), .A2(n18833), .B1(n18830), .B2(n18829), .ZN(
        P3_U3031) );
  NAND2_X1 U21946 ( .A1(n18972), .A2(n18833), .ZN(n18886) );
  CLKBUF_X1 U21947 ( .A(n18886), .Z(n18891) );
  OAI222_X1 U21948 ( .A1(n18942), .A2(n18895), .B1(n18834), .B2(n18972), .C1(
        n18835), .C2(n18891), .ZN(P3_U3032) );
  OAI222_X1 U21949 ( .A1(n18891), .A2(n18837), .B1(n18836), .B2(n18972), .C1(
        n18835), .C2(n18895), .ZN(P3_U3033) );
  OAI222_X1 U21950 ( .A1(n18891), .A2(n18839), .B1(n18838), .B2(n18972), .C1(
        n18837), .C2(n18895), .ZN(P3_U3034) );
  OAI222_X1 U21951 ( .A1(n18891), .A2(n18841), .B1(n18840), .B2(n18972), .C1(
        n18839), .C2(n18895), .ZN(P3_U3035) );
  OAI222_X1 U21952 ( .A1(n18891), .A2(n18843), .B1(n18842), .B2(n18972), .C1(
        n18841), .C2(n18895), .ZN(P3_U3036) );
  OAI222_X1 U21953 ( .A1(n18891), .A2(n18845), .B1(n18844), .B2(n18972), .C1(
        n18843), .C2(n18895), .ZN(P3_U3037) );
  OAI222_X1 U21954 ( .A1(n18891), .A2(n18848), .B1(n18846), .B2(n18972), .C1(
        n18845), .C2(n18895), .ZN(P3_U3038) );
  OAI222_X1 U21955 ( .A1(n18848), .A2(n18895), .B1(n18847), .B2(n18972), .C1(
        n18849), .C2(n18891), .ZN(P3_U3039) );
  OAI222_X1 U21956 ( .A1(n18891), .A2(n18851), .B1(n18850), .B2(n18972), .C1(
        n18849), .C2(n18895), .ZN(P3_U3040) );
  OAI222_X1 U21957 ( .A1(n18891), .A2(n18853), .B1(n18852), .B2(n18972), .C1(
        n18851), .C2(n18895), .ZN(P3_U3041) );
  OAI222_X1 U21958 ( .A1(n18891), .A2(n18855), .B1(n18854), .B2(n18972), .C1(
        n18853), .C2(n18895), .ZN(P3_U3042) );
  OAI222_X1 U21959 ( .A1(n18891), .A2(n21048), .B1(n18856), .B2(n18972), .C1(
        n18855), .C2(n18895), .ZN(P3_U3043) );
  OAI222_X1 U21960 ( .A1(n21048), .A2(n18895), .B1(n18857), .B2(n18972), .C1(
        n18859), .C2(n18891), .ZN(P3_U3044) );
  OAI222_X1 U21961 ( .A1(n18859), .A2(n18895), .B1(n18858), .B2(n18972), .C1(
        n18860), .C2(n18891), .ZN(P3_U3045) );
  INV_X1 U21962 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18862) );
  OAI222_X1 U21963 ( .A1(n18886), .A2(n18862), .B1(n18861), .B2(n18972), .C1(
        n18860), .C2(n18895), .ZN(P3_U3046) );
  OAI222_X1 U21964 ( .A1(n18886), .A2(n18865), .B1(n18863), .B2(n18972), .C1(
        n18862), .C2(n18895), .ZN(P3_U3047) );
  OAI222_X1 U21965 ( .A1(n18865), .A2(n18895), .B1(n18864), .B2(n18972), .C1(
        n18866), .C2(n18891), .ZN(P3_U3048) );
  OAI222_X1 U21966 ( .A1(n18886), .A2(n18868), .B1(n18867), .B2(n18972), .C1(
        n18866), .C2(n18895), .ZN(P3_U3049) );
  OAI222_X1 U21967 ( .A1(n18886), .A2(n18871), .B1(n18869), .B2(n18972), .C1(
        n18868), .C2(n18895), .ZN(P3_U3050) );
  OAI222_X1 U21968 ( .A1(n18871), .A2(n18895), .B1(n18870), .B2(n18972), .C1(
        n18872), .C2(n18891), .ZN(P3_U3051) );
  OAI222_X1 U21969 ( .A1(n18886), .A2(n18874), .B1(n18873), .B2(n18972), .C1(
        n18872), .C2(n18895), .ZN(P3_U3052) );
  OAI222_X1 U21970 ( .A1(n18886), .A2(n18876), .B1(n18875), .B2(n18972), .C1(
        n18874), .C2(n18895), .ZN(P3_U3053) );
  OAI222_X1 U21971 ( .A1(n18886), .A2(n18878), .B1(n18877), .B2(n18972), .C1(
        n18876), .C2(n18895), .ZN(P3_U3054) );
  OAI222_X1 U21972 ( .A1(n18886), .A2(n18880), .B1(n18879), .B2(n18972), .C1(
        n18878), .C2(n18895), .ZN(P3_U3055) );
  OAI222_X1 U21973 ( .A1(n18891), .A2(n18882), .B1(n18881), .B2(n18972), .C1(
        n18880), .C2(n18895), .ZN(P3_U3056) );
  OAI222_X1 U21974 ( .A1(n18891), .A2(n18884), .B1(n18883), .B2(n18972), .C1(
        n18882), .C2(n18895), .ZN(P3_U3057) );
  INV_X1 U21975 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18888) );
  OAI222_X1 U21976 ( .A1(n18886), .A2(n18888), .B1(n18885), .B2(n18972), .C1(
        n18884), .C2(n18895), .ZN(P3_U3058) );
  OAI222_X1 U21977 ( .A1(n18888), .A2(n18895), .B1(n18887), .B2(n18972), .C1(
        n18889), .C2(n18891), .ZN(P3_U3059) );
  OAI222_X1 U21978 ( .A1(n18891), .A2(n18894), .B1(n18890), .B2(n18972), .C1(
        n18889), .C2(n18895), .ZN(P3_U3060) );
  OAI222_X1 U21979 ( .A1(n18895), .A2(n18894), .B1(n18893), .B2(n18972), .C1(
        n18892), .C2(n18891), .ZN(P3_U3061) );
  INV_X1 U21980 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18896) );
  AOI22_X1 U21981 ( .A1(n18972), .A2(n18897), .B1(n18896), .B2(n18970), .ZN(
        P3_U3274) );
  INV_X1 U21982 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18944) );
  INV_X1 U21983 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18898) );
  AOI22_X1 U21984 ( .A1(n18972), .A2(n18944), .B1(n18898), .B2(n18970), .ZN(
        P3_U3275) );
  INV_X1 U21985 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18899) );
  AOI22_X1 U21986 ( .A1(n18972), .A2(n18900), .B1(n18899), .B2(n18970), .ZN(
        P3_U3276) );
  INV_X1 U21987 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18950) );
  INV_X1 U21988 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18901) );
  AOI22_X1 U21989 ( .A1(n18972), .A2(n18950), .B1(n18901), .B2(n18970), .ZN(
        P3_U3277) );
  INV_X1 U21990 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18903) );
  INV_X1 U21991 ( .A(n18905), .ZN(n18902) );
  AOI21_X1 U21992 ( .B1(n18904), .B2(n18903), .A(n18902), .ZN(P3_U3280) );
  OAI21_X1 U21993 ( .B1(n18907), .B2(n18906), .A(n18905), .ZN(P3_U3281) );
  NOR2_X1 U21994 ( .A1(n18908), .A2(n20997), .ZN(n18911) );
  OAI21_X1 U21995 ( .B1(n18911), .B2(n18910), .A(n18909), .ZN(P3_U3282) );
  INV_X1 U21996 ( .A(n18912), .ZN(n18916) );
  NOR2_X1 U21997 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18913), .ZN(
        n18915) );
  AOI22_X1 U21998 ( .A1(n18936), .A2(n18916), .B1(n18915), .B2(n18914), .ZN(
        n18920) );
  AOI21_X1 U21999 ( .B1(n18974), .B2(n18917), .A(n18941), .ZN(n18919) );
  OAI22_X1 U22000 ( .A1(n18941), .A2(n18920), .B1(n18919), .B2(n18918), .ZN(
        P3_U3285) );
  NOR2_X1 U22001 ( .A1(n18921), .A2(n18938), .ZN(n18929) );
  INV_X1 U22002 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18922) );
  AOI22_X1 U22003 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18923), .B2(n18922), .ZN(
        n18928) );
  AOI222_X1 U22004 ( .A1(n18925), .A2(n18974), .B1(n18929), .B2(n18928), .C1(
        n18936), .C2(n18924), .ZN(n18926) );
  AOI22_X1 U22005 ( .A1(n18941), .A2(n11534), .B1(n18926), .B2(n18939), .ZN(
        P3_U3288) );
  INV_X1 U22006 ( .A(n18927), .ZN(n18932) );
  INV_X1 U22007 ( .A(n18928), .ZN(n18930) );
  AOI222_X1 U22008 ( .A1(n18932), .A2(n18974), .B1(n18936), .B2(n18931), .C1(
        n18930), .C2(n18929), .ZN(n18933) );
  AOI22_X1 U22009 ( .A1(n18941), .A2(n18934), .B1(n18933), .B2(n18939), .ZN(
        P3_U3289) );
  INV_X1 U22010 ( .A(n18935), .ZN(n18937) );
  AOI222_X1 U22011 ( .A1(n18938), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18974), 
        .B2(n18937), .C1(n16981), .C2(n18936), .ZN(n18940) );
  AOI22_X1 U22012 ( .A1(n18941), .A2(n16981), .B1(n18940), .B2(n18939), .ZN(
        P3_U3290) );
  AOI21_X1 U22013 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18943) );
  AOI22_X1 U22014 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18943), .B2(n18942), .ZN(n18945) );
  AOI22_X1 U22015 ( .A1(n18946), .A2(n18945), .B1(n18944), .B2(n18949), .ZN(
        P3_U3292) );
  NOR2_X1 U22016 ( .A1(n18949), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18947) );
  AOI22_X1 U22017 ( .A1(n18950), .A2(n18949), .B1(n18948), .B2(n18947), .ZN(
        P3_U3293) );
  INV_X1 U22018 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18951) );
  AOI22_X1 U22019 ( .A1(n18972), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18951), 
        .B2(n18970), .ZN(P3_U3294) );
  NAND2_X1 U22020 ( .A1(n18954), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18952) );
  OAI21_X1 U22021 ( .B1(n18954), .B2(n18953), .A(n18952), .ZN(P3_U3295) );
  OAI22_X1 U22022 ( .A1(n18957), .A2(n18956), .B1(n18955), .B2(n20992), .ZN(
        n18958) );
  NOR2_X1 U22023 ( .A1(n18976), .A2(n18958), .ZN(n18969) );
  AOI21_X1 U22024 ( .B1(n18961), .B2(n18960), .A(n18959), .ZN(n18963) );
  OAI211_X1 U22025 ( .C1(n18964), .C2(n18963), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18962), .ZN(n18966) );
  AOI21_X1 U22026 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18966), .A(n18965), 
        .ZN(n18968) );
  NAND2_X1 U22027 ( .A1(n18969), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18967) );
  OAI21_X1 U22028 ( .B1(n18969), .B2(n18968), .A(n18967), .ZN(P3_U3296) );
  INV_X1 U22029 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18979) );
  INV_X1 U22030 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18971) );
  AOI22_X1 U22031 ( .A1(n18972), .A2(n18979), .B1(n18971), .B2(n18970), .ZN(
        P3_U3297) );
  AOI21_X1 U22032 ( .B1(n18974), .B2(n18973), .A(n18976), .ZN(n18980) );
  INV_X1 U22033 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18977) );
  AOI22_X1 U22034 ( .A1(n18980), .A2(n18977), .B1(n18976), .B2(n18975), .ZN(
        P3_U3298) );
  AOI21_X1 U22035 ( .B1(n18980), .B2(n18979), .A(n18978), .ZN(P3_U3299) );
  INV_X1 U22036 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18981) );
  INV_X1 U22037 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19884) );
  NAND2_X1 U22038 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19884), .ZN(n19877) );
  OR2_X1 U22039 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19873) );
  OAI21_X1 U22040 ( .B1(n19872), .B2(n19877), .A(n19873), .ZN(n19936) );
  INV_X1 U22041 ( .A(n19936), .ZN(n19866) );
  OAI21_X1 U22042 ( .B1(n19872), .B2(n18981), .A(n19866), .ZN(P2_U2815) );
  AOI22_X1 U22043 ( .A1(n20003), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19941), 
        .B2(n18982), .ZN(n18983) );
  INV_X1 U22044 ( .A(n18983), .ZN(P2_U2816) );
  AOI21_X1 U22045 ( .B1(n19872), .B2(n19884), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18984) );
  AOI22_X1 U22046 ( .A1(n20009), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18984), 
        .B2(n20007), .ZN(P2_U2817) );
  OAI21_X1 U22047 ( .B1(n19868), .B2(BS16), .A(n19936), .ZN(n19934) );
  OAI21_X1 U22048 ( .B1(n19936), .B2(n19781), .A(n19934), .ZN(P2_U2818) );
  NOR2_X1 U22049 ( .A1(n18986), .A2(n18985), .ZN(n19979) );
  OAI21_X1 U22050 ( .B1(n19979), .B2(n18988), .A(n18987), .ZN(P2_U2819) );
  NOR4_X1 U22051 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18992) );
  NOR4_X1 U22052 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18991) );
  NOR4_X1 U22053 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18990) );
  NOR4_X1 U22054 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18989) );
  NAND4_X1 U22055 ( .A1(n18992), .A2(n18991), .A3(n18990), .A4(n18989), .ZN(
        n18998) );
  NOR4_X1 U22056 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18996) );
  AOI211_X1 U22057 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_4__SCAN_IN), .B(
        P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(n18995) );
  NOR4_X1 U22058 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18994) );
  NOR4_X1 U22059 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18993) );
  NAND4_X1 U22060 ( .A1(n18996), .A2(n18995), .A3(n18994), .A4(n18993), .ZN(
        n18997) );
  NOR2_X1 U22061 ( .A1(n18998), .A2(n18997), .ZN(n19005) );
  INV_X1 U22062 ( .A(n19005), .ZN(n19004) );
  NOR2_X1 U22063 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19004), .ZN(n18999) );
  INV_X1 U22064 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U22065 ( .A1(n18999), .A2(n10421), .B1(n19004), .B2(n19932), .ZN(
        P2_U2820) );
  OR3_X1 U22066 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19003) );
  INV_X1 U22067 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19930) );
  AOI22_X1 U22068 ( .A1(n18999), .A2(n19003), .B1(n19004), .B2(n19930), .ZN(
        P2_U2821) );
  INV_X1 U22069 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19935) );
  NAND2_X1 U22070 ( .A1(n18999), .A2(n19935), .ZN(n19002) );
  OAI21_X1 U22071 ( .B1(n10439), .B2(n10421), .A(n19005), .ZN(n19000) );
  OAI21_X1 U22072 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19005), .A(n19000), 
        .ZN(n19001) );
  OAI221_X1 U22073 ( .B1(n19002), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19002), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19001), .ZN(P2_U2822) );
  INV_X1 U22074 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19928) );
  OAI221_X1 U22075 ( .B1(n19005), .B2(n19928), .C1(n19004), .C2(n19003), .A(
        n19002), .ZN(P2_U2823) );
  INV_X1 U22076 ( .A(n19006), .ZN(n19008) );
  AOI22_X1 U22077 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19167), .ZN(n19007) );
  OAI21_X1 U22078 ( .B1(n19008), .B2(n19201), .A(n19007), .ZN(n19012) );
  OAI22_X1 U22079 ( .A1(n19010), .A2(n19209), .B1(n15571), .B2(n19203), .ZN(
        n19011) );
  AOI211_X1 U22080 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n19207), .A(n19012), .B(
        n19011), .ZN(n19016) );
  OAI211_X1 U22081 ( .C1(n19014), .C2(n19017), .A(n19174), .B(n19013), .ZN(
        n19015) );
  OAI211_X1 U22082 ( .C1(n19017), .C2(n19091), .A(n19016), .B(n19015), .ZN(
        P2_U2835) );
  NAND2_X1 U22083 ( .A1(n9977), .A2(n19018), .ZN(n19019) );
  XOR2_X1 U22084 ( .A(n19020), .B(n19019), .Z(n19028) );
  OAI21_X1 U22085 ( .B1(n19906), .B2(n19204), .A(n19151), .ZN(n19024) );
  OAI22_X1 U22086 ( .A1(n19022), .A2(n19201), .B1(n19021), .B2(n19178), .ZN(
        n19023) );
  AOI211_X1 U22087 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19207), .A(n19024), .B(
        n19023), .ZN(n19027) );
  AOI22_X1 U22088 ( .A1(n19025), .A2(n19172), .B1(n10207), .B2(n19182), .ZN(
        n19026) );
  OAI211_X1 U22089 ( .C1(n19216), .C2(n19028), .A(n19027), .B(n19026), .ZN(
        P2_U2836) );
  AOI22_X1 U22090 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19207), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19213), .ZN(n19029) );
  OAI21_X1 U22091 ( .B1(n19030), .B2(n19201), .A(n19029), .ZN(n19031) );
  AOI211_X1 U22092 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19167), .A(n11352), 
        .B(n19031), .ZN(n19037) );
  NOR2_X1 U22093 ( .A1(n19192), .A2(n19039), .ZN(n19033) );
  XNOR2_X1 U22094 ( .A(n19033), .B(n19032), .ZN(n19034) );
  AOI22_X1 U22095 ( .A1(n19035), .A2(n19172), .B1(n19174), .B2(n19034), .ZN(
        n19036) );
  OAI211_X1 U22096 ( .C1(n19038), .C2(n19203), .A(n19037), .B(n19036), .ZN(
        P2_U2837) );
  AOI211_X1 U22097 ( .C1(n19041), .C2(n19040), .A(n19039), .B(n9883), .ZN(
        n19045) );
  AOI22_X1 U22098 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19167), .ZN(n19042) );
  OAI211_X1 U22099 ( .C1(n19043), .C2(n19201), .A(n19042), .B(n19151), .ZN(
        n19044) );
  AOI211_X1 U22100 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19207), .A(n19045), .B(
        n19044), .ZN(n19049) );
  AOI22_X1 U22101 ( .A1(n19047), .A2(n19182), .B1(n19046), .B2(n19172), .ZN(
        n19048) );
  OAI211_X1 U22102 ( .C1(n19050), .C2(n19091), .A(n19049), .B(n19048), .ZN(
        P2_U2838) );
  OAI22_X1 U22103 ( .A1(n19052), .A2(n19201), .B1(n19188), .B2(n19051), .ZN(
        n19053) );
  INV_X1 U22104 ( .A(n19053), .ZN(n19054) );
  OAI211_X1 U22105 ( .C1(n10870), .C2(n19204), .A(n19054), .B(n19151), .ZN(
        n19055) );
  AOI21_X1 U22106 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19213), .A(
        n19055), .ZN(n19062) );
  INV_X1 U22107 ( .A(n19056), .ZN(n19224) );
  NOR2_X1 U22108 ( .A1(n19192), .A2(n19057), .ZN(n19059) );
  XNOR2_X1 U22109 ( .A(n19059), .B(n19058), .ZN(n19060) );
  AOI22_X1 U22110 ( .A1(n19224), .A2(n19182), .B1(n19174), .B2(n19060), .ZN(
        n19061) );
  OAI211_X1 U22111 ( .C1(n19063), .C2(n19209), .A(n19062), .B(n19061), .ZN(
        P2_U2839) );
  NAND2_X1 U22112 ( .A1(n9977), .A2(n19064), .ZN(n19066) );
  XOR2_X1 U22113 ( .A(n19066), .B(n19065), .Z(n19074) );
  AOI22_X1 U22114 ( .A1(n19067), .A2(n19185), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19213), .ZN(n19068) );
  OAI211_X1 U22115 ( .C1(n19899), .C2(n19204), .A(n19068), .B(n19151), .ZN(
        n19072) );
  OAI22_X1 U22116 ( .A1(n19070), .A2(n19209), .B1(n19069), .B2(n19203), .ZN(
        n19071) );
  AOI211_X1 U22117 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19207), .A(n19072), .B(
        n19071), .ZN(n19073) );
  OAI21_X1 U22118 ( .B1(n19074), .B2(n19216), .A(n19073), .ZN(P2_U2840) );
  NOR2_X1 U22119 ( .A1(n19192), .A2(n19084), .ZN(n19076) );
  XOR2_X1 U22120 ( .A(n19076), .B(n19075), .Z(n19083) );
  AOI22_X1 U22121 ( .A1(n19077), .A2(n19185), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19207), .ZN(n19078) );
  OAI211_X1 U22122 ( .C1(n10855), .C2(n19204), .A(n19078), .B(n19151), .ZN(
        n19079) );
  AOI21_X1 U22123 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19213), .A(
        n19079), .ZN(n19082) );
  AOI22_X1 U22124 ( .A1(n19080), .A2(n19172), .B1(n19231), .B2(n19182), .ZN(
        n19081) );
  OAI211_X1 U22125 ( .C1(n19216), .C2(n19083), .A(n19082), .B(n19081), .ZN(
        P2_U2841) );
  AOI211_X1 U22126 ( .C1(n19093), .C2(n19085), .A(n19084), .B(n9883), .ZN(
        n19090) );
  INV_X1 U22127 ( .A(n19086), .ZN(n19088) );
  AOI22_X1 U22128 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19213), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19167), .ZN(n19087) );
  OAI211_X1 U22129 ( .C1(n19088), .C2(n19201), .A(n19087), .B(n19151), .ZN(
        n19089) );
  AOI211_X1 U22130 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n19207), .A(n19090), .B(
        n19089), .ZN(n19096) );
  INV_X1 U22131 ( .A(n19091), .ZN(n19092) );
  AOI22_X1 U22132 ( .A1(n19094), .A2(n19172), .B1(n19093), .B2(n19092), .ZN(
        n19095) );
  OAI211_X1 U22133 ( .C1(n19097), .C2(n19203), .A(n19096), .B(n19095), .ZN(
        P2_U2842) );
  INV_X1 U22134 ( .A(n19098), .ZN(n19100) );
  AOI22_X1 U22135 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n19207), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19213), .ZN(n19099) );
  OAI21_X1 U22136 ( .B1(n19100), .B2(n19201), .A(n19099), .ZN(n19101) );
  AOI211_X1 U22137 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19167), .A(n11352), 
        .B(n19101), .ZN(n19107) );
  NOR2_X1 U22138 ( .A1(n19192), .A2(n19102), .ZN(n19104) );
  XNOR2_X1 U22139 ( .A(n19104), .B(n19103), .ZN(n19105) );
  AOI22_X1 U22140 ( .A1(n19234), .A2(n19182), .B1(n19174), .B2(n19105), .ZN(
        n19106) );
  OAI211_X1 U22141 ( .C1(n19108), .C2(n19209), .A(n19107), .B(n19106), .ZN(
        P2_U2843) );
  AOI22_X1 U22142 ( .A1(n19109), .A2(n19185), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19213), .ZN(n19110) );
  OAI21_X1 U22143 ( .B1(n19188), .B2(n19111), .A(n19110), .ZN(n19112) );
  AOI211_X1 U22144 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19167), .A(n11352), 
        .B(n19112), .ZN(n19118) );
  NOR2_X1 U22145 ( .A1(n19192), .A2(n19113), .ZN(n19115) );
  XNOR2_X1 U22146 ( .A(n19115), .B(n19114), .ZN(n19116) );
  AOI22_X1 U22147 ( .A1(n19237), .A2(n19182), .B1(n19174), .B2(n19116), .ZN(
        n19117) );
  OAI211_X1 U22148 ( .C1(n19119), .C2(n19209), .A(n19118), .B(n19117), .ZN(
        P2_U2845) );
  OAI21_X1 U22149 ( .B1(n15464), .B2(n19204), .A(n19151), .ZN(n19122) );
  OAI22_X1 U22150 ( .A1(n19120), .A2(n19201), .B1(n10917), .B2(n19188), .ZN(
        n19121) );
  AOI211_X1 U22151 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19213), .A(
        n19122), .B(n19121), .ZN(n19129) );
  NAND2_X1 U22152 ( .A1(n9977), .A2(n19123), .ZN(n19124) );
  XNOR2_X1 U22153 ( .A(n19125), .B(n19124), .ZN(n19126) );
  AOI22_X1 U22154 ( .A1(n19127), .A2(n19172), .B1(n19174), .B2(n19126), .ZN(
        n19128) );
  OAI211_X1 U22155 ( .C1(n19242), .C2(n19203), .A(n19129), .B(n19128), .ZN(
        P2_U2846) );
  AOI22_X1 U22156 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19207), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19213), .ZN(n19130) );
  OAI21_X1 U22157 ( .B1(n19131), .B2(n19201), .A(n19130), .ZN(n19132) );
  AOI211_X1 U22158 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19167), .A(n11352), .B(
        n19132), .ZN(n19138) );
  NOR2_X1 U22159 ( .A1(n19192), .A2(n19133), .ZN(n19135) );
  XNOR2_X1 U22160 ( .A(n19135), .B(n19134), .ZN(n19136) );
  AOI22_X1 U22161 ( .A1(n19246), .A2(n19182), .B1(n19174), .B2(n19136), .ZN(
        n19137) );
  OAI211_X1 U22162 ( .C1(n19139), .C2(n19209), .A(n19138), .B(n19137), .ZN(
        P2_U2847) );
  NAND2_X1 U22163 ( .A1(n9977), .A2(n19140), .ZN(n19142) );
  XOR2_X1 U22164 ( .A(n19142), .B(n19141), .Z(n19150) );
  AOI22_X1 U22165 ( .A1(n19143), .A2(n19185), .B1(n19213), .B2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19144) );
  OAI211_X1 U22166 ( .C1(n10477), .C2(n19204), .A(n19144), .B(n19151), .ZN(
        n19148) );
  OAI22_X1 U22167 ( .A1(n19203), .A2(n19146), .B1(n19209), .B2(n19145), .ZN(
        n19147) );
  AOI211_X1 U22168 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19207), .A(n19148), .B(
        n19147), .ZN(n19149) );
  OAI21_X1 U22169 ( .B1(n19150), .B2(n19216), .A(n19149), .ZN(P2_U2848) );
  OAI21_X1 U22170 ( .B1(n10473), .B2(n19204), .A(n19151), .ZN(n19155) );
  INV_X1 U22171 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19152) );
  OAI22_X1 U22172 ( .A1(n19153), .A2(n19201), .B1(n19188), .B2(n19152), .ZN(
        n19154) );
  AOI211_X1 U22173 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19213), .A(
        n19155), .B(n19154), .ZN(n19162) );
  NOR2_X1 U22174 ( .A1(n19192), .A2(n19156), .ZN(n19158) );
  XNOR2_X1 U22175 ( .A(n19158), .B(n19157), .ZN(n19160) );
  AOI22_X1 U22176 ( .A1(n19174), .A2(n19160), .B1(n19172), .B2(n19159), .ZN(
        n19161) );
  OAI211_X1 U22177 ( .C1(n19203), .C2(n19163), .A(n19162), .B(n19161), .ZN(
        P2_U2849) );
  AOI22_X1 U22178 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n19207), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19213), .ZN(n19164) );
  OAI21_X1 U22179 ( .B1(n19165), .B2(n19201), .A(n19164), .ZN(n19166) );
  AOI211_X1 U22180 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19167), .A(n11352), .B(
        n19166), .ZN(n19176) );
  NAND2_X1 U22181 ( .A1(n9977), .A2(n19168), .ZN(n19169) );
  XNOR2_X1 U22182 ( .A(n19170), .B(n19169), .ZN(n19173) );
  AOI22_X1 U22183 ( .A1(n19174), .A2(n19173), .B1(n19172), .B2(n19171), .ZN(
        n19175) );
  OAI211_X1 U22184 ( .C1(n19203), .C2(n19177), .A(n19176), .B(n19175), .ZN(
        P2_U2850) );
  OAI21_X1 U22185 ( .B1(n19179), .B2(n19178), .A(n19151), .ZN(n19181) );
  NOR2_X1 U22186 ( .A1(n19204), .A2(n10694), .ZN(n19180) );
  AOI211_X1 U22187 ( .C1(n19183), .C2(n19182), .A(n19181), .B(n19180), .ZN(
        n19187) );
  NAND2_X1 U22188 ( .A1(n19185), .A2(n19184), .ZN(n19186) );
  OAI211_X1 U22189 ( .C1(n21133), .C2(n19188), .A(n19187), .B(n19186), .ZN(
        n19189) );
  AOI21_X1 U22190 ( .B1(n19190), .B2(n19211), .A(n19189), .ZN(n19197) );
  INV_X1 U22191 ( .A(n19293), .ZN(n19195) );
  NOR2_X1 U22192 ( .A1(n19192), .A2(n19191), .ZN(n19194) );
  AOI21_X1 U22193 ( .B1(n19195), .B2(n19194), .A(n19216), .ZN(n19193) );
  OAI21_X1 U22194 ( .B1(n19195), .B2(n19194), .A(n19193), .ZN(n19196) );
  OAI211_X1 U22195 ( .C1(n19288), .C2(n19209), .A(n19197), .B(n19196), .ZN(
        P2_U2851) );
  INV_X1 U22196 ( .A(n19199), .ZN(n19200) );
  OAI22_X1 U22197 ( .A1(n19203), .A2(n19202), .B1(n19201), .B2(n19200), .ZN(
        n19206) );
  NOR2_X1 U22198 ( .A1(n19204), .A2(n10421), .ZN(n19205) );
  AOI211_X1 U22199 ( .C1(P2_EBX_REG_0__SCAN_IN), .C2(n19207), .A(n19206), .B(
        n19205), .ZN(n19208) );
  OAI21_X1 U22200 ( .B1(n10072), .B2(n19209), .A(n19208), .ZN(n19210) );
  AOI21_X1 U22201 ( .B1(n19212), .B2(n19211), .A(n19210), .ZN(n19215) );
  NAND2_X1 U22202 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19213), .ZN(
        n19214) );
  OAI211_X1 U22203 ( .C1(n14260), .C2(n19216), .A(n19215), .B(n19214), .ZN(
        P2_U2855) );
  AOI22_X1 U22204 ( .A1(n19217), .A2(n13389), .B1(n19222), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U22205 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19239), .B1(n19223), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19218) );
  NAND2_X1 U22206 ( .A1(n19219), .A2(n19218), .ZN(P2_U2888) );
  AOI22_X1 U22207 ( .A1(n19221), .A2(n19220), .B1(n19239), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19229) );
  AOI22_X1 U22208 ( .A1(n19223), .A2(BUF1_REG_16__SCAN_IN), .B1(n19222), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19228) );
  AOI22_X1 U22209 ( .A1(n19226), .A2(n19225), .B1(n13389), .B2(n19224), .ZN(
        n19227) );
  NAND3_X1 U22210 ( .A1(n19229), .A2(n19228), .A3(n19227), .ZN(P2_U2903) );
  INV_X1 U22211 ( .A(n19243), .ZN(n19247) );
  AOI22_X1 U22212 ( .A1(n19247), .A2(n19231), .B1(n19245), .B2(n19230), .ZN(
        n19232) );
  OAI21_X1 U22213 ( .B1(n19249), .B2(n19253), .A(n19232), .ZN(P2_U2905) );
  AOI22_X1 U22214 ( .A1(n19247), .A2(n19234), .B1(n19245), .B2(n19233), .ZN(
        n19235) );
  OAI21_X1 U22215 ( .B1(n19249), .B2(n19257), .A(n19235), .ZN(P2_U2907) );
  AOI22_X1 U22216 ( .A1(n19237), .A2(n19247), .B1(n19245), .B2(n19236), .ZN(
        n19238) );
  OAI21_X1 U22217 ( .B1(n19249), .B2(n19261), .A(n19238), .ZN(P2_U2909) );
  AOI22_X1 U22218 ( .A1(n19245), .A2(n19240), .B1(n19239), .B2(
        P2_EAX_REG_9__SCAN_IN), .ZN(n19241) );
  OAI21_X1 U22219 ( .B1(n19243), .B2(n19242), .A(n19241), .ZN(P2_U2910) );
  AOI22_X1 U22220 ( .A1(n19247), .A2(n19246), .B1(n19245), .B2(n19244), .ZN(
        n19248) );
  OAI21_X1 U22221 ( .B1(n19249), .B2(n19265), .A(n19248), .ZN(P2_U2911) );
  AND2_X1 U22222 ( .A1(n19271), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22223 ( .A1(n19280), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19251) );
  OAI21_X1 U22224 ( .B1(n13526), .B2(n19282), .A(n19251), .ZN(P2_U2936) );
  AOI22_X1 U22225 ( .A1(n19280), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19252) );
  OAI21_X1 U22226 ( .B1(n19253), .B2(n19282), .A(n19252), .ZN(P2_U2937) );
  AOI22_X1 U22227 ( .A1(n19280), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19254) );
  OAI21_X1 U22228 ( .B1(n19255), .B2(n19282), .A(n19254), .ZN(P2_U2938) );
  AOI22_X1 U22229 ( .A1(n20002), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19256) );
  OAI21_X1 U22230 ( .B1(n19257), .B2(n19282), .A(n19256), .ZN(P2_U2939) );
  AOI22_X1 U22231 ( .A1(n20002), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19258) );
  OAI21_X1 U22232 ( .B1(n19259), .B2(n19282), .A(n19258), .ZN(P2_U2940) );
  AOI22_X1 U22233 ( .A1(n20002), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19260) );
  OAI21_X1 U22234 ( .B1(n19261), .B2(n19282), .A(n19260), .ZN(P2_U2941) );
  AOI22_X1 U22235 ( .A1(n20002), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19262) );
  OAI21_X1 U22236 ( .B1(n19263), .B2(n19282), .A(n19262), .ZN(P2_U2942) );
  AOI22_X1 U22237 ( .A1(n20002), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19264) );
  OAI21_X1 U22238 ( .B1(n19265), .B2(n19282), .A(n19264), .ZN(P2_U2943) );
  AOI22_X1 U22239 ( .A1(n20002), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19266) );
  OAI21_X1 U22240 ( .B1(n19267), .B2(n19282), .A(n19266), .ZN(P2_U2944) );
  AOI22_X1 U22241 ( .A1(n19280), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19268) );
  OAI21_X1 U22242 ( .B1(n19269), .B2(n19282), .A(n19268), .ZN(P2_U2945) );
  AOI22_X1 U22243 ( .A1(n19280), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19270) );
  OAI21_X1 U22244 ( .B1(n13919), .B2(n19282), .A(n19270), .ZN(P2_U2946) );
  AOI22_X1 U22245 ( .A1(n19280), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19271), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19272) );
  OAI21_X1 U22246 ( .B1(n13576), .B2(n19282), .A(n19272), .ZN(P2_U2947) );
  INV_X1 U22247 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19274) );
  AOI22_X1 U22248 ( .A1(n19280), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19273) );
  OAI21_X1 U22249 ( .B1(n19274), .B2(n19282), .A(n19273), .ZN(P2_U2948) );
  INV_X1 U22250 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19276) );
  AOI22_X1 U22251 ( .A1(n19280), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19275) );
  OAI21_X1 U22252 ( .B1(n19276), .B2(n19282), .A(n19275), .ZN(P2_U2949) );
  INV_X1 U22253 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19278) );
  AOI22_X1 U22254 ( .A1(n19280), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19277) );
  OAI21_X1 U22255 ( .B1(n19278), .B2(n19282), .A(n19277), .ZN(P2_U2950) );
  AOI22_X1 U22256 ( .A1(n19280), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19279), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19281) );
  OAI21_X1 U22257 ( .B1(n13529), .B2(n19282), .A(n19281), .ZN(P2_U2951) );
  AOI22_X1 U22258 ( .A1(n19296), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n11352), .ZN(n19292) );
  NAND2_X1 U22259 ( .A1(n19284), .A2(n19283), .ZN(n19287) );
  NAND2_X1 U22260 ( .A1(n19285), .A2(n19300), .ZN(n19286) );
  OAI211_X1 U22261 ( .C1(n19289), .C2(n19288), .A(n19287), .B(n19286), .ZN(
        n19290) );
  INV_X1 U22262 ( .A(n19290), .ZN(n19291) );
  OAI211_X1 U22263 ( .C1(n19294), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        P2_U3010) );
  NOR2_X1 U22264 ( .A1(n19296), .A2(n19295), .ZN(n19310) );
  INV_X1 U22265 ( .A(n19297), .ZN(n19298) );
  AOI21_X1 U22266 ( .B1(n19300), .B2(n19299), .A(n19298), .ZN(n19304) );
  NAND2_X1 U22267 ( .A1(n19302), .A2(n19301), .ZN(n19303) );
  OAI211_X1 U22268 ( .C1(n19306), .C2(n19305), .A(n19304), .B(n19303), .ZN(
        n19307) );
  INV_X1 U22269 ( .A(n19307), .ZN(n19308) );
  OAI21_X1 U22270 ( .B1(n19310), .B2(n19309), .A(n19308), .ZN(P2_U3014) );
  OR2_X1 U22271 ( .A1(n19312), .A2(n19311), .ZN(n19313) );
  AOI22_X1 U22272 ( .A1(n19316), .A2(n19315), .B1(n19314), .B2(n19313), .ZN(
        n19329) );
  NOR2_X1 U22273 ( .A1(n19317), .A2(n13670), .ZN(n19325) );
  NAND2_X1 U22274 ( .A1(n19319), .A2(n19318), .ZN(n19320) );
  OAI211_X1 U22275 ( .C1(n19323), .C2(n19322), .A(n19321), .B(n19320), .ZN(
        n19324) );
  AOI211_X1 U22276 ( .C1(n19327), .C2(n19326), .A(n19325), .B(n19324), .ZN(
        n19328) );
  OAI211_X1 U22277 ( .C1(n19331), .C2(n19330), .A(n19329), .B(n19328), .ZN(
        P2_U3044) );
  NAND2_X1 U22278 ( .A1(n19401), .A2(n19968), .ZN(n19378) );
  NOR2_X1 U22279 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19378), .ZN(
        n19369) );
  AOI22_X1 U22280 ( .A1(n19747), .A2(n19861), .B1(n19779), .B2(n19369), .ZN(
        n19343) );
  INV_X1 U22281 ( .A(n19400), .ZN(n19332) );
  NOR2_X1 U22282 ( .A1(n19861), .A2(n19332), .ZN(n19333) );
  OAI21_X1 U22283 ( .B1(n19333), .B2(n19781), .A(n19942), .ZN(n19341) );
  NOR2_X1 U22284 ( .A1(n19855), .A2(n19369), .ZN(n19340) );
  INV_X1 U22285 ( .A(n19340), .ZN(n19337) );
  INV_X1 U22286 ( .A(n19338), .ZN(n19335) );
  INV_X1 U22287 ( .A(n19369), .ZN(n19334) );
  INV_X1 U22288 ( .A(n19942), .ZN(n19703) );
  OAI211_X1 U22289 ( .C1(n19335), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19334), 
        .B(n19703), .ZN(n19336) );
  OAI211_X1 U22290 ( .C1(n19341), .C2(n19337), .A(n19738), .B(n19336), .ZN(
        n19372) );
  OAI21_X1 U22291 ( .B1(n19338), .B2(n19369), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19339) );
  OAI21_X1 U22292 ( .B1(n19341), .B2(n19340), .A(n19339), .ZN(n19371) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19372), .B1(
        n19790), .B2(n19371), .ZN(n19342) );
  OAI211_X1 U22294 ( .C1(n19710), .C2(n19400), .A(n19343), .B(n19342), .ZN(
        P2_U3048) );
  AOI22_X1 U22295 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19365), .ZN(n19819) );
  AOI22_X1 U22296 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19365), .ZN(n19754) );
  AOI22_X1 U22297 ( .A1(n19816), .A2(n19861), .B1(n19344), .B2(n19369), .ZN(
        n19347) );
  NOR2_X2 U22298 ( .A1(n19345), .A2(n19784), .ZN(n19815) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19372), .B1(
        n19815), .B2(n19371), .ZN(n19346) );
  OAI211_X1 U22300 ( .C1(n19819), .C2(n19400), .A(n19347), .B(n19346), .ZN(
        P2_U3049) );
  AOI22_X1 U22301 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19365), .ZN(n19798) );
  AOI22_X1 U22302 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19365), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19366), .ZN(n19676) );
  NOR2_X2 U22303 ( .A1(n10400), .A2(n19367), .ZN(n19820) );
  AOI22_X1 U22304 ( .A1(n19822), .A2(n19861), .B1(n19820), .B2(n19369), .ZN(
        n19350) );
  NOR2_X2 U22305 ( .A1(n19348), .A2(n19784), .ZN(n19821) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19372), .B1(
        n19821), .B2(n19371), .ZN(n19349) );
  OAI211_X1 U22307 ( .C1(n19798), .C2(n19400), .A(n19350), .B(n19349), .ZN(
        P2_U3050) );
  AOI22_X1 U22308 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19365), .ZN(n19832) );
  AOI22_X1 U22309 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19365), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19366), .ZN(n19679) );
  NOR2_X2 U22310 ( .A1(n10401), .A2(n19367), .ZN(n19827) );
  AOI22_X1 U22311 ( .A1(n19829), .A2(n19861), .B1(n19827), .B2(n19369), .ZN(
        n19354) );
  NOR2_X2 U22312 ( .A1(n19352), .A2(n19784), .ZN(n19828) );
  AOI22_X1 U22313 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19372), .B1(
        n19828), .B2(n19371), .ZN(n19353) );
  OAI211_X1 U22314 ( .C1(n19832), .C2(n19400), .A(n19354), .B(n19353), .ZN(
        P2_U3051) );
  AOI22_X1 U22315 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19365), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19366), .ZN(n19683) );
  NOR2_X2 U22316 ( .A1(n19355), .A2(n19367), .ZN(n19833) );
  AOI22_X1 U22317 ( .A1(n19835), .A2(n19861), .B1(n19833), .B2(n19369), .ZN(
        n19358) );
  NOR2_X2 U22318 ( .A1(n19356), .A2(n19784), .ZN(n19834) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19372), .B1(
        n19834), .B2(n19371), .ZN(n19357) );
  OAI211_X1 U22320 ( .C1(n19839), .C2(n19400), .A(n19358), .B(n19357), .ZN(
        P2_U3052) );
  AOI22_X1 U22321 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19365), .ZN(n19766) );
  AOI22_X1 U22322 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19365), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19366), .ZN(n19845) );
  INV_X1 U22323 ( .A(n19845), .ZN(n19763) );
  NOR2_X2 U22324 ( .A1(n10904), .A2(n19367), .ZN(n19840) );
  AOI22_X1 U22325 ( .A1(n19763), .A2(n19861), .B1(n19840), .B2(n19369), .ZN(
        n19361) );
  NOR2_X2 U22326 ( .A1(n19359), .A2(n19784), .ZN(n19841) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19372), .B1(
        n19841), .B2(n19371), .ZN(n19360) );
  OAI211_X1 U22328 ( .C1(n19766), .C2(n19400), .A(n19361), .B(n19360), .ZN(
        P2_U3053) );
  AOI22_X1 U22329 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19365), .ZN(n19723) );
  AOI22_X1 U22330 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19365), .ZN(n19853) );
  INV_X1 U22331 ( .A(n19853), .ZN(n19767) );
  NOR2_X2 U22332 ( .A1(n13541), .A2(n19367), .ZN(n19846) );
  AOI22_X1 U22333 ( .A1(n19767), .A2(n19861), .B1(n19846), .B2(n19369), .ZN(
        n19364) );
  NOR2_X2 U22334 ( .A1(n19362), .A2(n19784), .ZN(n19847) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19372), .B1(
        n19847), .B2(n19371), .ZN(n19363) );
  OAI211_X1 U22336 ( .C1(n19723), .C2(n19400), .A(n19364), .B(n19363), .ZN(
        P2_U3054) );
  AOI22_X1 U22337 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19365), .ZN(n19777) );
  AOI22_X1 U22338 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19366), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19365), .ZN(n19814) );
  INV_X1 U22339 ( .A(n19814), .ZN(n19858) );
  NOR2_X2 U22340 ( .A1(n19368), .A2(n19367), .ZN(n19854) );
  AOI22_X1 U22341 ( .A1(n19858), .A2(n19861), .B1(n19854), .B2(n19369), .ZN(
        n19374) );
  NOR2_X2 U22342 ( .A1(n19370), .A2(n19784), .ZN(n19856) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19372), .B1(
        n19856), .B2(n19371), .ZN(n19373) );
  OAI211_X1 U22344 ( .C1(n19777), .C2(n19400), .A(n19374), .B(n19373), .ZN(
        P2_U3055) );
  NAND2_X1 U22345 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19968), .ZN(
        n19600) );
  NOR2_X1 U22346 ( .A1(n19600), .A2(n19402), .ZN(n19395) );
  NOR3_X1 U22347 ( .A1(n19375), .A2(n19995), .A3(n19395), .ZN(n19377) );
  AOI211_X2 U22348 ( .C1(n19995), .C2(n19378), .A(n19510), .B(n19377), .ZN(
        n19396) );
  AOI22_X1 U22349 ( .A1(n19396), .A2(n19790), .B1(n19779), .B2(n19395), .ZN(
        n19382) );
  INV_X1 U22350 ( .A(n19538), .ZN(n19376) );
  NAND2_X1 U22351 ( .A1(n19376), .A2(n19599), .ZN(n19379) );
  AOI21_X1 U22352 ( .B1(n19379), .B2(n19378), .A(n19377), .ZN(n19380) );
  OAI211_X1 U22353 ( .C1(n19395), .C2(n20000), .A(n19380), .B(n19738), .ZN(
        n19397) );
  NAND2_X1 U22354 ( .A1(n19599), .A2(n19546), .ZN(n19419) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19780), .ZN(n19381) );
  OAI211_X1 U22356 ( .C1(n19793), .C2(n19400), .A(n19382), .B(n19381), .ZN(
        P2_U3056) );
  AOI22_X1 U22357 ( .A1(n19396), .A2(n19815), .B1(n19344), .B2(n19395), .ZN(
        n19384) );
  INV_X1 U22358 ( .A(n19819), .ZN(n19750) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19750), .ZN(n19383) );
  OAI211_X1 U22360 ( .C1(n19754), .C2(n19400), .A(n19384), .B(n19383), .ZN(
        P2_U3057) );
  AOI22_X1 U22361 ( .A1(n19396), .A2(n19821), .B1(n19820), .B2(n19395), .ZN(
        n19386) );
  INV_X1 U22362 ( .A(n19798), .ZN(n19823) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19823), .ZN(n19385) );
  OAI211_X1 U22364 ( .C1(n19676), .C2(n19400), .A(n19386), .B(n19385), .ZN(
        P2_U3058) );
  AOI22_X1 U22365 ( .A1(n19396), .A2(n19828), .B1(n19827), .B2(n19395), .ZN(
        n19388) );
  INV_X1 U22366 ( .A(n19832), .ZN(n19757) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19757), .ZN(n19387) );
  OAI211_X1 U22368 ( .C1(n19679), .C2(n19400), .A(n19388), .B(n19387), .ZN(
        P2_U3059) );
  AOI22_X1 U22369 ( .A1(n19396), .A2(n19834), .B1(n19833), .B2(n19395), .ZN(
        n19390) );
  INV_X1 U22370 ( .A(n19839), .ZN(n19680) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19680), .ZN(n19389) );
  OAI211_X1 U22372 ( .C1(n19683), .C2(n19400), .A(n19390), .B(n19389), .ZN(
        P2_U3060) );
  AOI22_X1 U22373 ( .A1(n19396), .A2(n19841), .B1(n19840), .B2(n19395), .ZN(
        n19392) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19842), .ZN(n19391) );
  OAI211_X1 U22375 ( .C1(n19845), .C2(n19400), .A(n19392), .B(n19391), .ZN(
        P2_U3061) );
  AOI22_X1 U22376 ( .A1(n19396), .A2(n19847), .B1(n19846), .B2(n19395), .ZN(
        n19394) );
  INV_X1 U22377 ( .A(n19723), .ZN(n19848) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19848), .ZN(n19393) );
  OAI211_X1 U22379 ( .C1(n19853), .C2(n19400), .A(n19394), .B(n19393), .ZN(
        P2_U3062) );
  AOI22_X1 U22380 ( .A1(n19396), .A2(n19856), .B1(n19854), .B2(n19395), .ZN(
        n19399) );
  INV_X1 U22381 ( .A(n19777), .ZN(n19860) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19397), .B1(
        n19428), .B2(n19860), .ZN(n19398) );
  OAI211_X1 U22383 ( .C1(n19814), .C2(n19400), .A(n19399), .B(n19398), .ZN(
        P2_U3063) );
  INV_X1 U22384 ( .A(n11079), .ZN(n19407) );
  NOR2_X1 U22385 ( .A1(n19968), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19632) );
  NAND2_X1 U22386 ( .A1(n19632), .A2(n19401), .ZN(n19406) );
  AOI21_X1 U22387 ( .B1(n19407), .B2(n19406), .A(n19995), .ZN(n19403) );
  NOR2_X1 U22388 ( .A1(n19402), .A2(n19634), .ZN(n19404) );
  OR2_X1 U22389 ( .A1(n19403), .A2(n19404), .ZN(n19427) );
  INV_X1 U22390 ( .A(n19406), .ZN(n19426) );
  AOI22_X1 U22391 ( .A1(n19427), .A2(n19790), .B1(n19779), .B2(n19426), .ZN(
        n19412) );
  AOI21_X1 U22392 ( .B1(n19442), .B2(n19419), .A(n19781), .ZN(n19405) );
  OR2_X1 U22393 ( .A1(n19405), .A2(n19404), .ZN(n19409) );
  OAI21_X1 U22394 ( .B1(n19407), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19406), 
        .ZN(n19408) );
  MUX2_X1 U22395 ( .A(n19409), .B(n19408), .S(n19703), .Z(n19410) );
  NAND2_X1 U22396 ( .A1(n19410), .A2(n19738), .ZN(n19429) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19429), .B1(
        n19428), .B2(n19747), .ZN(n19411) );
  OAI211_X1 U22398 ( .C1(n19710), .C2(n19442), .A(n19412), .B(n19411), .ZN(
        P2_U3064) );
  AOI22_X1 U22399 ( .A1(n19427), .A2(n19815), .B1(n19344), .B2(n19426), .ZN(
        n19414) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19429), .B1(
        n19428), .B2(n19816), .ZN(n19413) );
  OAI211_X1 U22401 ( .C1(n19819), .C2(n19442), .A(n19414), .B(n19413), .ZN(
        P2_U3065) );
  AOI22_X1 U22402 ( .A1(n19427), .A2(n19821), .B1(n19820), .B2(n19426), .ZN(
        n19416) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19429), .B1(
        n19428), .B2(n19822), .ZN(n19415) );
  OAI211_X1 U22404 ( .C1(n19798), .C2(n19442), .A(n19416), .B(n19415), .ZN(
        P2_U3066) );
  AOI22_X1 U22405 ( .A1(n19427), .A2(n19828), .B1(n19827), .B2(n19426), .ZN(
        n19418) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19429), .B1(
        n19446), .B2(n19757), .ZN(n19417) );
  OAI211_X1 U22407 ( .C1(n19679), .C2(n19419), .A(n19418), .B(n19417), .ZN(
        P2_U3067) );
  AOI22_X1 U22408 ( .A1(n19427), .A2(n19834), .B1(n19833), .B2(n19426), .ZN(
        n19421) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19429), .B1(
        n19428), .B2(n19835), .ZN(n19420) );
  OAI211_X1 U22410 ( .C1(n19839), .C2(n19442), .A(n19421), .B(n19420), .ZN(
        P2_U3068) );
  AOI22_X1 U22411 ( .A1(n19427), .A2(n19841), .B1(n19840), .B2(n19426), .ZN(
        n19423) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19429), .B1(
        n19428), .B2(n19763), .ZN(n19422) );
  OAI211_X1 U22413 ( .C1(n19766), .C2(n19442), .A(n19423), .B(n19422), .ZN(
        P2_U3069) );
  AOI22_X1 U22414 ( .A1(n19427), .A2(n19847), .B1(n19846), .B2(n19426), .ZN(
        n19425) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19429), .B1(
        n19428), .B2(n19767), .ZN(n19424) );
  OAI211_X1 U22416 ( .C1(n19723), .C2(n19442), .A(n19425), .B(n19424), .ZN(
        P2_U3070) );
  AOI22_X1 U22417 ( .A1(n19427), .A2(n19856), .B1(n19854), .B2(n19426), .ZN(
        n19431) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19429), .B1(
        n19428), .B2(n19858), .ZN(n19430) );
  OAI211_X1 U22419 ( .C1(n19777), .C2(n19442), .A(n19431), .B(n19430), .ZN(
        P2_U3071) );
  AOI22_X1 U22420 ( .A1(n19816), .A2(n19446), .B1(n19445), .B2(n19344), .ZN(
        n19433) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19448), .B1(
        n19815), .B2(n19447), .ZN(n19432) );
  OAI211_X1 U22422 ( .C1(n19819), .C2(n19481), .A(n19433), .B(n19432), .ZN(
        P2_U3073) );
  AOI22_X1 U22423 ( .A1(n19822), .A2(n19446), .B1(n19445), .B2(n19820), .ZN(
        n19435) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19448), .B1(
        n19821), .B2(n19447), .ZN(n19434) );
  OAI211_X1 U22425 ( .C1(n19798), .C2(n19481), .A(n19435), .B(n19434), .ZN(
        P2_U3074) );
  AOI22_X1 U22426 ( .A1(n19829), .A2(n19446), .B1(n19445), .B2(n19827), .ZN(
        n19437) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19448), .B1(
        n19828), .B2(n19447), .ZN(n19436) );
  OAI211_X1 U22428 ( .C1(n19832), .C2(n19481), .A(n19437), .B(n19436), .ZN(
        P2_U3075) );
  AOI22_X1 U22429 ( .A1(n19835), .A2(n19446), .B1(n19445), .B2(n19833), .ZN(
        n19439) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19448), .B1(
        n19834), .B2(n19447), .ZN(n19438) );
  OAI211_X1 U22431 ( .C1(n19839), .C2(n19481), .A(n19439), .B(n19438), .ZN(
        P2_U3076) );
  AOI22_X1 U22432 ( .A1(n19842), .A2(n19463), .B1(n19445), .B2(n19840), .ZN(
        n19441) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19448), .B1(
        n19841), .B2(n19447), .ZN(n19440) );
  OAI211_X1 U22434 ( .C1(n19845), .C2(n19442), .A(n19441), .B(n19440), .ZN(
        P2_U3077) );
  AOI22_X1 U22435 ( .A1(n19767), .A2(n19446), .B1(n19445), .B2(n19846), .ZN(
        n19444) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19448), .B1(
        n19847), .B2(n19447), .ZN(n19443) );
  OAI211_X1 U22437 ( .C1(n19723), .C2(n19481), .A(n19444), .B(n19443), .ZN(
        P2_U3078) );
  AOI22_X1 U22438 ( .A1(n19858), .A2(n19446), .B1(n19445), .B2(n19854), .ZN(
        n19450) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19448), .B1(
        n19856), .B2(n19447), .ZN(n19449) );
  OAI211_X1 U22440 ( .C1(n19777), .C2(n19481), .A(n19450), .B(n19449), .ZN(
        P2_U3079) );
  NAND3_X1 U22441 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19950), .A3(
        n19968), .ZN(n19487) );
  NOR2_X1 U22442 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19487), .ZN(
        n19476) );
  AOI22_X1 U22443 ( .A1(n19747), .A2(n19463), .B1(n19779), .B2(n19476), .ZN(
        n19462) );
  NOR2_X1 U22444 ( .A1(n19463), .A2(n19497), .ZN(n19451) );
  OAI21_X1 U22445 ( .B1(n19451), .B2(n19781), .A(n19942), .ZN(n19460) );
  INV_X1 U22446 ( .A(n19452), .ZN(n19697) );
  NAND2_X1 U22447 ( .A1(n19697), .A2(n19453), .ZN(n19702) );
  NOR2_X1 U22448 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19702), .ZN(
        n19457) );
  INV_X1 U22449 ( .A(n11125), .ZN(n19455) );
  INV_X1 U22450 ( .A(n19476), .ZN(n19454) );
  OAI211_X1 U22451 ( .C1(n19455), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19454), 
        .B(n19703), .ZN(n19456) );
  OAI211_X1 U22452 ( .C1(n19460), .C2(n19457), .A(n19738), .B(n19456), .ZN(
        n19478) );
  INV_X1 U22453 ( .A(n19457), .ZN(n19459) );
  OAI21_X1 U22454 ( .B1(n11125), .B2(n19476), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19458) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19478), .B1(
        n19790), .B2(n19477), .ZN(n19461) );
  OAI211_X1 U22456 ( .C1(n19710), .C2(n19509), .A(n19462), .B(n19461), .ZN(
        P2_U3080) );
  AOI22_X1 U22457 ( .A1(n19816), .A2(n19463), .B1(n19344), .B2(n19476), .ZN(
        n19465) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19478), .B1(
        n19815), .B2(n19477), .ZN(n19464) );
  OAI211_X1 U22459 ( .C1(n19819), .C2(n19509), .A(n19465), .B(n19464), .ZN(
        P2_U3081) );
  AOI22_X1 U22460 ( .A1(n19823), .A2(n19497), .B1(n19820), .B2(n19476), .ZN(
        n19467) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19478), .B1(
        n19821), .B2(n19477), .ZN(n19466) );
  OAI211_X1 U22462 ( .C1(n19676), .C2(n19481), .A(n19467), .B(n19466), .ZN(
        P2_U3082) );
  AOI22_X1 U22463 ( .A1(n19757), .A2(n19497), .B1(n19476), .B2(n19827), .ZN(
        n19469) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19478), .B1(
        n19828), .B2(n19477), .ZN(n19468) );
  OAI211_X1 U22465 ( .C1(n19679), .C2(n19481), .A(n19469), .B(n19468), .ZN(
        P2_U3083) );
  AOI22_X1 U22466 ( .A1(n19680), .A2(n19497), .B1(n19476), .B2(n19833), .ZN(
        n19471) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19478), .B1(
        n19834), .B2(n19477), .ZN(n19470) );
  OAI211_X1 U22468 ( .C1(n19683), .C2(n19481), .A(n19471), .B(n19470), .ZN(
        P2_U3084) );
  AOI22_X1 U22469 ( .A1(n19842), .A2(n19497), .B1(n19840), .B2(n19476), .ZN(
        n19473) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19478), .B1(
        n19841), .B2(n19477), .ZN(n19472) );
  OAI211_X1 U22471 ( .C1(n19845), .C2(n19481), .A(n19473), .B(n19472), .ZN(
        P2_U3085) );
  AOI22_X1 U22472 ( .A1(n19848), .A2(n19497), .B1(n19846), .B2(n19476), .ZN(
        n19475) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19478), .B1(
        n19847), .B2(n19477), .ZN(n19474) );
  OAI211_X1 U22474 ( .C1(n19853), .C2(n19481), .A(n19475), .B(n19474), .ZN(
        P2_U3086) );
  AOI22_X1 U22475 ( .A1(n19860), .A2(n19497), .B1(n19854), .B2(n19476), .ZN(
        n19480) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19478), .B1(
        n19856), .B2(n19477), .ZN(n19479) );
  OAI211_X1 U22477 ( .C1(n19814), .C2(n19481), .A(n19480), .B(n19479), .ZN(
        P2_U3087) );
  NOR2_X1 U22478 ( .A1(n19976), .A2(n19487), .ZN(n19514) );
  AOI22_X1 U22479 ( .A1(n19747), .A2(n19497), .B1(n19779), .B2(n19514), .ZN(
        n19490) );
  OAI21_X1 U22480 ( .B1(n19538), .B2(n19730), .A(n19942), .ZN(n19488) );
  INV_X1 U22481 ( .A(n19487), .ZN(n19485) );
  INV_X1 U22482 ( .A(n11111), .ZN(n19483) );
  INV_X1 U22483 ( .A(n19514), .ZN(n19482) );
  OAI211_X1 U22484 ( .C1(n19483), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19482), 
        .B(n19703), .ZN(n19484) );
  OAI211_X1 U22485 ( .C1(n19488), .C2(n19485), .A(n19738), .B(n19484), .ZN(
        n19506) );
  OAI21_X1 U22486 ( .B1(n11111), .B2(n19514), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19486) );
  OAI21_X1 U22487 ( .B1(n19488), .B2(n19487), .A(n19486), .ZN(n19505) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19506), .B1(
        n19790), .B2(n19505), .ZN(n19489) );
  OAI211_X1 U22489 ( .C1(n19710), .C2(n19537), .A(n19490), .B(n19489), .ZN(
        P2_U3088) );
  INV_X1 U22490 ( .A(n19537), .ZN(n19504) );
  AOI22_X1 U22491 ( .A1(n19750), .A2(n19504), .B1(n19344), .B2(n19514), .ZN(
        n19492) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19506), .B1(
        n19815), .B2(n19505), .ZN(n19491) );
  OAI211_X1 U22493 ( .C1(n19754), .C2(n19509), .A(n19492), .B(n19491), .ZN(
        P2_U3089) );
  AOI22_X1 U22494 ( .A1(n19822), .A2(n19497), .B1(n19514), .B2(n19820), .ZN(
        n19494) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19506), .B1(
        n19821), .B2(n19505), .ZN(n19493) );
  OAI211_X1 U22496 ( .C1(n19798), .C2(n19537), .A(n19494), .B(n19493), .ZN(
        P2_U3090) );
  AOI22_X1 U22497 ( .A1(n19829), .A2(n19497), .B1(n19514), .B2(n19827), .ZN(
        n19496) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19506), .B1(
        n19828), .B2(n19505), .ZN(n19495) );
  OAI211_X1 U22499 ( .C1(n19832), .C2(n19537), .A(n19496), .B(n19495), .ZN(
        P2_U3091) );
  AOI22_X1 U22500 ( .A1(n19835), .A2(n19497), .B1(n19514), .B2(n19833), .ZN(
        n19499) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19506), .B1(
        n19834), .B2(n19505), .ZN(n19498) );
  OAI211_X1 U22502 ( .C1(n19839), .C2(n19537), .A(n19499), .B(n19498), .ZN(
        P2_U3092) );
  AOI22_X1 U22503 ( .A1(n19842), .A2(n19504), .B1(n19514), .B2(n19840), .ZN(
        n19501) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19506), .B1(
        n19841), .B2(n19505), .ZN(n19500) );
  OAI211_X1 U22505 ( .C1(n19845), .C2(n19509), .A(n19501), .B(n19500), .ZN(
        P2_U3093) );
  AOI22_X1 U22506 ( .A1(n19848), .A2(n19504), .B1(n19514), .B2(n19846), .ZN(
        n19503) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19506), .B1(
        n19847), .B2(n19505), .ZN(n19502) );
  OAI211_X1 U22508 ( .C1(n19853), .C2(n19509), .A(n19503), .B(n19502), .ZN(
        P2_U3094) );
  AOI22_X1 U22509 ( .A1(n19860), .A2(n19504), .B1(n19514), .B2(n19854), .ZN(
        n19508) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19506), .B1(
        n19856), .B2(n19505), .ZN(n19507) );
  OAI211_X1 U22511 ( .C1(n19814), .C2(n19509), .A(n19508), .B(n19507), .ZN(
        P2_U3095) );
  NOR2_X1 U22512 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19544), .ZN(
        n19532) );
  NOR2_X1 U22513 ( .A1(n19514), .A2(n19532), .ZN(n19511) );
  NOR3_X1 U22514 ( .A1(n11114), .A2(n19995), .A3(n19532), .ZN(n19515) );
  AOI211_X2 U22515 ( .C1(n19995), .C2(n19511), .A(n19510), .B(n19515), .ZN(
        n19533) );
  AOI22_X1 U22516 ( .A1(n19533), .A2(n19790), .B1(n19779), .B2(n19532), .ZN(
        n19519) );
  NAND2_X1 U22517 ( .A1(n19545), .A2(n19512), .ZN(n19517) );
  AOI21_X1 U22518 ( .B1(n19537), .B2(n19517), .A(n19781), .ZN(n19513) );
  AOI221_X1 U22519 ( .B1(n20000), .B2(n19514), .C1(n20000), .C2(n19513), .A(
        n19532), .ZN(n19516) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19780), .ZN(n19518) );
  OAI211_X1 U22521 ( .C1(n19793), .C2(n19537), .A(n19519), .B(n19518), .ZN(
        P2_U3096) );
  AOI22_X1 U22522 ( .A1(n19533), .A2(n19815), .B1(n19344), .B2(n19532), .ZN(
        n19521) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19750), .ZN(n19520) );
  OAI211_X1 U22524 ( .C1(n19754), .C2(n19537), .A(n19521), .B(n19520), .ZN(
        P2_U3097) );
  AOI22_X1 U22525 ( .A1(n19533), .A2(n19821), .B1(n19820), .B2(n19532), .ZN(
        n19523) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19823), .ZN(n19522) );
  OAI211_X1 U22527 ( .C1(n19676), .C2(n19537), .A(n19523), .B(n19522), .ZN(
        P2_U3098) );
  AOI22_X1 U22528 ( .A1(n19533), .A2(n19828), .B1(n19827), .B2(n19532), .ZN(
        n19525) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19757), .ZN(n19524) );
  OAI211_X1 U22530 ( .C1(n19679), .C2(n19537), .A(n19525), .B(n19524), .ZN(
        P2_U3099) );
  AOI22_X1 U22531 ( .A1(n19533), .A2(n19834), .B1(n19833), .B2(n19532), .ZN(
        n19527) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19680), .ZN(n19526) );
  OAI211_X1 U22533 ( .C1(n19683), .C2(n19537), .A(n19527), .B(n19526), .ZN(
        P2_U3100) );
  AOI22_X1 U22534 ( .A1(n19533), .A2(n19841), .B1(n19840), .B2(n19532), .ZN(
        n19529) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19842), .ZN(n19528) );
  OAI211_X1 U22536 ( .C1(n19845), .C2(n19537), .A(n19529), .B(n19528), .ZN(
        P2_U3101) );
  AOI22_X1 U22537 ( .A1(n19533), .A2(n19847), .B1(n19846), .B2(n19532), .ZN(
        n19531) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19848), .ZN(n19530) );
  OAI211_X1 U22539 ( .C1(n19853), .C2(n19537), .A(n19531), .B(n19530), .ZN(
        P2_U3102) );
  AOI22_X1 U22540 ( .A1(n19533), .A2(n19856), .B1(n19854), .B2(n19532), .ZN(
        n19536) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19534), .B1(
        n19566), .B2(n19860), .ZN(n19535) );
  OAI211_X1 U22542 ( .C1(n19814), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3103) );
  OAI21_X1 U22543 ( .B1(n19538), .B2(n19937), .A(n19544), .ZN(n19542) );
  NAND2_X1 U22544 ( .A1(n11122), .A2(n20000), .ZN(n19540) );
  INV_X1 U22545 ( .A(n19574), .ZN(n19564) );
  NOR2_X1 U22546 ( .A1(n19942), .A2(n19564), .ZN(n19539) );
  AOI21_X1 U22547 ( .B1(n19540), .B2(n19539), .A(n19784), .ZN(n19541) );
  AND2_X1 U22548 ( .A1(n19542), .A2(n19541), .ZN(n19557) );
  INV_X1 U22549 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19549) );
  OAI21_X1 U22550 ( .B1(n11122), .B2(n19564), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19543) );
  OAI21_X1 U22551 ( .B1(n19544), .B2(n19703), .A(n19543), .ZN(n19565) );
  AOI22_X1 U22552 ( .A1(n19565), .A2(n19790), .B1(n19564), .B2(n19779), .ZN(
        n19548) );
  INV_X1 U22553 ( .A(n19598), .ZN(n19590) );
  AOI22_X1 U22554 ( .A1(n19590), .A2(n19780), .B1(n19566), .B2(n19747), .ZN(
        n19547) );
  OAI211_X1 U22555 ( .C1(n19557), .C2(n19549), .A(n19548), .B(n19547), .ZN(
        P2_U3104) );
  AOI22_X1 U22556 ( .A1(n19565), .A2(n19815), .B1(n19564), .B2(n19344), .ZN(
        n19551) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19816), .ZN(n19550) );
  OAI211_X1 U22558 ( .C1(n19819), .C2(n19598), .A(n19551), .B(n19550), .ZN(
        P2_U3105) );
  AOI22_X1 U22559 ( .A1(n19565), .A2(n19821), .B1(n19564), .B2(n19820), .ZN(
        n19553) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19822), .ZN(n19552) );
  OAI211_X1 U22561 ( .C1(n19798), .C2(n19598), .A(n19553), .B(n19552), .ZN(
        P2_U3106) );
  INV_X1 U22562 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n19556) );
  AOI22_X1 U22563 ( .A1(n19565), .A2(n19828), .B1(n19564), .B2(n19827), .ZN(
        n19555) );
  AOI22_X1 U22564 ( .A1(n19590), .A2(n19757), .B1(n19566), .B2(n19829), .ZN(
        n19554) );
  OAI211_X1 U22565 ( .C1(n19557), .C2(n19556), .A(n19555), .B(n19554), .ZN(
        P2_U3107) );
  AOI22_X1 U22566 ( .A1(n19565), .A2(n19834), .B1(n19564), .B2(n19833), .ZN(
        n19559) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19835), .ZN(n19558) );
  OAI211_X1 U22568 ( .C1(n19839), .C2(n19598), .A(n19559), .B(n19558), .ZN(
        P2_U3108) );
  AOI22_X1 U22569 ( .A1(n19565), .A2(n19841), .B1(n19564), .B2(n19840), .ZN(
        n19561) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19763), .ZN(n19560) );
  OAI211_X1 U22571 ( .C1(n19766), .C2(n19598), .A(n19561), .B(n19560), .ZN(
        P2_U3109) );
  AOI22_X1 U22572 ( .A1(n19565), .A2(n19847), .B1(n19564), .B2(n19846), .ZN(
        n19563) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19767), .ZN(n19562) );
  OAI211_X1 U22574 ( .C1(n19723), .C2(n19598), .A(n19563), .B(n19562), .ZN(
        P2_U3110) );
  AOI22_X1 U22575 ( .A1(n19565), .A2(n19856), .B1(n19564), .B2(n19854), .ZN(
        n19569) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19858), .ZN(n19568) );
  OAI211_X1 U22577 ( .C1(n19777), .C2(n19598), .A(n19569), .B(n19568), .ZN(
        P2_U3111) );
  NOR2_X1 U22578 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19950), .ZN(
        n19660) );
  NAND2_X1 U22579 ( .A1(n19660), .A2(n19968), .ZN(n19603) );
  NOR2_X1 U22580 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19603), .ZN(
        n19593) );
  AOI22_X1 U22581 ( .A1(n19747), .A2(n19590), .B1(n19779), .B2(n19593), .ZN(
        n19579) );
  NAND2_X1 U22582 ( .A1(n19625), .A2(n19598), .ZN(n19570) );
  AOI21_X1 U22583 ( .B1(n19570), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19703), 
        .ZN(n19573) );
  OAI21_X1 U22584 ( .B1(n11115), .B2(n19995), .A(n20000), .ZN(n19571) );
  AOI21_X1 U22585 ( .B1(n19573), .B2(n19574), .A(n19571), .ZN(n19572) );
  OAI21_X1 U22586 ( .B1(n19593), .B2(n19572), .A(n19738), .ZN(n19595) );
  NOR2_X1 U22587 ( .A1(n19573), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19577) );
  AOI21_X1 U22588 ( .B1(n11115), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19593), 
        .ZN(n19576) );
  INV_X1 U22589 ( .A(n19573), .ZN(n19575) );
  OAI22_X1 U22590 ( .A1(n19577), .A2(n19576), .B1(n19575), .B2(n19574), .ZN(
        n19594) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19595), .B1(
        n19790), .B2(n19594), .ZN(n19578) );
  OAI211_X1 U22592 ( .C1(n19710), .C2(n19625), .A(n19579), .B(n19578), .ZN(
        P2_U3112) );
  AOI22_X1 U22593 ( .A1(n19750), .A2(n19626), .B1(n19344), .B2(n19593), .ZN(
        n19581) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19815), .ZN(n19580) );
  OAI211_X1 U22595 ( .C1(n19754), .C2(n19598), .A(n19581), .B(n19580), .ZN(
        P2_U3113) );
  AOI22_X1 U22596 ( .A1(n19823), .A2(n19626), .B1(n19820), .B2(n19593), .ZN(
        n19583) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19821), .ZN(n19582) );
  OAI211_X1 U22598 ( .C1(n19676), .C2(n19598), .A(n19583), .B(n19582), .ZN(
        P2_U3114) );
  AOI22_X1 U22599 ( .A1(n19829), .A2(n19590), .B1(n19827), .B2(n19593), .ZN(
        n19585) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19828), .ZN(n19584) );
  OAI211_X1 U22601 ( .C1(n19832), .C2(n19625), .A(n19585), .B(n19584), .ZN(
        P2_U3115) );
  AOI22_X1 U22602 ( .A1(n19835), .A2(n19590), .B1(n19833), .B2(n19593), .ZN(
        n19587) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19834), .ZN(n19586) );
  OAI211_X1 U22604 ( .C1(n19839), .C2(n19625), .A(n19587), .B(n19586), .ZN(
        P2_U3116) );
  AOI22_X1 U22605 ( .A1(n19842), .A2(n19626), .B1(n19840), .B2(n19593), .ZN(
        n19589) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19841), .ZN(n19588) );
  OAI211_X1 U22607 ( .C1(n19845), .C2(n19598), .A(n19589), .B(n19588), .ZN(
        P2_U3117) );
  AOI22_X1 U22608 ( .A1(n19767), .A2(n19590), .B1(n19846), .B2(n19593), .ZN(
        n19592) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19847), .ZN(n19591) );
  OAI211_X1 U22610 ( .C1(n19723), .C2(n19625), .A(n19592), .B(n19591), .ZN(
        P2_U3118) );
  AOI22_X1 U22611 ( .A1(n19860), .A2(n19626), .B1(n19854), .B2(n19593), .ZN(
        n19597) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19856), .ZN(n19596) );
  OAI211_X1 U22613 ( .C1(n19814), .C2(n19598), .A(n19597), .B(n19596), .ZN(
        P2_U3119) );
  NOR2_X2 U22614 ( .A1(n19744), .A2(n19601), .ZN(n19656) );
  INV_X1 U22615 ( .A(n19656), .ZN(n19631) );
  INV_X1 U22616 ( .A(n19660), .ZN(n19662) );
  NOR2_X1 U22617 ( .A1(n19600), .A2(n19662), .ZN(n19635) );
  AOI22_X1 U22618 ( .A1(n19626), .A2(n19747), .B1(n19779), .B2(n19635), .ZN(
        n19612) );
  INV_X1 U22619 ( .A(n11116), .ZN(n19605) );
  INV_X1 U22620 ( .A(n19732), .ZN(n19602) );
  NOR2_X1 U22621 ( .A1(n19602), .A2(n19601), .ZN(n19610) );
  INV_X1 U22622 ( .A(n19603), .ZN(n19607) );
  NOR2_X1 U22623 ( .A1(n19610), .A2(n19607), .ZN(n19604) );
  AOI211_X1 U22624 ( .C1(n19605), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19604), .ZN(n19606) );
  OAI21_X1 U22625 ( .B1(n19635), .B2(n19606), .A(n19738), .ZN(n19628) );
  NAND2_X1 U22626 ( .A1(n19607), .A2(n19942), .ZN(n19609) );
  OAI21_X1 U22627 ( .B1(n11116), .B2(n19635), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19608) );
  OAI21_X1 U22628 ( .B1(n19610), .B2(n19609), .A(n19608), .ZN(n19627) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19628), .B1(
        n19790), .B2(n19627), .ZN(n19611) );
  OAI211_X1 U22630 ( .C1(n19710), .C2(n19631), .A(n19612), .B(n19611), .ZN(
        P2_U3120) );
  AOI22_X1 U22631 ( .A1(n19750), .A2(n19656), .B1(n19344), .B2(n19635), .ZN(
        n19614) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19628), .B1(
        n19815), .B2(n19627), .ZN(n19613) );
  OAI211_X1 U22633 ( .C1(n19754), .C2(n19625), .A(n19614), .B(n19613), .ZN(
        P2_U3121) );
  AOI22_X1 U22634 ( .A1(n19822), .A2(n19626), .B1(n19820), .B2(n19635), .ZN(
        n19616) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19628), .B1(
        n19821), .B2(n19627), .ZN(n19615) );
  OAI211_X1 U22636 ( .C1(n19798), .C2(n19631), .A(n19616), .B(n19615), .ZN(
        P2_U3122) );
  AOI22_X1 U22637 ( .A1(n19829), .A2(n19626), .B1(n19827), .B2(n19635), .ZN(
        n19618) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19628), .B1(
        n19828), .B2(n19627), .ZN(n19617) );
  OAI211_X1 U22639 ( .C1(n19832), .C2(n19631), .A(n19618), .B(n19617), .ZN(
        P2_U3123) );
  AOI22_X1 U22640 ( .A1(n19680), .A2(n19656), .B1(n19833), .B2(n19635), .ZN(
        n19620) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19628), .B1(
        n19834), .B2(n19627), .ZN(n19619) );
  OAI211_X1 U22642 ( .C1(n19683), .C2(n19625), .A(n19620), .B(n19619), .ZN(
        P2_U3124) );
  AOI22_X1 U22643 ( .A1(n19842), .A2(n19656), .B1(n19840), .B2(n19635), .ZN(
        n19622) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19628), .B1(
        n19841), .B2(n19627), .ZN(n19621) );
  OAI211_X1 U22645 ( .C1(n19845), .C2(n19625), .A(n19622), .B(n19621), .ZN(
        P2_U3125) );
  AOI22_X1 U22646 ( .A1(n19848), .A2(n19656), .B1(n19846), .B2(n19635), .ZN(
        n19624) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19628), .B1(
        n19847), .B2(n19627), .ZN(n19623) );
  OAI211_X1 U22648 ( .C1(n19853), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P2_U3126) );
  AOI22_X1 U22649 ( .A1(n19858), .A2(n19626), .B1(n19854), .B2(n19635), .ZN(
        n19630) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19628), .B1(
        n19856), .B2(n19627), .ZN(n19629) );
  OAI211_X1 U22651 ( .C1(n19777), .C2(n19631), .A(n19630), .B(n19629), .ZN(
        P2_U3127) );
  AND2_X1 U22652 ( .A1(n19632), .A2(n19660), .ZN(n19654) );
  OAI21_X1 U22653 ( .B1(n11126), .B2(n19654), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19633) );
  OAI21_X1 U22654 ( .B1(n19662), .B2(n19634), .A(n19633), .ZN(n19655) );
  AOI22_X1 U22655 ( .A1(n19655), .A2(n19790), .B1(n19779), .B2(n19654), .ZN(
        n19641) );
  NOR2_X1 U22656 ( .A1(n11126), .A2(n19995), .ZN(n19638) );
  INV_X1 U22657 ( .A(n19693), .ZN(n19636) );
  AOI221_X1 U22658 ( .B1(n19656), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19636), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19635), .ZN(n19637) );
  NOR3_X1 U22659 ( .A1(n19638), .A2(n19637), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19639) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19747), .ZN(n19640) );
  OAI211_X1 U22661 ( .C1(n19710), .C2(n19693), .A(n19641), .B(n19640), .ZN(
        P2_U3128) );
  AOI22_X1 U22662 ( .A1(n19655), .A2(n19815), .B1(n19344), .B2(n19654), .ZN(
        n19643) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19816), .ZN(n19642) );
  OAI211_X1 U22664 ( .C1(n19819), .C2(n19693), .A(n19643), .B(n19642), .ZN(
        P2_U3129) );
  AOI22_X1 U22665 ( .A1(n19655), .A2(n19821), .B1(n19820), .B2(n19654), .ZN(
        n19645) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19822), .ZN(n19644) );
  OAI211_X1 U22667 ( .C1(n19798), .C2(n19693), .A(n19645), .B(n19644), .ZN(
        P2_U3130) );
  AOI22_X1 U22668 ( .A1(n19655), .A2(n19828), .B1(n19827), .B2(n19654), .ZN(
        n19647) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19829), .ZN(n19646) );
  OAI211_X1 U22670 ( .C1(n19832), .C2(n19693), .A(n19647), .B(n19646), .ZN(
        P2_U3131) );
  AOI22_X1 U22671 ( .A1(n19655), .A2(n19834), .B1(n19833), .B2(n19654), .ZN(
        n19649) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19835), .ZN(n19648) );
  OAI211_X1 U22673 ( .C1(n19839), .C2(n19693), .A(n19649), .B(n19648), .ZN(
        P2_U3132) );
  AOI22_X1 U22674 ( .A1(n19655), .A2(n19841), .B1(n19840), .B2(n19654), .ZN(
        n19651) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19763), .ZN(n19650) );
  OAI211_X1 U22676 ( .C1(n19766), .C2(n19693), .A(n19651), .B(n19650), .ZN(
        P2_U3133) );
  AOI22_X1 U22677 ( .A1(n19655), .A2(n19847), .B1(n19846), .B2(n19654), .ZN(
        n19653) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19767), .ZN(n19652) );
  OAI211_X1 U22679 ( .C1(n19723), .C2(n19693), .A(n19653), .B(n19652), .ZN(
        P2_U3134) );
  AOI22_X1 U22680 ( .A1(n19655), .A2(n19856), .B1(n19854), .B2(n19654), .ZN(
        n19659) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19858), .ZN(n19658) );
  OAI211_X1 U22682 ( .C1(n19777), .C2(n19693), .A(n19659), .B(n19658), .ZN(
        P2_U3135) );
  NAND2_X1 U22683 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19660), .ZN(
        n19664) );
  OR2_X1 U22684 ( .A1(n19664), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19663) );
  NOR2_X1 U22685 ( .A1(n19662), .A2(n19661), .ZN(n19688) );
  NOR3_X1 U22686 ( .A1(n11121), .A2(n19995), .A3(n19688), .ZN(n19665) );
  AOI21_X1 U22687 ( .B1(n19995), .B2(n19663), .A(n19665), .ZN(n19689) );
  AOI22_X1 U22688 ( .A1(n19689), .A2(n19790), .B1(n19779), .B2(n19688), .ZN(
        n19671) );
  INV_X1 U22689 ( .A(n19664), .ZN(n19668) );
  INV_X1 U22690 ( .A(n19688), .ZN(n19666) );
  AOI211_X1 U22691 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19666), .A(n19784), 
        .B(n19665), .ZN(n19667) );
  OAI221_X1 U22692 ( .B1(n19668), .B2(n19940), .C1(n19668), .C2(n19732), .A(
        n19667), .ZN(n19690) );
  NOR2_X2 U22693 ( .A1(n19744), .A2(n19669), .ZN(n19726) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19780), .ZN(n19670) );
  OAI211_X1 U22695 ( .C1(n19793), .C2(n19693), .A(n19671), .B(n19670), .ZN(
        P2_U3136) );
  AOI22_X1 U22696 ( .A1(n19689), .A2(n19815), .B1(n19344), .B2(n19688), .ZN(
        n19673) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19750), .ZN(n19672) );
  OAI211_X1 U22698 ( .C1(n19754), .C2(n19693), .A(n19673), .B(n19672), .ZN(
        P2_U3137) );
  AOI22_X1 U22699 ( .A1(n19689), .A2(n19821), .B1(n19820), .B2(n19688), .ZN(
        n19675) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19823), .ZN(n19674) );
  OAI211_X1 U22701 ( .C1(n19676), .C2(n19693), .A(n19675), .B(n19674), .ZN(
        P2_U3138) );
  AOI22_X1 U22702 ( .A1(n19689), .A2(n19828), .B1(n19827), .B2(n19688), .ZN(
        n19678) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19757), .ZN(n19677) );
  OAI211_X1 U22704 ( .C1(n19679), .C2(n19693), .A(n19678), .B(n19677), .ZN(
        P2_U3139) );
  AOI22_X1 U22705 ( .A1(n19689), .A2(n19834), .B1(n19833), .B2(n19688), .ZN(
        n19682) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19680), .ZN(n19681) );
  OAI211_X1 U22707 ( .C1(n19683), .C2(n19693), .A(n19682), .B(n19681), .ZN(
        P2_U3140) );
  AOI22_X1 U22708 ( .A1(n19689), .A2(n19841), .B1(n19840), .B2(n19688), .ZN(
        n19685) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19842), .ZN(n19684) );
  OAI211_X1 U22710 ( .C1(n19845), .C2(n19693), .A(n19685), .B(n19684), .ZN(
        P2_U3141) );
  AOI22_X1 U22711 ( .A1(n19689), .A2(n19847), .B1(n19846), .B2(n19688), .ZN(
        n19687) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19848), .ZN(n19686) );
  OAI211_X1 U22713 ( .C1(n19853), .C2(n19693), .A(n19687), .B(n19686), .ZN(
        P2_U3142) );
  AOI22_X1 U22714 ( .A1(n19689), .A2(n19856), .B1(n19854), .B2(n19688), .ZN(
        n19692) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19690), .B1(
        n19726), .B2(n19860), .ZN(n19691) );
  OAI211_X1 U22716 ( .C1(n19814), .C2(n19693), .A(n19692), .B(n19691), .ZN(
        P2_U3143) );
  INV_X1 U22717 ( .A(n19694), .ZN(n19695) );
  NOR3_X1 U22718 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19958), .A3(
        n19950), .ZN(n19733) );
  INV_X1 U22719 ( .A(n19733), .ZN(n19741) );
  NOR2_X1 U22720 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19741), .ZN(
        n19724) );
  OAI21_X1 U22721 ( .B1(n11124), .B2(n19724), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19700) );
  NAND3_X1 U22722 ( .A1(n19698), .A2(n19697), .A3(n19696), .ZN(n19699) );
  NAND2_X1 U22723 ( .A1(n19700), .A2(n19699), .ZN(n19725) );
  AOI22_X1 U22724 ( .A1(n19725), .A2(n19790), .B1(n19779), .B2(n19724), .ZN(
        n19709) );
  OAI21_X1 U22725 ( .B1(n19773), .B2(n19726), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19701) );
  OAI21_X1 U22726 ( .B1(n19702), .B2(n19950), .A(n19701), .ZN(n19707) );
  INV_X1 U22727 ( .A(n11124), .ZN(n19705) );
  INV_X1 U22728 ( .A(n19724), .ZN(n19704) );
  OAI211_X1 U22729 ( .C1(n19705), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19704), 
        .B(n19703), .ZN(n19706) );
  NAND3_X1 U22730 ( .A1(n19707), .A2(n19738), .A3(n19706), .ZN(n19727) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19747), .ZN(n19708) );
  OAI211_X1 U22732 ( .C1(n19710), .C2(n19753), .A(n19709), .B(n19708), .ZN(
        P2_U3144) );
  AOI22_X1 U22733 ( .A1(n19725), .A2(n19815), .B1(n19344), .B2(n19724), .ZN(
        n19712) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19816), .ZN(n19711) );
  OAI211_X1 U22735 ( .C1(n19819), .C2(n19753), .A(n19712), .B(n19711), .ZN(
        P2_U3145) );
  AOI22_X1 U22736 ( .A1(n19725), .A2(n19821), .B1(n19820), .B2(n19724), .ZN(
        n19714) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19822), .ZN(n19713) );
  OAI211_X1 U22738 ( .C1(n19798), .C2(n19753), .A(n19714), .B(n19713), .ZN(
        P2_U3146) );
  AOI22_X1 U22739 ( .A1(n19725), .A2(n19828), .B1(n19827), .B2(n19724), .ZN(
        n19716) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19829), .ZN(n19715) );
  OAI211_X1 U22741 ( .C1(n19832), .C2(n19753), .A(n19716), .B(n19715), .ZN(
        P2_U3147) );
  AOI22_X1 U22742 ( .A1(n19725), .A2(n19834), .B1(n19833), .B2(n19724), .ZN(
        n19718) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19835), .ZN(n19717) );
  OAI211_X1 U22744 ( .C1(n19839), .C2(n19753), .A(n19718), .B(n19717), .ZN(
        P2_U3148) );
  AOI22_X1 U22745 ( .A1(n19725), .A2(n19841), .B1(n19840), .B2(n19724), .ZN(
        n19720) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19763), .ZN(n19719) );
  OAI211_X1 U22747 ( .C1(n19766), .C2(n19753), .A(n19720), .B(n19719), .ZN(
        P2_U3149) );
  AOI22_X1 U22748 ( .A1(n19725), .A2(n19847), .B1(n19846), .B2(n19724), .ZN(
        n19722) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19767), .ZN(n19721) );
  OAI211_X1 U22750 ( .C1(n19723), .C2(n19753), .A(n19722), .B(n19721), .ZN(
        P2_U3150) );
  AOI22_X1 U22751 ( .A1(n19725), .A2(n19856), .B1(n19854), .B2(n19724), .ZN(
        n19729) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n19858), .ZN(n19728) );
  OAI211_X1 U22753 ( .C1(n19777), .C2(n19753), .A(n19729), .B(n19728), .ZN(
        P2_U3151) );
  NOR2_X1 U22754 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19730), .ZN(n19731) );
  NAND2_X1 U22755 ( .A1(n19732), .A2(n19731), .ZN(n19735) );
  NAND2_X1 U22756 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19976), .ZN(n19969) );
  NAND2_X1 U22757 ( .A1(n19969), .A2(n19733), .ZN(n19734) );
  NAND2_X1 U22758 ( .A1(n19735), .A2(n19734), .ZN(n19740) );
  NOR2_X1 U22759 ( .A1(n19976), .A2(n19741), .ZN(n19786) );
  NOR2_X1 U22760 ( .A1(n19995), .A2(n19786), .ZN(n19736) );
  NAND2_X1 U22761 ( .A1(n19737), .A2(n19736), .ZN(n19743) );
  AND2_X1 U22762 ( .A1(n19743), .A2(n19738), .ZN(n19739) );
  OAI21_X1 U22763 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19741), .A(n19995), 
        .ZN(n19742) );
  AND2_X1 U22764 ( .A1(n19743), .A2(n19742), .ZN(n19772) );
  AOI22_X1 U22765 ( .A1(n19772), .A2(n19790), .B1(n19779), .B2(n19786), .ZN(
        n19749) );
  INV_X1 U22766 ( .A(n19744), .ZN(n19746) );
  AOI22_X1 U22767 ( .A1(n19773), .A2(n19747), .B1(n19801), .B2(n19780), .ZN(
        n19748) );
  OAI211_X1 U22768 ( .C1(n19771), .C2(n10604), .A(n19749), .B(n19748), .ZN(
        P2_U3152) );
  AOI22_X1 U22769 ( .A1(n19772), .A2(n19815), .B1(n19344), .B2(n19786), .ZN(
        n19752) );
  INV_X1 U22770 ( .A(n19771), .ZN(n19774) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19774), .B1(
        n19801), .B2(n19750), .ZN(n19751) );
  OAI211_X1 U22772 ( .C1(n19754), .C2(n19753), .A(n19752), .B(n19751), .ZN(
        P2_U3153) );
  AOI22_X1 U22773 ( .A1(n19772), .A2(n19821), .B1(n19820), .B2(n19786), .ZN(
        n19756) );
  AOI22_X1 U22774 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19774), .B1(
        n19773), .B2(n19822), .ZN(n19755) );
  OAI211_X1 U22775 ( .C1(n19798), .C2(n19813), .A(n19756), .B(n19755), .ZN(
        P2_U3154) );
  INV_X1 U22776 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U22777 ( .A1(n19772), .A2(n19828), .B1(n19827), .B2(n19786), .ZN(
        n19759) );
  AOI22_X1 U22778 ( .A1(n19773), .A2(n19829), .B1(n19801), .B2(n19757), .ZN(
        n19758) );
  OAI211_X1 U22779 ( .C1(n19771), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P2_U3155) );
  AOI22_X1 U22780 ( .A1(n19772), .A2(n19834), .B1(n19833), .B2(n19786), .ZN(
        n19762) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19774), .B1(
        n19773), .B2(n19835), .ZN(n19761) );
  OAI211_X1 U22782 ( .C1(n19839), .C2(n19813), .A(n19762), .B(n19761), .ZN(
        P2_U3156) );
  AOI22_X1 U22783 ( .A1(n19772), .A2(n19841), .B1(n19840), .B2(n19786), .ZN(
        n19765) );
  AOI22_X1 U22784 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19774), .B1(
        n19773), .B2(n19763), .ZN(n19764) );
  OAI211_X1 U22785 ( .C1(n19766), .C2(n19813), .A(n19765), .B(n19764), .ZN(
        P2_U3157) );
  AOI22_X1 U22786 ( .A1(n19772), .A2(n19847), .B1(n19846), .B2(n19786), .ZN(
        n19769) );
  AOI22_X1 U22787 ( .A1(n19773), .A2(n19767), .B1(n19801), .B2(n19848), .ZN(
        n19768) );
  OAI211_X1 U22788 ( .C1(n19771), .C2(n19770), .A(n19769), .B(n19768), .ZN(
        P2_U3158) );
  AOI22_X1 U22789 ( .A1(n19772), .A2(n19856), .B1(n19854), .B2(n19786), .ZN(
        n19776) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19774), .B1(
        n19773), .B2(n19858), .ZN(n19775) );
  OAI211_X1 U22791 ( .C1(n19777), .C2(n19813), .A(n19776), .B(n19775), .ZN(
        P2_U3159) );
  NOR2_X1 U22792 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19778), .ZN(
        n19808) );
  AOI22_X1 U22793 ( .A1(n19780), .A2(n19859), .B1(n19779), .B2(n19808), .ZN(
        n19792) );
  NOR3_X1 U22794 ( .A1(n11112), .A2(n19808), .A3(n19995), .ZN(n19785) );
  NOR2_X1 U22795 ( .A1(n19801), .A2(n19859), .ZN(n19782) );
  OAI21_X1 U22796 ( .B1(n19782), .B2(n19781), .A(n19942), .ZN(n19789) );
  AOI221_X1 U22797 ( .B1(n20000), .B2(n19789), .C1(n20000), .C2(n19786), .A(
        n19808), .ZN(n19783) );
  NOR2_X1 U22798 ( .A1(n19808), .A2(n19786), .ZN(n19788) );
  OAI21_X1 U22799 ( .B1(n11112), .B2(n19808), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19787) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19810), .B1(
        n19790), .B2(n19809), .ZN(n19791) );
  OAI211_X1 U22801 ( .C1(n19793), .C2(n19813), .A(n19792), .B(n19791), .ZN(
        P2_U3160) );
  AOI22_X1 U22802 ( .A1(n19816), .A2(n19801), .B1(n19344), .B2(n19808), .ZN(
        n19795) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19810), .B1(
        n19815), .B2(n19809), .ZN(n19794) );
  OAI211_X1 U22804 ( .C1(n19819), .C2(n19852), .A(n19795), .B(n19794), .ZN(
        P2_U3161) );
  AOI22_X1 U22805 ( .A1(n19822), .A2(n19801), .B1(n19820), .B2(n19808), .ZN(
        n19797) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19810), .B1(
        n19821), .B2(n19809), .ZN(n19796) );
  OAI211_X1 U22807 ( .C1(n19798), .C2(n19852), .A(n19797), .B(n19796), .ZN(
        P2_U3162) );
  AOI22_X1 U22808 ( .A1(n19829), .A2(n19801), .B1(n19827), .B2(n19808), .ZN(
        n19800) );
  AOI22_X1 U22809 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19810), .B1(
        n19828), .B2(n19809), .ZN(n19799) );
  OAI211_X1 U22810 ( .C1(n19832), .C2(n19852), .A(n19800), .B(n19799), .ZN(
        P2_U3163) );
  AOI22_X1 U22811 ( .A1(n19835), .A2(n19801), .B1(n19833), .B2(n19808), .ZN(
        n19803) );
  AOI22_X1 U22812 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19810), .B1(
        n19834), .B2(n19809), .ZN(n19802) );
  OAI211_X1 U22813 ( .C1(n19839), .C2(n19852), .A(n19803), .B(n19802), .ZN(
        P2_U3164) );
  AOI22_X1 U22814 ( .A1(n19842), .A2(n19859), .B1(n19840), .B2(n19808), .ZN(
        n19805) );
  AOI22_X1 U22815 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19810), .B1(
        n19841), .B2(n19809), .ZN(n19804) );
  OAI211_X1 U22816 ( .C1(n19845), .C2(n19813), .A(n19805), .B(n19804), .ZN(
        P2_U3165) );
  AOI22_X1 U22817 ( .A1(n19848), .A2(n19859), .B1(n19846), .B2(n19808), .ZN(
        n19807) );
  AOI22_X1 U22818 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19810), .B1(
        n19847), .B2(n19809), .ZN(n19806) );
  OAI211_X1 U22819 ( .C1(n19853), .C2(n19813), .A(n19807), .B(n19806), .ZN(
        P2_U3166) );
  AOI22_X1 U22820 ( .A1(n19860), .A2(n19859), .B1(n19854), .B2(n19808), .ZN(
        n19812) );
  AOI22_X1 U22821 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19810), .B1(
        n19856), .B2(n19809), .ZN(n19811) );
  OAI211_X1 U22822 ( .C1(n19814), .C2(n19813), .A(n19812), .B(n19811), .ZN(
        P2_U3167) );
  INV_X1 U22823 ( .A(n19861), .ZN(n19838) );
  AOI22_X1 U22824 ( .A1(n19857), .A2(n19815), .B1(n19855), .B2(n19344), .ZN(
        n19818) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19849), .B1(
        n19859), .B2(n19816), .ZN(n19817) );
  OAI211_X1 U22826 ( .C1(n19819), .C2(n19838), .A(n19818), .B(n19817), .ZN(
        P2_U3169) );
  INV_X1 U22827 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U22828 ( .A1(n19857), .A2(n19821), .B1(n19855), .B2(n19820), .ZN(
        n19825) );
  AOI22_X1 U22829 ( .A1(n19861), .A2(n19823), .B1(n19859), .B2(n19822), .ZN(
        n19824) );
  OAI211_X1 U22830 ( .C1(n19865), .C2(n19826), .A(n19825), .B(n19824), .ZN(
        P2_U3170) );
  AOI22_X1 U22831 ( .A1(n19857), .A2(n19828), .B1(n19855), .B2(n19827), .ZN(
        n19831) );
  AOI22_X1 U22832 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19849), .B1(
        n19859), .B2(n19829), .ZN(n19830) );
  OAI211_X1 U22833 ( .C1(n19832), .C2(n19838), .A(n19831), .B(n19830), .ZN(
        P2_U3171) );
  AOI22_X1 U22834 ( .A1(n19857), .A2(n19834), .B1(n19855), .B2(n19833), .ZN(
        n19837) );
  AOI22_X1 U22835 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19849), .B1(
        n19859), .B2(n19835), .ZN(n19836) );
  OAI211_X1 U22836 ( .C1(n19839), .C2(n19838), .A(n19837), .B(n19836), .ZN(
        P2_U3172) );
  AOI22_X1 U22837 ( .A1(n19857), .A2(n19841), .B1(n19855), .B2(n19840), .ZN(
        n19844) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19849), .B1(
        n19861), .B2(n19842), .ZN(n19843) );
  OAI211_X1 U22839 ( .C1(n19845), .C2(n19852), .A(n19844), .B(n19843), .ZN(
        P2_U3173) );
  AOI22_X1 U22840 ( .A1(n19857), .A2(n19847), .B1(n19855), .B2(n19846), .ZN(
        n19851) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19849), .B1(
        n19861), .B2(n19848), .ZN(n19850) );
  OAI211_X1 U22842 ( .C1(n19853), .C2(n19852), .A(n19851), .B(n19850), .ZN(
        P2_U3174) );
  INV_X1 U22843 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U22844 ( .A1(n19857), .A2(n19856), .B1(n19855), .B2(n19854), .ZN(
        n19863) );
  AOI22_X1 U22845 ( .A1(n19861), .A2(n19860), .B1(n19859), .B2(n19858), .ZN(
        n19862) );
  OAI211_X1 U22846 ( .C1(n19865), .C2(n19864), .A(n19863), .B(n19862), .ZN(
        P2_U3175) );
  AND2_X1 U22847 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19866), .ZN(
        P2_U3179) );
  AND2_X1 U22848 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19866), .ZN(
        P2_U3180) );
  AND2_X1 U22849 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19866), .ZN(
        P2_U3181) );
  AND2_X1 U22850 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19866), .ZN(
        P2_U3182) );
  AND2_X1 U22851 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19866), .ZN(
        P2_U3183) );
  AND2_X1 U22852 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19866), .ZN(
        P2_U3184) );
  AND2_X1 U22853 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19866), .ZN(
        P2_U3185) );
  AND2_X1 U22854 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19866), .ZN(
        P2_U3186) );
  AND2_X1 U22855 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19866), .ZN(
        P2_U3187) );
  AND2_X1 U22856 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19866), .ZN(
        P2_U3188) );
  AND2_X1 U22857 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19866), .ZN(
        P2_U3189) );
  AND2_X1 U22858 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19866), .ZN(
        P2_U3190) );
  AND2_X1 U22859 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19866), .ZN(
        P2_U3191) );
  AND2_X1 U22860 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19866), .ZN(
        P2_U3192) );
  AND2_X1 U22861 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19866), .ZN(
        P2_U3193) );
  AND2_X1 U22862 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19866), .ZN(
        P2_U3194) );
  AND2_X1 U22863 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19866), .ZN(
        P2_U3195) );
  AND2_X1 U22864 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19866), .ZN(
        P2_U3196) );
  AND2_X1 U22865 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19866), .ZN(
        P2_U3197) );
  AND2_X1 U22866 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19866), .ZN(
        P2_U3198) );
  AND2_X1 U22867 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19866), .ZN(
        P2_U3199) );
  AND2_X1 U22868 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19866), .ZN(
        P2_U3200) );
  AND2_X1 U22869 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19866), .ZN(P2_U3201) );
  AND2_X1 U22870 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19866), .ZN(P2_U3202) );
  AND2_X1 U22871 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19866), .ZN(P2_U3203) );
  AND2_X1 U22872 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19866), .ZN(P2_U3204) );
  AND2_X1 U22873 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19866), .ZN(P2_U3205) );
  AND2_X1 U22874 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19866), .ZN(P2_U3206) );
  AND2_X1 U22875 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19866), .ZN(P2_U3207) );
  AND2_X1 U22876 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19866), .ZN(P2_U3208) );
  INV_X1 U22877 ( .A(NA), .ZN(n19867) );
  OAI21_X1 U22878 ( .B1(n19867), .B2(n19873), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19883) );
  NAND2_X1 U22879 ( .A1(n19996), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19881) );
  NAND3_X1 U22880 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19881), .ZN(n19870) );
  AOI211_X1 U22881 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20902), .A(
        n20009), .B(n19868), .ZN(n19869) );
  AOI21_X1 U22882 ( .B1(n19883), .B2(n19870), .A(n19869), .ZN(n19871) );
  INV_X1 U22883 ( .A(n19871), .ZN(P2_U3209) );
  NOR2_X1 U22884 ( .A1(HOLD), .A2(n19872), .ZN(n19882) );
  OAI211_X1 U22885 ( .C1(n19882), .C2(n19884), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19873), .ZN(n19874) );
  AND3_X1 U22886 ( .A1(n19875), .A2(n19881), .A3(n19874), .ZN(n19876) );
  OAI21_X1 U22887 ( .B1(n20902), .B2(n19877), .A(n19876), .ZN(P2_U3210) );
  OAI22_X1 U22888 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19878), .B1(NA), 
        .B2(n19881), .ZN(n19879) );
  OAI211_X1 U22889 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19879), .ZN(n19880) );
  OAI221_X1 U22890 ( .B1(n19883), .B2(n19882), .C1(n19883), .C2(n19881), .A(
        n19880), .ZN(P2_U3211) );
  OAI222_X1 U22891 ( .A1(n19926), .A2(n19885), .B1(n21094), .B2(n20009), .C1(
        n10439), .C2(n19923), .ZN(P2_U3212) );
  OAI222_X1 U22892 ( .A1(n19926), .A2(n10663), .B1(n19886), .B2(n20009), .C1(
        n19885), .C2(n19923), .ZN(P2_U3213) );
  OAI222_X1 U22893 ( .A1(n19926), .A2(n10694), .B1(n19887), .B2(n20009), .C1(
        n10663), .C2(n19923), .ZN(P2_U3214) );
  OAI222_X1 U22894 ( .A1(n19926), .A2(n15751), .B1(n19888), .B2(n20009), .C1(
        n10694), .C2(n19923), .ZN(P2_U3215) );
  OAI222_X1 U22895 ( .A1(n19926), .A2(n10473), .B1(n19889), .B2(n20009), .C1(
        n15751), .C2(n19923), .ZN(P2_U3216) );
  OAI222_X1 U22896 ( .A1(n19926), .A2(n10477), .B1(n19890), .B2(n20009), .C1(
        n10473), .C2(n19923), .ZN(P2_U3217) );
  OAI222_X1 U22897 ( .A1(n19926), .A2(n10481), .B1(n19891), .B2(n20009), .C1(
        n10477), .C2(n19923), .ZN(P2_U3218) );
  OAI222_X1 U22898 ( .A1(n19926), .A2(n15464), .B1(n19892), .B2(n20009), .C1(
        n10481), .C2(n19923), .ZN(P2_U3219) );
  OAI222_X1 U22899 ( .A1(n19926), .A2(n10489), .B1(n19893), .B2(n20009), .C1(
        n15464), .C2(n19923), .ZN(P2_U3220) );
  OAI222_X1 U22900 ( .A1(n19926), .A2(n10808), .B1(n19894), .B2(n20009), .C1(
        n10489), .C2(n19923), .ZN(P2_U3221) );
  OAI222_X1 U22901 ( .A1(n19926), .A2(n10827), .B1(n19895), .B2(n20009), .C1(
        n10808), .C2(n19923), .ZN(P2_U3222) );
  OAI222_X1 U22902 ( .A1(n19926), .A2(n10842), .B1(n19896), .B2(n20009), .C1(
        n10827), .C2(n19923), .ZN(P2_U3223) );
  OAI222_X1 U22903 ( .A1(n19926), .A2(n10855), .B1(n19897), .B2(n20009), .C1(
        n10842), .C2(n19923), .ZN(P2_U3224) );
  OAI222_X1 U22904 ( .A1(n19926), .A2(n19899), .B1(n19898), .B2(n20009), .C1(
        n10855), .C2(n19923), .ZN(P2_U3225) );
  OAI222_X1 U22905 ( .A1(n19926), .A2(n10870), .B1(n19900), .B2(n20009), .C1(
        n19899), .C2(n19923), .ZN(P2_U3226) );
  OAI222_X1 U22906 ( .A1(n19926), .A2(n19902), .B1(n19901), .B2(n20009), .C1(
        n10870), .C2(n19923), .ZN(P2_U3227) );
  OAI222_X1 U22907 ( .A1(n19926), .A2(n19904), .B1(n19903), .B2(n20009), .C1(
        n19902), .C2(n19923), .ZN(P2_U3228) );
  OAI222_X1 U22908 ( .A1(n19926), .A2(n19906), .B1(n19905), .B2(n20009), .C1(
        n19904), .C2(n19923), .ZN(P2_U3229) );
  OAI222_X1 U22909 ( .A1(n19926), .A2(n19908), .B1(n19907), .B2(n20009), .C1(
        n19906), .C2(n19923), .ZN(P2_U3230) );
  OAI222_X1 U22910 ( .A1(n19926), .A2(n19910), .B1(n19909), .B2(n20009), .C1(
        n19908), .C2(n19923), .ZN(P2_U3231) );
  OAI222_X1 U22911 ( .A1(n19926), .A2(n15361), .B1(n19911), .B2(n20009), .C1(
        n19910), .C2(n19923), .ZN(P2_U3232) );
  OAI222_X1 U22912 ( .A1(n19926), .A2(n19913), .B1(n19912), .B2(n20009), .C1(
        n15361), .C2(n19923), .ZN(P2_U3233) );
  OAI222_X1 U22913 ( .A1(n19926), .A2(n15336), .B1(n19914), .B2(n20009), .C1(
        n19913), .C2(n19923), .ZN(P2_U3234) );
  OAI222_X1 U22914 ( .A1(n19926), .A2(n19916), .B1(n19915), .B2(n20009), .C1(
        n15336), .C2(n19923), .ZN(P2_U3235) );
  OAI222_X1 U22915 ( .A1(n19926), .A2(n19918), .B1(n19917), .B2(n20009), .C1(
        n19916), .C2(n19923), .ZN(P2_U3236) );
  OAI222_X1 U22916 ( .A1(n19926), .A2(n19919), .B1(n21027), .B2(n20009), .C1(
        n19918), .C2(n19923), .ZN(P2_U3237) );
  OAI222_X1 U22917 ( .A1(n19923), .A2(n19919), .B1(n21236), .B2(n20009), .C1(
        n10552), .C2(n19926), .ZN(P2_U3238) );
  OAI222_X1 U22918 ( .A1(n19926), .A2(n19921), .B1(n19920), .B2(n20009), .C1(
        n10552), .C2(n19923), .ZN(P2_U3239) );
  INV_X1 U22919 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19924) );
  OAI222_X1 U22920 ( .A1(n19926), .A2(n19924), .B1(n19922), .B2(n20009), .C1(
        n19921), .C2(n19923), .ZN(P2_U3240) );
  OAI222_X1 U22921 ( .A1(n19926), .A2(n16332), .B1(n19925), .B2(n20009), .C1(
        n19924), .C2(n19923), .ZN(P2_U3241) );
  INV_X1 U22922 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U22923 ( .A1(n20009), .A2(n19928), .B1(n19927), .B2(n20007), .ZN(
        P2_U3585) );
  MUX2_X1 U22924 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20009), .Z(P2_U3586) );
  INV_X1 U22925 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U22926 ( .A1(n20009), .A2(n19930), .B1(n19929), .B2(n20007), .ZN(
        P2_U3587) );
  INV_X1 U22927 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U22928 ( .A1(n20009), .A2(n19932), .B1(n19931), .B2(n20007), .ZN(
        P2_U3588) );
  OAI21_X1 U22929 ( .B1(n19936), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19934), 
        .ZN(n19933) );
  INV_X1 U22930 ( .A(n19933), .ZN(P2_U3591) );
  OAI21_X1 U22931 ( .B1(n19936), .B2(n19935), .A(n19934), .ZN(P2_U3592) );
  INV_X1 U22932 ( .A(n19944), .ZN(n19938) );
  AND2_X1 U22933 ( .A1(n19942), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19939) );
  INV_X1 U22934 ( .A(n19939), .ZN(n19964) );
  NOR3_X1 U22935 ( .A1(n19938), .A2(n19937), .A3(n19964), .ZN(n19947) );
  AND2_X1 U22936 ( .A1(n19940), .A2(n19939), .ZN(n19955) );
  INV_X1 U22937 ( .A(n19955), .ZN(n19945) );
  NAND2_X1 U22938 ( .A1(n19963), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19943) );
  AOI21_X1 U22939 ( .B1(n19943), .B2(n19942), .A(n19941), .ZN(n19952) );
  AOI21_X1 U22940 ( .B1(n19945), .B2(n19952), .A(n19944), .ZN(n19946) );
  AOI211_X1 U22941 ( .C1(n19948), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19947), 
        .B(n19946), .ZN(n19949) );
  AOI22_X1 U22942 ( .A1(n19977), .A2(n19950), .B1(n19949), .B2(n19974), .ZN(
        P2_U3602) );
  OAI22_X1 U22943 ( .A1(n19953), .A2(n19952), .B1(n19951), .B2(n20000), .ZN(
        n19954) );
  INV_X1 U22944 ( .A(n19954), .ZN(n19957) );
  NOR2_X1 U22945 ( .A1(n19977), .A2(n19955), .ZN(n19956) );
  AOI22_X1 U22946 ( .A1(n19958), .A2(n19977), .B1(n19957), .B2(n19956), .ZN(
        P2_U3603) );
  INV_X1 U22947 ( .A(n19959), .ZN(n19970) );
  OR3_X1 U22948 ( .A1(n19961), .A2(n19970), .A3(n19960), .ZN(n19962) );
  OAI21_X1 U22949 ( .B1(n19964), .B2(n19963), .A(n19962), .ZN(n19965) );
  AOI21_X1 U22950 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19966), .A(n19965), 
        .ZN(n19967) );
  AOI22_X1 U22951 ( .A1(n19977), .A2(n19968), .B1(n19967), .B2(n19974), .ZN(
        P2_U3604) );
  OAI21_X1 U22952 ( .B1(n19971), .B2(n19970), .A(n19969), .ZN(n19972) );
  AOI21_X1 U22953 ( .B1(n19973), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19972), 
        .ZN(n19975) );
  AOI22_X1 U22954 ( .A1(n19977), .A2(n19976), .B1(n19975), .B2(n19974), .ZN(
        P2_U3605) );
  INV_X1 U22955 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19978) );
  AOI22_X1 U22956 ( .A1(n20009), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19978), 
        .B2(n20007), .ZN(P2_U3608) );
  INV_X1 U22957 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19988) );
  INV_X1 U22958 ( .A(n19979), .ZN(n19987) );
  AOI22_X1 U22959 ( .A1(n19983), .A2(n19982), .B1(n19981), .B2(n19980), .ZN(
        n19986) );
  NOR2_X1 U22960 ( .A1(n19987), .A2(n19984), .ZN(n19985) );
  AOI22_X1 U22961 ( .A1(n19988), .A2(n19987), .B1(n19986), .B2(n19985), .ZN(
        P2_U3609) );
  OAI21_X1 U22962 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19990), .A(n19989), 
        .ZN(n19992) );
  NAND3_X1 U22963 ( .A1(n19992), .A2(n19991), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19998) );
  INV_X1 U22964 ( .A(n19993), .ZN(n19994) );
  OAI21_X1 U22965 ( .B1(n19996), .B2(n19995), .A(n19994), .ZN(n19997) );
  NAND2_X1 U22966 ( .A1(n19998), .A2(n19997), .ZN(n20006) );
  AOI22_X1 U22967 ( .A1(n20002), .A2(n20001), .B1(n20000), .B2(n19999), .ZN(
        n20004) );
  NAND2_X1 U22968 ( .A1(n20004), .A2(n20003), .ZN(n20005) );
  MUX2_X1 U22969 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n20006), .S(n20005), 
        .Z(P2_U3610) );
  INV_X1 U22970 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20008) );
  AOI22_X1 U22971 ( .A1(n20009), .A2(n21020), .B1(n20008), .B2(n20007), .ZN(
        P2_U3611) );
  AOI21_X1 U22972 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20905), .A(n20897), 
        .ZN(n20900) );
  INV_X1 U22973 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20010) );
  OR2_X1 U22974 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20894), .ZN(n20974) );
  INV_X2 U22975 ( .A(n20974), .ZN(n20988) );
  AOI21_X1 U22976 ( .B1(n20900), .B2(n20010), .A(n20988), .ZN(P1_U2802) );
  INV_X1 U22977 ( .A(n20011), .ZN(n20013) );
  OAI21_X1 U22978 ( .B1(n20013), .B2(n20012), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20014) );
  OAI21_X1 U22979 ( .B1(n20015), .B2(n20885), .A(n20014), .ZN(P1_U2803) );
  NOR2_X1 U22980 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20017) );
  OAI21_X1 U22981 ( .B1(n20017), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20974), .ZN(
        n20016) );
  OAI21_X1 U22982 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20974), .A(n20016), 
        .ZN(P1_U2804) );
  NOR2_X1 U22983 ( .A1(n20988), .A2(n20900), .ZN(n20965) );
  OAI21_X1 U22984 ( .B1(BS16), .B2(n20017), .A(n20965), .ZN(n20963) );
  OAI21_X1 U22985 ( .B1(n20965), .B2(n20789), .A(n20963), .ZN(P1_U2805) );
  INV_X1 U22986 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22987 ( .B1(n20019), .B2(n20018), .A(n20198), .ZN(P1_U2806) );
  NOR4_X1 U22988 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20023) );
  NOR4_X1 U22989 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20022) );
  NOR4_X1 U22990 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20021) );
  NOR4_X1 U22991 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20020) );
  NAND4_X1 U22992 ( .A1(n20023), .A2(n20022), .A3(n20021), .A4(n20020), .ZN(
        n20029) );
  NOR4_X1 U22993 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20027) );
  AOI211_X1 U22994 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_9__SCAN_IN), .B(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20026) );
  NOR4_X1 U22995 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20025) );
  NOR4_X1 U22996 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20024) );
  NAND4_X1 U22997 ( .A1(n20027), .A2(n20026), .A3(n20025), .A4(n20024), .ZN(
        n20028) );
  NOR2_X1 U22998 ( .A1(n20029), .A2(n20028), .ZN(n20970) );
  INV_X1 U22999 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20958) );
  NOR3_X1 U23000 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20031) );
  OAI21_X1 U23001 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20031), .A(n20970), .ZN(
        n20030) );
  OAI21_X1 U23002 ( .B1(n20970), .B2(n20958), .A(n20030), .ZN(P1_U2807) );
  INV_X1 U23003 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20964) );
  AOI21_X1 U23004 ( .B1(n20966), .B2(n20964), .A(n20031), .ZN(n20032) );
  INV_X1 U23005 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20955) );
  INV_X1 U23006 ( .A(n20970), .ZN(n20972) );
  AOI22_X1 U23007 ( .A1(n20970), .A2(n20032), .B1(n20955), .B2(n20972), .ZN(
        P1_U2808) );
  AOI22_X1 U23008 ( .A1(n20033), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20071), 
        .B2(P1_EBX_REG_9__SCAN_IN), .ZN(n20034) );
  OAI21_X1 U23009 ( .B1(n20061), .B2(n20035), .A(n20034), .ZN(n20036) );
  AOI211_X1 U23010 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20050), .B(n20036), .ZN(n20044) );
  INV_X1 U23011 ( .A(n20037), .ZN(n20040) );
  AOI22_X1 U23012 ( .A1(n20040), .A2(n20066), .B1(n20039), .B2(n20038), .ZN(
        n20043) );
  INV_X1 U23013 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21146) );
  NAND3_X1 U23014 ( .A1(n20041), .A2(n20074), .A3(n21146), .ZN(n20042) );
  NAND3_X1 U23015 ( .A1(n20044), .A2(n20043), .A3(n20042), .ZN(P1_U2831) );
  INV_X1 U23016 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21198) );
  INV_X1 U23017 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20914) );
  NOR2_X1 U23018 ( .A1(n21198), .A2(n20914), .ZN(n20053) );
  OAI21_X1 U23019 ( .B1(n20046), .B2(n20053), .A(n20045), .ZN(n20067) );
  AOI22_X1 U23020 ( .A1(n20067), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20071), 
        .B2(P1_EBX_REG_7__SCAN_IN), .ZN(n20047) );
  OAI21_X1 U23021 ( .B1(n20061), .B2(n20048), .A(n20047), .ZN(n20049) );
  AOI211_X1 U23022 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20050), .B(n20049), .ZN(n20058) );
  INV_X1 U23023 ( .A(n20052), .ZN(n20056) );
  INV_X1 U23024 ( .A(n20053), .ZN(n20054) );
  NOR2_X1 U23025 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20054), .ZN(n20055) );
  AOI22_X1 U23026 ( .A1(n20056), .A2(n20066), .B1(n20074), .B2(n20055), .ZN(
        n20057) );
  OAI211_X1 U23027 ( .C1(n20059), .C2(n20107), .A(n20058), .B(n20057), .ZN(
        P1_U2833) );
  NOR2_X1 U23028 ( .A1(n20061), .A2(n20060), .ZN(n20065) );
  NAND2_X1 U23029 ( .A1(n20071), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n20062) );
  OAI211_X1 U23030 ( .C1(n20093), .C2(n20063), .A(n20062), .B(n20091), .ZN(
        n20064) );
  AOI211_X1 U23031 ( .C1(n20109), .C2(n20066), .A(n20065), .B(n20064), .ZN(
        n20069) );
  NOR2_X1 U23032 ( .A1(n20103), .A2(n21198), .ZN(n20075) );
  OAI21_X1 U23033 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20075), .A(n20067), .ZN(
        n20068) );
  OAI211_X1 U23034 ( .C1(n20107), .C2(n20070), .A(n20069), .B(n20068), .ZN(
        P1_U2834) );
  NAND2_X1 U23035 ( .A1(n20071), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20072) );
  OAI211_X1 U23036 ( .C1(n20093), .C2(n20073), .A(n20072), .B(n20091), .ZN(
        n20078) );
  INV_X1 U23037 ( .A(n20074), .ZN(n20076) );
  AOI21_X1 U23038 ( .B1(n20076), .B2(n21198), .A(n20075), .ZN(n20077) );
  AOI211_X1 U23039 ( .C1(n20099), .C2(n20079), .A(n20078), .B(n20077), .ZN(
        n20080) );
  INV_X1 U23040 ( .A(n20080), .ZN(n20081) );
  AOI21_X1 U23041 ( .B1(n20104), .B2(n20082), .A(n20081), .ZN(n20083) );
  OAI21_X1 U23042 ( .B1(n20084), .B2(n20107), .A(n20083), .ZN(P1_U2835) );
  NAND2_X1 U23043 ( .A1(n20086), .A2(n20085), .ZN(n20089) );
  INV_X1 U23044 ( .A(n20087), .ZN(n20088) );
  NAND2_X1 U23045 ( .A1(n20089), .A2(n20088), .ZN(n20090) );
  AND2_X1 U23046 ( .A1(n20090), .A2(n13990), .ZN(n20203) );
  OAI21_X1 U23047 ( .B1(n20093), .B2(n20092), .A(n20091), .ZN(n20098) );
  OAI22_X1 U23048 ( .A1(n20096), .A2(n20095), .B1(n21063), .B2(n20094), .ZN(
        n20097) );
  AOI211_X1 U23049 ( .C1(n20099), .C2(n20203), .A(n20098), .B(n20097), .ZN(
        n20106) );
  OAI21_X1 U23050 ( .B1(n20101), .B2(n20100), .A(n20910), .ZN(n20102) );
  AOI22_X1 U23051 ( .A1(n20104), .A2(n20175), .B1(n20103), .B2(n20102), .ZN(
        n20105) );
  OAI211_X1 U23052 ( .C1(n20178), .C2(n20107), .A(n20106), .B(n20105), .ZN(
        P1_U2836) );
  AOI22_X1 U23053 ( .A1(n20109), .A2(n20113), .B1(n20112), .B2(n20108), .ZN(
        n20110) );
  OAI21_X1 U23054 ( .B1(n20115), .B2(n20111), .A(n20110), .ZN(P1_U2866) );
  AOI22_X1 U23055 ( .A1(n20175), .A2(n20113), .B1(n20112), .B2(n20203), .ZN(
        n20114) );
  OAI21_X1 U23056 ( .B1(n20115), .B2(n21063), .A(n20114), .ZN(P1_U2868) );
  AOI22_X1 U23057 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20119), .B1(n20132), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20116) );
  OAI21_X1 U23058 ( .B1(n20118), .B2(n20117), .A(n20116), .ZN(P1_U2921) );
  AOI22_X1 U23059 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20120) );
  OAI21_X1 U23060 ( .B1(n14845), .B2(n20142), .A(n20120), .ZN(P1_U2922) );
  INV_X1 U23061 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U23062 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U23063 ( .B1(n20122), .B2(n20142), .A(n20121), .ZN(P1_U2923) );
  AOI22_X1 U23064 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20123) );
  OAI21_X1 U23065 ( .B1(n14855), .B2(n20142), .A(n20123), .ZN(P1_U2924) );
  AOI22_X1 U23066 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20124) );
  OAI21_X1 U23067 ( .B1(n21189), .B2(n20142), .A(n20124), .ZN(P1_U2925) );
  AOI22_X1 U23068 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20125) );
  OAI21_X1 U23069 ( .B1(n14862), .B2(n20142), .A(n20125), .ZN(P1_U2926) );
  AOI22_X1 U23070 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20126) );
  OAI21_X1 U23071 ( .B1(n14240), .B2(n20142), .A(n20126), .ZN(P1_U2927) );
  AOI22_X1 U23072 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20127) );
  OAI21_X1 U23073 ( .B1(n14232), .B2(n20142), .A(n20127), .ZN(P1_U2928) );
  AOI22_X1 U23074 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20128) );
  OAI21_X1 U23075 ( .B1(n12102), .B2(n20142), .A(n20128), .ZN(P1_U2929) );
  AOI22_X1 U23076 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20129) );
  OAI21_X1 U23077 ( .B1(n14235), .B2(n20142), .A(n20129), .ZN(P1_U2930) );
  AOI22_X1 U23078 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20130) );
  OAI21_X1 U23079 ( .B1(n20131), .B2(n20142), .A(n20130), .ZN(P1_U2931) );
  AOI22_X1 U23080 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20979), .B1(n20132), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20133) );
  OAI21_X1 U23081 ( .B1(n14141), .B2(n20142), .A(n20133), .ZN(P1_U2932) );
  AOI22_X1 U23082 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20134) );
  OAI21_X1 U23083 ( .B1(n20135), .B2(n20142), .A(n20134), .ZN(P1_U2933) );
  AOI22_X1 U23084 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20136) );
  OAI21_X1 U23085 ( .B1(n20137), .B2(n20142), .A(n20136), .ZN(P1_U2934) );
  AOI22_X1 U23086 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20138) );
  OAI21_X1 U23087 ( .B1(n20139), .B2(n20142), .A(n20138), .ZN(P1_U2935) );
  AOI22_X1 U23088 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20979), .B1(n20140), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20141) );
  OAI21_X1 U23089 ( .B1(n20143), .B2(n20142), .A(n20141), .ZN(P1_U2936) );
  AOI22_X1 U23090 ( .A1(n20168), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20144), .ZN(n20147) );
  INV_X1 U23091 ( .A(n20145), .ZN(n20146) );
  NAND2_X1 U23092 ( .A1(n20155), .A2(n20146), .ZN(n20157) );
  NAND2_X1 U23093 ( .A1(n20147), .A2(n20157), .ZN(P1_U2945) );
  AOI22_X1 U23094 ( .A1(n20168), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20167), .ZN(n20150) );
  INV_X1 U23095 ( .A(n20148), .ZN(n20149) );
  NAND2_X1 U23096 ( .A1(n20155), .A2(n20149), .ZN(n20163) );
  NAND2_X1 U23097 ( .A1(n20150), .A2(n20163), .ZN(P1_U2949) );
  AOI22_X1 U23098 ( .A1(n20168), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20167), .ZN(n20152) );
  NAND2_X1 U23099 ( .A1(n20155), .A2(n20151), .ZN(n20165) );
  NAND2_X1 U23100 ( .A1(n20152), .A2(n20165), .ZN(P1_U2950) );
  AOI22_X1 U23101 ( .A1(n20168), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20167), .ZN(n20156) );
  INV_X1 U23102 ( .A(n20153), .ZN(n20154) );
  NAND2_X1 U23103 ( .A1(n20155), .A2(n20154), .ZN(n20169) );
  NAND2_X1 U23104 ( .A1(n20156), .A2(n20169), .ZN(P1_U2951) );
  AOI22_X1 U23105 ( .A1(n20168), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20144), .ZN(n20158) );
  NAND2_X1 U23106 ( .A1(n20158), .A2(n20157), .ZN(P1_U2960) );
  AOI22_X1 U23107 ( .A1(n20168), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20167), .ZN(n20160) );
  NAND2_X1 U23108 ( .A1(n20160), .A2(n20159), .ZN(P1_U2961) );
  AOI22_X1 U23109 ( .A1(n20168), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20144), .ZN(n20162) );
  NAND2_X1 U23110 ( .A1(n20162), .A2(n20161), .ZN(P1_U2962) );
  AOI22_X1 U23111 ( .A1(n20168), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20167), .ZN(n20164) );
  NAND2_X1 U23112 ( .A1(n20164), .A2(n20163), .ZN(P1_U2964) );
  AOI22_X1 U23113 ( .A1(n20168), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20144), .ZN(n20166) );
  NAND2_X1 U23114 ( .A1(n20166), .A2(n20165), .ZN(P1_U2965) );
  AOI22_X1 U23115 ( .A1(n20168), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20167), .ZN(n20170) );
  NAND2_X1 U23116 ( .A1(n20170), .A2(n20169), .ZN(P1_U2966) );
  AOI22_X1 U23117 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20177) );
  OAI21_X1 U23118 ( .B1(n20173), .B2(n20172), .A(n9810), .ZN(n20174) );
  INV_X1 U23119 ( .A(n20174), .ZN(n20206) );
  AOI22_X1 U23120 ( .A1(n20206), .A2(n20186), .B1(n20194), .B2(n20175), .ZN(
        n20176) );
  OAI211_X1 U23121 ( .C1(n20179), .C2(n20178), .A(n20177), .B(n20176), .ZN(
        P1_U2995) );
  AOI22_X1 U23122 ( .A1(n20180), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20236), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20188) );
  OAI21_X1 U23123 ( .B1(n20182), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20181), .ZN(n20183) );
  INV_X1 U23124 ( .A(n20183), .ZN(n20244) );
  INV_X1 U23125 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20184) );
  AOI22_X1 U23126 ( .A1(n20244), .A2(n20186), .B1(n20185), .B2(n20184), .ZN(
        n20187) );
  OAI211_X1 U23127 ( .C1(n20258), .C2(n20189), .A(n20188), .B(n20187), .ZN(
        P1_U2998) );
  NAND2_X1 U23128 ( .A1(n20191), .A2(n20190), .ZN(n20192) );
  AOI22_X1 U23129 ( .A1(n20194), .A2(n20193), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20192), .ZN(n20196) );
  OAI211_X1 U23130 ( .C1(n20198), .C2(n20197), .A(n20196), .B(n20195), .ZN(
        P1_U2999) );
  AOI21_X1 U23131 ( .B1(n20201), .B2(n20200), .A(n20199), .ZN(n20202) );
  INV_X1 U23132 ( .A(n20202), .ZN(n20209) );
  AOI22_X1 U23133 ( .A1(n20236), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n20238), 
        .B2(n20203), .ZN(n20208) );
  OAI21_X1 U23134 ( .B1(n20223), .B2(n20205), .A(n20204), .ZN(n20213) );
  AOI22_X1 U23135 ( .A1(n20206), .A2(n20243), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20213), .ZN(n20207) );
  OAI211_X1 U23136 ( .C1(n20216), .C2(n20209), .A(n20208), .B(n20207), .ZN(
        P1_U3027) );
  AOI22_X1 U23137 ( .A1(n20236), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20238), 
        .B2(n20210), .ZN(n20215) );
  INV_X1 U23138 ( .A(n20211), .ZN(n20212) );
  AOI22_X1 U23139 ( .A1(n20213), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20212), .B2(n20243), .ZN(n20214) );
  OAI211_X1 U23140 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20216), .A(
        n20215), .B(n20214), .ZN(P1_U3028) );
  NAND2_X1 U23141 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20217), .ZN(
        n20234) );
  AOI21_X1 U23142 ( .B1(n20247), .B2(n20219), .A(n20218), .ZN(n20233) );
  INV_X1 U23143 ( .A(n20220), .ZN(n20229) );
  NAND3_X1 U23144 ( .A1(n20221), .A2(n13794), .A3(n20243), .ZN(n20228) );
  AND2_X1 U23145 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20222) );
  NAND2_X1 U23146 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20222), .ZN(
        n20224) );
  NAND2_X1 U23147 ( .A1(n20224), .A2(n20223), .ZN(n20225) );
  AOI22_X1 U23148 ( .A1(n20226), .A2(n20225), .B1(n20236), .B2(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20227) );
  OAI211_X1 U23149 ( .C1(n20230), .C2(n20229), .A(n20228), .B(n20227), .ZN(
        n20231) );
  INV_X1 U23150 ( .A(n20231), .ZN(n20232) );
  OAI221_X1 U23151 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20234), .C1(
        n21112), .C2(n20233), .A(n20232), .ZN(P1_U3029) );
  INV_X1 U23152 ( .A(n20235), .ZN(n20237) );
  AOI22_X1 U23153 ( .A1(n20238), .A2(n20237), .B1(n20236), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20246) );
  AOI211_X1 U23154 ( .C1(n20241), .C2(n20240), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n20239), .ZN(n20242) );
  AOI21_X1 U23155 ( .B1(n20244), .B2(n20243), .A(n20242), .ZN(n20245) );
  OAI211_X1 U23156 ( .C1(n20248), .C2(n20247), .A(n20246), .B(n20245), .ZN(
        P1_U3030) );
  NOR2_X1 U23157 ( .A1(n20250), .A2(n20249), .ZN(P1_U3032) );
  INV_X1 U23158 ( .A(n20608), .ZN(n20552) );
  OR2_X1 U23159 ( .A1(n20551), .A2(n20552), .ZN(n20429) );
  NAND2_X1 U23160 ( .A1(n20265), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20788) );
  NAND2_X1 U23161 ( .A1(n20324), .A2(n20788), .ZN(n20555) );
  INV_X1 U23162 ( .A(n13828), .ZN(n20251) );
  OR2_X1 U23163 ( .A1(n13831), .A2(n12686), .ZN(n20548) );
  OAI21_X1 U23164 ( .B1(n20345), .B2(n20862), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20253) );
  NAND2_X1 U23165 ( .A1(n20253), .A2(n20829), .ZN(n20267) );
  INV_X1 U23166 ( .A(n20690), .ZN(n20254) );
  OR2_X1 U23167 ( .A1(n20549), .A2(n20254), .ZN(n20392) );
  OR2_X1 U23168 ( .A1(n20392), .A2(n20791), .ZN(n20266) );
  INV_X1 U23169 ( .A(n20266), .ZN(n20255) );
  NAND3_X1 U23170 ( .A1(n20652), .A2(n20611), .A3(n20693), .ZN(n20323) );
  NOR2_X1 U23171 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20323), .ZN(
        n20262) );
  OAI22_X1 U23172 ( .A1(n20267), .A2(n20255), .B1(n20262), .B2(n20701), .ZN(
        n20256) );
  AOI211_X2 U23173 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20429), .A(n20555), 
        .B(n20256), .ZN(n20315) );
  NOR2_X2 U23174 ( .A1(n20258), .A2(n20257), .ZN(n20310) );
  NOR2_X2 U23175 ( .A1(n20259), .A2(n20258), .ZN(n20311) );
  AOI22_X1 U23176 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20310), .B1(DATAI_24_), 
        .B2(n20311), .ZN(n20387) );
  NAND2_X1 U23177 ( .A1(n20312), .A2(n20261), .ZN(n20694) );
  INV_X1 U23178 ( .A(n20262), .ZN(n20313) );
  OAI22_X1 U23179 ( .A1(n20882), .A2(n20387), .B1(n20694), .B2(n20313), .ZN(
        n20263) );
  INV_X1 U23180 ( .A(n20263), .ZN(n20270) );
  NOR2_X2 U23181 ( .A1(n20264), .A2(n20432), .ZN(n20820) );
  NOR2_X1 U23182 ( .A1(n20265), .A2(n20888), .ZN(n20610) );
  INV_X1 U23183 ( .A(n20610), .ZN(n20554) );
  OAI22_X1 U23184 ( .A1(n20267), .A2(n20266), .B1(n20554), .B2(n20429), .ZN(
        n20317) );
  INV_X1 U23185 ( .A(n20834), .ZN(n20268) );
  AOI22_X1 U23186 ( .A1(n20820), .A2(n20317), .B1(n20345), .B2(n20268), .ZN(
        n20269) );
  OAI211_X1 U23187 ( .C1(n20315), .C2(n20271), .A(n20270), .B(n20269), .ZN(
        P1_U3033) );
  NAND2_X1 U23188 ( .A1(n20312), .A2(n20272), .ZN(n20706) );
  OAI22_X1 U23189 ( .A1(n20882), .A2(n20840), .B1(n20706), .B2(n20313), .ZN(
        n20273) );
  INV_X1 U23190 ( .A(n20273), .ZN(n20277) );
  NOR2_X2 U23191 ( .A1(n20274), .A2(n20432), .ZN(n20836) );
  INV_X1 U23192 ( .A(DATAI_17_), .ZN(n21017) );
  INV_X1 U23193 ( .A(n20311), .ZN(n20298) );
  INV_X1 U23194 ( .A(n20310), .ZN(n20300) );
  AOI22_X1 U23195 ( .A1(n20836), .A2(n20317), .B1(n20345), .B2(n20837), .ZN(
        n20276) );
  OAI211_X1 U23196 ( .C1(n20315), .C2(n12124), .A(n20277), .B(n20276), .ZN(
        P1_U3034) );
  NAND2_X1 U23197 ( .A1(n20312), .A2(n20278), .ZN(n20713) );
  OAI22_X1 U23198 ( .A1(n20882), .A2(n20846), .B1(n20713), .B2(n20313), .ZN(
        n20279) );
  INV_X1 U23199 ( .A(n20279), .ZN(n20282) );
  NOR2_X2 U23200 ( .A1(n20280), .A2(n20432), .ZN(n20842) );
  AOI22_X1 U23201 ( .A1(DATAI_18_), .A2(n20311), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20310), .ZN(n20714) );
  INV_X1 U23202 ( .A(n20714), .ZN(n20843) );
  AOI22_X1 U23203 ( .A1(n20842), .A2(n20317), .B1(n20345), .B2(n20843), .ZN(
        n20281) );
  OAI211_X1 U23204 ( .C1(n20315), .C2(n20283), .A(n20282), .B(n20281), .ZN(
        P1_U3035) );
  NAND2_X1 U23205 ( .A1(n20312), .A2(n20284), .ZN(n20720) );
  OAI22_X1 U23206 ( .A1(n20882), .A2(n20852), .B1(n20720), .B2(n20313), .ZN(
        n20285) );
  INV_X1 U23207 ( .A(n20285), .ZN(n20288) );
  NOR2_X2 U23208 ( .A1(n20286), .A2(n20432), .ZN(n20848) );
  AOI22_X1 U23209 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20310), .B1(DATAI_19_), 
        .B2(n20311), .ZN(n20721) );
  INV_X1 U23210 ( .A(n20721), .ZN(n20849) );
  AOI22_X1 U23211 ( .A1(n20848), .A2(n20317), .B1(n20345), .B2(n20849), .ZN(
        n20287) );
  OAI211_X1 U23212 ( .C1(n20315), .C2(n12167), .A(n20288), .B(n20287), .ZN(
        P1_U3036) );
  INV_X1 U23213 ( .A(DATAI_28_), .ZN(n20289) );
  INV_X1 U23214 ( .A(n20855), .ZN(n20631) );
  NAND2_X1 U23215 ( .A1(n20312), .A2(n11823), .ZN(n20727) );
  OAI22_X1 U23216 ( .A1(n20882), .A2(n20631), .B1(n20727), .B2(n20313), .ZN(
        n20291) );
  INV_X1 U23217 ( .A(n20291), .ZN(n20294) );
  NOR2_X2 U23218 ( .A1(n20292), .A2(n20432), .ZN(n20854) );
  INV_X1 U23219 ( .A(n20858), .ZN(n20633) );
  AOI22_X1 U23220 ( .A1(n20854), .A2(n20317), .B1(n20345), .B2(n20633), .ZN(
        n20293) );
  OAI211_X1 U23221 ( .C1(n20315), .C2(n20295), .A(n20294), .B(n20293), .ZN(
        P1_U3037) );
  OAI22_X1 U23222 ( .A1(n20882), .A2(n20866), .B1(n20732), .B2(n20313), .ZN(
        n20296) );
  INV_X1 U23223 ( .A(n20296), .ZN(n20303) );
  NOR2_X2 U23224 ( .A1(n20297), .A2(n20432), .ZN(n20860) );
  INV_X1 U23225 ( .A(DATAI_21_), .ZN(n20299) );
  AOI22_X1 U23226 ( .A1(n20860), .A2(n20317), .B1(n20345), .B2(n20861), .ZN(
        n20302) );
  OAI211_X1 U23227 ( .C1(n20315), .C2(n20304), .A(n20303), .B(n20302), .ZN(
        P1_U3038) );
  AOI22_X1 U23228 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20310), .B1(DATAI_30_), 
        .B2(n20311), .ZN(n20678) );
  NAND2_X1 U23229 ( .A1(n20312), .A2(n11826), .ZN(n20739) );
  OAI22_X1 U23230 ( .A1(n20882), .A2(n20678), .B1(n20739), .B2(n20313), .ZN(
        n20305) );
  INV_X1 U23231 ( .A(n20305), .ZN(n20308) );
  NOR2_X2 U23232 ( .A1(n20306), .A2(n20432), .ZN(n20868) );
  AOI22_X1 U23233 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20310), .B1(DATAI_22_), 
        .B2(n20311), .ZN(n20872) );
  INV_X1 U23234 ( .A(n20872), .ZN(n20675) );
  AOI22_X1 U23235 ( .A1(n20868), .A2(n20317), .B1(n20345), .B2(n20675), .ZN(
        n20307) );
  OAI211_X1 U23236 ( .C1(n20315), .C2(n20309), .A(n20308), .B(n20307), .ZN(
        P1_U3039) );
  AOI22_X1 U23237 ( .A1(DATAI_31_), .A2(n20311), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20310), .ZN(n20784) );
  NAND2_X1 U23238 ( .A1(n20312), .A2(n11827), .ZN(n20745) );
  OAI22_X1 U23239 ( .A1(n20882), .A2(n20784), .B1(n20745), .B2(n20313), .ZN(
        n20314) );
  INV_X1 U23240 ( .A(n20314), .ZN(n20320) );
  INV_X1 U23241 ( .A(n20315), .ZN(n20318) );
  NOR2_X2 U23242 ( .A1(n20316), .A2(n20432), .ZN(n20876) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20318), .B1(
        n20876), .B2(n20317), .ZN(n20319) );
  OAI211_X1 U23244 ( .C1(n20883), .C2(n20342), .A(n20320), .B(n20319), .ZN(
        P1_U3040) );
  OR2_X1 U23245 ( .A1(n13831), .A2(n20349), .ZN(n20580) );
  INV_X1 U23246 ( .A(n20392), .ZN(n20322) );
  INV_X1 U23247 ( .A(n20321), .ZN(n20756) );
  NOR2_X1 U23248 ( .A1(n20755), .A2(n20323), .ZN(n20343) );
  AOI21_X1 U23249 ( .B1(n20322), .B2(n20756), .A(n20343), .ZN(n20325) );
  OAI22_X1 U23250 ( .A1(n20325), .A2(n20822), .B1(n20323), .B2(n20888), .ZN(
        n20344) );
  AOI22_X1 U23251 ( .A1(n20820), .A2(n20344), .B1(n20819), .B2(n20343), .ZN(
        n20329) );
  INV_X1 U23252 ( .A(n20323), .ZN(n20327) );
  OAI21_X1 U23253 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20701), .A(
        n20324), .ZN(n20394) );
  OAI211_X1 U23254 ( .C1(n20389), .C2(n20789), .A(n20325), .B(n20829), .ZN(
        n20326) );
  OAI211_X1 U23255 ( .C1(n20829), .C2(n20327), .A(n20828), .B(n20326), .ZN(
        n20346) );
  INV_X1 U23256 ( .A(n20387), .ZN(n20831) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20831), .ZN(n20328) );
  OAI211_X1 U23258 ( .C1(n20834), .C2(n20379), .A(n20329), .B(n20328), .ZN(
        P1_U3041) );
  AOI22_X1 U23259 ( .A1(n20836), .A2(n20344), .B1(n20835), .B2(n20343), .ZN(
        n20331) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20346), .B1(
        n20351), .B2(n20837), .ZN(n20330) );
  OAI211_X1 U23261 ( .C1(n20840), .C2(n20342), .A(n20331), .B(n20330), .ZN(
        P1_U3042) );
  AOI22_X1 U23262 ( .A1(n20842), .A2(n20344), .B1(n20841), .B2(n20343), .ZN(
        n20333) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20346), .B1(
        n20351), .B2(n20843), .ZN(n20332) );
  OAI211_X1 U23264 ( .C1(n20846), .C2(n20342), .A(n20333), .B(n20332), .ZN(
        P1_U3043) );
  AOI22_X1 U23265 ( .A1(n20848), .A2(n20344), .B1(n20847), .B2(n20343), .ZN(
        n20335) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20346), .B1(
        n20351), .B2(n20849), .ZN(n20334) );
  OAI211_X1 U23267 ( .C1(n20852), .C2(n20342), .A(n20335), .B(n20334), .ZN(
        P1_U3044) );
  AOI22_X1 U23268 ( .A1(n20854), .A2(n20344), .B1(n20853), .B2(n20343), .ZN(
        n20337) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20855), .ZN(n20336) );
  OAI211_X1 U23270 ( .C1(n20858), .C2(n20379), .A(n20337), .B(n20336), .ZN(
        P1_U3045) );
  AOI22_X1 U23271 ( .A1(n20860), .A2(n20344), .B1(n20859), .B2(n20343), .ZN(
        n20339) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20346), .B1(
        n20351), .B2(n20861), .ZN(n20338) );
  OAI211_X1 U23273 ( .C1(n20866), .C2(n20342), .A(n20339), .B(n20338), .ZN(
        P1_U3046) );
  AOI22_X1 U23274 ( .A1(n20868), .A2(n20344), .B1(n20867), .B2(n20343), .ZN(
        n20341) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20346), .B1(
        n20351), .B2(n20675), .ZN(n20340) );
  OAI211_X1 U23276 ( .C1(n20678), .C2(n20342), .A(n20341), .B(n20340), .ZN(
        P1_U3047) );
  AOI22_X1 U23277 ( .A1(n20876), .A2(n20344), .B1(n20874), .B2(n20343), .ZN(
        n20348) );
  INV_X1 U23278 ( .A(n20784), .ZN(n20877) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20877), .ZN(n20347) );
  OAI211_X1 U23280 ( .C1(n20883), .C2(n20379), .A(n20348), .B(n20347), .ZN(
        P1_U3048) );
  NAND3_X1 U23281 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20652), .A3(
        n20611), .ZN(n20397) );
  OR2_X1 U23282 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20397), .ZN(
        n20378) );
  OAI22_X1 U23283 ( .A1(n20379), .A2(n20387), .B1(n20378), .B2(n20694), .ZN(
        n20350) );
  INV_X1 U23284 ( .A(n20350), .ZN(n20359) );
  INV_X1 U23285 ( .A(n20426), .ZN(n20352) );
  OAI21_X1 U23286 ( .B1(n20352), .B2(n20351), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20353) );
  NAND2_X1 U23287 ( .A1(n20353), .A2(n20829), .ZN(n20357) );
  NOR2_X1 U23288 ( .A1(n20392), .A2(n20550), .ZN(n20355) );
  OR2_X1 U23289 ( .A1(n20608), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20482) );
  AND2_X1 U23290 ( .A1(n20482), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20486) );
  AOI211_X1 U23291 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20378), .A(n20486), 
        .B(n20555), .ZN(n20354) );
  INV_X1 U23292 ( .A(n20355), .ZN(n20356) );
  OAI22_X1 U23293 ( .A1(n20357), .A2(n20356), .B1(n20554), .B2(n20482), .ZN(
        n20381) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20382), .B1(
        n20820), .B2(n20381), .ZN(n20358) );
  OAI211_X1 U23295 ( .C1(n20834), .C2(n20426), .A(n20359), .B(n20358), .ZN(
        P1_U3049) );
  INV_X1 U23296 ( .A(n20837), .ZN(n20707) );
  OAI22_X1 U23297 ( .A1(n20426), .A2(n20707), .B1(n20706), .B2(n20378), .ZN(
        n20360) );
  INV_X1 U23298 ( .A(n20360), .ZN(n20362) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20382), .B1(
        n20836), .B2(n20381), .ZN(n20361) );
  OAI211_X1 U23300 ( .C1(n20840), .C2(n20379), .A(n20362), .B(n20361), .ZN(
        P1_U3050) );
  OAI22_X1 U23301 ( .A1(n20426), .A2(n20714), .B1(n20378), .B2(n20713), .ZN(
        n20363) );
  INV_X1 U23302 ( .A(n20363), .ZN(n20365) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20382), .B1(
        n20842), .B2(n20381), .ZN(n20364) );
  OAI211_X1 U23304 ( .C1(n20846), .C2(n20379), .A(n20365), .B(n20364), .ZN(
        P1_U3051) );
  OAI22_X1 U23305 ( .A1(n20426), .A2(n20721), .B1(n20378), .B2(n20720), .ZN(
        n20366) );
  INV_X1 U23306 ( .A(n20366), .ZN(n20368) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20382), .B1(
        n20848), .B2(n20381), .ZN(n20367) );
  OAI211_X1 U23308 ( .C1(n20852), .C2(n20379), .A(n20368), .B(n20367), .ZN(
        P1_U3052) );
  OAI22_X1 U23309 ( .A1(n20379), .A2(n20631), .B1(n20378), .B2(n20727), .ZN(
        n20369) );
  INV_X1 U23310 ( .A(n20369), .ZN(n20371) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20382), .B1(
        n20854), .B2(n20381), .ZN(n20370) );
  OAI211_X1 U23312 ( .C1(n20858), .C2(n20426), .A(n20371), .B(n20370), .ZN(
        P1_U3053) );
  INV_X1 U23313 ( .A(n20861), .ZN(n20733) );
  OAI22_X1 U23314 ( .A1(n20426), .A2(n20733), .B1(n20378), .B2(n20732), .ZN(
        n20372) );
  INV_X1 U23315 ( .A(n20372), .ZN(n20374) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20382), .B1(
        n20860), .B2(n20381), .ZN(n20373) );
  OAI211_X1 U23317 ( .C1(n20866), .C2(n20379), .A(n20374), .B(n20373), .ZN(
        P1_U3054) );
  OAI22_X1 U23318 ( .A1(n20379), .A2(n20678), .B1(n20378), .B2(n20739), .ZN(
        n20375) );
  INV_X1 U23319 ( .A(n20375), .ZN(n20377) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20382), .B1(
        n20868), .B2(n20381), .ZN(n20376) );
  OAI211_X1 U23321 ( .C1(n20872), .C2(n20426), .A(n20377), .B(n20376), .ZN(
        P1_U3055) );
  OAI22_X1 U23322 ( .A1(n20379), .A2(n20784), .B1(n20378), .B2(n20745), .ZN(
        n20380) );
  INV_X1 U23323 ( .A(n20380), .ZN(n20384) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20382), .B1(
        n20876), .B2(n20381), .ZN(n20383) );
  OAI211_X1 U23325 ( .C1(n20883), .C2(n20426), .A(n20384), .B(n20383), .ZN(
        P1_U3056) );
  INV_X1 U23326 ( .A(n20653), .ZN(n20386) );
  NAND2_X1 U23327 ( .A1(n20386), .A2(n20652), .ZN(n20420) );
  OAI22_X1 U23328 ( .A1(n20426), .A2(n20387), .B1(n20694), .B2(n20420), .ZN(
        n20388) );
  INV_X1 U23329 ( .A(n20388), .ZN(n20401) );
  AOI21_X1 U23330 ( .B1(n20389), .B2(n20829), .A(n20825), .ZN(n20399) );
  AND2_X1 U23331 ( .A1(n9785), .A2(n20390), .ZN(n20817) );
  INV_X1 U23332 ( .A(n20817), .ZN(n20391) );
  OR2_X1 U23333 ( .A1(n20392), .A2(n20391), .ZN(n20393) );
  AND2_X1 U23334 ( .A1(n20393), .A2(n20420), .ZN(n20398) );
  INV_X1 U23335 ( .A(n20398), .ZN(n20396) );
  AOI21_X1 U23336 ( .B1(n20822), .B2(n20397), .A(n20394), .ZN(n20395) );
  OAI21_X1 U23337 ( .B1(n20399), .B2(n20396), .A(n20395), .ZN(n20423) );
  OAI22_X1 U23338 ( .A1(n20399), .A2(n20398), .B1(n20888), .B2(n20397), .ZN(
        n20422) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20423), .B1(
        n20820), .B2(n20422), .ZN(n20400) );
  OAI211_X1 U23340 ( .C1(n20834), .C2(n20446), .A(n20401), .B(n20400), .ZN(
        P1_U3057) );
  OAI22_X1 U23341 ( .A1(n20446), .A2(n20707), .B1(n20706), .B2(n20420), .ZN(
        n20402) );
  INV_X1 U23342 ( .A(n20402), .ZN(n20404) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20423), .B1(
        n20836), .B2(n20422), .ZN(n20403) );
  OAI211_X1 U23344 ( .C1(n20840), .C2(n20426), .A(n20404), .B(n20403), .ZN(
        P1_U3058) );
  OAI22_X1 U23345 ( .A1(n20426), .A2(n20846), .B1(n20713), .B2(n20420), .ZN(
        n20405) );
  INV_X1 U23346 ( .A(n20405), .ZN(n20407) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20423), .B1(
        n20842), .B2(n20422), .ZN(n20406) );
  OAI211_X1 U23348 ( .C1(n20714), .C2(n20446), .A(n20407), .B(n20406), .ZN(
        P1_U3059) );
  OAI22_X1 U23349 ( .A1(n20426), .A2(n20852), .B1(n20720), .B2(n20420), .ZN(
        n20408) );
  INV_X1 U23350 ( .A(n20408), .ZN(n20410) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20423), .B1(
        n20848), .B2(n20422), .ZN(n20409) );
  OAI211_X1 U23352 ( .C1(n20721), .C2(n20446), .A(n20410), .B(n20409), .ZN(
        P1_U3060) );
  OAI22_X1 U23353 ( .A1(n20426), .A2(n20631), .B1(n20420), .B2(n20727), .ZN(
        n20411) );
  INV_X1 U23354 ( .A(n20411), .ZN(n20413) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20423), .B1(
        n20854), .B2(n20422), .ZN(n20412) );
  OAI211_X1 U23356 ( .C1(n20858), .C2(n20446), .A(n20413), .B(n20412), .ZN(
        P1_U3061) );
  OAI22_X1 U23357 ( .A1(n20446), .A2(n20733), .B1(n20732), .B2(n20420), .ZN(
        n20414) );
  INV_X1 U23358 ( .A(n20414), .ZN(n20416) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20423), .B1(
        n20860), .B2(n20422), .ZN(n20415) );
  OAI211_X1 U23360 ( .C1(n20866), .C2(n20426), .A(n20416), .B(n20415), .ZN(
        P1_U3062) );
  OAI22_X1 U23361 ( .A1(n20446), .A2(n20872), .B1(n20420), .B2(n20739), .ZN(
        n20417) );
  INV_X1 U23362 ( .A(n20417), .ZN(n20419) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20423), .B1(
        n20868), .B2(n20422), .ZN(n20418) );
  OAI211_X1 U23364 ( .C1(n20678), .C2(n20426), .A(n20419), .B(n20418), .ZN(
        P1_U3063) );
  OAI22_X1 U23365 ( .A1(n20446), .A2(n20883), .B1(n20420), .B2(n20745), .ZN(
        n20421) );
  INV_X1 U23366 ( .A(n20421), .ZN(n20425) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20423), .B1(
        n20876), .B2(n20422), .ZN(n20424) );
  OAI211_X1 U23368 ( .C1(n20784), .C2(n20426), .A(n20425), .B(n20424), .ZN(
        P1_U3064) );
  NOR2_X1 U23369 ( .A1(n20690), .A2(n20427), .ZN(n20520) );
  NAND3_X1 U23370 ( .A1(n20520), .A2(n20550), .A3(n20829), .ZN(n20428) );
  OAI21_X1 U23371 ( .B1(n20788), .B2(n20429), .A(n20428), .ZN(n20450) );
  NAND3_X1 U23372 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20652), .A3(
        n20693), .ZN(n20455) );
  NOR2_X1 U23373 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20455), .ZN(
        n20449) );
  AOI22_X1 U23374 ( .A1(n20820), .A2(n20450), .B1(n20819), .B2(n20449), .ZN(
        n20435) );
  AOI21_X1 U23375 ( .B1(n20446), .B2(n20480), .A(n20789), .ZN(n20430) );
  AOI21_X1 U23376 ( .B1(n20520), .B2(n20550), .A(n20430), .ZN(n20431) );
  NOR2_X1 U23377 ( .A1(n20431), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20433) );
  NOR2_X1 U23378 ( .A1(n20610), .A2(n20432), .ZN(n20794) );
  INV_X1 U23379 ( .A(n20446), .ZN(n20451) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20831), .ZN(n20434) );
  OAI211_X1 U23381 ( .C1(n20834), .C2(n20480), .A(n20435), .B(n20434), .ZN(
        P1_U3065) );
  AOI22_X1 U23382 ( .A1(n20836), .A2(n20450), .B1(n20835), .B2(n20449), .ZN(
        n20437) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20837), .ZN(n20436) );
  OAI211_X1 U23384 ( .C1(n20840), .C2(n20446), .A(n20437), .B(n20436), .ZN(
        P1_U3066) );
  AOI22_X1 U23385 ( .A1(n20842), .A2(n20450), .B1(n20841), .B2(n20449), .ZN(
        n20439) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20843), .ZN(n20438) );
  OAI211_X1 U23387 ( .C1(n20846), .C2(n20446), .A(n20439), .B(n20438), .ZN(
        P1_U3067) );
  AOI22_X1 U23388 ( .A1(n20848), .A2(n20450), .B1(n20847), .B2(n20449), .ZN(
        n20441) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20849), .ZN(n20440) );
  OAI211_X1 U23390 ( .C1(n20852), .C2(n20446), .A(n20441), .B(n20440), .ZN(
        P1_U3068) );
  AOI22_X1 U23391 ( .A1(n20854), .A2(n20450), .B1(n20853), .B2(n20449), .ZN(
        n20443) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20855), .ZN(n20442) );
  OAI211_X1 U23393 ( .C1(n20858), .C2(n20480), .A(n20443), .B(n20442), .ZN(
        P1_U3069) );
  AOI22_X1 U23394 ( .A1(n20860), .A2(n20450), .B1(n20859), .B2(n20449), .ZN(
        n20445) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20861), .ZN(n20444) );
  OAI211_X1 U23396 ( .C1(n20866), .C2(n20446), .A(n20445), .B(n20444), .ZN(
        P1_U3070) );
  AOI22_X1 U23397 ( .A1(n20868), .A2(n20450), .B1(n20867), .B2(n20449), .ZN(
        n20448) );
  INV_X1 U23398 ( .A(n20678), .ZN(n20869) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20869), .ZN(n20447) );
  OAI211_X1 U23400 ( .C1(n20872), .C2(n20480), .A(n20448), .B(n20447), .ZN(
        P1_U3071) );
  AOI22_X1 U23401 ( .A1(n20876), .A2(n20450), .B1(n20874), .B2(n20449), .ZN(
        n20454) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20877), .ZN(n20453) );
  OAI211_X1 U23403 ( .C1(n20883), .C2(n20480), .A(n20454), .B(n20453), .ZN(
        P1_U3072) );
  NOR2_X1 U23404 ( .A1(n20755), .A2(n20455), .ZN(n20475) );
  AOI21_X1 U23405 ( .B1(n20520), .B2(n20756), .A(n20475), .ZN(n20456) );
  OAI22_X1 U23406 ( .A1(n20456), .A2(n20822), .B1(n20455), .B2(n20888), .ZN(
        n20476) );
  AOI22_X1 U23407 ( .A1(n20820), .A2(n20476), .B1(n20819), .B2(n20475), .ZN(
        n20461) );
  INV_X1 U23408 ( .A(n20455), .ZN(n20459) );
  OAI211_X1 U23409 ( .C1(n20457), .C2(n20789), .A(n20456), .B(n20829), .ZN(
        n20458) );
  OAI211_X1 U23410 ( .C1(n20829), .C2(n20459), .A(n20828), .B(n20458), .ZN(
        n20477) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20477), .B1(
        n20468), .B2(n20831), .ZN(n20460) );
  OAI211_X1 U23412 ( .C1(n20834), .C2(n20513), .A(n20461), .B(n20460), .ZN(
        P1_U3073) );
  AOI22_X1 U23413 ( .A1(n20836), .A2(n20476), .B1(n20835), .B2(n20475), .ZN(
        n20463) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20477), .B1(
        n20509), .B2(n20837), .ZN(n20462) );
  OAI211_X1 U23415 ( .C1(n20840), .C2(n20480), .A(n20463), .B(n20462), .ZN(
        P1_U3074) );
  AOI22_X1 U23416 ( .A1(n20842), .A2(n20476), .B1(n20841), .B2(n20475), .ZN(
        n20465) );
  INV_X1 U23417 ( .A(n20846), .ZN(n20716) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20477), .B1(
        n20468), .B2(n20716), .ZN(n20464) );
  OAI211_X1 U23419 ( .C1(n20714), .C2(n20513), .A(n20465), .B(n20464), .ZN(
        P1_U3075) );
  AOI22_X1 U23420 ( .A1(n20848), .A2(n20476), .B1(n20847), .B2(n20475), .ZN(
        n20467) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20477), .B1(
        n20509), .B2(n20849), .ZN(n20466) );
  OAI211_X1 U23422 ( .C1(n20852), .C2(n20480), .A(n20467), .B(n20466), .ZN(
        P1_U3076) );
  AOI22_X1 U23423 ( .A1(n20854), .A2(n20476), .B1(n20853), .B2(n20475), .ZN(
        n20470) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20477), .B1(
        n20468), .B2(n20855), .ZN(n20469) );
  OAI211_X1 U23425 ( .C1(n20858), .C2(n20513), .A(n20470), .B(n20469), .ZN(
        P1_U3077) );
  AOI22_X1 U23426 ( .A1(n20860), .A2(n20476), .B1(n20859), .B2(n20475), .ZN(
        n20472) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20477), .B1(
        n20509), .B2(n20861), .ZN(n20471) );
  OAI211_X1 U23428 ( .C1(n20866), .C2(n20480), .A(n20472), .B(n20471), .ZN(
        P1_U3078) );
  AOI22_X1 U23429 ( .A1(n20868), .A2(n20476), .B1(n20867), .B2(n20475), .ZN(
        n20474) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20477), .B1(
        n20509), .B2(n20675), .ZN(n20473) );
  OAI211_X1 U23431 ( .C1(n20678), .C2(n20480), .A(n20474), .B(n20473), .ZN(
        P1_U3079) );
  AOI22_X1 U23432 ( .A1(n20876), .A2(n20476), .B1(n20874), .B2(n20475), .ZN(
        n20479) );
  INV_X1 U23433 ( .A(n20883), .ZN(n20779) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20477), .B1(
        n20509), .B2(n20779), .ZN(n20478) );
  OAI211_X1 U23435 ( .C1(n20784), .C2(n20480), .A(n20479), .B(n20478), .ZN(
        P1_U3080) );
  NAND3_X1 U23436 ( .A1(n20541), .A2(n20513), .A3(n20829), .ZN(n20481) );
  NAND2_X1 U23437 ( .A1(n20481), .A2(n20687), .ZN(n20488) );
  AND2_X1 U23438 ( .A1(n20520), .A2(n20791), .ZN(n20485) );
  INV_X1 U23439 ( .A(n20482), .ZN(n20483) );
  INV_X1 U23440 ( .A(n20788), .ZN(n20692) );
  AOI22_X1 U23441 ( .A1(n20488), .A2(n20485), .B1(n20483), .B2(n20692), .ZN(
        n20518) );
  INV_X1 U23442 ( .A(n20820), .ZN(n20705) );
  INV_X1 U23443 ( .A(n20526), .ZN(n20521) );
  NOR2_X1 U23444 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20521), .ZN(
        n20490) );
  INV_X1 U23445 ( .A(n20490), .ZN(n20512) );
  OAI22_X1 U23446 ( .A1(n20541), .A2(n20834), .B1(n20694), .B2(n20512), .ZN(
        n20484) );
  INV_X1 U23447 ( .A(n20484), .ZN(n20492) );
  INV_X1 U23448 ( .A(n20485), .ZN(n20487) );
  AOI21_X1 U23449 ( .B1(n20488), .B2(n20487), .A(n20486), .ZN(n20489) );
  OAI211_X1 U23450 ( .C1(n20490), .C2(n20701), .A(n20794), .B(n20489), .ZN(
        n20515) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20515), .B1(
        n20509), .B2(n20831), .ZN(n20491) );
  OAI211_X1 U23452 ( .C1(n20518), .C2(n20705), .A(n20492), .B(n20491), .ZN(
        P1_U3081) );
  INV_X1 U23453 ( .A(n20836), .ZN(n20712) );
  OAI22_X1 U23454 ( .A1(n20513), .A2(n20840), .B1(n20706), .B2(n20512), .ZN(
        n20493) );
  INV_X1 U23455 ( .A(n20493), .ZN(n20495) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20515), .B1(
        n20544), .B2(n20837), .ZN(n20494) );
  OAI211_X1 U23457 ( .C1(n20518), .C2(n20712), .A(n20495), .B(n20494), .ZN(
        P1_U3082) );
  INV_X1 U23458 ( .A(n20842), .ZN(n20719) );
  OAI22_X1 U23459 ( .A1(n20513), .A2(n20846), .B1(n20713), .B2(n20512), .ZN(
        n20496) );
  INV_X1 U23460 ( .A(n20496), .ZN(n20498) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20515), .B1(
        n20544), .B2(n20843), .ZN(n20497) );
  OAI211_X1 U23462 ( .C1(n20518), .C2(n20719), .A(n20498), .B(n20497), .ZN(
        P1_U3083) );
  INV_X1 U23463 ( .A(n20848), .ZN(n20726) );
  OAI22_X1 U23464 ( .A1(n20513), .A2(n20852), .B1(n20720), .B2(n20512), .ZN(
        n20499) );
  INV_X1 U23465 ( .A(n20499), .ZN(n20501) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20515), .B1(
        n20544), .B2(n20849), .ZN(n20500) );
  OAI211_X1 U23467 ( .C1(n20518), .C2(n20726), .A(n20501), .B(n20500), .ZN(
        P1_U3084) );
  INV_X1 U23468 ( .A(n20854), .ZN(n20731) );
  OAI22_X1 U23469 ( .A1(n20513), .A2(n20631), .B1(n20727), .B2(n20512), .ZN(
        n20502) );
  INV_X1 U23470 ( .A(n20502), .ZN(n20504) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20515), .B1(
        n20544), .B2(n20633), .ZN(n20503) );
  OAI211_X1 U23472 ( .C1(n20518), .C2(n20731), .A(n20504), .B(n20503), .ZN(
        P1_U3085) );
  INV_X1 U23473 ( .A(n20860), .ZN(n20738) );
  OAI22_X1 U23474 ( .A1(n20541), .A2(n20733), .B1(n20732), .B2(n20512), .ZN(
        n20505) );
  INV_X1 U23475 ( .A(n20505), .ZN(n20507) );
  INV_X1 U23476 ( .A(n20866), .ZN(n20735) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20515), .B1(
        n20509), .B2(n20735), .ZN(n20506) );
  OAI211_X1 U23478 ( .C1(n20518), .C2(n20738), .A(n20507), .B(n20506), .ZN(
        P1_U3086) );
  INV_X1 U23479 ( .A(n20868), .ZN(n20743) );
  OAI22_X1 U23480 ( .A1(n20541), .A2(n20872), .B1(n20739), .B2(n20512), .ZN(
        n20508) );
  INV_X1 U23481 ( .A(n20508), .ZN(n20511) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20515), .B1(
        n20509), .B2(n20869), .ZN(n20510) );
  OAI211_X1 U23483 ( .C1(n20518), .C2(n20743), .A(n20511), .B(n20510), .ZN(
        P1_U3087) );
  INV_X1 U23484 ( .A(n20876), .ZN(n20751) );
  OAI22_X1 U23485 ( .A1(n20513), .A2(n20784), .B1(n20745), .B2(n20512), .ZN(
        n20514) );
  INV_X1 U23486 ( .A(n20514), .ZN(n20517) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20515), .B1(
        n20544), .B2(n20779), .ZN(n20516) );
  OAI211_X1 U23488 ( .C1(n20518), .C2(n20751), .A(n20517), .B(n20516), .ZN(
        P1_U3088) );
  NAND2_X1 U23489 ( .A1(n20522), .A2(n20650), .ZN(n20571) );
  INV_X1 U23490 ( .A(n20519), .ZN(n20542) );
  AOI21_X1 U23491 ( .B1(n20520), .B2(n20817), .A(n20542), .ZN(n20523) );
  OAI22_X1 U23492 ( .A1(n20523), .A2(n20822), .B1(n20521), .B2(n20888), .ZN(
        n20543) );
  AOI22_X1 U23493 ( .A1(n20820), .A2(n20543), .B1(n20819), .B2(n20542), .ZN(
        n20528) );
  NOR2_X1 U23494 ( .A1(n20522), .A2(n20822), .ZN(n20524) );
  OAI21_X1 U23495 ( .B1(n20524), .B2(n20825), .A(n20523), .ZN(n20525) );
  OAI211_X1 U23496 ( .C1(n20526), .C2(n20829), .A(n20828), .B(n20525), .ZN(
        n20545) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20831), .ZN(n20527) );
  OAI211_X1 U23498 ( .C1(n20834), .C2(n20571), .A(n20528), .B(n20527), .ZN(
        P1_U3089) );
  AOI22_X1 U23499 ( .A1(n20836), .A2(n20543), .B1(n20835), .B2(n20542), .ZN(
        n20530) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20545), .B1(
        n20576), .B2(n20837), .ZN(n20529) );
  OAI211_X1 U23501 ( .C1(n20840), .C2(n20541), .A(n20530), .B(n20529), .ZN(
        P1_U3090) );
  AOI22_X1 U23502 ( .A1(n20842), .A2(n20543), .B1(n20841), .B2(n20542), .ZN(
        n20532) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20545), .B1(
        n20576), .B2(n20843), .ZN(n20531) );
  OAI211_X1 U23504 ( .C1(n20846), .C2(n20541), .A(n20532), .B(n20531), .ZN(
        P1_U3091) );
  AOI22_X1 U23505 ( .A1(n20848), .A2(n20543), .B1(n20847), .B2(n20542), .ZN(
        n20534) );
  INV_X1 U23506 ( .A(n20852), .ZN(n20723) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20723), .ZN(n20533) );
  OAI211_X1 U23508 ( .C1(n20721), .C2(n20571), .A(n20534), .B(n20533), .ZN(
        P1_U3092) );
  AOI22_X1 U23509 ( .A1(n20854), .A2(n20543), .B1(n20853), .B2(n20542), .ZN(
        n20536) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20855), .ZN(n20535) );
  OAI211_X1 U23511 ( .C1(n20858), .C2(n20571), .A(n20536), .B(n20535), .ZN(
        P1_U3093) );
  AOI22_X1 U23512 ( .A1(n20860), .A2(n20543), .B1(n20859), .B2(n20542), .ZN(
        n20538) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20545), .B1(
        n20576), .B2(n20861), .ZN(n20537) );
  OAI211_X1 U23514 ( .C1(n20866), .C2(n20541), .A(n20538), .B(n20537), .ZN(
        P1_U3094) );
  AOI22_X1 U23515 ( .A1(n20868), .A2(n20543), .B1(n20867), .B2(n20542), .ZN(
        n20540) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20545), .B1(
        n20576), .B2(n20675), .ZN(n20539) );
  OAI211_X1 U23517 ( .C1(n20678), .C2(n20541), .A(n20540), .B(n20539), .ZN(
        P1_U3095) );
  AOI22_X1 U23518 ( .A1(n20876), .A2(n20543), .B1(n20874), .B2(n20542), .ZN(
        n20547) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20877), .ZN(n20546) );
  OAI211_X1 U23520 ( .C1(n20883), .C2(n20571), .A(n20547), .B(n20546), .ZN(
        P1_U3096) );
  AND2_X1 U23521 ( .A1(n20549), .A2(n20690), .ZN(n20654) );
  NAND3_X1 U23522 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20611), .A3(
        n20693), .ZN(n20581) );
  NOR2_X1 U23523 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20581), .ZN(
        n20574) );
  AOI21_X1 U23524 ( .B1(n20654), .B2(n20550), .A(n20574), .ZN(n20556) );
  INV_X1 U23525 ( .A(n20551), .ZN(n20553) );
  NOR2_X1 U23526 ( .A1(n20553), .A2(n20552), .ZN(n20691) );
  INV_X1 U23527 ( .A(n20691), .ZN(n20697) );
  OAI22_X1 U23528 ( .A1(n20556), .A2(n20822), .B1(n20697), .B2(n20554), .ZN(
        n20575) );
  AOI22_X1 U23529 ( .A1(n20820), .A2(n20575), .B1(n20819), .B2(n20574), .ZN(
        n20560) );
  INV_X1 U23530 ( .A(n20555), .ZN(n20614) );
  OAI21_X1 U23531 ( .B1(n20602), .B2(n20576), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20557) );
  NAND2_X1 U23532 ( .A1(n20557), .A2(n20556), .ZN(n20558) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20577), .B1(
        n20576), .B2(n20831), .ZN(n20559) );
  OAI211_X1 U23534 ( .C1(n20834), .C2(n20599), .A(n20560), .B(n20559), .ZN(
        P1_U3097) );
  AOI22_X1 U23535 ( .A1(n20836), .A2(n20575), .B1(n20835), .B2(n20574), .ZN(
        n20562) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20577), .B1(
        n20602), .B2(n20837), .ZN(n20561) );
  OAI211_X1 U23537 ( .C1(n20840), .C2(n20571), .A(n20562), .B(n20561), .ZN(
        P1_U3098) );
  AOI22_X1 U23538 ( .A1(n20842), .A2(n20575), .B1(n20841), .B2(n20574), .ZN(
        n20564) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20577), .B1(
        n20576), .B2(n20716), .ZN(n20563) );
  OAI211_X1 U23540 ( .C1(n20714), .C2(n20599), .A(n20564), .B(n20563), .ZN(
        P1_U3099) );
  AOI22_X1 U23541 ( .A1(n20848), .A2(n20575), .B1(n20847), .B2(n20574), .ZN(
        n20566) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20577), .B1(
        n20576), .B2(n20723), .ZN(n20565) );
  OAI211_X1 U23543 ( .C1(n20721), .C2(n20599), .A(n20566), .B(n20565), .ZN(
        P1_U3100) );
  AOI22_X1 U23544 ( .A1(n20854), .A2(n20575), .B1(n20853), .B2(n20574), .ZN(
        n20568) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20577), .B1(
        n20576), .B2(n20855), .ZN(n20567) );
  OAI211_X1 U23546 ( .C1(n20858), .C2(n20599), .A(n20568), .B(n20567), .ZN(
        P1_U3101) );
  AOI22_X1 U23547 ( .A1(n20860), .A2(n20575), .B1(n20859), .B2(n20574), .ZN(
        n20570) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20577), .B1(
        n20602), .B2(n20861), .ZN(n20569) );
  OAI211_X1 U23549 ( .C1(n20866), .C2(n20571), .A(n20570), .B(n20569), .ZN(
        P1_U3102) );
  AOI22_X1 U23550 ( .A1(n20868), .A2(n20575), .B1(n20867), .B2(n20574), .ZN(
        n20573) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20577), .B1(
        n20576), .B2(n20869), .ZN(n20572) );
  OAI211_X1 U23552 ( .C1(n20872), .C2(n20599), .A(n20573), .B(n20572), .ZN(
        P1_U3103) );
  AOI22_X1 U23553 ( .A1(n20876), .A2(n20575), .B1(n20874), .B2(n20574), .ZN(
        n20579) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20577), .B1(
        n20576), .B2(n20877), .ZN(n20578) );
  OAI211_X1 U23555 ( .C1(n20883), .C2(n20599), .A(n20579), .B(n20578), .ZN(
        P1_U3104) );
  NOR2_X1 U23556 ( .A1(n20755), .A2(n20581), .ZN(n20600) );
  AOI21_X1 U23557 ( .B1(n20654), .B2(n20756), .A(n20600), .ZN(n20582) );
  OAI22_X1 U23558 ( .A1(n20582), .A2(n20822), .B1(n20581), .B2(n20888), .ZN(
        n20601) );
  AOI22_X1 U23559 ( .A1(n20820), .A2(n20601), .B1(n20819), .B2(n20600), .ZN(
        n20586) );
  INV_X1 U23560 ( .A(n20581), .ZN(n20584) );
  OAI211_X1 U23561 ( .C1(n20656), .C2(n20789), .A(n20582), .B(n20829), .ZN(
        n20583) );
  OAI211_X1 U23562 ( .C1(n20829), .C2(n20584), .A(n20828), .B(n20583), .ZN(
        n20603) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20831), .ZN(n20585) );
  OAI211_X1 U23564 ( .C1(n20834), .C2(n20639), .A(n20586), .B(n20585), .ZN(
        P1_U3105) );
  AOI22_X1 U23565 ( .A1(n20836), .A2(n20601), .B1(n20835), .B2(n20600), .ZN(
        n20588) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20603), .B1(
        n20645), .B2(n20837), .ZN(n20587) );
  OAI211_X1 U23567 ( .C1(n20840), .C2(n20599), .A(n20588), .B(n20587), .ZN(
        P1_U3106) );
  AOI22_X1 U23568 ( .A1(n20842), .A2(n20601), .B1(n20841), .B2(n20600), .ZN(
        n20590) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20603), .B1(
        n20645), .B2(n20843), .ZN(n20589) );
  OAI211_X1 U23570 ( .C1(n20846), .C2(n20599), .A(n20590), .B(n20589), .ZN(
        P1_U3107) );
  AOI22_X1 U23571 ( .A1(n20848), .A2(n20601), .B1(n20847), .B2(n20600), .ZN(
        n20592) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20723), .ZN(n20591) );
  OAI211_X1 U23573 ( .C1(n20721), .C2(n20639), .A(n20592), .B(n20591), .ZN(
        P1_U3108) );
  AOI22_X1 U23574 ( .A1(n20854), .A2(n20601), .B1(n20853), .B2(n20600), .ZN(
        n20594) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20855), .ZN(n20593) );
  OAI211_X1 U23576 ( .C1(n20858), .C2(n20639), .A(n20594), .B(n20593), .ZN(
        P1_U3109) );
  AOI22_X1 U23577 ( .A1(n20860), .A2(n20601), .B1(n20859), .B2(n20600), .ZN(
        n20596) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20603), .B1(
        n20645), .B2(n20861), .ZN(n20595) );
  OAI211_X1 U23579 ( .C1(n20866), .C2(n20599), .A(n20596), .B(n20595), .ZN(
        P1_U3110) );
  AOI22_X1 U23580 ( .A1(n20868), .A2(n20601), .B1(n20867), .B2(n20600), .ZN(
        n20598) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20603), .B1(
        n20645), .B2(n20675), .ZN(n20597) );
  OAI211_X1 U23582 ( .C1(n20678), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        P1_U3111) );
  AOI22_X1 U23583 ( .A1(n20876), .A2(n20601), .B1(n20874), .B2(n20600), .ZN(
        n20605) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20877), .ZN(n20604) );
  OAI211_X1 U23585 ( .C1(n20883), .C2(n20639), .A(n20605), .B(n20604), .ZN(
        P1_U3112) );
  INV_X1 U23586 ( .A(n20785), .ZN(n20606) );
  NAND3_X1 U23587 ( .A1(n20684), .A2(n20639), .A3(n20829), .ZN(n20607) );
  NAND2_X1 U23588 ( .A1(n20607), .A2(n20687), .ZN(n20618) );
  AND2_X1 U23589 ( .A1(n20654), .A2(n20791), .ZN(n20613) );
  OR2_X1 U23590 ( .A1(n20608), .A2(n20652), .ZN(n20787) );
  INV_X1 U23591 ( .A(n20787), .ZN(n20609) );
  AOI22_X1 U23592 ( .A1(n20618), .A2(n20613), .B1(n20610), .B2(n20609), .ZN(
        n20649) );
  NAND3_X1 U23593 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20611), .ZN(n20655) );
  NOR2_X1 U23594 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20655), .ZN(
        n20615) );
  INV_X1 U23595 ( .A(n20615), .ZN(n20643) );
  OAI22_X1 U23596 ( .A1(n20684), .A2(n20834), .B1(n20694), .B2(n20643), .ZN(
        n20612) );
  INV_X1 U23597 ( .A(n20612), .ZN(n20621) );
  INV_X1 U23598 ( .A(n20613), .ZN(n20617) );
  NAND2_X1 U23599 ( .A1(n20787), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20793) );
  OAI211_X1 U23600 ( .C1(n20701), .C2(n20615), .A(n20793), .B(n20614), .ZN(
        n20616) );
  AOI21_X1 U23601 ( .B1(n20618), .B2(n20617), .A(n20616), .ZN(n20619) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20831), .ZN(n20620) );
  OAI211_X1 U23603 ( .C1(n20649), .C2(n20705), .A(n20621), .B(n20620), .ZN(
        P1_U3113) );
  OAI22_X1 U23604 ( .A1(n20684), .A2(n20707), .B1(n20706), .B2(n20643), .ZN(
        n20622) );
  INV_X1 U23605 ( .A(n20622), .ZN(n20624) );
  INV_X1 U23606 ( .A(n20840), .ZN(n20709) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20709), .ZN(n20623) );
  OAI211_X1 U23608 ( .C1(n20649), .C2(n20712), .A(n20624), .B(n20623), .ZN(
        P1_U3114) );
  OAI22_X1 U23609 ( .A1(n20639), .A2(n20846), .B1(n20713), .B2(n20643), .ZN(
        n20625) );
  INV_X1 U23610 ( .A(n20625), .ZN(n20627) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20646), .B1(
        n20670), .B2(n20843), .ZN(n20626) );
  OAI211_X1 U23612 ( .C1(n20649), .C2(n20719), .A(n20627), .B(n20626), .ZN(
        P1_U3115) );
  OAI22_X1 U23613 ( .A1(n20639), .A2(n20852), .B1(n20720), .B2(n20643), .ZN(
        n20628) );
  INV_X1 U23614 ( .A(n20628), .ZN(n20630) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20646), .B1(
        n20670), .B2(n20849), .ZN(n20629) );
  OAI211_X1 U23616 ( .C1(n20649), .C2(n20726), .A(n20630), .B(n20629), .ZN(
        P1_U3116) );
  OAI22_X1 U23617 ( .A1(n20639), .A2(n20631), .B1(n20727), .B2(n20643), .ZN(
        n20632) );
  INV_X1 U23618 ( .A(n20632), .ZN(n20635) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20646), .B1(
        n20670), .B2(n20633), .ZN(n20634) );
  OAI211_X1 U23620 ( .C1(n20649), .C2(n20731), .A(n20635), .B(n20634), .ZN(
        P1_U3117) );
  OAI22_X1 U23621 ( .A1(n20684), .A2(n20733), .B1(n20732), .B2(n20643), .ZN(
        n20636) );
  INV_X1 U23622 ( .A(n20636), .ZN(n20638) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20735), .ZN(n20637) );
  OAI211_X1 U23624 ( .C1(n20649), .C2(n20738), .A(n20638), .B(n20637), .ZN(
        P1_U3118) );
  OAI22_X1 U23625 ( .A1(n20639), .A2(n20678), .B1(n20643), .B2(n20739), .ZN(
        n20640) );
  INV_X1 U23626 ( .A(n20640), .ZN(n20642) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20646), .B1(
        n20670), .B2(n20675), .ZN(n20641) );
  OAI211_X1 U23628 ( .C1(n20649), .C2(n20743), .A(n20642), .B(n20641), .ZN(
        P1_U3119) );
  OAI22_X1 U23629 ( .A1(n20684), .A2(n20883), .B1(n20643), .B2(n20745), .ZN(
        n20644) );
  INV_X1 U23630 ( .A(n20644), .ZN(n20648) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20646), .B1(
        n20645), .B2(n20877), .ZN(n20647) );
  OAI211_X1 U23632 ( .C1(n20649), .C2(n20751), .A(n20648), .B(n20647), .ZN(
        P1_U3120) );
  INV_X1 U23633 ( .A(n20650), .ZN(n20651) );
  NOR2_X1 U23634 ( .A1(n20653), .A2(n20652), .ZN(n20679) );
  AOI21_X1 U23635 ( .B1(n20654), .B2(n20817), .A(n20679), .ZN(n20658) );
  OAI22_X1 U23636 ( .A1(n20658), .A2(n20822), .B1(n20655), .B2(n20888), .ZN(
        n20680) );
  AOI22_X1 U23637 ( .A1(n20820), .A2(n20680), .B1(n20819), .B2(n20679), .ZN(
        n20663) );
  INV_X1 U23638 ( .A(n20655), .ZN(n20661) );
  INV_X1 U23639 ( .A(n20656), .ZN(n20657) );
  NOR2_X1 U23640 ( .A1(n20657), .A2(n20822), .ZN(n20659) );
  OAI21_X1 U23641 ( .B1(n20659), .B2(n20825), .A(n20658), .ZN(n20660) );
  OAI211_X1 U23642 ( .C1(n20829), .C2(n20661), .A(n20828), .B(n20660), .ZN(
        n20681) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20681), .B1(
        n20670), .B2(n20831), .ZN(n20662) );
  OAI211_X1 U23644 ( .C1(n20834), .C2(n20686), .A(n20663), .B(n20662), .ZN(
        P1_U3121) );
  AOI22_X1 U23645 ( .A1(n20836), .A2(n20680), .B1(n20835), .B2(n20679), .ZN(
        n20665) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20681), .B1(
        n20747), .B2(n20837), .ZN(n20664) );
  OAI211_X1 U23647 ( .C1(n20840), .C2(n20684), .A(n20665), .B(n20664), .ZN(
        P1_U3122) );
  AOI22_X1 U23648 ( .A1(n20842), .A2(n20680), .B1(n20841), .B2(n20679), .ZN(
        n20667) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20681), .B1(
        n20670), .B2(n20716), .ZN(n20666) );
  OAI211_X1 U23650 ( .C1(n20714), .C2(n20686), .A(n20667), .B(n20666), .ZN(
        P1_U3123) );
  AOI22_X1 U23651 ( .A1(n20848), .A2(n20680), .B1(n20847), .B2(n20679), .ZN(
        n20669) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20681), .B1(
        n20747), .B2(n20849), .ZN(n20668) );
  OAI211_X1 U23653 ( .C1(n20852), .C2(n20684), .A(n20669), .B(n20668), .ZN(
        P1_U3124) );
  AOI22_X1 U23654 ( .A1(n20854), .A2(n20680), .B1(n20853), .B2(n20679), .ZN(
        n20672) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20681), .B1(
        n20670), .B2(n20855), .ZN(n20671) );
  OAI211_X1 U23656 ( .C1(n20858), .C2(n20686), .A(n20672), .B(n20671), .ZN(
        P1_U3125) );
  AOI22_X1 U23657 ( .A1(n20860), .A2(n20680), .B1(n20859), .B2(n20679), .ZN(
        n20674) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20681), .B1(
        n20747), .B2(n20861), .ZN(n20673) );
  OAI211_X1 U23659 ( .C1(n20866), .C2(n20684), .A(n20674), .B(n20673), .ZN(
        P1_U3126) );
  AOI22_X1 U23660 ( .A1(n20868), .A2(n20680), .B1(n20867), .B2(n20679), .ZN(
        n20677) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20681), .B1(
        n20747), .B2(n20675), .ZN(n20676) );
  OAI211_X1 U23662 ( .C1(n20678), .C2(n20684), .A(n20677), .B(n20676), .ZN(
        P1_U3127) );
  AOI22_X1 U23663 ( .A1(n20876), .A2(n20680), .B1(n20874), .B2(n20679), .ZN(
        n20683) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20681), .B1(
        n20747), .B2(n20779), .ZN(n20682) );
  OAI211_X1 U23665 ( .C1(n20784), .C2(n20684), .A(n20683), .B(n20682), .ZN(
        P1_U3128) );
  NAND3_X1 U23666 ( .A1(n20686), .A2(n20829), .A3(n20783), .ZN(n20688) );
  NAND2_X1 U23667 ( .A1(n20688), .A2(n20687), .ZN(n20699) );
  OR2_X1 U23668 ( .A1(n20690), .A2(n20689), .ZN(n20754) );
  NOR2_X1 U23669 ( .A1(n20754), .A2(n20791), .ZN(n20696) );
  AOI22_X1 U23670 ( .A1(n20699), .A2(n20696), .B1(n20692), .B2(n20691), .ZN(
        n20752) );
  NAND3_X1 U23671 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20693), .ZN(n20757) );
  NOR2_X1 U23672 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20757), .ZN(
        n20702) );
  INV_X1 U23673 ( .A(n20702), .ZN(n20744) );
  OAI22_X1 U23674 ( .A1(n20783), .A2(n20834), .B1(n20694), .B2(n20744), .ZN(
        n20695) );
  INV_X1 U23675 ( .A(n20695), .ZN(n20704) );
  INV_X1 U23676 ( .A(n20696), .ZN(n20698) );
  AOI22_X1 U23677 ( .A1(n20699), .A2(n20698), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20697), .ZN(n20700) );
  OAI211_X1 U23678 ( .C1(n20702), .C2(n20701), .A(n20794), .B(n20700), .ZN(
        n20748) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20831), .ZN(n20703) );
  OAI211_X1 U23680 ( .C1(n20752), .C2(n20705), .A(n20704), .B(n20703), .ZN(
        P1_U3129) );
  OAI22_X1 U23681 ( .A1(n20783), .A2(n20707), .B1(n20706), .B2(n20744), .ZN(
        n20708) );
  INV_X1 U23682 ( .A(n20708), .ZN(n20711) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20709), .ZN(n20710) );
  OAI211_X1 U23684 ( .C1(n20752), .C2(n20712), .A(n20711), .B(n20710), .ZN(
        P1_U3130) );
  OAI22_X1 U23685 ( .A1(n20783), .A2(n20714), .B1(n20713), .B2(n20744), .ZN(
        n20715) );
  INV_X1 U23686 ( .A(n20715), .ZN(n20718) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20716), .ZN(n20717) );
  OAI211_X1 U23688 ( .C1(n20752), .C2(n20719), .A(n20718), .B(n20717), .ZN(
        P1_U3131) );
  OAI22_X1 U23689 ( .A1(n20783), .A2(n20721), .B1(n20720), .B2(n20744), .ZN(
        n20722) );
  INV_X1 U23690 ( .A(n20722), .ZN(n20725) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20723), .ZN(n20724) );
  OAI211_X1 U23692 ( .C1(n20752), .C2(n20726), .A(n20725), .B(n20724), .ZN(
        P1_U3132) );
  OAI22_X1 U23693 ( .A1(n20783), .A2(n20858), .B1(n20727), .B2(n20744), .ZN(
        n20728) );
  INV_X1 U23694 ( .A(n20728), .ZN(n20730) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20855), .ZN(n20729) );
  OAI211_X1 U23696 ( .C1(n20752), .C2(n20731), .A(n20730), .B(n20729), .ZN(
        P1_U3133) );
  OAI22_X1 U23697 ( .A1(n20783), .A2(n20733), .B1(n20732), .B2(n20744), .ZN(
        n20734) );
  INV_X1 U23698 ( .A(n20734), .ZN(n20737) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20735), .ZN(n20736) );
  OAI211_X1 U23700 ( .C1(n20752), .C2(n20738), .A(n20737), .B(n20736), .ZN(
        P1_U3134) );
  OAI22_X1 U23701 ( .A1(n20783), .A2(n20872), .B1(n20739), .B2(n20744), .ZN(
        n20740) );
  INV_X1 U23702 ( .A(n20740), .ZN(n20742) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20869), .ZN(n20741) );
  OAI211_X1 U23704 ( .C1(n20752), .C2(n20743), .A(n20742), .B(n20741), .ZN(
        P1_U3135) );
  OAI22_X1 U23705 ( .A1(n20783), .A2(n20883), .B1(n20745), .B2(n20744), .ZN(
        n20746) );
  INV_X1 U23706 ( .A(n20746), .ZN(n20750) );
  AOI22_X1 U23707 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20877), .ZN(n20749) );
  OAI211_X1 U23708 ( .C1(n20752), .C2(n20751), .A(n20750), .B(n20749), .ZN(
        P1_U3136) );
  INV_X1 U23709 ( .A(n20754), .ZN(n20818) );
  NOR2_X1 U23710 ( .A1(n20755), .A2(n20757), .ZN(n20777) );
  AOI21_X1 U23711 ( .B1(n20818), .B2(n20756), .A(n20777), .ZN(n20758) );
  OAI22_X1 U23712 ( .A1(n20758), .A2(n20822), .B1(n20757), .B2(n20888), .ZN(
        n20778) );
  AOI22_X1 U23713 ( .A1(n20820), .A2(n20778), .B1(n20819), .B2(n20777), .ZN(
        n20763) );
  INV_X1 U23714 ( .A(n20757), .ZN(n20761) );
  OAI211_X1 U23715 ( .C1(n20759), .C2(n20789), .A(n20758), .B(n20829), .ZN(
        n20760) );
  OAI211_X1 U23716 ( .C1(n20829), .C2(n20761), .A(n20828), .B(n20760), .ZN(
        n20780) );
  INV_X1 U23717 ( .A(n20783), .ZN(n20774) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20780), .B1(
        n20774), .B2(n20831), .ZN(n20762) );
  OAI211_X1 U23719 ( .C1(n20834), .C2(n20808), .A(n20763), .B(n20762), .ZN(
        P1_U3137) );
  AOI22_X1 U23720 ( .A1(n20836), .A2(n20778), .B1(n20835), .B2(n20777), .ZN(
        n20765) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20780), .B1(
        n20813), .B2(n20837), .ZN(n20764) );
  OAI211_X1 U23722 ( .C1(n20840), .C2(n20783), .A(n20765), .B(n20764), .ZN(
        P1_U3138) );
  AOI22_X1 U23723 ( .A1(n20842), .A2(n20778), .B1(n20841), .B2(n20777), .ZN(
        n20767) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20780), .B1(
        n20813), .B2(n20843), .ZN(n20766) );
  OAI211_X1 U23725 ( .C1(n20846), .C2(n20783), .A(n20767), .B(n20766), .ZN(
        P1_U3139) );
  AOI22_X1 U23726 ( .A1(n20848), .A2(n20778), .B1(n20847), .B2(n20777), .ZN(
        n20769) );
  AOI22_X1 U23727 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20780), .B1(
        n20813), .B2(n20849), .ZN(n20768) );
  OAI211_X1 U23728 ( .C1(n20852), .C2(n20783), .A(n20769), .B(n20768), .ZN(
        P1_U3140) );
  AOI22_X1 U23729 ( .A1(n20854), .A2(n20778), .B1(n20853), .B2(n20777), .ZN(
        n20771) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20780), .B1(
        n20774), .B2(n20855), .ZN(n20770) );
  OAI211_X1 U23731 ( .C1(n20858), .C2(n20808), .A(n20771), .B(n20770), .ZN(
        P1_U3141) );
  AOI22_X1 U23732 ( .A1(n20860), .A2(n20778), .B1(n20859), .B2(n20777), .ZN(
        n20773) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20780), .B1(
        n20813), .B2(n20861), .ZN(n20772) );
  OAI211_X1 U23734 ( .C1(n20866), .C2(n20783), .A(n20773), .B(n20772), .ZN(
        P1_U3142) );
  AOI22_X1 U23735 ( .A1(n20868), .A2(n20778), .B1(n20867), .B2(n20777), .ZN(
        n20776) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20780), .B1(
        n20774), .B2(n20869), .ZN(n20775) );
  OAI211_X1 U23737 ( .C1(n20872), .C2(n20808), .A(n20776), .B(n20775), .ZN(
        P1_U3143) );
  AOI22_X1 U23738 ( .A1(n20876), .A2(n20778), .B1(n20874), .B2(n20777), .ZN(
        n20782) );
  AOI22_X1 U23739 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20780), .B1(
        n20813), .B2(n20779), .ZN(n20781) );
  OAI211_X1 U23740 ( .C1(n20784), .C2(n20783), .A(n20782), .B(n20781), .ZN(
        P1_U3144) );
  NAND3_X1 U23741 ( .A1(n20818), .A2(n20791), .A3(n20829), .ZN(n20786) );
  OAI21_X1 U23742 ( .B1(n20788), .B2(n20787), .A(n20786), .ZN(n20812) );
  NOR2_X1 U23743 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20821), .ZN(
        n20811) );
  AOI22_X1 U23744 ( .A1(n20820), .A2(n20812), .B1(n20819), .B2(n20811), .ZN(
        n20797) );
  AOI21_X1 U23745 ( .B1(n20865), .B2(n20808), .A(n20789), .ZN(n20790) );
  AOI21_X1 U23746 ( .B1(n20818), .B2(n20791), .A(n20790), .ZN(n20792) );
  NOR2_X1 U23747 ( .A1(n20792), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20795) );
  AOI22_X1 U23748 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20814), .B1(
        n20813), .B2(n20831), .ZN(n20796) );
  OAI211_X1 U23749 ( .C1(n20834), .C2(n20865), .A(n20797), .B(n20796), .ZN(
        P1_U3145) );
  AOI22_X1 U23750 ( .A1(n20836), .A2(n20812), .B1(n20835), .B2(n20811), .ZN(
        n20799) );
  AOI22_X1 U23751 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20814), .B1(
        n20878), .B2(n20837), .ZN(n20798) );
  OAI211_X1 U23752 ( .C1(n20840), .C2(n20808), .A(n20799), .B(n20798), .ZN(
        P1_U3146) );
  AOI22_X1 U23753 ( .A1(n20842), .A2(n20812), .B1(n20841), .B2(n20811), .ZN(
        n20801) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20814), .B1(
        n20878), .B2(n20843), .ZN(n20800) );
  OAI211_X1 U23755 ( .C1(n20846), .C2(n20808), .A(n20801), .B(n20800), .ZN(
        P1_U3147) );
  AOI22_X1 U23756 ( .A1(n20848), .A2(n20812), .B1(n20847), .B2(n20811), .ZN(
        n20803) );
  AOI22_X1 U23757 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20814), .B1(
        n20878), .B2(n20849), .ZN(n20802) );
  OAI211_X1 U23758 ( .C1(n20852), .C2(n20808), .A(n20803), .B(n20802), .ZN(
        P1_U3148) );
  AOI22_X1 U23759 ( .A1(n20854), .A2(n20812), .B1(n20853), .B2(n20811), .ZN(
        n20805) );
  AOI22_X1 U23760 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20814), .B1(
        n20813), .B2(n20855), .ZN(n20804) );
  OAI211_X1 U23761 ( .C1(n20858), .C2(n20865), .A(n20805), .B(n20804), .ZN(
        P1_U3149) );
  AOI22_X1 U23762 ( .A1(n20860), .A2(n20812), .B1(n20859), .B2(n20811), .ZN(
        n20807) );
  AOI22_X1 U23763 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20814), .B1(
        n20878), .B2(n20861), .ZN(n20806) );
  OAI211_X1 U23764 ( .C1(n20866), .C2(n20808), .A(n20807), .B(n20806), .ZN(
        P1_U3150) );
  AOI22_X1 U23765 ( .A1(n20868), .A2(n20812), .B1(n20867), .B2(n20811), .ZN(
        n20810) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20814), .B1(
        n20813), .B2(n20869), .ZN(n20809) );
  OAI211_X1 U23767 ( .C1(n20872), .C2(n20865), .A(n20810), .B(n20809), .ZN(
        P1_U3151) );
  AOI22_X1 U23768 ( .A1(n20876), .A2(n20812), .B1(n20874), .B2(n20811), .ZN(
        n20816) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20814), .B1(
        n20813), .B2(n20877), .ZN(n20815) );
  OAI211_X1 U23770 ( .C1(n20883), .C2(n20865), .A(n20816), .B(n20815), .ZN(
        P1_U3152) );
  AOI21_X1 U23771 ( .B1(n20818), .B2(n20817), .A(n20873), .ZN(n20824) );
  OAI22_X1 U23772 ( .A1(n20824), .A2(n20822), .B1(n20821), .B2(n20888), .ZN(
        n20875) );
  AOI22_X1 U23773 ( .A1(n20820), .A2(n20875), .B1(n20819), .B2(n20873), .ZN(
        n20833) );
  INV_X1 U23774 ( .A(n20821), .ZN(n20830) );
  NOR2_X1 U23775 ( .A1(n20823), .A2(n20822), .ZN(n20826) );
  OAI21_X1 U23776 ( .B1(n20826), .B2(n20825), .A(n20824), .ZN(n20827) );
  OAI211_X1 U23777 ( .C1(n20830), .C2(n20829), .A(n20828), .B(n20827), .ZN(
        n20879) );
  AOI22_X1 U23778 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20879), .B1(
        n20878), .B2(n20831), .ZN(n20832) );
  OAI211_X1 U23779 ( .C1(n20834), .C2(n20882), .A(n20833), .B(n20832), .ZN(
        P1_U3153) );
  AOI22_X1 U23780 ( .A1(n20836), .A2(n20875), .B1(n20835), .B2(n20873), .ZN(
        n20839) );
  AOI22_X1 U23781 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20879), .B1(
        n20862), .B2(n20837), .ZN(n20838) );
  OAI211_X1 U23782 ( .C1(n20840), .C2(n20865), .A(n20839), .B(n20838), .ZN(
        P1_U3154) );
  AOI22_X1 U23783 ( .A1(n20842), .A2(n20875), .B1(n20841), .B2(n20873), .ZN(
        n20845) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20879), .B1(
        n20862), .B2(n20843), .ZN(n20844) );
  OAI211_X1 U23785 ( .C1(n20846), .C2(n20865), .A(n20845), .B(n20844), .ZN(
        P1_U3155) );
  AOI22_X1 U23786 ( .A1(n20848), .A2(n20875), .B1(n20847), .B2(n20873), .ZN(
        n20851) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20879), .B1(
        n20862), .B2(n20849), .ZN(n20850) );
  OAI211_X1 U23788 ( .C1(n20852), .C2(n20865), .A(n20851), .B(n20850), .ZN(
        P1_U3156) );
  AOI22_X1 U23789 ( .A1(n20854), .A2(n20875), .B1(n20853), .B2(n20873), .ZN(
        n20857) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20879), .B1(
        n20878), .B2(n20855), .ZN(n20856) );
  OAI211_X1 U23791 ( .C1(n20858), .C2(n20882), .A(n20857), .B(n20856), .ZN(
        P1_U3157) );
  AOI22_X1 U23792 ( .A1(n20860), .A2(n20875), .B1(n20859), .B2(n20873), .ZN(
        n20864) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20879), .B1(
        n20862), .B2(n20861), .ZN(n20863) );
  OAI211_X1 U23794 ( .C1(n20866), .C2(n20865), .A(n20864), .B(n20863), .ZN(
        P1_U3158) );
  AOI22_X1 U23795 ( .A1(n20868), .A2(n20875), .B1(n20867), .B2(n20873), .ZN(
        n20871) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20879), .B1(
        n20878), .B2(n20869), .ZN(n20870) );
  OAI211_X1 U23797 ( .C1(n20872), .C2(n20882), .A(n20871), .B(n20870), .ZN(
        P1_U3159) );
  AOI22_X1 U23798 ( .A1(n20876), .A2(n20875), .B1(n20874), .B2(n20873), .ZN(
        n20881) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20879), .B1(
        n20878), .B2(n20877), .ZN(n20880) );
  OAI211_X1 U23800 ( .C1(n20883), .C2(n20882), .A(n20881), .B(n20880), .ZN(
        P1_U3160) );
  NOR2_X1 U23801 ( .A1(n20885), .A2(n20884), .ZN(n20889) );
  INV_X1 U23802 ( .A(n20886), .ZN(n20887) );
  OAI21_X1 U23803 ( .B1(n20889), .B2(n20888), .A(n20887), .ZN(P1_U3163) );
  INV_X1 U23804 ( .A(n20965), .ZN(n20961) );
  AND2_X1 U23805 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20961), .ZN(
        P1_U3164) );
  AND2_X1 U23806 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20961), .ZN(
        P1_U3165) );
  AND2_X1 U23807 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20961), .ZN(
        P1_U3166) );
  AND2_X1 U23808 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20961), .ZN(
        P1_U3167) );
  AND2_X1 U23809 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20961), .ZN(
        P1_U3168) );
  AND2_X1 U23810 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20961), .ZN(
        P1_U3169) );
  AND2_X1 U23811 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20961), .ZN(
        P1_U3170) );
  AND2_X1 U23812 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20961), .ZN(
        P1_U3171) );
  AND2_X1 U23813 ( .A1(n20961), .A2(P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(
        P1_U3172) );
  AND2_X1 U23814 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20961), .ZN(
        P1_U3173) );
  AND2_X1 U23815 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20961), .ZN(
        P1_U3174) );
  AND2_X1 U23816 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20961), .ZN(
        P1_U3175) );
  AND2_X1 U23817 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20961), .ZN(
        P1_U3176) );
  AND2_X1 U23818 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20961), .ZN(
        P1_U3177) );
  AND2_X1 U23819 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20961), .ZN(
        P1_U3178) );
  AND2_X1 U23820 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20961), .ZN(
        P1_U3179) );
  AND2_X1 U23821 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20961), .ZN(
        P1_U3180) );
  AND2_X1 U23822 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20961), .ZN(
        P1_U3181) );
  AND2_X1 U23823 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20961), .ZN(
        P1_U3182) );
  AND2_X1 U23824 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20961), .ZN(
        P1_U3183) );
  AND2_X1 U23825 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20961), .ZN(
        P1_U3184) );
  AND2_X1 U23826 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20961), .ZN(
        P1_U3185) );
  AND2_X1 U23827 ( .A1(n20961), .A2(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(P1_U3186) );
  AND2_X1 U23828 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20961), .ZN(P1_U3187) );
  AND2_X1 U23829 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20961), .ZN(P1_U3188) );
  AND2_X1 U23830 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20961), .ZN(P1_U3189) );
  AND2_X1 U23831 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20961), .ZN(P1_U3190) );
  AND2_X1 U23832 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20961), .ZN(P1_U3191) );
  AND2_X1 U23833 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20961), .ZN(P1_U3192) );
  AND2_X1 U23834 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20961), .ZN(P1_U3193) );
  AOI21_X1 U23835 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20890), .A(n20897), 
        .ZN(n20904) );
  NOR2_X1 U23836 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20891) );
  NOR2_X1 U23837 ( .A1(n20891), .A2(n20902), .ZN(n20892) );
  AOI211_X1 U23838 ( .C1(NA), .C2(n20897), .A(n20892), .B(n20898), .ZN(n20893)
         );
  OAI22_X1 U23839 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20904), .B1(n20988), 
        .B2(n20893), .ZN(P1_U3194) );
  NOR2_X1 U23840 ( .A1(NA), .A2(n20898), .ZN(n20896) );
  AOI21_X1 U23841 ( .B1(NA), .B2(n20894), .A(n20905), .ZN(n20895) );
  AOI21_X1 U23842 ( .B1(n20896), .B2(P1_STATE_REG_0__SCAN_IN), .A(n20895), 
        .ZN(n20903) );
  NOR3_X1 U23843 ( .A1(NA), .A2(n20897), .A3(n20978), .ZN(n20899) );
  OAI22_X1 U23844 ( .A1(n20900), .A2(n20899), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20898), .ZN(n20901) );
  OAI22_X1 U23845 ( .A1(n20904), .A2(n20903), .B1(n20902), .B2(n20901), .ZN(
        P1_U3196) );
  NAND2_X1 U23846 ( .A1(n20988), .A2(n20905), .ZN(n20950) );
  INV_X1 U23847 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20906) );
  NAND2_X1 U23848 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20988), .ZN(n20953) );
  OAI222_X1 U23849 ( .A1(n20950), .A2(n20908), .B1(n20906), .B2(n20988), .C1(
        n20966), .C2(n20953), .ZN(P1_U3197) );
  INV_X1 U23850 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20907) );
  OAI222_X1 U23851 ( .A1(n20953), .A2(n20908), .B1(n20907), .B2(n20988), .C1(
        n14655), .C2(n20950), .ZN(P1_U3198) );
  OAI222_X1 U23852 ( .A1(n20953), .A2(n14655), .B1(n20909), .B2(n20988), .C1(
        n20910), .C2(n20950), .ZN(P1_U3199) );
  INV_X1 U23853 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20911) );
  OAI222_X1 U23854 ( .A1(n20950), .A2(n21198), .B1(n20911), .B2(n20988), .C1(
        n20910), .C2(n20953), .ZN(P1_U3200) );
  INV_X1 U23855 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20912) );
  OAI222_X1 U23856 ( .A1(n20950), .A2(n20914), .B1(n20912), .B2(n20988), .C1(
        n21198), .C2(n20953), .ZN(P1_U3201) );
  INV_X1 U23857 ( .A(n20950), .ZN(n20942) );
  AOI22_X1 U23858 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20974), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20942), .ZN(n20913) );
  OAI21_X1 U23859 ( .B1(n20914), .B2(n20953), .A(n20913), .ZN(P1_U3202) );
  INV_X1 U23860 ( .A(n20953), .ZN(n20945) );
  AOI22_X1 U23861 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20974), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20945), .ZN(n20915) );
  OAI21_X1 U23862 ( .B1(n20917), .B2(n20950), .A(n20915), .ZN(P1_U3203) );
  INV_X1 U23863 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20916) );
  OAI222_X1 U23864 ( .A1(n20953), .A2(n20917), .B1(n20916), .B2(n20988), .C1(
        n21146), .C2(n20950), .ZN(P1_U3204) );
  AOI222_X1 U23865 ( .A1(n20945), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20974), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20942), .ZN(n20918) );
  INV_X1 U23866 ( .A(n20918), .ZN(P1_U3205) );
  AOI222_X1 U23867 ( .A1(n20945), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20974), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20942), .ZN(n20919) );
  INV_X1 U23868 ( .A(n20919), .ZN(P1_U3206) );
  AOI222_X1 U23869 ( .A1(n20942), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20974), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20945), .ZN(n20920) );
  INV_X1 U23870 ( .A(n20920), .ZN(P1_U3207) );
  AOI222_X1 U23871 ( .A1(n20942), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20974), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20945), .ZN(n20921) );
  INV_X1 U23872 ( .A(n20921), .ZN(P1_U3208) );
  INV_X1 U23873 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20922) );
  OAI222_X1 U23874 ( .A1(n20953), .A2(n20923), .B1(n20922), .B2(n20988), .C1(
        n20924), .C2(n20950), .ZN(P1_U3209) );
  INV_X1 U23875 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20925) );
  OAI222_X1 U23876 ( .A1(n20950), .A2(n20927), .B1(n20925), .B2(n20988), .C1(
        n20924), .C2(n20953), .ZN(P1_U3210) );
  AOI22_X1 U23877 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20974), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20942), .ZN(n20926) );
  OAI21_X1 U23878 ( .B1(n20927), .B2(n20953), .A(n20926), .ZN(P1_U3211) );
  AOI22_X1 U23879 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20974), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20945), .ZN(n20928) );
  OAI21_X1 U23880 ( .B1(n20929), .B2(n20950), .A(n20928), .ZN(P1_U3212) );
  INV_X1 U23881 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20930) );
  OAI222_X1 U23882 ( .A1(n20950), .A2(n20932), .B1(n20930), .B2(n20988), .C1(
        n20929), .C2(n20953), .ZN(P1_U3213) );
  AOI22_X1 U23883 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20974), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20942), .ZN(n20931) );
  OAI21_X1 U23884 ( .B1(n20932), .B2(n20953), .A(n20931), .ZN(P1_U3214) );
  INV_X1 U23885 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20935) );
  AOI22_X1 U23886 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20974), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20945), .ZN(n20933) );
  OAI21_X1 U23887 ( .B1(n20935), .B2(n20950), .A(n20933), .ZN(P1_U3215) );
  INV_X1 U23888 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20934) );
  OAI222_X1 U23889 ( .A1(n20953), .A2(n20935), .B1(n20934), .B2(n20988), .C1(
        n20937), .C2(n20950), .ZN(P1_U3216) );
  INV_X1 U23890 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20936) );
  OAI222_X1 U23891 ( .A1(n20953), .A2(n20937), .B1(n20936), .B2(n20988), .C1(
        n21230), .C2(n20950), .ZN(P1_U3217) );
  INV_X1 U23892 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20938) );
  INV_X1 U23893 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21170) );
  OAI222_X1 U23894 ( .A1(n20953), .A2(n21230), .B1(n20938), .B2(n20988), .C1(
        n21170), .C2(n20950), .ZN(P1_U3218) );
  AOI222_X1 U23895 ( .A1(n20945), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20974), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20942), .ZN(n20939) );
  INV_X1 U23896 ( .A(n20939), .ZN(P1_U3219) );
  AOI222_X1 U23897 ( .A1(n20945), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20974), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20942), .ZN(n20940) );
  INV_X1 U23898 ( .A(n20940), .ZN(P1_U3220) );
  INV_X1 U23899 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20941) );
  OAI222_X1 U23900 ( .A1(n20953), .A2(n21204), .B1(n20941), .B2(n20988), .C1(
        n20944), .C2(n20950), .ZN(P1_U3221) );
  AOI22_X1 U23901 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20942), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20974), .ZN(n20943) );
  OAI21_X1 U23902 ( .B1(n20944), .B2(n20953), .A(n20943), .ZN(P1_U3222) );
  AOI22_X1 U23903 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20945), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20974), .ZN(n20946) );
  OAI21_X1 U23904 ( .B1(n20948), .B2(n20950), .A(n20946), .ZN(P1_U3223) );
  INV_X1 U23905 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20947) );
  OAI222_X1 U23906 ( .A1(n20953), .A2(n20948), .B1(n20947), .B2(n20988), .C1(
        n21143), .C2(n20950), .ZN(P1_U3224) );
  INV_X1 U23907 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20949) );
  OAI222_X1 U23908 ( .A1(n20950), .A2(n21043), .B1(n20949), .B2(n20988), .C1(
        n21143), .C2(n20953), .ZN(P1_U3225) );
  INV_X1 U23909 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20952) );
  OAI222_X1 U23910 ( .A1(n20953), .A2(n21043), .B1(n20952), .B2(n20988), .C1(
        n20951), .C2(n20950), .ZN(P1_U3226) );
  INV_X1 U23911 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20954) );
  AOI22_X1 U23912 ( .A1(n20988), .A2(n20955), .B1(n20954), .B2(n20974), .ZN(
        P1_U3458) );
  INV_X1 U23913 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20968) );
  INV_X1 U23914 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20956) );
  AOI22_X1 U23915 ( .A1(n20988), .A2(n20968), .B1(n20956), .B2(n20974), .ZN(
        P1_U3459) );
  INV_X1 U23916 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20957) );
  AOI22_X1 U23917 ( .A1(n20988), .A2(n20958), .B1(n20957), .B2(n20974), .ZN(
        P1_U3460) );
  INV_X1 U23918 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20973) );
  INV_X1 U23919 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20959) );
  AOI22_X1 U23920 ( .A1(n20988), .A2(n20973), .B1(n20959), .B2(n20974), .ZN(
        P1_U3461) );
  INV_X1 U23921 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20962) );
  INV_X1 U23922 ( .A(n20963), .ZN(n20960) );
  AOI21_X1 U23923 ( .B1(n20962), .B2(n20961), .A(n20960), .ZN(P1_U3464) );
  OAI21_X1 U23924 ( .B1(n20965), .B2(n20964), .A(n20963), .ZN(P1_U3465) );
  AOI21_X1 U23925 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20967) );
  AOI22_X1 U23926 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20967), .B2(n20966), .ZN(n20969) );
  AOI22_X1 U23927 ( .A1(n20970), .A2(n20969), .B1(n20968), .B2(n20972), .ZN(
        P1_U3481) );
  NOR2_X1 U23928 ( .A1(n20972), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20971) );
  AOI22_X1 U23929 ( .A1(n20973), .A2(n20972), .B1(n13803), .B2(n20971), .ZN(
        P1_U3482) );
  AOI22_X1 U23930 ( .A1(n20988), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20975), 
        .B2(n20974), .ZN(P1_U3483) );
  AOI211_X1 U23931 ( .C1(n20979), .C2(n20978), .A(n20977), .B(n20976), .ZN(
        n20987) );
  INV_X1 U23932 ( .A(n20980), .ZN(n20981) );
  OAI211_X1 U23933 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20982), .A(n20981), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20984) );
  AOI21_X1 U23934 ( .B1(n20984), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20983), 
        .ZN(n20986) );
  NAND2_X1 U23935 ( .A1(n20987), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20985) );
  OAI21_X1 U23936 ( .B1(n20987), .B2(n20986), .A(n20985), .ZN(P1_U3485) );
  MUX2_X1 U23937 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20988), .Z(P1_U3486) );
  NAND2_X1 U23938 ( .A1(n20990), .A2(n20989), .ZN(n20994) );
  AOI21_X1 U23939 ( .B1(n20992), .B2(n20995), .A(n20991), .ZN(n20993) );
  AOI21_X1 U23940 ( .B1(n20995), .B2(n20994), .A(n20993), .ZN(n21308) );
  AOI22_X1 U23941 ( .A1(n10916), .A2(keyinput113), .B1(keyinput93), .B2(n20997), .ZN(n20996) );
  OAI221_X1 U23942 ( .B1(n10916), .B2(keyinput113), .C1(n20997), .C2(
        keyinput93), .A(n20996), .ZN(n21009) );
  AOI22_X1 U23943 ( .A1(n20999), .A2(keyinput49), .B1(keyinput12), .B2(n13697), 
        .ZN(n20998) );
  OAI221_X1 U23944 ( .B1(n20999), .B2(keyinput49), .C1(n13697), .C2(keyinput12), .A(n20998), .ZN(n21008) );
  INV_X1 U23945 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n21002) );
  INV_X1 U23946 ( .A(keyinput10), .ZN(n21001) );
  AOI22_X1 U23947 ( .A1(n21002), .A2(keyinput7), .B1(
        P2_DATAWIDTH_REG_2__SCAN_IN), .B2(n21001), .ZN(n21000) );
  OAI221_X1 U23948 ( .B1(n21002), .B2(keyinput7), .C1(n21001), .C2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A(n21000), .ZN(n21007) );
  INV_X1 U23949 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n21005) );
  INV_X1 U23950 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n21004) );
  AOI22_X1 U23951 ( .A1(n21005), .A2(keyinput87), .B1(keyinput52), .B2(n21004), 
        .ZN(n21003) );
  OAI221_X1 U23952 ( .B1(n21005), .B2(keyinput87), .C1(n21004), .C2(keyinput52), .A(n21003), .ZN(n21006) );
  NOR4_X1 U23953 ( .A1(n21009), .A2(n21008), .A3(n21007), .A4(n21006), .ZN(
        n21057) );
  INV_X1 U23954 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U23955 ( .A1(n21012), .A2(keyinput16), .B1(n21011), .B2(keyinput78), 
        .ZN(n21010) );
  OAI221_X1 U23956 ( .B1(n21012), .B2(keyinput16), .C1(n21011), .C2(keyinput78), .A(n21010), .ZN(n21025) );
  INV_X1 U23957 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21014) );
  AOI22_X1 U23958 ( .A1(n21015), .A2(keyinput71), .B1(keyinput104), .B2(n21014), .ZN(n21013) );
  OAI221_X1 U23959 ( .B1(n21015), .B2(keyinput71), .C1(n21014), .C2(
        keyinput104), .A(n21013), .ZN(n21024) );
  AOI22_X1 U23960 ( .A1(n21018), .A2(keyinput26), .B1(keyinput116), .B2(n21017), .ZN(n21016) );
  OAI221_X1 U23961 ( .B1(n21018), .B2(keyinput26), .C1(n21017), .C2(
        keyinput116), .A(n21016), .ZN(n21023) );
  INV_X1 U23962 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n21021) );
  AOI22_X1 U23963 ( .A1(n21021), .A2(keyinput82), .B1(keyinput38), .B2(n21020), 
        .ZN(n21019) );
  OAI221_X1 U23964 ( .B1(n21021), .B2(keyinput82), .C1(n21020), .C2(keyinput38), .A(n21019), .ZN(n21022) );
  NOR4_X1 U23965 ( .A1(n21025), .A2(n21024), .A3(n21023), .A4(n21022), .ZN(
        n21056) );
  AOI22_X1 U23966 ( .A1(n13499), .A2(keyinput101), .B1(n21027), .B2(
        keyinput127), .ZN(n21026) );
  OAI221_X1 U23967 ( .B1(n13499), .B2(keyinput101), .C1(n21027), .C2(
        keyinput127), .A(n21026), .ZN(n21038) );
  AOI22_X1 U23968 ( .A1(n21029), .A2(keyinput108), .B1(keyinput80), .B2(n13529), .ZN(n21028) );
  OAI221_X1 U23969 ( .B1(n21029), .B2(keyinput108), .C1(n13529), .C2(
        keyinput80), .A(n21028), .ZN(n21037) );
  INV_X1 U23970 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n21032) );
  INV_X1 U23971 ( .A(DATAI_22_), .ZN(n21031) );
  AOI22_X1 U23972 ( .A1(n21032), .A2(keyinput123), .B1(keyinput124), .B2(
        n21031), .ZN(n21030) );
  OAI221_X1 U23973 ( .B1(n21032), .B2(keyinput123), .C1(n21031), .C2(
        keyinput124), .A(n21030), .ZN(n21036) );
  XNOR2_X1 U23974 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput110), 
        .ZN(n21034) );
  XNOR2_X1 U23975 ( .A(keyinput11), .B(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n21033) );
  NAND2_X1 U23976 ( .A1(n21034), .A2(n21033), .ZN(n21035) );
  NOR4_X1 U23977 ( .A1(n21038), .A2(n21037), .A3(n21036), .A4(n21035), .ZN(
        n21055) );
  INV_X1 U23978 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n21040) );
  AOI22_X1 U23979 ( .A1(n21041), .A2(keyinput79), .B1(n21040), .B2(keyinput19), 
        .ZN(n21039) );
  OAI221_X1 U23980 ( .B1(n21041), .B2(keyinput79), .C1(n21040), .C2(keyinput19), .A(n21039), .ZN(n21053) );
  AOI22_X1 U23981 ( .A1(n21043), .A2(keyinput31), .B1(n12775), .B2(keyinput83), 
        .ZN(n21042) );
  OAI221_X1 U23982 ( .B1(n21043), .B2(keyinput31), .C1(n12775), .C2(keyinput83), .A(n21042), .ZN(n21052) );
  INV_X1 U23983 ( .A(DATAI_26_), .ZN(n21045) );
  AOI22_X1 U23984 ( .A1(n21046), .A2(keyinput23), .B1(keyinput56), .B2(n21045), 
        .ZN(n21044) );
  OAI221_X1 U23985 ( .B1(n21046), .B2(keyinput23), .C1(n21045), .C2(keyinput56), .A(n21044), .ZN(n21051) );
  AOI22_X1 U23986 ( .A1(n21049), .A2(keyinput65), .B1(n21048), .B2(keyinput46), 
        .ZN(n21047) );
  OAI221_X1 U23987 ( .B1(n21049), .B2(keyinput65), .C1(n21048), .C2(keyinput46), .A(n21047), .ZN(n21050) );
  NOR4_X1 U23988 ( .A1(n21053), .A2(n21052), .A3(n21051), .A4(n21050), .ZN(
        n21054) );
  NAND4_X1 U23989 ( .A1(n21057), .A2(n21056), .A3(n21055), .A4(n21054), .ZN(
        n21306) );
  INV_X1 U23990 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n21060) );
  INV_X1 U23991 ( .A(keyinput119), .ZN(n21059) );
  AOI22_X1 U23992 ( .A1(n21060), .A2(keyinput2), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n21059), .ZN(n21058) );
  OAI221_X1 U23993 ( .B1(n21060), .B2(keyinput2), .C1(n21059), .C2(
        P3_ADDRESS_REG_21__SCAN_IN), .A(n21058), .ZN(n21073) );
  AOI22_X1 U23994 ( .A1(n21063), .A2(keyinput100), .B1(keyinput47), .B2(n21062), .ZN(n21061) );
  OAI221_X1 U23995 ( .B1(n21063), .B2(keyinput100), .C1(n21062), .C2(
        keyinput47), .A(n21061), .ZN(n21072) );
  INV_X1 U23996 ( .A(DATAI_7_), .ZN(n21065) );
  AOI22_X1 U23997 ( .A1(n21066), .A2(keyinput55), .B1(n21065), .B2(keyinput35), 
        .ZN(n21064) );
  OAI221_X1 U23998 ( .B1(n21066), .B2(keyinput55), .C1(n21065), .C2(keyinput35), .A(n21064), .ZN(n21071) );
  INV_X1 U23999 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n21069) );
  INV_X1 U24000 ( .A(keyinput32), .ZN(n21068) );
  AOI22_X1 U24001 ( .A1(n21069), .A2(keyinput94), .B1(HOLD), .B2(n21068), .ZN(
        n21067) );
  OAI221_X1 U24002 ( .B1(n21069), .B2(keyinput94), .C1(n21068), .C2(HOLD), .A(
        n21067), .ZN(n21070) );
  NOR4_X1 U24003 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        n21122) );
  INV_X1 U24004 ( .A(DATAI_23_), .ZN(n21076) );
  INV_X1 U24005 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21075) );
  AOI22_X1 U24006 ( .A1(n21076), .A2(keyinput76), .B1(n21075), .B2(keyinput98), 
        .ZN(n21074) );
  OAI221_X1 U24007 ( .B1(n21076), .B2(keyinput76), .C1(n21075), .C2(keyinput98), .A(n21074), .ZN(n21089) );
  INV_X1 U24008 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n21079) );
  AOI22_X1 U24009 ( .A1(n21079), .A2(keyinput60), .B1(keyinput75), .B2(n21078), 
        .ZN(n21077) );
  OAI221_X1 U24010 ( .B1(n21079), .B2(keyinput60), .C1(n21078), .C2(keyinput75), .A(n21077), .ZN(n21088) );
  INV_X1 U24011 ( .A(keyinput111), .ZN(n21081) );
  AOI22_X1 U24012 ( .A1(n21082), .A2(keyinput1), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n21081), .ZN(n21080) );
  OAI221_X1 U24013 ( .B1(n21082), .B2(keyinput1), .C1(n21081), .C2(
        P3_ADDRESS_REG_20__SCAN_IN), .A(n21080), .ZN(n21087) );
  INV_X1 U24014 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n21085) );
  INV_X1 U24015 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n21084) );
  AOI22_X1 U24016 ( .A1(n21085), .A2(keyinput20), .B1(keyinput29), .B2(n21084), 
        .ZN(n21083) );
  OAI221_X1 U24017 ( .B1(n21085), .B2(keyinput20), .C1(n21084), .C2(keyinput29), .A(n21083), .ZN(n21086) );
  NOR4_X1 U24018 ( .A1(n21089), .A2(n21088), .A3(n21087), .A4(n21086), .ZN(
        n21121) );
  INV_X1 U24019 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n21091) );
  AOI22_X1 U24020 ( .A1(n10922), .A2(keyinput125), .B1(keyinput8), .B2(n21091), 
        .ZN(n21090) );
  OAI221_X1 U24021 ( .B1(n10922), .B2(keyinput125), .C1(n21091), .C2(keyinput8), .A(n21090), .ZN(n21104) );
  INV_X1 U24022 ( .A(keyinput43), .ZN(n21093) );
  AOI22_X1 U24023 ( .A1(n21094), .A2(keyinput6), .B1(
        P2_DATAWIDTH_REG_24__SCAN_IN), .B2(n21093), .ZN(n21092) );
  OAI221_X1 U24024 ( .B1(n21094), .B2(keyinput6), .C1(n21093), .C2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A(n21092), .ZN(n21103) );
  AOI22_X1 U24025 ( .A1(n21097), .A2(keyinput51), .B1(n21096), .B2(keyinput117), .ZN(n21095) );
  OAI221_X1 U24026 ( .B1(n21097), .B2(keyinput51), .C1(n21096), .C2(
        keyinput117), .A(n21095), .ZN(n21102) );
  INV_X1 U24027 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n21100) );
  AOI22_X1 U24028 ( .A1(n21100), .A2(keyinput88), .B1(keyinput14), .B2(n21099), 
        .ZN(n21098) );
  OAI221_X1 U24029 ( .B1(n21100), .B2(keyinput88), .C1(n21099), .C2(keyinput14), .A(n21098), .ZN(n21101) );
  NOR4_X1 U24030 ( .A1(n21104), .A2(n21103), .A3(n21102), .A4(n21101), .ZN(
        n21120) );
  INV_X1 U24031 ( .A(keyinput90), .ZN(n21106) );
  AOI22_X1 U24032 ( .A1(n12162), .A2(keyinput66), .B1(
        P3_DATAWIDTH_REG_13__SCAN_IN), .B2(n21106), .ZN(n21105) );
  OAI221_X1 U24033 ( .B1(n12162), .B2(keyinput66), .C1(n21106), .C2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A(n21105), .ZN(n21118) );
  INV_X1 U24034 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n21109) );
  INV_X1 U24035 ( .A(keyinput50), .ZN(n21108) );
  AOI22_X1 U24036 ( .A1(n21109), .A2(keyinput13), .B1(P3_DATAO_REG_3__SCAN_IN), 
        .B2(n21108), .ZN(n21107) );
  OAI221_X1 U24037 ( .B1(n21109), .B2(keyinput13), .C1(n21108), .C2(
        P3_DATAO_REG_3__SCAN_IN), .A(n21107), .ZN(n21117) );
  AOI22_X1 U24038 ( .A1(n21112), .A2(keyinput39), .B1(keyinput28), .B2(n21111), 
        .ZN(n21110) );
  OAI221_X1 U24039 ( .B1(n21112), .B2(keyinput39), .C1(n21111), .C2(keyinput28), .A(n21110), .ZN(n21116) );
  INV_X1 U24040 ( .A(keyinput120), .ZN(n21114) );
  AOI22_X1 U24041 ( .A1(n9910), .A2(keyinput42), .B1(
        P1_DATAWIDTH_REG_23__SCAN_IN), .B2(n21114), .ZN(n21113) );
  OAI221_X1 U24042 ( .B1(n9910), .B2(keyinput42), .C1(n21114), .C2(
        P1_DATAWIDTH_REG_23__SCAN_IN), .A(n21113), .ZN(n21115) );
  NOR4_X1 U24043 ( .A1(n21118), .A2(n21117), .A3(n21116), .A4(n21115), .ZN(
        n21119) );
  NAND4_X1 U24044 ( .A1(n21122), .A2(n21121), .A3(n21120), .A4(n21119), .ZN(
        n21305) );
  INV_X1 U24045 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n21124) );
  AOI22_X1 U24046 ( .A1(n21125), .A2(keyinput27), .B1(n21124), .B2(keyinput22), 
        .ZN(n21123) );
  OAI221_X1 U24047 ( .B1(n21125), .B2(keyinput27), .C1(n21124), .C2(keyinput22), .A(n21123), .ZN(n21138) );
  INV_X1 U24048 ( .A(READY12_REG_SCAN_IN), .ZN(n21128) );
  AOI22_X1 U24049 ( .A1(n21128), .A2(keyinput96), .B1(keyinput81), .B2(n21127), 
        .ZN(n21126) );
  OAI221_X1 U24050 ( .B1(n21128), .B2(keyinput96), .C1(n21127), .C2(keyinput81), .A(n21126), .ZN(n21137) );
  INV_X1 U24051 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n21131) );
  INV_X1 U24052 ( .A(keyinput85), .ZN(n21130) );
  AOI22_X1 U24053 ( .A1(n21131), .A2(keyinput17), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n21130), .ZN(n21129) );
  OAI221_X1 U24054 ( .B1(n21131), .B2(keyinput17), .C1(n21130), .C2(
        P3_ADDRESS_REG_0__SCAN_IN), .A(n21129), .ZN(n21136) );
  AOI22_X1 U24055 ( .A1(n21134), .A2(keyinput33), .B1(n21133), .B2(keyinput59), 
        .ZN(n21132) );
  OAI221_X1 U24056 ( .B1(n21134), .B2(keyinput33), .C1(n21133), .C2(keyinput59), .A(n21132), .ZN(n21135) );
  NOR4_X1 U24057 ( .A1(n21138), .A2(n21137), .A3(n21136), .A4(n21135), .ZN(
        n21187) );
  AOI22_X1 U24058 ( .A1(n10917), .A2(keyinput73), .B1(keyinput92), .B2(n21140), 
        .ZN(n21139) );
  OAI221_X1 U24059 ( .B1(n10917), .B2(keyinput73), .C1(n21140), .C2(keyinput92), .A(n21139), .ZN(n21152) );
  AOI22_X1 U24060 ( .A1(n21143), .A2(keyinput36), .B1(n21142), .B2(keyinput77), 
        .ZN(n21141) );
  OAI221_X1 U24061 ( .B1(n21143), .B2(keyinput36), .C1(n21142), .C2(keyinput77), .A(n21141), .ZN(n21151) );
  AOI22_X1 U24062 ( .A1(n21146), .A2(keyinput74), .B1(keyinput0), .B2(n21145), 
        .ZN(n21144) );
  OAI221_X1 U24063 ( .B1(n21146), .B2(keyinput74), .C1(n21145), .C2(keyinput0), 
        .A(n21144), .ZN(n21150) );
  AOI22_X1 U24064 ( .A1(n12284), .A2(keyinput18), .B1(keyinput121), .B2(n21148), .ZN(n21147) );
  OAI221_X1 U24065 ( .B1(n12284), .B2(keyinput18), .C1(n21148), .C2(
        keyinput121), .A(n21147), .ZN(n21149) );
  NOR4_X1 U24066 ( .A1(n21152), .A2(n21151), .A3(n21150), .A4(n21149), .ZN(
        n21186) );
  INV_X1 U24067 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n21155) );
  INV_X1 U24068 ( .A(keyinput40), .ZN(n21154) );
  AOI22_X1 U24069 ( .A1(n21155), .A2(keyinput105), .B1(
        P2_DATAWIDTH_REG_4__SCAN_IN), .B2(n21154), .ZN(n21153) );
  OAI221_X1 U24070 ( .B1(n21155), .B2(keyinput105), .C1(n21154), .C2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A(n21153), .ZN(n21167) );
  INV_X1 U24071 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n21157) );
  AOI22_X1 U24072 ( .A1(n21158), .A2(keyinput4), .B1(keyinput91), .B2(n21157), 
        .ZN(n21156) );
  OAI221_X1 U24073 ( .B1(n21158), .B2(keyinput4), .C1(n21157), .C2(keyinput91), 
        .A(n21156), .ZN(n21166) );
  INV_X1 U24074 ( .A(keyinput44), .ZN(n21160) );
  AOI22_X1 U24075 ( .A1(n21161), .A2(keyinput5), .B1(
        P3_DATAWIDTH_REG_20__SCAN_IN), .B2(n21160), .ZN(n21159) );
  OAI221_X1 U24076 ( .B1(n21161), .B2(keyinput5), .C1(n21160), .C2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A(n21159), .ZN(n21165) );
  INV_X1 U24077 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n21163) );
  AOI22_X1 U24078 ( .A1(n21163), .A2(keyinput107), .B1(keyinput109), .B2(
        n13492), .ZN(n21162) );
  OAI221_X1 U24079 ( .B1(n21163), .B2(keyinput107), .C1(n13492), .C2(
        keyinput109), .A(n21162), .ZN(n21164) );
  NOR4_X1 U24080 ( .A1(n21167), .A2(n21166), .A3(n21165), .A4(n21164), .ZN(
        n21185) );
  INV_X1 U24081 ( .A(keyinput21), .ZN(n21169) );
  AOI22_X1 U24082 ( .A1(n21170), .A2(keyinput25), .B1(P3_DATAO_REG_20__SCAN_IN), .B2(n21169), .ZN(n21168) );
  OAI221_X1 U24083 ( .B1(n21170), .B2(keyinput25), .C1(n21169), .C2(
        P3_DATAO_REG_20__SCAN_IN), .A(n21168), .ZN(n21183) );
  INV_X1 U24084 ( .A(DATAI_27_), .ZN(n21173) );
  INV_X1 U24085 ( .A(keyinput45), .ZN(n21172) );
  AOI22_X1 U24086 ( .A1(n21173), .A2(keyinput64), .B1(
        P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n21172), .ZN(n21171) );
  OAI221_X1 U24087 ( .B1(n21173), .B2(keyinput64), .C1(n21172), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(n21171), .ZN(n21182) );
  INV_X1 U24088 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n21176) );
  INV_X1 U24089 ( .A(keyinput48), .ZN(n21175) );
  AOI22_X1 U24090 ( .A1(n21176), .A2(keyinput122), .B1(
        P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n21175), .ZN(n21174) );
  OAI221_X1 U24091 ( .B1(n21176), .B2(keyinput122), .C1(n21175), .C2(
        P3_BYTEENABLE_REG_3__SCAN_IN), .A(n21174), .ZN(n21181) );
  INV_X1 U24092 ( .A(keyinput57), .ZN(n21178) );
  AOI22_X1 U24093 ( .A1(n21179), .A2(keyinput24), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n21178), .ZN(n21177) );
  OAI221_X1 U24094 ( .B1(n21179), .B2(keyinput24), .C1(n21178), .C2(
        P3_ADDRESS_REG_13__SCAN_IN), .A(n21177), .ZN(n21180) );
  NOR4_X1 U24095 ( .A1(n21183), .A2(n21182), .A3(n21181), .A4(n21180), .ZN(
        n21184) );
  NAND4_X1 U24096 ( .A1(n21187), .A2(n21186), .A3(n21185), .A4(n21184), .ZN(
        n21304) );
  AOI22_X1 U24097 ( .A1(n21190), .A2(keyinput61), .B1(n21189), .B2(keyinput84), 
        .ZN(n21188) );
  OAI221_X1 U24098 ( .B1(n21190), .B2(keyinput61), .C1(n21189), .C2(keyinput84), .A(n21188), .ZN(n21202) );
  INV_X1 U24099 ( .A(keyinput3), .ZN(n21192) );
  AOI22_X1 U24100 ( .A1(n14796), .A2(keyinput114), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n21192), .ZN(n21191) );
  OAI221_X1 U24101 ( .B1(n14796), .B2(keyinput114), .C1(n21192), .C2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .A(n21191), .ZN(n21201) );
  AOI22_X1 U24102 ( .A1(n21195), .A2(keyinput106), .B1(n21194), .B2(keyinput69), .ZN(n21193) );
  OAI221_X1 U24103 ( .B1(n21195), .B2(keyinput106), .C1(n21194), .C2(
        keyinput69), .A(n21193), .ZN(n21200) );
  AOI22_X1 U24104 ( .A1(n21198), .A2(keyinput67), .B1(n21197), .B2(keyinput54), 
        .ZN(n21196) );
  OAI221_X1 U24105 ( .B1(n21198), .B2(keyinput67), .C1(n21197), .C2(keyinput54), .A(n21196), .ZN(n21199) );
  NOR4_X1 U24106 ( .A1(n21202), .A2(n21201), .A3(n21200), .A4(n21199), .ZN(
        n21302) );
  INV_X1 U24107 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n21205) );
  AOI22_X1 U24108 ( .A1(n21205), .A2(keyinput9), .B1(n21204), .B2(keyinput89), 
        .ZN(n21203) );
  OAI221_X1 U24109 ( .B1(n21205), .B2(keyinput9), .C1(n21204), .C2(keyinput89), 
        .A(n21203), .ZN(n21216) );
  INV_X1 U24110 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n21208) );
  AOI22_X1 U24111 ( .A1(n21208), .A2(keyinput86), .B1(keyinput126), .B2(n21207), .ZN(n21206) );
  OAI221_X1 U24112 ( .B1(n21208), .B2(keyinput86), .C1(n21207), .C2(
        keyinput126), .A(n21206), .ZN(n21215) );
  AOI22_X1 U24113 ( .A1(n11722), .A2(keyinput112), .B1(keyinput115), .B2(
        n21210), .ZN(n21209) );
  OAI221_X1 U24114 ( .B1(n11722), .B2(keyinput112), .C1(n21210), .C2(
        keyinput115), .A(n21209), .ZN(n21214) );
  AOI22_X1 U24115 ( .A1(n12514), .A2(keyinput70), .B1(keyinput68), .B2(n21212), 
        .ZN(n21211) );
  OAI221_X1 U24116 ( .B1(n12514), .B2(keyinput70), .C1(n21212), .C2(keyinput68), .A(n21211), .ZN(n21213) );
  NOR4_X1 U24117 ( .A1(n21216), .A2(n21215), .A3(n21214), .A4(n21213), .ZN(
        n21301) );
  INV_X1 U24118 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n21218) );
  AOI22_X1 U24119 ( .A1(n21219), .A2(keyinput102), .B1(keyinput63), .B2(n21218), .ZN(n21217) );
  OAI221_X1 U24120 ( .B1(n21219), .B2(keyinput102), .C1(n21218), .C2(
        keyinput63), .A(n21217), .ZN(n21247) );
  INV_X1 U24121 ( .A(keyinput58), .ZN(n21221) );
  AOI22_X1 U24122 ( .A1(n11730), .A2(keyinput37), .B1(
        P1_DATAWIDTH_REG_9__SCAN_IN), .B2(n21221), .ZN(n21220) );
  OAI221_X1 U24123 ( .B1(n11730), .B2(keyinput37), .C1(n21221), .C2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A(n21220), .ZN(n21246) );
  XOR2_X1 U24124 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput62), .Z(n21226) );
  AOI22_X1 U24125 ( .A1(n21224), .A2(keyinput103), .B1(keyinput72), .B2(n21223), .ZN(n21222) );
  OAI221_X1 U24126 ( .B1(n21224), .B2(keyinput103), .C1(n21223), .C2(
        keyinput72), .A(n21222), .ZN(n21225) );
  AOI211_X1 U24127 ( .C1(n21228), .C2(keyinput99), .A(n21226), .B(n21225), 
        .ZN(n21227) );
  OAI21_X1 U24128 ( .B1(n21228), .B2(keyinput99), .A(n21227), .ZN(n21245) );
  OAI22_X1 U24129 ( .A1(n14771), .A2(keyinput97), .B1(n21230), .B2(keyinput15), 
        .ZN(n21229) );
  AOI221_X1 U24130 ( .B1(n14771), .B2(keyinput97), .C1(keyinput15), .C2(n21230), .A(n21229), .ZN(n21243) );
  INV_X1 U24131 ( .A(keyinput95), .ZN(n21232) );
  OAI22_X1 U24132 ( .A1(n21233), .A2(keyinput34), .B1(n21232), .B2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21231) );
  AOI221_X1 U24133 ( .B1(n21233), .B2(keyinput34), .C1(
        P2_DATAWIDTH_REG_13__SCAN_IN), .C2(n21232), .A(n21231), .ZN(n21242) );
  INV_X1 U24134 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n21235) );
  OAI22_X1 U24135 ( .A1(n21236), .A2(keyinput41), .B1(n21235), .B2(keyinput53), 
        .ZN(n21234) );
  AOI221_X1 U24136 ( .B1(n21236), .B2(keyinput41), .C1(keyinput53), .C2(n21235), .A(n21234), .ZN(n21241) );
  INV_X1 U24137 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21239) );
  OAI22_X1 U24138 ( .A1(n21239), .A2(keyinput118), .B1(n21238), .B2(keyinput30), .ZN(n21237) );
  AOI221_X1 U24139 ( .B1(n21239), .B2(keyinput118), .C1(keyinput30), .C2(
        n21238), .A(n21237), .ZN(n21240) );
  NAND4_X1 U24140 ( .A1(n21243), .A2(n21242), .A3(n21241), .A4(n21240), .ZN(
        n21244) );
  NOR4_X1 U24141 ( .A1(n21247), .A2(n21246), .A3(n21245), .A4(n21244), .ZN(
        n21300) );
  NAND2_X1 U24142 ( .A1(keyinput25), .A2(keyinput45), .ZN(n21248) );
  NOR3_X1 U24143 ( .A1(keyinput21), .A2(keyinput64), .A3(n21248), .ZN(n21249)
         );
  NAND3_X1 U24144 ( .A1(keyinput24), .A2(keyinput57), .A3(n21249), .ZN(n21262)
         );
  NAND2_X1 U24145 ( .A1(keyinput17), .A2(keyinput22), .ZN(n21250) );
  NOR3_X1 U24146 ( .A1(keyinput27), .A2(keyinput85), .A3(n21250), .ZN(n21260)
         );
  NOR4_X1 U24147 ( .A1(keyinput96), .A2(keyinput81), .A3(keyinput33), .A4(
        keyinput59), .ZN(n21259) );
  NAND4_X1 U24148 ( .A1(keyinput18), .A2(keyinput121), .A3(keyinput74), .A4(
        keyinput0), .ZN(n21257) );
  INV_X1 U24149 ( .A(keyinput73), .ZN(n21251) );
  NAND4_X1 U24150 ( .A1(keyinput77), .A2(keyinput36), .A3(keyinput92), .A4(
        n21251), .ZN(n21256) );
  NOR2_X1 U24151 ( .A1(keyinput44), .A2(keyinput109), .ZN(n21252) );
  NAND3_X1 U24152 ( .A1(keyinput107), .A2(keyinput5), .A3(n21252), .ZN(n21255)
         );
  INV_X1 U24153 ( .A(keyinput4), .ZN(n21253) );
  NAND4_X1 U24154 ( .A1(keyinput91), .A2(keyinput105), .A3(keyinput40), .A4(
        n21253), .ZN(n21254) );
  NOR4_X1 U24155 ( .A1(n21257), .A2(n21256), .A3(n21255), .A4(n21254), .ZN(
        n21258) );
  NAND3_X1 U24156 ( .A1(n21260), .A2(n21259), .A3(n21258), .ZN(n21261) );
  NOR4_X1 U24157 ( .A1(keyinput122), .A2(keyinput48), .A3(n21262), .A4(n21261), 
        .ZN(n21298) );
  NAND4_X1 U24158 ( .A1(keyinput9), .A2(keyinput12), .A3(keyinput56), .A4(
        keyinput68), .ZN(n21266) );
  NAND4_X1 U24159 ( .A1(keyinput19), .A2(keyinput7), .A3(keyinput10), .A4(
        keyinput49), .ZN(n21265) );
  NAND4_X1 U24160 ( .A1(keyinput89), .A2(keyinput116), .A3(keyinput84), .A4(
        keyinput80), .ZN(n21264) );
  NAND4_X1 U24161 ( .A1(keyinput52), .A2(keyinput113), .A3(keyinput93), .A4(
        keyinput69), .ZN(n21263) );
  NOR4_X1 U24162 ( .A1(n21266), .A2(n21265), .A3(n21264), .A4(n21263), .ZN(
        n21297) );
  NAND4_X1 U24163 ( .A1(keyinput83), .A2(keyinput82), .A3(keyinput79), .A4(
        keyinput78), .ZN(n21270) );
  NAND4_X1 U24164 ( .A1(keyinput127), .A2(keyinput115), .A3(keyinput126), .A4(
        keyinput99), .ZN(n21269) );
  NAND4_X1 U24165 ( .A1(keyinput38), .A2(keyinput23), .A3(keyinput26), .A4(
        keyinput15), .ZN(n21268) );
  NAND4_X1 U24166 ( .A1(keyinput67), .A2(keyinput54), .A3(keyinput46), .A4(
        keyinput34), .ZN(n21267) );
  NOR4_X1 U24167 ( .A1(n21270), .A2(n21269), .A3(n21268), .A4(n21267), .ZN(
        n21296) );
  NAND2_X1 U24168 ( .A1(keyinput120), .A2(keyinput90), .ZN(n21271) );
  NOR3_X1 U24169 ( .A1(keyinput42), .A2(keyinput66), .A3(n21271), .ZN(n21275)
         );
  NOR4_X1 U24170 ( .A1(keyinput50), .A2(keyinput13), .A3(keyinput39), .A4(
        keyinput28), .ZN(n21274) );
  NOR4_X1 U24171 ( .A1(keyinput125), .A2(keyinput8), .A3(keyinput88), .A4(
        keyinput14), .ZN(n21273) );
  AND4_X1 U24172 ( .A1(keyinput6), .A2(keyinput43), .A3(keyinput51), .A4(
        keyinput117), .ZN(n21272) );
  NAND4_X1 U24173 ( .A1(n21275), .A2(n21274), .A3(n21273), .A4(n21272), .ZN(
        n21294) );
  INV_X1 U24174 ( .A(keyinput1), .ZN(n21276) );
  NOR4_X1 U24175 ( .A1(keyinput76), .A2(keyinput98), .A3(keyinput111), .A4(
        n21276), .ZN(n21282) );
  AND4_X1 U24176 ( .A1(keyinput60), .A2(keyinput75), .A3(keyinput20), .A4(
        keyinput29), .ZN(n21281) );
  INV_X1 U24177 ( .A(keyinput55), .ZN(n21277) );
  NOR4_X1 U24178 ( .A1(keyinput94), .A2(keyinput32), .A3(keyinput35), .A4(
        n21277), .ZN(n21280) );
  NAND2_X1 U24179 ( .A1(keyinput2), .A2(keyinput100), .ZN(n21278) );
  NOR3_X1 U24180 ( .A1(keyinput47), .A2(keyinput119), .A3(n21278), .ZN(n21279)
         );
  NAND4_X1 U24181 ( .A1(n21282), .A2(n21281), .A3(n21280), .A4(n21279), .ZN(
        n21293) );
  NOR4_X1 U24182 ( .A1(keyinput37), .A2(keyinput61), .A3(keyinput53), .A4(
        keyinput16), .ZN(n21286) );
  NOR4_X1 U24183 ( .A1(keyinput30), .A2(keyinput31), .A3(keyinput11), .A4(
        keyinput41), .ZN(n21285) );
  NOR4_X1 U24184 ( .A1(keyinput104), .A2(keyinput112), .A3(keyinput72), .A4(
        keyinput108), .ZN(n21284) );
  NOR4_X1 U24185 ( .A1(keyinput101), .A2(keyinput97), .A3(keyinput65), .A4(
        keyinput124), .ZN(n21283) );
  NAND4_X1 U24186 ( .A1(n21286), .A2(n21285), .A3(n21284), .A4(n21283), .ZN(
        n21292) );
  NOR4_X1 U24187 ( .A1(keyinput110), .A2(keyinput106), .A3(keyinput102), .A4(
        keyinput103), .ZN(n21290) );
  NOR4_X1 U24188 ( .A1(keyinput3), .A2(keyinput123), .A3(keyinput118), .A4(
        keyinput114), .ZN(n21289) );
  NOR4_X1 U24189 ( .A1(keyinput71), .A2(keyinput62), .A3(keyinput63), .A4(
        keyinput58), .ZN(n21288) );
  NOR4_X1 U24190 ( .A1(keyinput95), .A2(keyinput86), .A3(keyinput87), .A4(
        keyinput70), .ZN(n21287) );
  NAND4_X1 U24191 ( .A1(n21290), .A2(n21289), .A3(n21288), .A4(n21287), .ZN(
        n21291) );
  NOR4_X1 U24192 ( .A1(n21294), .A2(n21293), .A3(n21292), .A4(n21291), .ZN(
        n21295) );
  NAND4_X1 U24193 ( .A1(n21298), .A2(n21297), .A3(n21296), .A4(n21295), .ZN(
        n21299) );
  NAND4_X1 U24194 ( .A1(n21302), .A2(n21301), .A3(n21300), .A4(n21299), .ZN(
        n21303) );
  NOR4_X1 U24195 ( .A1(n21306), .A2(n21305), .A3(n21304), .A4(n21303), .ZN(
        n21307) );
  XNOR2_X1 U24196 ( .A(n21308), .B(n21307), .ZN(P3_U2863) );
  NOR2_X2 U12205 ( .A1(n16734), .A2(n17660), .ZN(n16733) );
  NOR2_X2 U16705 ( .A1(n17699), .A2(n16763), .ZN(n16762) );
  NOR2_X2 U12219 ( .A1(n13419), .A2(n17653), .ZN(n13420) );
  NOR2_X2 U19899 ( .A1(n16695), .A2(n16696), .ZN(n16694) );
  XNOR2_X2 U11300 ( .A(n12696), .B(n12697), .ZN(n20182) );
  NAND2_X1 U11484 ( .A1(n9998), .A2(n11836), .ZN(n11923) );
  NAND2_X1 U11620 ( .A1(n13952), .A2(n12713), .ZN(n20173) );
  OR2_X2 U11327 ( .A1(n11965), .A2(n11964), .ZN(n11966) );
  OR2_X4 U11518 ( .A1(n11818), .A2(n11817), .ZN(n20272) );
  AND2_X4 U11550 ( .A1(n11705), .A2(n10161), .ZN(n11955) );
  AND2_X4 U11649 ( .A1(n14593), .A2(n14742), .ZN(n14578) );
  NOR2_X4 U11650 ( .A1(n14591), .A2(n14594), .ZN(n14593) );
  AND2_X2 U11320 ( .A1(n14522), .A2(n14703), .ZN(n14506) );
  OR2_X2 U11369 ( .A1(n14790), .A2(n20258), .ZN(n13049) );
  OR2_X4 U11281 ( .A1(n11802), .A2(n11801), .ZN(n20261) );
  AND2_X2 U11822 ( .A1(n12677), .A2(n12676), .ZN(n13646) );
  NAND2_X2 U11520 ( .A1(n9824), .A2(n9820), .ZN(n11826) );
  NAND2_X2 U15003 ( .A1(n11943), .A2(n20321), .ZN(n14677) );
  NOR2_X2 U11561 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11693), .ZN(
        n11706) );
  AND2_X2 U11569 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13621) );
  AND2_X2 U11563 ( .A1(n11693), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10161) );
  INV_X2 U12745 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10119) );
  INV_X2 U14780 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12011) );
  AND2_X2 U11547 ( .A1(n10161), .A2(n11708), .ZN(n11812) );
  INV_X1 U11562 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13655) );
  AND2_X1 U12832 ( .A1(n11704), .A2(n11707), .ZN(n10222) );
  AND2_X1 U11523 ( .A1(n11765), .A2(n11763), .ZN(n10124) );
  AND4_X1 U11526 ( .A1(n11733), .A2(n11736), .A3(n11734), .A4(n11738), .ZN(
        n9824) );
  OR2_X1 U14830 ( .A1(n11753), .A2(n11752), .ZN(n11823) );
  INV_X2 U11233 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11534) );
  CLKBUF_X1 U14984 ( .A(n11955), .Z(n12577) );
  AND2_X1 U11218 ( .A1(n10373), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10664) );
  NAND2_X1 U11210 ( .A1(n12759), .A2(n11992), .ZN(n12640) );
  NOR2_X1 U11715 ( .A1(n10160), .A2(n13829), .ZN(n12037) );
  AND2_X1 U14035 ( .A1(n11059), .A2(n11063), .ZN(n11122) );
  CLKBUF_X2 U11200 ( .A(n20252), .Z(n9752) );
  AND2_X1 U11692 ( .A1(n12841), .A2(n14132), .ZN(n12963) );
  NOR2_X1 U11328 ( .A1(n20226), .A2(n14277), .ZN(n13801) );
  AND2_X1 U14782 ( .A1(n11704), .A2(n11706), .ZN(n11853) );
  AND2_X1 U12761 ( .A1(n11704), .A2(n10161), .ZN(n11860) );
  AND4_X1 U11296 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n9799) );
  CLKBUF_X2 U11229 ( .A(n11946), .Z(n12580) );
  CLKBUF_X2 U14951 ( .A(n11896), .Z(n12490) );
  OR2_X1 U11197 ( .A1(n12648), .A2(n11824), .ZN(n12667) );
  OR2_X1 U11221 ( .A1(n11912), .A2(n11911), .ZN(n11929) );
  CLKBUF_X2 U11228 ( .A(n11847), .Z(n12582) );
  CLKBUF_X2 U11248 ( .A(n11812), .Z(n12595) );
  CLKBUF_X2 U11249 ( .A(n11862), .Z(n12581) );
  CLKBUF_X2 U11259 ( .A(n12001), .Z(n11901) );
  NAND2_X1 U11277 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11694) );
  NOR2_X2 U11292 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11709) );
  INV_X1 U11340 ( .A(n12064), .ZN(n12062) );
  INV_X2 U11351 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11693) );
  OAI22_X1 U11354 ( .A1(n13654), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12706), 
        .B2(n12759), .ZN(n9999) );
  AND2_X1 U11358 ( .A1(n11708), .A2(n11707), .ZN(n11861) );
  INV_X1 U11361 ( .A(n20261), .ZN(n14197) );
  BUF_X1 U11366 ( .A(n9812), .Z(n12624) );
  NOR2_X1 U11383 ( .A1(n16121), .A2(n12765), .ZN(n12767) );
  AND2_X1 U11413 ( .A1(n11819), .A2(n9803), .ZN(n11825) );
  AND3_X1 U11458 ( .A1(n11755), .A2(n11756), .A3(n11764), .ZN(n10123) );
  CLKBUF_X1 U11504 ( .A(n10464), .Z(n10556) );
  INV_X1 U11533 ( .A(n11821), .ZN(n11767) );
  CLKBUF_X1 U11544 ( .A(n14887), .Z(n9779) );
  NAND2_X1 U11570 ( .A1(n11824), .A2(n20261), .ZN(n20982) );
  OAI21_X1 U11571 ( .B1(n14988), .B2(n14997), .A(n14998), .ZN(n14993) );
  NOR2_X1 U11577 ( .A1(n14708), .A2(n14515), .ZN(n9906) );
  AOI21_X1 U11599 ( .B1(n16263), .B2(n16194), .A(n16191), .ZN(n16185) );
  CLKBUF_X1 U11610 ( .A(n14929), .Z(n16133) );
  NOR2_X1 U11617 ( .A1(n15999), .A2(n12961), .ZN(n20239) );
  CLKBUF_X1 U11622 ( .A(n11830), .Z(n15030) );
  CLKBUF_X1 U11633 ( .A(n15680), .Z(n15681) );
  NOR2_X1 U11642 ( .A1(n17614), .A2(n16714), .ZN(n16713) );
  OR2_X1 U11654 ( .A1(n9913), .A2(n9912), .ZN(n9911) );
  NOR2_X1 U11792 ( .A1(n13412), .A2(n9927), .ZN(n17638) );
  OR2_X1 U11954 ( .A1(n9915), .A2(n9914), .ZN(n17749) );
  NOR2_X1 U11989 ( .A1(n17832), .A2(n17896), .ZN(n17863) );
  NOR2_X2 U12095 ( .A1(n20272), .A2(n20261), .ZN(n13480) );
  CLKBUF_X1 U12203 ( .A(n14911), .Z(n14920) );
  OR2_X1 U12208 ( .A1(n14281), .A2(n14280), .ZN(n16179) );
  CLKBUF_X1 U12225 ( .A(n19280), .Z(n20002) );
  INV_X2 U12259 ( .A(n19990), .ZN(n10625) );
  XNOR2_X1 U12327 ( .A(n14344), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14357) );
  NAND2_X1 U12386 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17922) );
  AND2_X1 U12413 ( .A1(n13049), .A2(n13048), .ZN(n13050) );
  INV_X1 U12673 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13684) );
  CLKBUF_X1 U12683 ( .A(n19279), .Z(n19271) );
endmodule

