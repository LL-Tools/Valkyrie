

module b14_C_AntiSAT_k_128_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758;

  CLKBUF_X2 U2289 ( .A(n2477), .Z(n3629) );
  NAND3_X2 U2290 ( .A1(n2198), .A2(n4360), .A3(n2197), .ZN(n2864) );
  INV_X1 U2291 ( .A(n2782), .ZN(n2797) );
  AND2_X1 U2292 ( .A1(n2885), .A2(n2336), .ZN(n2467) );
  XNOR2_X2 U2293 ( .A(n2334), .B(IR_REG_30__SCAN_IN), .ZN(n2885) );
  NAND2_X2 U2294 ( .A1(n2882), .A2(IR_REG_31__SCAN_IN), .ZN(n2334) );
  NAND2_X2 U2295 ( .A1(n2440), .A2(n2439), .ZN(n2447) );
  XNOR2_X2 U2296 ( .A(n3395), .B(n3421), .ZN(n3445) );
  AOI22_X2 U2297 ( .A1(n3865), .A2(n3872), .B1(n3868), .B2(n3895), .ZN(n3395)
         );
  AND2_X1 U2298 ( .A1(n2271), .A2(n3308), .ZN(n2268) );
  NAND4_X1 U2299 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n3770)
         );
  NAND4_X2 U2300 ( .A1(n2408), .A2(n2409), .A3(n2407), .A4(n2410), .ZN(n3773)
         );
  CLKBUF_X2 U2301 ( .A(n2406), .Z(n2134) );
  XNOR2_X1 U2302 ( .A(n2331), .B(IR_REG_29__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U2303 ( .A1(n2152), .A2(n2151), .ZN(n2579) );
  MUX2_X1 U2304 ( .A(n4214), .B(n4292), .S(n4568), .Z(n4215) );
  MUX2_X1 U2305 ( .A(n4293), .B(n4292), .S(n4756), .Z(n4294) );
  NAND2_X1 U2306 ( .A1(n3391), .A2(n3390), .ZN(n3882) );
  AOI21_X1 U2307 ( .B1(n3501), .B2(n2221), .A(n2224), .ZN(n2220) );
  NAND2_X1 U2308 ( .A1(n3551), .A2(n3552), .ZN(n3550) );
  OAI22_X1 U2309 ( .A1(n3472), .A2(n3471), .B1(n2688), .B2(n2687), .ZN(n3551)
         );
  NAND2_X1 U2310 ( .A1(n3842), .A2(n3843), .ZN(n3854) );
  INV_X1 U2311 ( .A(n2189), .ZN(n3583) );
  NAND2_X1 U2312 ( .A1(n4135), .A2(n2295), .ZN(n4116) );
  NAND2_X1 U2313 ( .A1(n4137), .A2(n4136), .ZN(n4135) );
  AND2_X1 U2314 ( .A1(n2212), .A2(n2211), .ZN(n4458) );
  NOR2_X1 U2315 ( .A1(n3378), .A2(n2296), .ZN(n4137) );
  OAI21_X1 U2316 ( .B1(n2641), .B2(n2187), .A(n2185), .ZN(n2188) );
  NAND2_X1 U2317 ( .A1(n4426), .A2(n3836), .ZN(n4436) );
  AOI21_X1 U2318 ( .B1(n2264), .B2(n2265), .A(n2070), .ZN(n2261) );
  NAND2_X1 U2319 ( .A1(n3030), .A2(n3072), .ZN(n3142) );
  AND2_X1 U2320 ( .A1(n3653), .A2(n3656), .ZN(n3027) );
  NOR2_X2 U2321 ( .A1(n2932), .A2(n2931), .ZN(n4457) );
  NAND2_X2 U2322 ( .A1(n2474), .A2(n2473), .ZN(n3771) );
  NOR2_X1 U2323 ( .A1(n3003), .A2(n3002), .ZN(n4496) );
  INV_X4 U2324 ( .A(n2848), .ZN(n3424) );
  AND2_X1 U2325 ( .A1(n2333), .A2(n2336), .ZN(n2454) );
  NAND2_X2 U2326 ( .A1(n3035), .A2(n2837), .ZN(n2782) );
  MUX2_X1 U2327 ( .A(IR_REG_31__SCAN_IN), .B(n2349), .S(IR_REG_25__SCAN_IN), 
        .Z(n2351) );
  NAND2_X1 U2328 ( .A1(n2821), .A2(IR_REG_31__SCAN_IN), .ZN(n2120) );
  XNOR2_X1 U2329 ( .A(n2354), .B(IR_REG_26__SCAN_IN), .ZN(n4360) );
  INV_X1 U2330 ( .A(n2579), .ZN(n2125) );
  AND3_X1 U2331 ( .A1(n2318), .A2(n2316), .A3(n2317), .ZN(n2319) );
  AND2_X1 U2332 ( .A1(n2106), .A2(n2105), .ZN(n2104) );
  INV_X1 U2333 ( .A(IR_REG_14__SCAN_IN), .ZN(n4595) );
  INV_X1 U2334 ( .A(IR_REG_9__SCAN_IN), .ZN(n2151) );
  INV_X1 U2335 ( .A(n2567), .ZN(n2152) );
  XNOR2_X1 U2336 ( .A(n2917), .B(n4390), .ZN(n4382) );
  NAND2_X1 U2337 ( .A1(n3530), .A2(n2441), .ZN(n2744) );
  NOR2_X1 U2338 ( .A1(n2237), .A2(n2717), .ZN(n2236) );
  INV_X1 U2339 ( .A(n3554), .ZN(n2237) );
  INV_X1 U2340 ( .A(IR_REG_30__SCAN_IN), .ZN(n2329) );
  NOR2_X1 U2341 ( .A1(n4458), .A2(n2210), .ZN(n3840) );
  AND2_X1 U2342 ( .A1(n3839), .A2(REG2_REG_15__SCAN_IN), .ZN(n2210) );
  NAND2_X1 U2343 ( .A1(n2374), .A2(n3652), .ZN(n3035) );
  NAND2_X1 U2344 ( .A1(n2288), .A2(n3389), .ZN(n2287) );
  NAND2_X1 U2345 ( .A1(n2293), .A2(n2289), .ZN(n2288) );
  NOR2_X1 U2346 ( .A1(n2290), .A2(n2283), .ZN(n2282) );
  INV_X1 U2347 ( .A(n3386), .ZN(n2283) );
  INV_X1 U2348 ( .A(n2293), .ZN(n2290) );
  NAND2_X1 U2349 ( .A1(n2308), .A2(n2307), .ZN(n2306) );
  INV_X1 U2350 ( .A(IR_REG_25__SCAN_IN), .ZN(n2307) );
  INV_X1 U2351 ( .A(IR_REG_20__SCAN_IN), .ZN(n2345) );
  INV_X1 U2352 ( .A(IR_REG_17__SCAN_IN), .ZN(n2357) );
  NOR2_X1 U2353 ( .A1(n2343), .A2(IR_REG_13__SCAN_IN), .ZN(n2249) );
  INV_X1 U2354 ( .A(n2626), .ZN(n2342) );
  NAND2_X1 U2355 ( .A1(n2125), .A2(n2302), .ZN(n2626) );
  OR2_X1 U2356 ( .A1(n2879), .A2(IR_REG_27__SCAN_IN), .ZN(n2200) );
  NAND2_X1 U2357 ( .A1(n2879), .A2(IR_REG_28__SCAN_IN), .ZN(n2199) );
  OR2_X1 U2358 ( .A1(n2484), .A2(n2119), .ZN(n2117) );
  INV_X1 U2359 ( .A(n2454), .ZN(n2848) );
  NAND2_X1 U2360 ( .A1(n2180), .A2(n3791), .ZN(n3792) );
  NAND2_X1 U2361 ( .A1(n2170), .A2(n2080), .ZN(n2169) );
  INV_X1 U2362 ( .A(n2971), .ZN(n2170) );
  AND3_X1 U2363 ( .A1(n2174), .A2(n2097), .A3(n2175), .ZN(n3817) );
  AND2_X1 U2364 ( .A1(n2376), .A2(n2375), .ZN(n3085) );
  OAI21_X1 U2365 ( .B1(n3000), .B2(D_REG_0__SCAN_IN), .A(n2888), .ZN(n3031) );
  NAND2_X1 U2366 ( .A1(n3866), .A2(n3705), .ZN(n4196) );
  AND2_X1 U2367 ( .A1(n2064), .A2(n3387), .ZN(n2291) );
  AND2_X1 U2368 ( .A1(n3996), .A2(n3975), .ZN(n3960) );
  AOI21_X1 U2369 ( .B1(n4116), .B2(n3379), .A(n2312), .ZN(n4101) );
  NAND2_X1 U2370 ( .A1(n2374), .A2(n3085), .ZN(n4530) );
  NOR2_X1 U2371 ( .A1(n2323), .A2(n2299), .ZN(n2298) );
  NAND2_X1 U2372 ( .A1(n2302), .A2(n2324), .ZN(n2299) );
  NAND2_X1 U2373 ( .A1(n3525), .A2(n2194), .ZN(n3501) );
  NAND2_X1 U2374 ( .A1(n2124), .A2(n2123), .ZN(n2194) );
  INV_X1 U2375 ( .A(n3528), .ZN(n2123) );
  NAND2_X1 U2376 ( .A1(n3935), .A2(n2682), .ZN(n2766) );
  INV_X1 U2377 ( .A(n3590), .ZN(n2229) );
  AOI21_X1 U2378 ( .B1(n3837), .B2(REG1_REG_13__SCAN_IN), .A(n4430), .ZN(n3816) );
  INV_X1 U2379 ( .A(n2291), .ZN(n2289) );
  NOR2_X1 U2380 ( .A1(n2157), .A2(n4123), .ZN(n2156) );
  INV_X1 U2381 ( .A(n3686), .ZN(n2157) );
  INV_X1 U2382 ( .A(n3617), .ZN(n2271) );
  NAND2_X1 U2383 ( .A1(n3767), .A2(n3466), .ZN(n2272) );
  NAND2_X1 U2384 ( .A1(n3106), .A2(n3544), .ZN(n3659) );
  NAND2_X1 U2385 ( .A1(n3771), .A2(n3117), .ZN(n3661) );
  NAND2_X1 U2386 ( .A1(n3025), .A2(n3043), .ZN(n3653) );
  NOR2_X1 U2387 ( .A1(n4177), .A2(n4148), .ZN(n4117) );
  NOR2_X1 U2388 ( .A1(n2306), .A2(IR_REG_22__SCAN_IN), .ZN(n2208) );
  AND2_X1 U2389 ( .A1(n2322), .A2(n2303), .ZN(n2302) );
  INV_X1 U2390 ( .A(IR_REG_10__SCAN_IN), .ZN(n2303) );
  NOR2_X1 U2391 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2322)
         );
  NOR2_X1 U2392 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2310)
         );
  INV_X1 U2393 ( .A(IR_REG_2__SCAN_IN), .ZN(n2318) );
  INV_X1 U2394 ( .A(IR_REG_1__SCAN_IN), .ZN(n2317) );
  NOR2_X1 U2395 ( .A1(n2634), .A2(n2245), .ZN(n2244) );
  INV_X1 U2396 ( .A(n3274), .ZN(n2245) );
  INV_X1 U2397 ( .A(n2233), .ZN(n2232) );
  NOR2_X1 U2398 ( .A1(n2239), .A2(n2069), .ZN(n2230) );
  XNOR2_X1 U2399 ( .A(n2466), .B(n2782), .ZN(n2481) );
  NAND2_X1 U2400 ( .A1(n2229), .A2(n2226), .ZN(n2225) );
  NAND2_X1 U2401 ( .A1(n3589), .A2(n2227), .ZN(n2226) );
  NAND2_X1 U2402 ( .A1(n2229), .A2(n3498), .ZN(n2228) );
  INV_X1 U2403 ( .A(n2225), .ZN(n2224) );
  INV_X1 U2404 ( .A(n3256), .ZN(n3248) );
  NAND2_X1 U2405 ( .A1(n2238), .A2(n2195), .ZN(n2124) );
  NOR2_X1 U2406 ( .A1(n2748), .A2(n2747), .ZN(n2195) );
  AOI22_X1 U2407 ( .A1(n3773), .A2(n2785), .B1(n2682), .B2(n3483), .ZN(n2430)
         );
  NAND2_X1 U2408 ( .A1(n2414), .A2(n2413), .ZN(n2415) );
  NAND2_X1 U2409 ( .A1(n2355), .A2(n2864), .ZN(n2840) );
  AND2_X1 U2410 ( .A1(n2795), .A2(n2794), .ZN(n3394) );
  OR2_X1 U2411 ( .A1(n3869), .A2(n2790), .ZN(n2795) );
  OR2_X1 U2412 ( .A1(n4104), .A2(n2790), .ZN(n2382) );
  INV_X1 U2413 ( .A(n3545), .ZN(n2135) );
  NAND2_X1 U2414 ( .A1(n2468), .A2(n2059), .ZN(n2469) );
  AND2_X1 U2415 ( .A1(n2333), .A2(n2332), .ZN(n2455) );
  XNOR2_X1 U2416 ( .A(n4365), .B(n3047), .ZN(n3788) );
  NAND2_X1 U2417 ( .A1(n3792), .A2(n2912), .ZN(n2913) );
  AND2_X1 U2418 ( .A1(n2218), .A2(n2217), .ZN(n2949) );
  NAND2_X1 U2419 ( .A1(n2929), .A2(REG2_REG_5__SCAN_IN), .ZN(n2217) );
  XNOR2_X1 U2420 ( .A(n3810), .B(n3828), .ZN(n2966) );
  NAND2_X1 U2421 ( .A1(n3809), .A2(n2171), .ZN(n3811) );
  OR2_X1 U2422 ( .A1(n3810), .A2(n3828), .ZN(n2171) );
  NAND2_X1 U2423 ( .A1(n2099), .A2(n2066), .ZN(n2212) );
  OR2_X1 U2424 ( .A1(n4441), .A2(n2176), .ZN(n2174) );
  OR2_X1 U2425 ( .A1(n4454), .A2(n4442), .ZN(n2176) );
  OR2_X1 U2426 ( .A1(n2056), .A2(n4454), .ZN(n2175) );
  OR2_X1 U2427 ( .A1(n4441), .A2(n4442), .ZN(n2177) );
  NAND2_X1 U2428 ( .A1(n3854), .A2(n2095), .ZN(n4484) );
  NAND2_X1 U2429 ( .A1(n3849), .A2(n2094), .ZN(n4477) );
  NOR2_X1 U2430 ( .A1(n4484), .A2(n4485), .ZN(n4483) );
  AOI21_X1 U2431 ( .B1(n3871), .B2(n3711), .A(n3710), .ZN(n3422) );
  NOR2_X1 U2432 ( .A1(n2057), .A2(n2289), .ZN(n2286) );
  AND2_X1 U2433 ( .A1(n3388), .A2(n2063), .ZN(n2293) );
  AOI21_X1 U2434 ( .B1(n4083), .B2(n3383), .A(n3382), .ZN(n4063) );
  AND2_X1 U2435 ( .A1(n4111), .A2(n4090), .ZN(n3382) );
  AND2_X1 U2436 ( .A1(n4142), .A2(n4165), .ZN(n2296) );
  NAND2_X1 U2437 ( .A1(n3246), .A2(n3241), .ZN(n2297) );
  NAND2_X1 U2438 ( .A1(n2275), .A2(n2274), .ZN(n2273) );
  NAND2_X1 U2439 ( .A1(n3150), .A2(n2048), .ZN(n2276) );
  AND2_X1 U2440 ( .A1(n3228), .A2(n3667), .ZN(n3665) );
  INV_X1 U2441 ( .A(n3197), .ZN(n3191) );
  INV_X1 U2442 ( .A(n4169), .ZN(n4143) );
  OR2_X1 U2443 ( .A1(n4531), .A2(n3652), .ZN(n3003) );
  AND2_X1 U2444 ( .A1(n3960), .A2(n2092), .ZN(n3885) );
  AND2_X1 U2445 ( .A1(n3885), .A2(n3876), .ZN(n3866) );
  NAND2_X1 U2446 ( .A1(n2281), .A2(n2068), .ZN(n3391) );
  AND2_X1 U2447 ( .A1(n3960), .A2(n3951), .ZN(n3953) );
  AND2_X1 U2448 ( .A1(n4367), .A2(n2988), .ZN(n4166) );
  NAND2_X1 U2449 ( .A1(n3749), .A2(n2991), .ZN(n4172) );
  OR2_X1 U2450 ( .A1(n4367), .A2(n2987), .ZN(n4169) );
  OR2_X1 U2451 ( .A1(n3090), .A2(n3756), .ZN(n4531) );
  NAND2_X1 U2452 ( .A1(n2803), .A2(n4360), .ZN(n3000) );
  NAND2_X1 U2453 ( .A1(n2305), .A2(n2326), .ZN(n2304) );
  INV_X1 U2454 ( .A(n2306), .ZN(n2305) );
  AND2_X1 U2455 ( .A1(n2370), .A2(n2208), .ZN(n2362) );
  NAND2_X1 U2456 ( .A1(n2821), .A2(n2820), .ZN(n2922) );
  NAND2_X1 U2457 ( .A1(n2309), .A2(n2058), .ZN(n2323) );
  AND4_X1 U2458 ( .A1(n2368), .A2(n2386), .A3(n2248), .A4(n2387), .ZN(n2309)
         );
  INV_X1 U2459 ( .A(n2302), .ZN(n2300) );
  INV_X1 U2460 ( .A(IR_REG_19__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U2461 ( .A1(n2247), .A2(IR_REG_31__SCAN_IN), .ZN(n2369) );
  AND2_X1 U2462 ( .A1(n2402), .A2(n2401), .ZN(n3839) );
  INV_X1 U2463 ( .A(IR_REG_7__SCAN_IN), .ZN(n2548) );
  OR2_X1 U2464 ( .A1(n2525), .A2(n2259), .ZN(n2549) );
  INV_X1 U2465 ( .A(IR_REG_6__SCAN_IN), .ZN(n2523) );
  INV_X1 U2466 ( .A(IR_REG_3__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U2467 ( .A1(n2317), .A2(n2259), .ZN(n2258) );
  OAI21_X1 U2468 ( .B1(n3501), .B2(n2224), .A(n2222), .ZN(n2860) );
  AND2_X1 U2469 ( .A1(n3446), .A2(n2223), .ZN(n2222) );
  NAND2_X1 U2470 ( .A1(n2228), .A2(n2225), .ZN(n2223) );
  OAI21_X1 U2471 ( .B1(n2477), .B2(n3778), .A(n2412), .ZN(n3483) );
  NAND2_X1 U2472 ( .A1(n2477), .A2(DATAI_1_), .ZN(n2412) );
  NAND2_X1 U2473 ( .A1(n2126), .A2(n2191), .ZN(n3519) );
  NAND2_X1 U2474 ( .A1(n2193), .A2(n2192), .ZN(n2191) );
  OAI211_X1 U2475 ( .C1(n3598), .C2(n3599), .A(n3510), .B(n3596), .ZN(n2126)
         );
  INV_X1 U2476 ( .A(n2661), .ZN(n2192) );
  NAND2_X1 U2477 ( .A1(n2559), .A2(n2558), .ZN(n3265) );
  OAI21_X1 U2478 ( .B1(n2116), .B2(n2088), .A(n2108), .ZN(n2107) );
  NAND2_X1 U2479 ( .A1(n3501), .A2(n2065), .ZN(n2110) );
  OR2_X1 U2480 ( .A1(n3501), .A2(n2112), .ZN(n2111) );
  INV_X1 U2481 ( .A(n3577), .ZN(n3609) );
  OAI211_X1 U2482 ( .C1(n3502), .C2(n2790), .A(n2752), .B(n2751), .ZN(n3946)
         );
  OAI211_X1 U2483 ( .C1(n3949), .C2(n2790), .A(n2743), .B(n2742), .ZN(n3973)
         );
  NAND4_X1 U2484 ( .A1(n2733), .A2(n2732), .A3(n2731), .A4(n2730), .ZN(n3987)
         );
  OAI22_X1 U2485 ( .A1(n4382), .A2(n2252), .B1(n2918), .B2(n2251), .ZN(n2971)
         );
  NAND2_X1 U2486 ( .A1(n2919), .A2(REG1_REG_4__SCAN_IN), .ZN(n2252) );
  INV_X1 U2487 ( .A(n2919), .ZN(n2251) );
  XOR2_X1 U2488 ( .A(n4363), .B(n2949), .Z(n2950) );
  XNOR2_X1 U2489 ( .A(n3827), .B(n3828), .ZN(n3826) );
  NAND2_X1 U2490 ( .A1(n2102), .A2(n2100), .ZN(n4399) );
  NAND2_X1 U2491 ( .A1(n3827), .A2(n2101), .ZN(n2100) );
  NAND2_X1 U2492 ( .A1(n3826), .A2(REG2_REG_8__SCAN_IN), .ZN(n2102) );
  INV_X1 U2493 ( .A(n3828), .ZN(n2101) );
  XNOR2_X1 U2494 ( .A(n3831), .B(n4520), .ZN(n4409) );
  NAND2_X1 U2495 ( .A1(n4409), .A2(REG2_REG_10__SCAN_IN), .ZN(n4408) );
  OR2_X1 U2496 ( .A1(n4380), .A2(n3799), .ZN(n4490) );
  INV_X1 U2497 ( .A(n4443), .ZN(n4487) );
  OR2_X1 U2498 ( .A1(n2773), .A2(n2760), .ZN(n3912) );
  AND2_X1 U2499 ( .A1(n4066), .A2(n2093), .ZN(n3996) );
  NAND2_X1 U2500 ( .A1(n2166), .A2(n2084), .ZN(n3436) );
  INV_X1 U2501 ( .A(n3442), .ZN(n2166) );
  NAND2_X1 U2502 ( .A1(n3987), .A2(n2441), .ZN(n2735) );
  INV_X1 U2503 ( .A(n2236), .ZN(n2231) );
  NAND2_X1 U2504 ( .A1(n2241), .A2(n2240), .ZN(n2239) );
  INV_X1 U2505 ( .A(n3455), .ZN(n2240) );
  INV_X1 U2506 ( .A(n3454), .ZN(n2241) );
  NAND2_X1 U2507 ( .A1(n3946), .A2(n2682), .ZN(n2754) );
  NAND2_X1 U2508 ( .A1(n4091), .A2(n2682), .ZN(n2672) );
  NAND2_X1 U2509 ( .A1(n3159), .A2(n2682), .ZN(n2512) );
  INV_X1 U2510 ( .A(n2186), .ZN(n2185) );
  OAI21_X1 U2511 ( .B1(n2640), .B2(n2187), .A(n3337), .ZN(n2186) );
  NAND2_X1 U2512 ( .A1(n2963), .A2(n2962), .ZN(n2965) );
  NAND2_X1 U2513 ( .A1(n3420), .A2(n3706), .ZN(n3890) );
  NAND2_X1 U2514 ( .A1(n2129), .A2(n2127), .ZN(n3929) );
  AOI21_X1 U2515 ( .B1(n2130), .B2(n3732), .A(n2128), .ZN(n2127) );
  NOR2_X1 U2516 ( .A1(n2133), .A2(n2131), .ZN(n2130) );
  AND2_X1 U2517 ( .A1(n3410), .A2(n2132), .ZN(n2131) );
  INV_X1 U2518 ( .A(n3731), .ZN(n2133) );
  NAND2_X1 U2519 ( .A1(n4134), .A2(n3406), .ZN(n2158) );
  AOI21_X1 U2520 ( .B1(n2270), .B2(n2267), .A(n2049), .ZN(n2264) );
  INV_X1 U2521 ( .A(n2267), .ZN(n2265) );
  INV_X1 U2522 ( .A(n3027), .ZN(n3614) );
  AND2_X1 U2523 ( .A1(n2833), .A2(n2988), .ZN(n3001) );
  AND2_X1 U2524 ( .A1(n4044), .A2(n4035), .ZN(n2206) );
  NAND2_X1 U2525 ( .A1(n2196), .A2(n2308), .ZN(n2348) );
  INV_X1 U2526 ( .A(n2352), .ZN(n2196) );
  INV_X1 U2527 ( .A(IR_REG_23__SCAN_IN), .ZN(n2818) );
  INV_X1 U2528 ( .A(IR_REG_15__SCAN_IN), .ZN(n2386) );
  NOR2_X1 U2529 ( .A1(n2579), .A2(IR_REG_10__SCAN_IN), .ZN(n2596) );
  NOR2_X1 U2530 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2106)
         );
  NOR2_X1 U2531 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2105)
         );
  INV_X1 U2532 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U2533 ( .A1(n4073), .A2(n2441), .ZN(n2684) );
  INV_X1 U2534 ( .A(n2785), .ZN(n2799) );
  INV_X1 U2535 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U2536 ( .A1(n3763), .A2(n2682), .ZN(n2712) );
  NAND2_X1 U2537 ( .A1(n2441), .A2(n4009), .ZN(n2714) );
  INV_X1 U2538 ( .A(n2660), .ZN(n2193) );
  NAND2_X1 U2539 ( .A1(n3015), .A2(n2484), .ZN(n3539) );
  AND2_X1 U2540 ( .A1(n3056), .A2(n3033), .ZN(n2852) );
  NAND2_X1 U2541 ( .A1(n2676), .A2(REG3_REG_19__SCAN_IN), .ZN(n2689) );
  NAND2_X1 U2542 ( .A1(n4054), .A2(n2682), .ZN(n2696) );
  NAND2_X1 U2543 ( .A1(n2682), .A2(n3558), .ZN(n2698) );
  OR2_X1 U2544 ( .A1(n2620), .A2(n3355), .ZN(n2643) );
  NOR2_X1 U2545 ( .A1(n3566), .A2(n2234), .ZN(n2233) );
  INV_X1 U2546 ( .A(n2242), .ZN(n2234) );
  NAND2_X1 U2547 ( .A1(n3489), .A2(n2716), .ZN(n2242) );
  NAND2_X1 U2548 ( .A1(n3550), .A2(n2236), .ZN(n2235) );
  INV_X1 U2549 ( .A(n2852), .ZN(n2854) );
  NOR2_X1 U2550 ( .A1(n2502), .A2(n2933), .ZN(n2517) );
  NAND2_X1 U2551 ( .A1(n3592), .A2(n2227), .ZN(n2112) );
  NAND2_X1 U2552 ( .A1(n2116), .A2(n2227), .ZN(n2108) );
  OR2_X1 U2553 ( .A1(n3962), .A2(n2790), .ZN(n2733) );
  INV_X1 U2554 ( .A(n4120), .ZN(n2146) );
  INV_X1 U2555 ( .A(n4152), .ZN(n2145) );
  INV_X1 U2556 ( .A(n4181), .ZN(n2143) );
  INV_X1 U2557 ( .A(n3331), .ZN(n2144) );
  INV_X1 U2558 ( .A(n3316), .ZN(n2137) );
  INV_X1 U2559 ( .A(n3258), .ZN(n2142) );
  INV_X1 U2560 ( .A(n3186), .ZN(n2138) );
  INV_X1 U2561 ( .A(n3167), .ZN(n2139) );
  NAND2_X1 U2562 ( .A1(n2406), .A2(REG3_REG_0__SCAN_IN), .ZN(n2419) );
  AOI21_X1 U2563 ( .B1(n2219), .B2(n2216), .A(n2976), .ZN(n2213) );
  INV_X1 U2564 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2216) );
  NOR2_X1 U2565 ( .A1(n4393), .A2(n2089), .ZN(n3812) );
  AOI21_X1 U2566 ( .B1(n3824), .B2(REG1_REG_11__SCAN_IN), .A(n4412), .ZN(n3814) );
  OAI21_X1 U2567 ( .B1(n4422), .B2(n2254), .A(n2253), .ZN(n4430) );
  NAND2_X1 U2568 ( .A1(n2255), .A2(REG1_REG_12__SCAN_IN), .ZN(n2254) );
  NAND2_X1 U2569 ( .A1(n3815), .A2(n2255), .ZN(n2253) );
  INV_X1 U2570 ( .A(n4431), .ZN(n2255) );
  INV_X1 U2571 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U2572 ( .A1(n2342), .A2(n2341), .ZN(n2650) );
  OAI22_X1 U2573 ( .A1(n4436), .A2(n4434), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3837), .ZN(n3838) );
  NAND2_X1 U2574 ( .A1(n4465), .A2(n3841), .ZN(n3842) );
  NAND2_X1 U2575 ( .A1(n4467), .A2(n3818), .ZN(n3819) );
  NAND2_X1 U2576 ( .A1(n3819), .A2(n3820), .ZN(n3849) );
  INV_X1 U2577 ( .A(n3868), .ZN(n3876) );
  OAI21_X1 U2578 ( .B1(n3890), .B2(n3889), .A(n3736), .ZN(n3871) );
  NOR2_X1 U2579 ( .A1(n2749), .A2(n3503), .ZN(n2759) );
  OR2_X1 U2580 ( .A1(n2740), .A2(n3533), .ZN(n2749) );
  AND4_X1 U2581 ( .A1(n2723), .A2(n2722), .A3(n2721), .A4(n2720), .ZN(n4002)
         );
  NAND2_X1 U2582 ( .A1(n4066), .A2(n2055), .ZN(n4011) );
  AND2_X1 U2583 ( .A1(n2664), .A2(REG3_REG_18__SCAN_IN), .ZN(n2676) );
  INV_X1 U2584 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2378) );
  OR2_X1 U2585 ( .A1(n2394), .A2(n2378), .ZN(n2380) );
  AOI21_X1 U2586 ( .B1(n4136), .B2(n2156), .A(n2154), .ZN(n2153) );
  INV_X1 U2587 ( .A(n2156), .ZN(n2155) );
  INV_X1 U2588 ( .A(n3675), .ZN(n2154) );
  NAND2_X1 U2589 ( .A1(n2644), .A2(REG3_REG_15__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U2590 ( .A1(n2158), .A2(n2156), .ZN(n4124) );
  INV_X1 U2591 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2604) );
  AND2_X1 U2592 ( .A1(n2572), .A2(REG3_REG_10__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U2593 ( .A1(n2590), .A2(REG3_REG_11__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U2594 ( .A1(n2266), .A2(n2272), .ZN(n3328) );
  OR2_X1 U2595 ( .A1(n3361), .A2(n3308), .ZN(n2266) );
  INV_X1 U2596 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2560) );
  NOR2_X1 U2597 ( .A1(n2561), .A2(n2560), .ZN(n2572) );
  AOI21_X1 U2598 ( .B1(n2162), .B2(n2161), .A(n2160), .ZN(n2159) );
  INV_X1 U2599 ( .A(n3667), .ZN(n2161) );
  INV_X1 U2600 ( .A(n3668), .ZN(n2160) );
  INV_X1 U2601 ( .A(n3239), .ZN(n3137) );
  OAI21_X1 U2602 ( .B1(n3132), .B2(n3131), .A(n3661), .ZN(n3196) );
  OR2_X1 U2603 ( .A1(n3116), .A2(n3544), .ZN(n3190) );
  NAND2_X1 U2604 ( .A1(n3110), .A2(n3658), .ZN(n3132) );
  AND2_X1 U2605 ( .A1(n3659), .A2(n3661), .ZN(n3616) );
  NAND2_X1 U2606 ( .A1(n3074), .A2(n3612), .ZN(n3110) );
  NAND2_X1 U2607 ( .A1(n2148), .A2(n3027), .ZN(n3073) );
  NAND2_X1 U2608 ( .A1(n3038), .A2(n3037), .ZN(n2148) );
  NAND2_X1 U2609 ( .A1(n2150), .A2(n2149), .ZN(n3038) );
  INV_X1 U2610 ( .A(n2985), .ZN(n2149) );
  INV_X1 U2611 ( .A(n3483), .ZN(n2996) );
  NOR2_X1 U2612 ( .A1(n4196), .A2(n4197), .ZN(n4195) );
  AND2_X1 U2613 ( .A1(n3629), .A2(DATAI_28_), .ZN(n3868) );
  NAND2_X1 U2614 ( .A1(n3960), .A2(n2054), .ZN(n3915) );
  NAND2_X1 U2615 ( .A1(n3960), .A2(n2053), .ZN(n3921) );
  AOI21_X1 U2616 ( .B1(n4006), .B2(n3385), .A(n2277), .ZN(n3983) );
  AND2_X1 U2617 ( .A1(n4021), .A2(n3416), .ZN(n2277) );
  NAND2_X1 U2618 ( .A1(n2278), .A2(n3635), .ZN(n4006) );
  OAI21_X1 U2619 ( .B1(n4043), .B2(n4018), .A(n2279), .ZN(n2278) );
  AND2_X1 U2620 ( .A1(n3634), .A2(n4019), .ZN(n2279) );
  AND2_X1 U2621 ( .A1(n3615), .A2(n3968), .ZN(n4005) );
  NAND2_X1 U2622 ( .A1(n4066), .A2(n2206), .ZN(n4034) );
  INV_X1 U2623 ( .A(n4053), .ZN(n4044) );
  AND2_X1 U2624 ( .A1(n4084), .A2(n4065), .ZN(n4066) );
  NAND2_X1 U2625 ( .A1(n4066), .A2(n4044), .ZN(n4046) );
  NAND2_X1 U2626 ( .A1(n4062), .A2(n2280), .ZN(n4043) );
  OR2_X1 U2627 ( .A1(n4091), .A2(n4072), .ZN(n2280) );
  NAND2_X1 U2628 ( .A1(n4107), .A2(n3694), .ZN(n4088) );
  INV_X1 U2629 ( .A(n3411), .ZN(n4090) );
  OR2_X1 U2630 ( .A1(n4118), .A2(n4110), .ZN(n4103) );
  NOR2_X1 U2631 ( .A1(n4103), .A2(n4090), .ZN(n4084) );
  NAND2_X1 U2632 ( .A1(n4127), .A2(n4110), .ZN(n3381) );
  OR2_X1 U2633 ( .A1(n4167), .A2(n4148), .ZN(n2295) );
  NAND2_X1 U2634 ( .A1(n3367), .A2(n2086), .ZN(n4177) );
  NAND2_X1 U2635 ( .A1(n3367), .A2(n2052), .ZN(n4176) );
  INV_X1 U2636 ( .A(n3309), .ZN(n3326) );
  NAND2_X1 U2637 ( .A1(n3367), .A2(n2051), .ZN(n3329) );
  NOR2_X1 U2638 ( .A1(n3255), .A2(n3303), .ZN(n3367) );
  AND2_X1 U2639 ( .A1(n3367), .A2(n3315), .ZN(n3368) );
  OR2_X1 U2640 ( .A1(n3254), .A2(n3248), .ZN(n3255) );
  NOR2_X1 U2641 ( .A1(n3190), .A2(n3191), .ZN(n3189) );
  AND2_X1 U2642 ( .A1(n3189), .A2(n2274), .ZN(n3166) );
  NOR2_X1 U2643 ( .A1(n3044), .A2(n3043), .ZN(n3079) );
  NAND2_X1 U2644 ( .A1(n2363), .A2(IR_REG_31__SCAN_IN), .ZN(n2879) );
  AND2_X1 U2645 ( .A1(n2208), .A2(n2361), .ZN(n2207) );
  NAND2_X1 U2646 ( .A1(n2819), .A2(n2818), .ZN(n2821) );
  NAND2_X1 U2647 ( .A1(n2344), .A2(IR_REG_31__SCAN_IN), .ZN(n2346) );
  AND2_X1 U2648 ( .A1(n2342), .A2(n2249), .ZN(n2356) );
  INV_X1 U2649 ( .A(IR_REG_16__SCAN_IN), .ZN(n2387) );
  INV_X1 U2650 ( .A(n2220), .ZN(n3447) );
  INV_X1 U2651 ( .A(n2228), .ZN(n2221) );
  INV_X1 U2652 ( .A(n3102), .ZN(n3103) );
  AOI21_X1 U2653 ( .B1(n3174), .B2(n2531), .A(n2540), .ZN(n3213) );
  NAND2_X1 U2654 ( .A1(n3550), .A2(n3554), .ZN(n3491) );
  NAND2_X1 U2655 ( .A1(n3629), .A2(DATAI_25_), .ZN(n3926) );
  NAND2_X1 U2656 ( .A1(n3539), .A2(n2488), .ZN(n3064) );
  INV_X1 U2657 ( .A(n2124), .ZN(n3527) );
  INV_X1 U2658 ( .A(n3570), .ZN(n3604) );
  INV_X1 U2659 ( .A(n3773), .ZN(n3089) );
  AND2_X1 U2660 ( .A1(n2235), .A2(n2233), .ZN(n3564) );
  NAND2_X1 U2661 ( .A1(n2235), .A2(n2242), .ZN(n3565) );
  NAND2_X1 U2662 ( .A1(n2122), .A2(n2121), .ZN(n3276) );
  AOI21_X1 U2663 ( .B1(n2586), .B2(n3266), .A(n2067), .ZN(n2121) );
  NAND2_X1 U2664 ( .A1(n2429), .A2(n2431), .ZN(n2432) );
  INV_X1 U2665 ( .A(n2430), .ZN(n2431) );
  OAI21_X1 U2666 ( .B1(n3519), .B2(n2081), .A(n2190), .ZN(n2189) );
  NAND2_X1 U2667 ( .A1(n2663), .A2(n3516), .ZN(n2190) );
  NOR2_X1 U2668 ( .A1(n3433), .A2(n2243), .ZN(n2657) );
  OR2_X1 U2669 ( .A1(n2840), .A2(n2839), .ZN(n3755) );
  OAI21_X1 U2670 ( .B1(n3912), .B2(n2790), .A(n2764), .ZN(n3935) );
  NOR2_X1 U2671 ( .A1(n2314), .A2(n2469), .ZN(n2474) );
  NAND3_X1 U2672 ( .A1(n2459), .A2(n2458), .A3(n2457), .ZN(n3543) );
  NAND2_X1 U2673 ( .A1(n2467), .A2(REG2_REG_3__SCAN_IN), .ZN(n2457) );
  OR2_X2 U2674 ( .A1(n2864), .A2(n2863), .ZN(n3772) );
  INV_X1 U2675 ( .A(n2215), .ZN(n2977) );
  OAI21_X1 U2676 ( .B1(n4383), .B2(n2216), .A(n2219), .ZN(n2215) );
  OR2_X1 U2677 ( .A1(n4382), .A2(n2916), .ZN(n2250) );
  XNOR2_X1 U2678 ( .A(n2169), .B(n2948), .ZN(n2946) );
  NAND2_X1 U2679 ( .A1(n2954), .A2(n2209), .ZN(n2959) );
  INV_X1 U2680 ( .A(n2952), .ZN(n2209) );
  AND2_X1 U2681 ( .A1(n2168), .A2(n2167), .ZN(n2963) );
  NAND2_X1 U2682 ( .A1(n2169), .A2(n4363), .ZN(n2167) );
  NAND2_X1 U2683 ( .A1(n2946), .A2(REG1_REG_6__SCAN_IN), .ZN(n2168) );
  OR2_X1 U2684 ( .A1(n2966), .A2(n3286), .ZN(n3809) );
  AND2_X1 U2685 ( .A1(n3811), .A2(n2256), .ZN(n4393) );
  INV_X1 U2686 ( .A(n4394), .ZN(n2256) );
  INV_X1 U2687 ( .A(n3811), .ZN(n4395) );
  XNOR2_X1 U2688 ( .A(n3812), .B(n4520), .ZN(n4404) );
  NOR2_X1 U2689 ( .A1(n4404), .A2(n4405), .ZN(n4403) );
  NAND2_X1 U2690 ( .A1(n4408), .A2(n3832), .ZN(n4417) );
  OAI21_X1 U2691 ( .B1(n4404), .B2(n2182), .A(n2181), .ZN(n4412) );
  NAND2_X1 U2692 ( .A1(n2183), .A2(REG1_REG_10__SCAN_IN), .ZN(n2182) );
  NAND2_X1 U2693 ( .A1(n3813), .A2(n2183), .ZN(n2181) );
  INV_X1 U2694 ( .A(n4413), .ZN(n2183) );
  XNOR2_X1 U2695 ( .A(n3835), .B(n4516), .ZN(n4427) );
  XNOR2_X1 U2696 ( .A(n3814), .B(n4516), .ZN(n4422) );
  NOR2_X1 U2697 ( .A1(n4422), .A2(n4423), .ZN(n4421) );
  NAND2_X1 U2698 ( .A1(n4427), .A2(REG2_REG_12__SCAN_IN), .ZN(n4426) );
  INV_X1 U2699 ( .A(n4460), .ZN(n2211) );
  INV_X1 U2700 ( .A(n2212), .ZN(n4459) );
  NAND2_X1 U2701 ( .A1(n2174), .A2(n2175), .ZN(n4453) );
  XNOR2_X1 U2702 ( .A(n3817), .B(n2389), .ZN(n4469) );
  NAND2_X1 U2703 ( .A1(n4469), .A2(n4468), .ZN(n4467) );
  XNOR2_X1 U2704 ( .A(n2103), .B(n3857), .ZN(n3862) );
  NOR2_X1 U2705 ( .A1(n4483), .A2(n2098), .ZN(n2103) );
  AND2_X1 U2706 ( .A1(n2173), .A2(n2172), .ZN(n3852) );
  NAND2_X1 U2707 ( .A1(n3856), .A2(REG1_REG_18__SCAN_IN), .ZN(n2172) );
  OR2_X1 U2708 ( .A1(n4380), .A2(n4377), .ZN(n4475) );
  NAND2_X1 U2709 ( .A1(n4196), .A2(n3435), .ZN(n3438) );
  NAND2_X1 U2710 ( .A1(n3432), .A2(n3431), .ZN(n3442) );
  NAND2_X1 U2711 ( .A1(n2285), .A2(n2284), .ZN(n3900) );
  OR2_X1 U2712 ( .A1(n2057), .A2(n2293), .ZN(n2284) );
  NAND2_X1 U2713 ( .A1(n2292), .A2(n2286), .ZN(n2285) );
  AND2_X1 U2714 ( .A1(n2292), .A2(n2064), .ZN(n3939) );
  NAND2_X1 U2715 ( .A1(n2263), .A2(n2267), .ZN(n3375) );
  NAND2_X1 U2716 ( .A1(n3361), .A2(n2269), .ZN(n2263) );
  NAND2_X1 U2717 ( .A1(n2297), .A2(n3242), .ZN(n3302) );
  NAND2_X1 U2718 ( .A1(n2276), .A2(n2273), .ZN(n3152) );
  NAND2_X1 U2719 ( .A1(n3150), .A2(n3149), .ZN(n3157) );
  INV_X1 U2720 ( .A(n3860), .ZN(n3850) );
  INV_X1 U2721 ( .A(n4496), .ZN(n4180) );
  AND2_X1 U2722 ( .A1(n4080), .A2(n4551), .ZN(n4498) );
  INV_X1 U2723 ( .A(n4498), .ZN(n4151) );
  INV_X1 U2724 ( .A(n4188), .ZN(n4499) );
  NAND2_X1 U2725 ( .A1(n4556), .A2(REG0_REG_29__SCAN_IN), .ZN(n2204) );
  AND2_X1 U2726 ( .A1(n2294), .A2(n2063), .ZN(n3920) );
  NAND2_X1 U2727 ( .A1(n2292), .A2(n2291), .ZN(n2294) );
  OR2_X1 U2728 ( .A1(n3953), .A2(n3952), .ZN(n4304) );
  INV_X1 U2729 ( .A(n4330), .ZN(n4358) );
  XNOR2_X1 U2730 ( .A(n2844), .B(n4596), .ZN(n4367) );
  OR2_X1 U2731 ( .A1(n2362), .A2(n2259), .ZN(n2354) );
  AND2_X1 U2732 ( .A1(n2922), .A2(STATE_REG_SCAN_IN), .ZN(n4506) );
  XNOR2_X1 U2733 ( .A(n2372), .B(IR_REG_22__SCAN_IN), .ZN(n3756) );
  XNOR2_X1 U2734 ( .A(n2347), .B(IR_REG_21__SCAN_IN), .ZN(n3652) );
  NOR2_X1 U2735 ( .A1(n2300), .A2(n2323), .ZN(n2301) );
  XNOR2_X1 U2736 ( .A(n2369), .B(n2368), .ZN(n3860) );
  INV_X1 U2737 ( .A(IR_REG_8__SCAN_IN), .ZN(n2320) );
  INV_X1 U2738 ( .A(IR_REG_5__SCAN_IN), .ZN(n2321) );
  XNOR2_X1 U2739 ( .A(n2476), .B(IR_REG_4__SCAN_IN), .ZN(n4390) );
  AND2_X1 U2740 ( .A1(n2475), .A2(n2463), .ZN(n4364) );
  OR2_X1 U2741 ( .A1(n2442), .A2(n2259), .ZN(n2443) );
  AND2_X1 U2742 ( .A1(n2260), .A2(n2258), .ZN(n2257) );
  INV_X1 U2743 ( .A(IR_REG_0__SCAN_IN), .ZN(n2316) );
  OR2_X1 U2744 ( .A1(n2860), .A2(n2825), .ZN(n2862) );
  INV_X1 U2745 ( .A(n3595), .ZN(n2113) );
  AOI21_X1 U2746 ( .B1(n4482), .B2(n2173), .A(n4481), .ZN(n4489) );
  OAI21_X1 U2747 ( .B1(n3436), .B2(n4565), .A(n2165), .ZN(n3437) );
  OR2_X1 U2748 ( .A1(n4568), .A2(REG1_REG_29__SCAN_IN), .ZN(n2165) );
  NAND2_X1 U2749 ( .A1(n2205), .A2(n2202), .ZN(U3515) );
  NAND2_X1 U2750 ( .A1(n3436), .A2(n4756), .ZN(n2205) );
  INV_X1 U2751 ( .A(n2203), .ZN(n2202) );
  OAI21_X1 U2752 ( .B1(n3445), .B2(n4341), .A(n2204), .ZN(n2203) );
  INV_X1 U2753 ( .A(IR_REG_31__SCAN_IN), .ZN(n2259) );
  INV_X1 U2754 ( .A(n3466), .ZN(n3315) );
  AND2_X1 U2755 ( .A1(n3966), .A2(n3702), .ZN(n3410) );
  AND2_X1 U2756 ( .A1(n2311), .A2(n2830), .ZN(n2047) );
  AND2_X1 U2757 ( .A1(n2073), .A2(n3149), .ZN(n2048) );
  NOR2_X1 U2758 ( .A1(n4170), .A2(n3374), .ZN(n2049) );
  OR2_X1 U2759 ( .A1(n3440), .A2(n2790), .ZN(n2050) );
  NAND2_X1 U2760 ( .A1(n2959), .A2(n2085), .ZN(n3827) );
  INV_X1 U2761 ( .A(n3159), .ZN(n2274) );
  INV_X1 U2762 ( .A(n3499), .ZN(n2227) );
  AND2_X1 U2763 ( .A1(n3315), .A2(n3326), .ZN(n2051) );
  AND2_X1 U2764 ( .A1(n2051), .A2(n3374), .ZN(n2052) );
  AND2_X1 U2765 ( .A1(n3926), .A2(n3951), .ZN(n2053) );
  AND2_X1 U2766 ( .A1(n2053), .A2(n3905), .ZN(n2054) );
  AND2_X1 U2767 ( .A1(n2206), .A2(n3416), .ZN(n2055) );
  INV_X1 U2768 ( .A(n2840), .ZN(n2441) );
  OR2_X1 U2769 ( .A1(n3816), .A2(n4513), .ZN(n2056) );
  XNOR2_X1 U2770 ( .A(n2346), .B(n2345), .ZN(n2374) );
  NAND2_X1 U2771 ( .A1(n2319), .A2(n2310), .ZN(n2495) );
  NOR2_X1 U2772 ( .A1(n3906), .A2(n3926), .ZN(n2057) );
  INV_X1 U2773 ( .A(n2416), .ZN(n2796) );
  AND4_X1 U2774 ( .A1(n2357), .A2(n4595), .A3(n2341), .A4(n2345), .ZN(n2058)
         );
  NAND2_X1 U2775 ( .A1(n2467), .A2(REG2_REG_4__SCAN_IN), .ZN(n2059) );
  NAND2_X1 U2776 ( .A1(n3768), .A2(n3303), .ZN(n2060) );
  AND2_X1 U2777 ( .A1(n2249), .A2(n2357), .ZN(n2061) );
  NAND2_X1 U2778 ( .A1(n2534), .A2(n2535), .ZN(n2062) );
  OR2_X1 U2779 ( .A1(n3973), .A2(n3530), .ZN(n2063) );
  NAND2_X1 U2780 ( .A1(n3987), .A2(n3961), .ZN(n2064) );
  AND2_X1 U2781 ( .A1(n2116), .A2(n3498), .ZN(n2065) );
  OR2_X1 U2782 ( .A1(n4513), .A2(n3838), .ZN(n2066) );
  INV_X1 U2783 ( .A(n2319), .ZN(n2460) );
  AND2_X1 U2784 ( .A1(n2589), .A2(n2588), .ZN(n2067) );
  NOR2_X1 U2785 ( .A1(n2057), .A2(n2287), .ZN(n2068) );
  OR2_X1 U2786 ( .A1(n4477), .A2(n4476), .ZN(n2173) );
  AND2_X1 U2787 ( .A1(n2231), .A2(n2233), .ZN(n2069) );
  NOR2_X1 U2788 ( .A1(n3765), .A2(n3376), .ZN(n2070) );
  INV_X1 U2789 ( .A(n2238), .ZN(n3453) );
  OAI21_X1 U2790 ( .B1(n3550), .B2(n2232), .A(n2230), .ZN(n2238) );
  AND2_X1 U2791 ( .A1(n3327), .A2(n3326), .ZN(n2071) );
  NAND2_X1 U2792 ( .A1(n2125), .A2(n2301), .ZN(n2072) );
  INV_X1 U2793 ( .A(IR_REG_22__SCAN_IN), .ZN(n2325) );
  INV_X1 U2794 ( .A(IR_REG_13__SCAN_IN), .ZN(n2341) );
  XNOR2_X1 U2795 ( .A(n2415), .B(n2782), .ZN(n2429) );
  INV_X1 U2796 ( .A(n2270), .ZN(n2269) );
  NAND2_X1 U2797 ( .A1(n2272), .A2(n2271), .ZN(n2270) );
  NAND2_X1 U2798 ( .A1(n3183), .A2(n3159), .ZN(n2073) );
  OR2_X1 U2799 ( .A1(n2859), .A2(n2858), .ZN(n2074) );
  AND2_X1 U2800 ( .A1(n3242), .A2(n2060), .ZN(n2075) );
  AND2_X1 U2801 ( .A1(n2454), .A2(REG0_REG_3__SCAN_IN), .ZN(n2076) );
  AND2_X1 U2802 ( .A1(n3151), .A2(n2273), .ZN(n2077) );
  INV_X1 U2803 ( .A(n2488), .ZN(n2119) );
  AND2_X1 U2804 ( .A1(n2177), .A2(n2056), .ZN(n2078) );
  AND2_X1 U2805 ( .A1(n2061), .A2(n2248), .ZN(n2079) );
  INV_X1 U2806 ( .A(n2163), .ZN(n2162) );
  INV_X1 U2807 ( .A(IR_REG_18__SCAN_IN), .ZN(n2248) );
  NAND4_X1 U2808 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2313), .ZN(n2984)
         );
  NAND2_X1 U2809 ( .A1(n2885), .A2(n2332), .ZN(n2434) );
  NAND2_X1 U2810 ( .A1(n2246), .A2(n3274), .ZN(n3292) );
  NAND4_X1 U2811 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n3183)
         );
  INV_X1 U2812 ( .A(n2198), .ZN(n2804) );
  XNOR2_X1 U2813 ( .A(n2120), .B(IR_REG_24__SCAN_IN), .ZN(n2198) );
  NAND2_X1 U2814 ( .A1(n2411), .A2(n2257), .ZN(n3778) );
  OR2_X1 U2815 ( .A1(n2974), .A2(n2920), .ZN(n2080) );
  NAND2_X1 U2816 ( .A1(n2262), .A2(n2261), .ZN(n4158) );
  INV_X1 U2817 ( .A(n3498), .ZN(n2109) );
  NAND2_X1 U2818 ( .A1(n2641), .A2(n2640), .ZN(n3336) );
  INV_X1 U2819 ( .A(n3694), .ZN(n2132) );
  INV_X1 U2820 ( .A(IR_REG_24__SCAN_IN), .ZN(n2353) );
  AND2_X1 U2821 ( .A1(n3517), .A2(n2662), .ZN(n2081) );
  INV_X1 U2822 ( .A(n3338), .ZN(n2187) );
  INV_X1 U2823 ( .A(n4178), .ZN(n4165) );
  NOR2_X1 U2824 ( .A1(n4421), .A2(n3815), .ZN(n2082) );
  INV_X1 U2825 ( .A(n3374), .ZN(n3376) );
  NOR2_X1 U2826 ( .A1(n3328), .A2(n3617), .ZN(n2083) );
  NAND2_X1 U2827 ( .A1(n2990), .A2(n2989), .ZN(n3649) );
  INV_X1 U2828 ( .A(n3649), .ZN(n2150) );
  OR2_X1 U2829 ( .A1(n3438), .A2(n4530), .ZN(n2084) );
  OR2_X1 U2830 ( .A1(n2960), .A2(n2951), .ZN(n2085) );
  AND2_X1 U2831 ( .A1(n2052), .A2(n4178), .ZN(n2086) );
  AND2_X1 U2832 ( .A1(n2158), .A2(n3686), .ZN(n2087) );
  INV_X1 U2833 ( .A(n3734), .ZN(n2128) );
  INV_X1 U2834 ( .A(IR_REG_28__SCAN_IN), .ZN(n4596) );
  AND2_X1 U2835 ( .A1(n2227), .A2(n2109), .ZN(n2088) );
  NAND2_X1 U2836 ( .A1(n2342), .A2(n2061), .ZN(n2359) );
  INV_X1 U2837 ( .A(n3834), .ZN(n4516) );
  OR2_X1 U2838 ( .A1(n3265), .A2(n3266), .ZN(n3263) );
  NAND2_X1 U2839 ( .A1(n3016), .A2(n3017), .ZN(n3015) );
  INV_X1 U2840 ( .A(n3558), .ZN(n4035) );
  AND2_X1 U2841 ( .A1(n3825), .A2(REG1_REG_9__SCAN_IN), .ZN(n2089) );
  NAND2_X1 U2842 ( .A1(n3263), .A2(n2586), .ZN(n3462) );
  INV_X1 U2843 ( .A(n3893), .ZN(n3883) );
  INV_X1 U2844 ( .A(n3416), .ZN(n4009) );
  NOR2_X1 U2845 ( .A1(n4403), .A2(n3813), .ZN(n2090) );
  AND2_X1 U2846 ( .A1(n3629), .A2(DATAI_22_), .ZN(n3990) );
  INV_X1 U2847 ( .A(n3990), .ZN(n3569) );
  INV_X1 U2848 ( .A(n2455), .ZN(n2489) );
  OR2_X1 U2849 ( .A1(n4522), .A2(n3237), .ZN(n2091) );
  AND2_X1 U2850 ( .A1(n2054), .A2(n3893), .ZN(n2092) );
  AND2_X1 U2851 ( .A1(n2055), .A2(n3569), .ZN(n2093) );
  INV_X2 U2852 ( .A(n4556), .ZN(n4756) );
  INV_X2 U2853 ( .A(n4565), .ZN(n4568) );
  OR2_X1 U2854 ( .A1(n3057), .A2(n3031), .ZN(n4565) );
  OR2_X1 U2855 ( .A1(n3855), .A2(REG1_REG_17__SCAN_IN), .ZN(n2094) );
  OR2_X1 U2856 ( .A1(n3855), .A2(REG2_REG_17__SCAN_IN), .ZN(n2095) );
  AND2_X1 U2857 ( .A1(n2250), .A2(n2918), .ZN(n2096) );
  INV_X1 U2858 ( .A(n4047), .ZN(n2147) );
  NAND2_X1 U2859 ( .A1(n3839), .A2(REG1_REG_15__SCAN_IN), .ZN(n2097) );
  AND2_X1 U2860 ( .A1(n3856), .A2(REG2_REG_18__SCAN_IN), .ZN(n2098) );
  INV_X1 U2861 ( .A(n4495), .ZN(n2140) );
  INV_X1 U2862 ( .A(n3269), .ZN(n2141) );
  NAND2_X1 U2863 ( .A1(n2351), .A2(n2350), .ZN(n2876) );
  INV_X1 U2864 ( .A(n2876), .ZN(n2197) );
  INV_X1 U2865 ( .A(IR_REG_29__SCAN_IN), .ZN(n2327) );
  INV_X1 U2866 ( .A(n3205), .ZN(n2136) );
  INV_X1 U2867 ( .A(DATAI_0_), .ZN(n2201) );
  NAND2_X1 U2868 ( .A1(n4398), .A2(n2091), .ZN(n3831) );
  NAND2_X1 U2869 ( .A1(n4416), .A2(n3833), .ZN(n3835) );
  XNOR2_X1 U2870 ( .A(n3840), .B(n2389), .ZN(n4466) );
  INV_X1 U2871 ( .A(n4444), .ZN(n2099) );
  NAND3_X1 U2872 ( .A1(n2319), .A2(n2310), .A3(n2104), .ZN(n2567) );
  NAND3_X1 U2873 ( .A1(n2111), .A2(n2110), .A3(n2107), .ZN(n2115) );
  NAND2_X1 U2874 ( .A1(n2114), .A2(n2113), .ZN(U3237) );
  NAND2_X1 U2875 ( .A1(n2115), .A2(n3609), .ZN(n2114) );
  INV_X1 U2876 ( .A(n3592), .ZN(n2116) );
  NAND3_X1 U2877 ( .A1(n2118), .A2(n2117), .A3(n3063), .ZN(n3174) );
  NAND3_X1 U2878 ( .A1(n3016), .A2(n2488), .A3(n3017), .ZN(n2118) );
  NAND2_X1 U2879 ( .A1(n3265), .A2(n2586), .ZN(n2122) );
  NAND2_X2 U2880 ( .A1(n2370), .A2(n2325), .ZN(n2352) );
  AND2_X2 U2881 ( .A1(n2125), .A2(n2298), .ZN(n2370) );
  OAI21_X1 U2882 ( .B1(n4107), .B2(n3732), .A(n2130), .ZN(n3941) );
  NAND2_X1 U2883 ( .A1(n4107), .A2(n2130), .ZN(n2129) );
  NAND2_X1 U2884 ( .A1(n2134), .A2(n2135), .ZN(n2473) );
  NAND2_X1 U2885 ( .A1(n2134), .A2(n2136), .ZN(n2492) );
  NAND2_X1 U2886 ( .A1(n2134), .A2(n2137), .ZN(n2593) );
  NAND2_X1 U2887 ( .A1(n2134), .A2(n2138), .ZN(n2520) );
  NAND2_X1 U2888 ( .A1(n2134), .A2(n2139), .ZN(n2505) );
  NAND2_X1 U2889 ( .A1(n2134), .A2(n2140), .ZN(n2576) );
  NAND2_X1 U2890 ( .A1(n2134), .A2(n2141), .ZN(n2564) );
  NAND2_X1 U2891 ( .A1(n2134), .A2(n2142), .ZN(n2545) );
  NAND2_X1 U2892 ( .A1(n2134), .A2(n2143), .ZN(n2623) );
  NAND2_X1 U2893 ( .A1(n2134), .A2(n2144), .ZN(n2608) );
  NAND2_X1 U2894 ( .A1(n2145), .A2(n2134), .ZN(n2647) );
  NAND2_X1 U2895 ( .A1(n2146), .A2(n2134), .ZN(n2396) );
  NAND2_X1 U2896 ( .A1(n2147), .A2(n2134), .ZN(n2679) );
  NAND2_X2 U2897 ( .A1(n3037), .A2(n3650), .ZN(n2985) );
  NOR2_X2 U2898 ( .A1(n2352), .A2(n2304), .ZN(n2843) );
  OAI21_X1 U2899 ( .B1(n4134), .B2(n2155), .A(n2153), .ZN(n4109) );
  OAI21_X1 U2900 ( .B1(n3230), .B2(n2163), .A(n2159), .ZN(n3299) );
  OAI21_X1 U2901 ( .B1(n3230), .B2(n3229), .A(n3667), .ZN(n3247) );
  NAND2_X1 U2902 ( .A1(n3669), .A2(n2164), .ZN(n2163) );
  NAND2_X1 U2903 ( .A1(n3229), .A2(n3667), .ZN(n2164) );
  INV_X1 U2904 ( .A(n2177), .ZN(n4440) );
  OR2_X1 U2905 ( .A1(n4365), .A2(n2910), .ZN(n2179) );
  XNOR2_X2 U2906 ( .A(n2443), .B(IR_REG_2__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U2907 ( .A1(n2179), .A2(n2178), .ZN(n2180) );
  NAND2_X1 U2908 ( .A1(n4365), .A2(n2910), .ZN(n2178) );
  NAND2_X1 U2909 ( .A1(n2184), .A2(n2903), .ZN(n2428) );
  XNOR2_X1 U2910 ( .A(n2184), .B(n2903), .ZN(n3800) );
  NAND2_X1 U2911 ( .A1(n2424), .A2(n2425), .ZN(n2184) );
  OAI21_X1 U2912 ( .B1(n3338), .B2(n3336), .A(n2188), .ZN(n2659) );
  INV_X1 U2913 ( .A(n3087), .ZN(n2989) );
  MUX2_X1 U2914 ( .A(n2316), .B(n2201), .S(n2477), .Z(n3087) );
  NAND3_X1 U2915 ( .A1(n2200), .A2(n2199), .A3(n2364), .ZN(n2477) );
  NAND2_X1 U2916 ( .A1(n2370), .A2(n2207), .ZN(n2363) );
  NAND2_X1 U2917 ( .A1(n2214), .A2(n2213), .ZN(n2218) );
  NAND2_X1 U2918 ( .A1(n4383), .A2(n2219), .ZN(n2214) );
  INV_X1 U2919 ( .A(n2218), .ZN(n2975) );
  NAND2_X1 U2920 ( .A1(n2927), .A2(n4390), .ZN(n2219) );
  XOR2_X1 U2921 ( .A(n4448), .B(n3838), .Z(n4445) );
  NAND2_X1 U2922 ( .A1(n2682), .A2(n2984), .ZN(n2421) );
  CLKBUF_X1 U2923 ( .A(n2840), .Z(n2243) );
  NAND2_X1 U2924 ( .A1(n3276), .A2(n3273), .ZN(n2246) );
  NAND2_X1 U2925 ( .A1(n2246), .A2(n2244), .ZN(n2641) );
  NAND2_X1 U2926 ( .A1(n2342), .A2(n2079), .ZN(n2247) );
  NAND3_X1 U2927 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_31__SCAN_IN), .ZN(n2260) );
  NAND2_X1 U2928 ( .A1(n3026), .A2(n3614), .ZN(n3030) );
  NAND2_X1 U2929 ( .A1(n3361), .A2(n2264), .ZN(n2262) );
  AOI21_X2 U2930 ( .B1(n2272), .B2(n2268), .A(n2071), .ZN(n2267) );
  NAND2_X1 U2931 ( .A1(n2276), .A2(n2077), .ZN(n4544) );
  INV_X1 U2932 ( .A(n3183), .ZN(n2275) );
  NAND2_X1 U2933 ( .A1(n3959), .A2(n3386), .ZN(n2292) );
  NAND2_X1 U2934 ( .A1(n3959), .A2(n2282), .ZN(n2281) );
  NAND2_X1 U2935 ( .A1(n2297), .A2(n2075), .ZN(n3306) );
  NAND2_X1 U2936 ( .A1(n3089), .A2(n3483), .ZN(n3037) );
  NAND2_X1 U2937 ( .A1(n3773), .A2(n2996), .ZN(n3650) );
  AOI21_X1 U2938 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n4482) );
  NAND2_X1 U2939 ( .A1(n2467), .A2(REG2_REG_2__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U2940 ( .A1(n2467), .A2(REG2_REG_1__SCAN_IN), .ZN(n2408) );
  NOR2_X1 U2941 ( .A1(n2434), .A2(n3046), .ZN(n2438) );
  NAND2_X1 U2942 ( .A1(n2406), .A2(n2456), .ZN(n2458) );
  NAND2_X1 U2943 ( .A1(n3008), .A2(n2453), .ZN(n3016) );
  INV_X1 U2944 ( .A(n2332), .ZN(n2336) );
  NAND2_X1 U2945 ( .A1(n2330), .A2(IR_REG_31__SCAN_IN), .ZN(n2331) );
  OAI21_X1 U2946 ( .B1(n4002), .B2(n3569), .A(n3982), .ZN(n3959) );
  OAI21_X2 U2947 ( .B1(n3882), .B2(n3393), .A(n3392), .ZN(n3865) );
  AND2_X1 U2948 ( .A1(n2818), .A2(n2353), .ZN(n2308) );
  INV_X1 U2949 ( .A(n4127), .ZN(n4094) );
  AND2_X1 U2950 ( .A1(n2829), .A2(n3609), .ZN(n2311) );
  AND2_X1 U2951 ( .A1(n4140), .A2(n3433), .ZN(n2312) );
  NAND2_X1 U2952 ( .A1(n2467), .A2(REG2_REG_0__SCAN_IN), .ZN(n2313) );
  AND2_X1 U2953 ( .A1(n2454), .A2(REG0_REG_4__SCAN_IN), .ZN(n2314) );
  AND2_X1 U2954 ( .A1(n2455), .A2(REG1_REG_3__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2955 ( .A1(n4180), .A2(n3034), .ZN(n4373) );
  INV_X1 U2956 ( .A(IR_REG_21__SCAN_IN), .ZN(n2324) );
  AND2_X1 U2957 ( .A1(n3632), .A2(n3940), .ZN(n3734) );
  AND2_X1 U2958 ( .A1(n3419), .A2(n3418), .ZN(n3731) );
  INV_X1 U2959 ( .A(n2486), .ZN(n2487) );
  INV_X1 U2960 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3556) );
  INV_X1 U2961 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2933) );
  INV_X1 U2962 ( .A(n3543), .ZN(n3104) );
  NAND2_X1 U2963 ( .A1(n2485), .A2(n2487), .ZN(n2488) );
  AND2_X1 U2964 ( .A1(n2619), .A2(n2618), .ZN(n3349) );
  NOR2_X1 U2965 ( .A1(n2705), .A2(n2704), .ZN(n2718) );
  AND2_X1 U2966 ( .A1(n2773), .A2(REG3_REG_27__SCAN_IN), .ZN(n2786) );
  AND2_X1 U2967 ( .A1(n3756), .A2(n3652), .ZN(n2988) );
  OR2_X1 U2968 ( .A1(n2689), .A2(n3556), .ZN(n2705) );
  NOR2_X1 U2969 ( .A1(n2380), .A2(n4610), .ZN(n2664) );
  NOR2_X1 U2970 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  OR2_X1 U2971 ( .A1(n2605), .A2(n2604), .ZN(n2620) );
  OR2_X1 U2972 ( .A1(n2542), .A2(n2541), .ZN(n2561) );
  AND2_X1 U2973 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2490) );
  INV_X1 U2974 ( .A(n3713), .ZN(n3705) );
  INV_X1 U2975 ( .A(n4072), .ZN(n4065) );
  INV_X1 U2976 ( .A(n4126), .ZN(n3433) );
  AND2_X1 U2977 ( .A1(n3658), .A2(n3655), .ZN(n3612) );
  AND2_X1 U2978 ( .A1(n2984), .A2(n2989), .ZN(n2986) );
  OR2_X1 U2979 ( .A1(n2728), .A2(n2727), .ZN(n2740) );
  INV_X1 U2980 ( .A(n3987), .ZN(n3944) );
  AND2_X1 U2981 ( .A1(n2855), .A2(n4180), .ZN(n3570) );
  AND2_X1 U2982 ( .A1(n2759), .A2(REG3_REG_26__SCAN_IN), .ZN(n2773) );
  INV_X1 U2983 ( .A(n3792), .ZN(n3793) );
  INV_X1 U2984 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4610) );
  OR2_X1 U2985 ( .A1(n2786), .A2(n2774), .ZN(n3887) );
  INV_X1 U2986 ( .A(n3764), .ZN(n4140) );
  INV_X1 U2987 ( .A(n4172), .ZN(n4147) );
  AND2_X1 U2988 ( .A1(n3400), .A2(n3397), .ZN(n3617) );
  INV_X1 U2989 ( .A(n3665), .ZN(n3151) );
  OR2_X1 U2990 ( .A1(n3147), .A2(n3146), .ZN(n3192) );
  NAND2_X1 U2991 ( .A1(n4361), .A2(n3085), .ZN(n4200) );
  INV_X1 U2992 ( .A(n3905), .ZN(n3913) );
  AND2_X1 U2993 ( .A1(n3629), .A2(DATAI_20_), .ZN(n3558) );
  INV_X1 U2994 ( .A(n4530), .ZN(n4551) );
  NAND2_X1 U2995 ( .A1(n2983), .A2(n3860), .ZN(n4175) );
  NAND2_X1 U2996 ( .A1(n2864), .A2(n4506), .ZN(n3002) );
  AND2_X1 U2997 ( .A1(n2842), .A2(n2905), .ZN(n3607) );
  INV_X1 U2998 ( .A(n2406), .ZN(n2790) );
  INV_X1 U2999 ( .A(n4475), .ZN(n4471) );
  INV_X1 U3000 ( .A(n4200), .ZN(n4192) );
  AND2_X1 U3001 ( .A1(n4373), .A2(n3860), .ZN(n4080) );
  INV_X1 U3002 ( .A(n4368), .ZN(n4183) );
  AND2_X1 U3003 ( .A1(n4568), .A2(n4551), .ZN(n4248) );
  NAND2_X1 U3004 ( .A1(n4101), .A2(n4100), .ZN(n4099) );
  NAND2_X1 U3005 ( .A1(n4175), .A2(n4531), .ZN(n4549) );
  AND2_X1 U3006 ( .A1(n4756), .A2(n4551), .ZN(n4330) );
  INV_X1 U3007 ( .A(n4531), .ZN(n4540) );
  OR2_X1 U3008 ( .A1(n2854), .A2(n2823), .ZN(n3577) );
  INV_X1 U3009 ( .A(n3394), .ZN(n3895) );
  NAND4_X1 U3010 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .ZN(n4054)
         );
  OR2_X1 U3011 ( .A1(n4380), .A2(n3802), .ZN(n4443) );
  NAND2_X1 U3012 ( .A1(n4183), .A2(n3154), .ZN(n4133) );
  NAND2_X1 U3013 ( .A1(n4183), .A2(n3036), .ZN(n4188) );
  NAND2_X1 U3014 ( .A1(n4568), .A2(n4549), .ZN(n4257) );
  INV_X1 U3015 ( .A(n4248), .ZN(n4276) );
  NAND2_X1 U3016 ( .A1(n4756), .A2(n4549), .ZN(n4341) );
  AND3_X1 U3017 ( .A1(n4555), .A2(n4554), .A3(n4553), .ZN(n4567) );
  OR2_X1 U3018 ( .A1(n3057), .A2(n3056), .ZN(n4556) );
  NAND2_X1 U3019 ( .A1(n2904), .A2(n3000), .ZN(n4505) );
  INV_X1 U3020 ( .A(n3837), .ZN(n4514) );
  XNOR2_X1 U3021 ( .A(n2549), .B(IR_REG_7__SCAN_IN), .ZN(n4362) );
  INV_X1 U3022 ( .A(n3772), .ZN(U4043) );
  INV_X2 U3023 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U3024 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2326)
         );
  NAND2_X1 U3025 ( .A1(n2843), .A2(n4596), .ZN(n2330) );
  INV_X1 U3026 ( .A(n2330), .ZN(n2328) );
  NAND2_X1 U3027 ( .A1(n2328), .A2(n2327), .ZN(n2882) );
  XNOR2_X1 U3028 ( .A(n2334), .B(n2329), .ZN(n2333) );
  NAND2_X1 U3029 ( .A1(n3424), .A2(REG0_REG_17__SCAN_IN), .ZN(n2340) );
  INV_X4 U3030 ( .A(n2489), .ZN(n2775) );
  NAND2_X1 U3031 ( .A1(n2775), .A2(REG1_REG_17__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U3032 ( .A1(n2490), .A2(REG3_REG_5__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U3033 ( .A1(n2517), .A2(REG3_REG_7__SCAN_IN), .ZN(n2542) );
  AND2_X1 U3034 ( .A1(n2380), .A2(n4610), .ZN(n2335) );
  OR2_X1 U3035 ( .A1(n2335), .A2(n2664), .ZN(n4085) );
  OR2_X1 U3036 ( .A1(n2790), .A2(n4085), .ZN(n2338) );
  INV_X2 U3037 ( .A(n2467), .ZN(n2895) );
  INV_X1 U3038 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4096) );
  OR2_X1 U3039 ( .A1(n2895), .A2(n4096), .ZN(n2337) );
  NAND4_X1 U3040 ( .A1(n2340), .A2(n2339), .A3(n2338), .A4(n2337), .ZN(n4111)
         );
  NAND3_X1 U3041 ( .A1(n4595), .A2(n2386), .A3(n2387), .ZN(n2343) );
  NAND2_X1 U3042 ( .A1(n2369), .A2(n2368), .ZN(n2344) );
  NAND2_X1 U3043 ( .A1(n2072), .A2(IR_REG_31__SCAN_IN), .ZN(n2347) );
  INV_X1 U3044 ( .A(n3035), .ZN(n2355) );
  NAND2_X1 U3045 ( .A1(n2348), .A2(IR_REG_31__SCAN_IN), .ZN(n2349) );
  INV_X1 U3046 ( .A(n2362), .ZN(n2350) );
  NAND2_X1 U3047 ( .A1(n2352), .A2(IR_REG_31__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U3048 ( .A1(n4111), .A2(n2682), .ZN(n2367) );
  OR2_X1 U3049 ( .A1(n2356), .A2(n2259), .ZN(n2358) );
  MUX2_X1 U3050 ( .A(n2358), .B(IR_REG_31__SCAN_IN), .S(n2357), .Z(n2360) );
  NAND2_X1 U3051 ( .A1(n2360), .A2(n2359), .ZN(n3823) );
  INV_X1 U3052 ( .A(DATAI_17_), .ZN(n2365) );
  INV_X1 U3053 ( .A(IR_REG_26__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3054 ( .A1(n4596), .A2(IR_REG_27__SCAN_IN), .ZN(n2364) );
  MUX2_X1 U3055 ( .A(n3823), .B(n2365), .S(n3629), .Z(n3411) );
  AND2_X2 U3056 ( .A1(n2864), .A2(n3035), .ZN(n2416) );
  NAND2_X1 U3057 ( .A1(n4090), .A2(n2416), .ZN(n2366) );
  NAND2_X1 U3058 ( .A1(n2367), .A2(n2366), .ZN(n2373) );
  INV_X1 U3059 ( .A(n2370), .ZN(n2371) );
  NAND2_X1 U3060 ( .A1(n2371), .A2(IR_REG_31__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U3061 ( .A1(n3860), .A2(n3756), .ZN(n2837) );
  XNOR2_X1 U3062 ( .A(n2373), .B(n2797), .ZN(n3517) );
  INV_X1 U3063 ( .A(n3517), .ZN(n2663) );
  INV_X1 U3064 ( .A(n3756), .ZN(n2376) );
  INV_X1 U3065 ( .A(n3652), .ZN(n2375) );
  AND2_X4 U3066 ( .A1(n2416), .A2(n4530), .ZN(n2785) );
  NOR2_X1 U3067 ( .A1(n3411), .A2(n2243), .ZN(n2377) );
  AOI21_X1 U3068 ( .B1(n4111), .B2(n2785), .A(n2377), .ZN(n2662) );
  INV_X1 U3069 ( .A(n2662), .ZN(n3516) );
  NAND2_X1 U3070 ( .A1(n3424), .A2(REG0_REG_16__SCAN_IN), .ZN(n2384) );
  NAND2_X1 U3071 ( .A1(n2775), .A2(REG1_REG_16__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U3072 ( .A1(n2394), .A2(n2378), .ZN(n2379) );
  NAND2_X1 U3073 ( .A1(n2380), .A2(n2379), .ZN(n4104) );
  INV_X1 U3074 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4105) );
  OR2_X1 U3075 ( .A1(n2895), .A2(n4105), .ZN(n2381) );
  NAND4_X1 U3076 ( .A1(n2384), .A2(n2383), .A3(n2382), .A4(n2381), .ZN(n4127)
         );
  OR2_X1 U3077 ( .A1(n2650), .A2(IR_REG_14__SCAN_IN), .ZN(n2385) );
  NAND2_X1 U3078 ( .A1(n2385), .A2(IR_REG_31__SCAN_IN), .ZN(n2399) );
  NAND2_X1 U3079 ( .A1(n2399), .A2(n2386), .ZN(n2401) );
  NAND2_X1 U3080 ( .A1(n2401), .A2(IR_REG_31__SCAN_IN), .ZN(n2388) );
  XNOR2_X1 U3081 ( .A(n2388), .B(n2387), .ZN(n4510) );
  INV_X1 U3082 ( .A(n4510), .ZN(n2389) );
  MUX2_X1 U3083 ( .A(n2389), .B(DATAI_16_), .S(n3629), .Z(n4110) );
  INV_X1 U3084 ( .A(n4110), .ZN(n3380) );
  OAI22_X1 U3085 ( .A1(n4094), .A2(n2799), .B1(n2243), .B2(n3380), .ZN(n2661)
         );
  NAND2_X1 U3086 ( .A1(n4127), .A2(n2682), .ZN(n2391) );
  NAND2_X1 U3087 ( .A1(n4110), .A2(n2416), .ZN(n2390) );
  NAND2_X1 U3088 ( .A1(n2391), .A2(n2390), .ZN(n2392) );
  XNOR2_X1 U3089 ( .A(n2392), .B(n2782), .ZN(n2660) );
  NAND2_X1 U3090 ( .A1(n3424), .A2(REG0_REG_15__SCAN_IN), .ZN(n2398) );
  NAND2_X1 U3091 ( .A1(n2775), .A2(REG1_REG_15__SCAN_IN), .ZN(n2397) );
  OR2_X1 U3092 ( .A1(n2644), .A2(REG3_REG_15__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3093 ( .A1(n2394), .A2(n2393), .ZN(n4120) );
  INV_X1 U3094 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4121) );
  OR2_X1 U3095 ( .A1(n2895), .A2(n4121), .ZN(n2395) );
  NAND4_X1 U3096 ( .A1(n2398), .A2(n2397), .A3(n2396), .A4(n2395), .ZN(n3764)
         );
  NAND2_X1 U3097 ( .A1(n3764), .A2(n2682), .ZN(n2404) );
  INV_X1 U3098 ( .A(n2399), .ZN(n2400) );
  NAND2_X1 U3099 ( .A1(n2400), .A2(IR_REG_15__SCAN_IN), .ZN(n2402) );
  MUX2_X1 U3100 ( .A(n3839), .B(DATAI_15_), .S(n3629), .Z(n4126) );
  NAND2_X1 U3101 ( .A1(n4126), .A2(n2416), .ZN(n2403) );
  NAND2_X1 U3102 ( .A1(n2404), .A2(n2403), .ZN(n2405) );
  XNOR2_X1 U3103 ( .A(n2405), .B(n2782), .ZN(n2658) );
  NAND2_X1 U3104 ( .A1(n2455), .A2(REG1_REG_1__SCAN_IN), .ZN(n2410) );
  INV_X1 U3105 ( .A(n2434), .ZN(n2406) );
  NAND2_X1 U3106 ( .A1(n2406), .A2(REG3_REG_1__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3107 ( .A1(n2454), .A2(REG0_REG_1__SCAN_IN), .ZN(n2407) );
  INV_X2 U3108 ( .A(n2840), .ZN(n2682) );
  NOR2_X1 U3109 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2442)
         );
  INV_X1 U3110 ( .A(n2442), .ZN(n2411) );
  INV_X1 U3111 ( .A(n3778), .ZN(n3777) );
  NAND2_X1 U3112 ( .A1(n3773), .A2(n2441), .ZN(n2414) );
  NAND2_X1 U3113 ( .A1(n3483), .A2(n2416), .ZN(n2413) );
  XNOR2_X1 U3114 ( .A(n2430), .B(n2429), .ZN(n3479) );
  INV_X1 U3115 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U3116 ( .A1(n2989), .A2(n2416), .ZN(n2426) );
  OAI21_X1 U3117 ( .B1(n2864), .B2(n4558), .A(n2426), .ZN(n2417) );
  INV_X1 U3118 ( .A(n2417), .ZN(n2422) );
  NAND2_X1 U3119 ( .A1(n2455), .A2(REG1_REG_0__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3120 ( .A1(n2454), .A2(REG0_REG_0__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3121 ( .A1(n2422), .A2(n2421), .ZN(n2903) );
  NAND2_X1 U3122 ( .A1(n2984), .A2(n2785), .ZN(n2425) );
  NOR2_X1 U3123 ( .A1(n2864), .A2(n2316), .ZN(n2423) );
  AOI21_X1 U3124 ( .B1(n2989), .B2(n2682), .A(n2423), .ZN(n2424) );
  NAND2_X1 U3125 ( .A1(n2426), .A2(n2797), .ZN(n2427) );
  NAND2_X1 U3126 ( .A1(n2428), .A2(n2427), .ZN(n3480) );
  NAND2_X1 U3127 ( .A1(n3479), .A2(n3480), .ZN(n2433) );
  NAND2_X1 U3128 ( .A1(n2433), .A2(n2432), .ZN(n3007) );
  INV_X1 U3129 ( .A(n3007), .ZN(n2452) );
  INV_X1 U3130 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3046) );
  NAND2_X1 U3131 ( .A1(n2455), .A2(REG1_REG_2__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U3132 ( .A1(n2454), .A2(REG0_REG_2__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U3133 ( .A1(n2436), .A2(n2435), .ZN(n2437) );
  NOR2_X1 U3134 ( .A1(n2438), .A2(n2437), .ZN(n2440) );
  NAND2_X1 U3135 ( .A1(n2447), .A2(n2441), .ZN(n2445) );
  MUX2_X1 U3136 ( .A(n4365), .B(DATAI_2_), .S(n2477), .Z(n3043) );
  NAND2_X1 U3137 ( .A1(n3043), .A2(n2416), .ZN(n2444) );
  NAND2_X1 U3138 ( .A1(n2445), .A2(n2444), .ZN(n2446) );
  XNOR2_X1 U3139 ( .A(n2446), .B(n2797), .ZN(n2449) );
  AOI22_X1 U3140 ( .A1(n2447), .A2(n2785), .B1(n2682), .B2(n3043), .ZN(n2448)
         );
  NAND2_X1 U3141 ( .A1(n2449), .A2(n2448), .ZN(n2453) );
  OR2_X1 U3142 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  NAND2_X1 U3143 ( .A1(n2453), .A2(n2450), .ZN(n3010) );
  INV_X1 U3144 ( .A(n3010), .ZN(n2451) );
  NAND2_X1 U3145 ( .A1(n2452), .A2(n2451), .ZN(n3008) );
  NOR2_X1 U3146 ( .A1(n2076), .A2(n2315), .ZN(n2459) );
  INV_X1 U3147 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U31480 ( .A1(n3543), .A2(n2682), .ZN(n2465) );
  NAND2_X1 U31490 ( .A1(n2460), .A2(IR_REG_31__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U3150 ( .A1(n2462), .A2(n2461), .ZN(n2475) );
  OR2_X1 U3151 ( .A1(n2462), .A2(n2461), .ZN(n2463) );
  MUX2_X1 U3152 ( .A(n4364), .B(DATAI_3_), .S(n2477), .Z(n3102) );
  NAND2_X1 U3153 ( .A1(n3102), .A2(n2416), .ZN(n2464) );
  NAND2_X1 U3154 ( .A1(n2465), .A2(n2464), .ZN(n2466) );
  AOI22_X1 U3155 ( .A1(n3543), .A2(n2785), .B1(n2682), .B2(n3102), .ZN(n2482)
         );
  XNOR2_X1 U3156 ( .A(n2481), .B(n2482), .ZN(n3017) );
  NAND2_X1 U3157 ( .A1(n2455), .A2(REG1_REG_4__SCAN_IN), .ZN(n2468) );
  INV_X1 U3158 ( .A(n2490), .ZN(n2472) );
  INV_X1 U3159 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3160 ( .A1(n2456), .A2(n2470), .ZN(n2471) );
  NAND2_X1 U3161 ( .A1(n2472), .A2(n2471), .ZN(n3545) );
  NAND2_X1 U3162 ( .A1(n3771), .A2(n2682), .ZN(n2479) );
  NAND2_X1 U3163 ( .A1(n2475), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  MUX2_X1 U3164 ( .A(n4390), .B(DATAI_4_), .S(n2477), .Z(n3544) );
  NAND2_X1 U3165 ( .A1(n3544), .A2(n2416), .ZN(n2478) );
  NAND2_X1 U3166 ( .A1(n2479), .A2(n2478), .ZN(n2480) );
  XNOR2_X1 U3167 ( .A(n2480), .B(n2782), .ZN(n2485) );
  AOI22_X1 U3168 ( .A1(n3771), .A2(n2785), .B1(n2682), .B2(n3544), .ZN(n2486)
         );
  XNOR2_X1 U3169 ( .A(n2485), .B(n2486), .ZN(n3540) );
  INV_X1 U3170 ( .A(n2481), .ZN(n2483) );
  NAND2_X1 U3171 ( .A1(n2483), .A2(n2482), .ZN(n3538) );
  AND2_X1 U3172 ( .A1(n3540), .A2(n3538), .ZN(n2484) );
  NAND2_X1 U3173 ( .A1(n3424), .A2(REG0_REG_5__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U3174 ( .A1(n2775), .A2(REG1_REG_5__SCAN_IN), .ZN(n2493) );
  OAI21_X1 U3175 ( .B1(n2490), .B2(REG3_REG_5__SCAN_IN), .A(n2502), .ZN(n3205)
         );
  OR2_X1 U3176 ( .A1(n2895), .A2(n2928), .ZN(n2491) );
  NAND4_X1 U3177 ( .A1(n2494), .A2(n2493), .A3(n2492), .A4(n2491), .ZN(n3542)
         );
  NAND2_X1 U3178 ( .A1(n3542), .A2(n2682), .ZN(n2499) );
  NAND2_X1 U3179 ( .A1(n2495), .A2(IR_REG_31__SCAN_IN), .ZN(n2496) );
  XNOR2_X1 U3180 ( .A(n2496), .B(n2321), .ZN(n2974) );
  INV_X1 U3181 ( .A(DATAI_5_), .ZN(n2497) );
  MUX2_X1 U3182 ( .A(n2974), .B(n2497), .S(n3629), .Z(n3197) );
  NAND2_X1 U3183 ( .A1(n3191), .A2(n2416), .ZN(n2498) );
  NAND2_X1 U3184 ( .A1(n2499), .A2(n2498), .ZN(n2500) );
  XNOR2_X1 U3185 ( .A(n2500), .B(n2782), .ZN(n2516) );
  NOR2_X1 U3186 ( .A1(n3197), .A2(n2243), .ZN(n2501) );
  AOI21_X1 U3187 ( .B1(n3542), .B2(n2785), .A(n2501), .ZN(n2514) );
  XNOR2_X1 U3188 ( .A(n2516), .B(n2514), .ZN(n3063) );
  NAND2_X1 U3189 ( .A1(n3424), .A2(REG0_REG_6__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3190 ( .A1(n2775), .A2(REG1_REG_6__SCAN_IN), .ZN(n2506) );
  AND2_X1 U3191 ( .A1(n2502), .A2(n2933), .ZN(n2503) );
  OR2_X1 U3192 ( .A1(n2503), .A2(n2517), .ZN(n3167) );
  INV_X1 U3193 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3168) );
  OR2_X1 U3194 ( .A1(n2895), .A2(n3168), .ZN(n2504) );
  NAND2_X1 U3195 ( .A1(n3183), .A2(n2441), .ZN(n2510) );
  NOR2_X1 U3196 ( .A1(n2495), .A2(IR_REG_5__SCAN_IN), .ZN(n2524) );
  OR2_X1 U3197 ( .A1(n2524), .A2(n2259), .ZN(n2508) );
  XNOR2_X1 U3198 ( .A(n2508), .B(IR_REG_6__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U3199 ( .A(n4363), .B(DATAI_6_), .S(n3629), .Z(n3159) );
  NAND2_X1 U3200 ( .A1(n3159), .A2(n2416), .ZN(n2509) );
  NAND2_X1 U3201 ( .A1(n2510), .A2(n2509), .ZN(n2511) );
  XNOR2_X1 U3202 ( .A(n2511), .B(n2782), .ZN(n2534) );
  NAND2_X1 U3203 ( .A1(n3183), .A2(n2785), .ZN(n2513) );
  NAND2_X1 U3204 ( .A1(n2513), .A2(n2512), .ZN(n2535) );
  INV_X1 U3205 ( .A(n2514), .ZN(n2515) );
  NAND2_X1 U3206 ( .A1(n2516), .A2(n2515), .ZN(n3122) );
  AND2_X1 U3207 ( .A1(n2062), .A2(n3122), .ZN(n3173) );
  NAND2_X1 U3208 ( .A1(n3424), .A2(REG0_REG_7__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3209 ( .A1(n2775), .A2(REG1_REG_7__SCAN_IN), .ZN(n2521) );
  OR2_X1 U32100 ( .A1(n2517), .A2(REG3_REG_7__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32110 ( .A1(n2542), .A2(n2518), .ZN(n3186) );
  INV_X1 U32120 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2951) );
  OR2_X1 U32130 ( .A1(n2895), .A2(n2951), .ZN(n2519) );
  NAND2_X1 U32140 ( .A1(n3770), .A2(n2682), .ZN(n2527) );
  AND2_X1 U32150 ( .A1(n2524), .A2(n2523), .ZN(n2525) );
  MUX2_X1 U32160 ( .A(n4362), .B(DATAI_7_), .S(n3629), .Z(n3239) );
  NAND2_X1 U32170 ( .A1(n3239), .A2(n2416), .ZN(n2526) );
  NAND2_X1 U32180 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  XNOR2_X1 U32190 ( .A(n2528), .B(n2797), .ZN(n2533) );
  INV_X1 U32200 ( .A(n2533), .ZN(n2530) );
  AOI22_X1 U32210 ( .A1(n3770), .A2(n2785), .B1(n2682), .B2(n3239), .ZN(n2532)
         );
  INV_X1 U32220 ( .A(n2532), .ZN(n2529) );
  NAND2_X1 U32230 ( .A1(n2530), .A2(n2529), .ZN(n2539) );
  AND2_X1 U32240 ( .A1(n3173), .A2(n2539), .ZN(n2531) );
  XNOR2_X1 U32250 ( .A(n2533), .B(n2532), .ZN(n3181) );
  INV_X1 U32260 ( .A(n3181), .ZN(n2538) );
  INV_X1 U32270 ( .A(n2534), .ZN(n2537) );
  INV_X1 U32280 ( .A(n2535), .ZN(n2536) );
  NAND2_X1 U32290 ( .A1(n2537), .A2(n2536), .ZN(n3175) );
  NAND2_X1 U32300 ( .A1(n2538), .A2(n3175), .ZN(n3177) );
  AND2_X1 U32310 ( .A1(n2539), .A2(n3177), .ZN(n2540) );
  NAND2_X1 U32320 ( .A1(n3424), .A2(REG0_REG_8__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32330 ( .A1(n2775), .A2(REG1_REG_8__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32340 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  NAND2_X1 U32350 ( .A1(n2561), .A2(n2543), .ZN(n3258) );
  INV_X1 U32360 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3829) );
  OR2_X1 U32370 ( .A1(n2895), .A2(n3829), .ZN(n2544) );
  NAND4_X1 U32380 ( .A1(n2547), .A2(n2546), .A3(n2545), .A4(n2544), .ZN(n3769)
         );
  NAND2_X1 U32390 ( .A1(n3769), .A2(n2785), .ZN(n2554) );
  NAND2_X1 U32400 ( .A1(n2549), .A2(n2548), .ZN(n2550) );
  NAND2_X1 U32410 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2551) );
  XNOR2_X1 U32420 ( .A(n2551), .B(n2320), .ZN(n3828) );
  INV_X1 U32430 ( .A(DATAI_8_), .ZN(n2552) );
  MUX2_X1 U32440 ( .A(n3828), .B(n2552), .S(n3629), .Z(n3256) );
  NAND2_X1 U32450 ( .A1(n3248), .A2(n2682), .ZN(n2553) );
  NAND2_X1 U32460 ( .A1(n2554), .A2(n2553), .ZN(n3210) );
  NAND2_X1 U32470 ( .A1(n3769), .A2(n2682), .ZN(n2556) );
  NAND2_X1 U32480 ( .A1(n3248), .A2(n2416), .ZN(n2555) );
  NAND2_X1 U32490 ( .A1(n2556), .A2(n2555), .ZN(n2557) );
  XNOR2_X1 U32500 ( .A(n2557), .B(n2782), .ZN(n3211) );
  OAI21_X1 U32510 ( .B1(n3213), .B2(n3210), .A(n3211), .ZN(n2559) );
  NAND2_X1 U32520 ( .A1(n3213), .A2(n3210), .ZN(n2558) );
  NAND2_X1 U32530 ( .A1(n3424), .A2(REG0_REG_9__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U32540 ( .A1(n2775), .A2(REG1_REG_9__SCAN_IN), .ZN(n2565) );
  AND2_X1 U32550 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  OR2_X1 U32560 ( .A1(n2562), .A2(n2572), .ZN(n3269) );
  INV_X1 U32570 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3237) );
  OR2_X1 U32580 ( .A1(n2895), .A2(n3237), .ZN(n2563) );
  NAND4_X1 U32590 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n3768)
         );
  NAND2_X1 U32600 ( .A1(n3768), .A2(n2441), .ZN(n2570) );
  NAND2_X1 U32610 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  XNOR2_X1 U32620 ( .A(n2568), .B(IR_REG_9__SCAN_IN), .ZN(n3825) );
  MUX2_X1 U32630 ( .A(n3825), .B(DATAI_9_), .S(n3629), .Z(n3303) );
  NAND2_X1 U32640 ( .A1(n3303), .A2(n2416), .ZN(n2569) );
  NAND2_X1 U32650 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  XNOR2_X1 U32660 ( .A(n2571), .B(n2797), .ZN(n2585) );
  AOI22_X1 U32670 ( .A1(n3768), .A2(n2785), .B1(n2682), .B2(n3303), .ZN(n2584)
         );
  XNOR2_X1 U32680 ( .A(n2585), .B(n2584), .ZN(n3266) );
  NAND2_X1 U32690 ( .A1(n2775), .A2(REG1_REG_10__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32700 ( .A1(n3424), .A2(REG0_REG_10__SCAN_IN), .ZN(n2577) );
  NOR2_X1 U32710 ( .A1(n2572), .A2(REG3_REG_10__SCAN_IN), .ZN(n2573) );
  OR2_X1 U32720 ( .A1(n2590), .A2(n2573), .ZN(n4495) );
  INV_X1 U32730 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2574) );
  OR2_X1 U32740 ( .A1(n2895), .A2(n2574), .ZN(n2575) );
  NAND4_X1 U32750 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(n3767)
         );
  NAND2_X1 U32760 ( .A1(n3767), .A2(n2682), .ZN(n2582) );
  NAND2_X1 U32770 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2580) );
  XNOR2_X1 U32780 ( .A(n2580), .B(IR_REG_10__SCAN_IN), .ZN(n3830) );
  MUX2_X1 U32790 ( .A(n3830), .B(DATAI_10_), .S(n3629), .Z(n3466) );
  NAND2_X1 U32800 ( .A1(n3466), .A2(n2416), .ZN(n2581) );
  NAND2_X1 U32810 ( .A1(n2582), .A2(n2581), .ZN(n2583) );
  XNOR2_X1 U32820 ( .A(n2583), .B(n2782), .ZN(n2589) );
  AOI22_X1 U32830 ( .A1(n3767), .A2(n2785), .B1(n2682), .B2(n3466), .ZN(n2587)
         );
  XNOR2_X1 U32840 ( .A(n2589), .B(n2587), .ZN(n3463) );
  NAND2_X1 U32850 ( .A1(n2585), .A2(n2584), .ZN(n3461) );
  AND2_X1 U32860 ( .A1(n3463), .A2(n3461), .ZN(n2586) );
  INV_X1 U32870 ( .A(n2587), .ZN(n2588) );
  NAND2_X1 U32880 ( .A1(n3424), .A2(REG0_REG_11__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U32890 ( .A1(n2775), .A2(REG1_REG_11__SCAN_IN), .ZN(n2594) );
  OR2_X1 U32900 ( .A1(n2590), .A2(REG3_REG_11__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U32910 ( .A1(n2605), .A2(n2591), .ZN(n3316) );
  INV_X1 U32920 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3317) );
  OR2_X1 U32930 ( .A1(n2895), .A2(n3317), .ZN(n2592) );
  NAND4_X1 U32940 ( .A1(n2595), .A2(n2594), .A3(n2593), .A4(n2592), .ZN(n3766)
         );
  NAND2_X1 U32950 ( .A1(n3766), .A2(n2441), .ZN(n2598) );
  OR2_X1 U32960 ( .A1(n2596), .A2(n2259), .ZN(n2612) );
  XNOR2_X1 U32970 ( .A(n2612), .B(IR_REG_11__SCAN_IN), .ZN(n3824) );
  MUX2_X1 U32980 ( .A(n3824), .B(DATAI_11_), .S(n3629), .Z(n3309) );
  NAND2_X1 U32990 ( .A1(n3309), .A2(n2416), .ZN(n2597) );
  NAND2_X1 U33000 ( .A1(n2598), .A2(n2597), .ZN(n2599) );
  XNOR2_X1 U33010 ( .A(n2599), .B(n2797), .ZN(n2600) );
  AOI22_X1 U33020 ( .A1(n3766), .A2(n2785), .B1(n2682), .B2(n3309), .ZN(n2601)
         );
  NAND2_X1 U33030 ( .A1(n2600), .A2(n2601), .ZN(n3273) );
  INV_X1 U33040 ( .A(n2600), .ZN(n2603) );
  INV_X1 U33050 ( .A(n2601), .ZN(n2602) );
  NAND2_X1 U33060 ( .A1(n2603), .A2(n2602), .ZN(n3274) );
  NAND2_X1 U33070 ( .A1(n3424), .A2(REG0_REG_12__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U33080 ( .A1(n2775), .A2(REG1_REG_12__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U33090 ( .A1(n2605), .A2(n2604), .ZN(n2606) );
  NAND2_X1 U33100 ( .A1(n2620), .A2(n2606), .ZN(n3331) );
  INV_X1 U33110 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3332) );
  OR2_X1 U33120 ( .A1(n2895), .A2(n3332), .ZN(n2607) );
  NAND4_X1 U33130 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(n3765)
         );
  NAND2_X1 U33140 ( .A1(n3765), .A2(n2682), .ZN(n2616) );
  INV_X1 U33150 ( .A(IR_REG_11__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U33160 ( .A1(n2612), .A2(n2611), .ZN(n2613) );
  NAND2_X1 U33170 ( .A1(n2613), .A2(IR_REG_31__SCAN_IN), .ZN(n2614) );
  XNOR2_X1 U33180 ( .A(n2614), .B(IR_REG_12__SCAN_IN), .ZN(n3834) );
  INV_X1 U33190 ( .A(DATAI_12_), .ZN(n4515) );
  MUX2_X1 U33200 ( .A(n4516), .B(n4515), .S(n3629), .Z(n3374) );
  NAND2_X1 U33210 ( .A1(n3376), .A2(n2416), .ZN(n2615) );
  NAND2_X1 U33220 ( .A1(n2616), .A2(n2615), .ZN(n2617) );
  XNOR2_X1 U33230 ( .A(n2617), .B(n2797), .ZN(n3347) );
  NAND2_X1 U33240 ( .A1(n3765), .A2(n2785), .ZN(n2619) );
  NAND2_X1 U33250 ( .A1(n3376), .A2(n2682), .ZN(n2618) );
  NAND2_X1 U33260 ( .A1(n3424), .A2(REG0_REG_13__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U33270 ( .A1(n2775), .A2(REG1_REG_13__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U33280 ( .A1(n2620), .A2(n3355), .ZN(n2621) );
  NAND2_X1 U33290 ( .A1(n2643), .A2(n2621), .ZN(n4181) );
  INV_X1 U33300 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4182) );
  OR2_X1 U33310 ( .A1(n2895), .A2(n4182), .ZN(n2622) );
  NAND4_X1 U33320 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n4142)
         );
  NAND2_X1 U33330 ( .A1(n4142), .A2(n2682), .ZN(n2630) );
  NAND2_X1 U33340 ( .A1(n2626), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  XNOR2_X1 U33350 ( .A(n2627), .B(IR_REG_13__SCAN_IN), .ZN(n3837) );
  INV_X1 U33360 ( .A(DATAI_13_), .ZN(n2628) );
  MUX2_X1 U33370 ( .A(n4514), .B(n2628), .S(n3629), .Z(n4178) );
  NAND2_X1 U33380 ( .A1(n4165), .A2(n2416), .ZN(n2629) );
  NAND2_X1 U33390 ( .A1(n2630), .A2(n2629), .ZN(n2631) );
  XNOR2_X1 U33400 ( .A(n2631), .B(n2782), .ZN(n2635) );
  NAND2_X1 U33410 ( .A1(n4142), .A2(n2785), .ZN(n2633) );
  NAND2_X1 U33420 ( .A1(n4165), .A2(n2682), .ZN(n2632) );
  NAND2_X1 U33430 ( .A1(n2633), .A2(n2632), .ZN(n2636) );
  NAND2_X1 U33440 ( .A1(n2635), .A2(n2636), .ZN(n3352) );
  OAI21_X1 U33450 ( .B1(n3347), .B2(n3349), .A(n3352), .ZN(n2634) );
  NAND3_X1 U33460 ( .A1(n3352), .A2(n3349), .A3(n3347), .ZN(n2639) );
  INV_X1 U33470 ( .A(n2635), .ZN(n2638) );
  INV_X1 U33480 ( .A(n2636), .ZN(n2637) );
  NAND2_X1 U33490 ( .A1(n2638), .A2(n2637), .ZN(n3351) );
  AND2_X1 U33500 ( .A1(n2639), .A2(n3351), .ZN(n2640) );
  NAND2_X1 U33510 ( .A1(n3424), .A2(REG0_REG_14__SCAN_IN), .ZN(n2649) );
  NAND2_X1 U33520 ( .A1(n2775), .A2(REG1_REG_14__SCAN_IN), .ZN(n2648) );
  AND2_X1 U3353 ( .A1(n2643), .A2(n2642), .ZN(n2645) );
  OR2_X1 U33540 ( .A1(n2645), .A2(n2644), .ZN(n4152) );
  INV_X1 U3355 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4153) );
  OR2_X1 U3356 ( .A1(n2895), .A2(n4153), .ZN(n2646) );
  NAND4_X1 U3357 ( .A1(n2649), .A2(n2648), .A3(n2647), .A4(n2646), .ZN(n4167)
         );
  NAND2_X1 U3358 ( .A1(n4167), .A2(n2441), .ZN(n2653) );
  NAND2_X1 U3359 ( .A1(n2650), .A2(IR_REG_31__SCAN_IN), .ZN(n2651) );
  XNOR2_X1 U3360 ( .A(n2651), .B(IR_REG_14__SCAN_IN), .ZN(n4448) );
  MUX2_X1 U3361 ( .A(n4448), .B(DATAI_14_), .S(n3629), .Z(n4148) );
  NAND2_X1 U3362 ( .A1(n4148), .A2(n2416), .ZN(n2652) );
  NAND2_X1 U3363 ( .A1(n2653), .A2(n2652), .ZN(n2654) );
  XNOR2_X1 U3364 ( .A(n2654), .B(n2797), .ZN(n3338) );
  NAND2_X1 U3365 ( .A1(n4167), .A2(n2785), .ZN(n2656) );
  NAND2_X1 U3366 ( .A1(n4148), .A2(n2441), .ZN(n2655) );
  NAND2_X1 U3367 ( .A1(n2656), .A2(n2655), .ZN(n3337) );
  NOR2_X1 U3368 ( .A1(n2658), .A2(n2659), .ZN(n3598) );
  AOI21_X1 U3369 ( .B1(n3764), .B2(n2785), .A(n2657), .ZN(n3599) );
  XOR2_X1 U3370 ( .A(n2661), .B(n2660), .Z(n3510) );
  NAND2_X1 U3371 ( .A1(n2659), .A2(n2658), .ZN(n3596) );
  NAND2_X1 U3372 ( .A1(n3424), .A2(REG0_REG_18__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3373 ( .A1(n2775), .A2(REG1_REG_18__SCAN_IN), .ZN(n2668) );
  NOR2_X1 U3374 ( .A1(n2664), .A2(REG3_REG_18__SCAN_IN), .ZN(n2665) );
  OR2_X1 U3375 ( .A1(n2676), .A2(n2665), .ZN(n4068) );
  OR2_X1 U3376 ( .A1(n2790), .A2(n4068), .ZN(n2667) );
  INV_X1 U3377 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4069) );
  OR2_X1 U3378 ( .A1(n2895), .A2(n4069), .ZN(n2666) );
  NAND4_X1 U3379 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .ZN(n4091)
         );
  NAND2_X1 U3380 ( .A1(n2359), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  XNOR2_X1 U3381 ( .A(n2670), .B(IR_REG_18__SCAN_IN), .ZN(n3856) );
  MUX2_X1 U3382 ( .A(n3856), .B(DATAI_18_), .S(n3629), .Z(n4072) );
  NAND2_X1 U3383 ( .A1(n4072), .A2(n2416), .ZN(n2671) );
  NAND2_X1 U3384 ( .A1(n2672), .A2(n2671), .ZN(n2673) );
  XNOR2_X1 U3385 ( .A(n2673), .B(n2797), .ZN(n2675) );
  AOI22_X1 U3386 ( .A1(n4091), .A2(n2785), .B1(n2682), .B2(n4072), .ZN(n2674)
         );
  OR2_X1 U3387 ( .A1(n2675), .A2(n2674), .ZN(n3579) );
  AND2_X1 U3388 ( .A1(n2675), .A2(n2674), .ZN(n3580) );
  AOI21_X1 U3389 ( .B1(n3583), .B2(n3579), .A(n3580), .ZN(n3472) );
  NAND2_X1 U3390 ( .A1(n3424), .A2(REG0_REG_19__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3391 ( .A1(n2775), .A2(REG1_REG_19__SCAN_IN), .ZN(n2680) );
  OR2_X1 U3392 ( .A1(n2676), .A2(REG3_REG_19__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3393 ( .A1(n2689), .A2(n2677), .ZN(n4047) );
  INV_X1 U3394 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4059) );
  OR2_X1 U3395 ( .A1(n2895), .A2(n4059), .ZN(n2678) );
  NAND4_X1 U3396 ( .A1(n2681), .A2(n2680), .A3(n2679), .A4(n2678), .ZN(n4073)
         );
  MUX2_X1 U3397 ( .A(n3850), .B(DATAI_19_), .S(n3629), .Z(n4053) );
  AOI22_X1 U3398 ( .A1(n4073), .A2(n2785), .B1(n2682), .B2(n4053), .ZN(n2686)
         );
  NAND2_X1 U3399 ( .A1(n4053), .A2(n2416), .ZN(n2683) );
  NAND2_X1 U3400 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  XNOR2_X1 U3401 ( .A(n2685), .B(n2782), .ZN(n2688) );
  XOR2_X1 U3402 ( .A(n2686), .B(n2688), .Z(n3471) );
  INV_X1 U3403 ( .A(n2686), .ZN(n2687) );
  NAND2_X1 U3404 ( .A1(n3424), .A2(REG0_REG_20__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3405 ( .A1(n2775), .A2(REG1_REG_20__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3406 ( .A1(n2689), .A2(n3556), .ZN(n2690) );
  NAND2_X1 U3407 ( .A1(n2705), .A2(n2690), .ZN(n4037) );
  OR2_X1 U3408 ( .A1(n2790), .A2(n4037), .ZN(n2692) );
  INV_X1 U3409 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4038) );
  OR2_X1 U3410 ( .A1(n2895), .A2(n4038), .ZN(n2691) );
  NAND2_X1 U3411 ( .A1(n3558), .A2(n2416), .ZN(n2695) );
  NAND2_X1 U3412 ( .A1(n2696), .A2(n2695), .ZN(n2697) );
  XNOR2_X1 U3413 ( .A(n2697), .B(n2782), .ZN(n2700) );
  NAND2_X1 U3414 ( .A1(n4054), .A2(n2785), .ZN(n2699) );
  NAND2_X1 U3415 ( .A1(n2699), .A2(n2698), .ZN(n2701) );
  NAND2_X1 U3416 ( .A1(n2700), .A2(n2701), .ZN(n3552) );
  INV_X1 U3417 ( .A(n2700), .ZN(n2703) );
  INV_X1 U3418 ( .A(n2701), .ZN(n2702) );
  NAND2_X1 U3419 ( .A1(n2703), .A2(n2702), .ZN(n3554) );
  INV_X1 U3420 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2704) );
  AND2_X1 U3421 ( .A1(n2705), .A2(n2704), .ZN(n2706) );
  NOR2_X1 U3422 ( .A1(n2718), .A2(n2706), .ZN(n3492) );
  NAND2_X1 U3423 ( .A1(n2406), .A2(n3492), .ZN(n2710) );
  NAND2_X1 U3424 ( .A1(n3424), .A2(REG0_REG_21__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U3425 ( .A1(n2775), .A2(REG1_REG_21__SCAN_IN), .ZN(n2708) );
  INV_X1 U3426 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4013) );
  OR2_X1 U3427 ( .A1(n2895), .A2(n4013), .ZN(n2707) );
  NAND4_X1 U3428 ( .A1(n2710), .A2(n2709), .A3(n2708), .A4(n2707), .ZN(n3763)
         );
  NAND2_X1 U3429 ( .A1(n3629), .A2(DATAI_21_), .ZN(n3416) );
  NAND2_X1 U3430 ( .A1(n4009), .A2(n2416), .ZN(n2711) );
  NAND2_X1 U3431 ( .A1(n2712), .A2(n2711), .ZN(n2713) );
  XNOR2_X1 U3432 ( .A(n2713), .B(n2782), .ZN(n3489) );
  NAND2_X1 U3433 ( .A1(n3763), .A2(n2785), .ZN(n2715) );
  NAND2_X1 U3434 ( .A1(n2715), .A2(n2714), .ZN(n2716) );
  NOR2_X1 U3435 ( .A1(n3489), .A2(n2716), .ZN(n2717) );
  INV_X1 U3436 ( .A(n2716), .ZN(n3488) );
  NAND2_X1 U3437 ( .A1(n2775), .A2(REG1_REG_22__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3438 ( .A1(n3424), .A2(REG0_REG_22__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U3439 ( .A1(n2718), .A2(REG3_REG_22__SCAN_IN), .ZN(n2728) );
  OR2_X1 U3440 ( .A1(n2718), .A2(REG3_REG_22__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U3441 ( .A1(n2728), .A2(n2719), .ZN(n3991) );
  OR2_X1 U3442 ( .A1(n3991), .A2(n2790), .ZN(n2721) );
  INV_X1 U3443 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3992) );
  OR2_X1 U3444 ( .A1(n2895), .A2(n3992), .ZN(n2720) );
  OAI22_X1 U3445 ( .A1(n4002), .A2(n2243), .B1(n2796), .B2(n3569), .ZN(n2724)
         );
  XNOR2_X1 U3446 ( .A(n2724), .B(n2782), .ZN(n2726) );
  OAI22_X1 U3447 ( .A1(n4002), .A2(n2799), .B1(n2243), .B2(n3569), .ZN(n2725)
         );
  XNOR2_X1 U3448 ( .A(n2726), .B(n2725), .ZN(n3566) );
  NOR2_X1 U3449 ( .A1(n2726), .A2(n2725), .ZN(n3455) );
  INV_X1 U3450 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U3451 ( .A1(n2728), .A2(n2727), .ZN(n2729) );
  NAND2_X1 U3452 ( .A1(n2740), .A2(n2729), .ZN(n3962) );
  NAND2_X1 U3453 ( .A1(n3424), .A2(REG0_REG_23__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U3454 ( .A1(n2775), .A2(REG1_REG_23__SCAN_IN), .ZN(n2731) );
  INV_X1 U3455 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3979) );
  OR2_X1 U3456 ( .A1(n2895), .A2(n3979), .ZN(n2730) );
  NAND2_X1 U3457 ( .A1(n3629), .A2(DATAI_23_), .ZN(n3975) );
  INV_X1 U34580 ( .A(n3975), .ZN(n3961) );
  NAND2_X1 U34590 ( .A1(n3961), .A2(n2416), .ZN(n2734) );
  NAND2_X1 U3460 ( .A1(n2735), .A2(n2734), .ZN(n2736) );
  XNOR2_X1 U3461 ( .A(n2736), .B(n2797), .ZN(n2739) );
  NOR2_X1 U3462 ( .A1(n3975), .A2(n2243), .ZN(n2737) );
  AOI21_X1 U3463 ( .B1(n3987), .B2(n2785), .A(n2737), .ZN(n2738) );
  XNOR2_X1 U3464 ( .A(n2739), .B(n2738), .ZN(n3454) );
  NOR2_X1 U3465 ( .A1(n2739), .A2(n2738), .ZN(n2748) );
  INV_X1 U3466 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U34670 ( .A1(n2740), .A2(n3533), .ZN(n2741) );
  NAND2_X1 U3468 ( .A1(n2749), .A2(n2741), .ZN(n3949) );
  AOI22_X1 U34690 ( .A1(n3424), .A2(REG0_REG_24__SCAN_IN), .B1(n2775), .B2(
        REG1_REG_24__SCAN_IN), .ZN(n2743) );
  INV_X1 U3470 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3950) );
  OR2_X1 U34710 ( .A1(n2895), .A2(n3950), .ZN(n2742) );
  NAND2_X1 U3472 ( .A1(n3973), .A2(n2785), .ZN(n2745) );
  NAND2_X1 U34730 ( .A1(n3629), .A2(DATAI_24_), .ZN(n3951) );
  INV_X1 U3474 ( .A(n3951), .ZN(n3530) );
  NAND2_X1 U34750 ( .A1(n2745), .A2(n2744), .ZN(n2747) );
  AOI22_X1 U3476 ( .A1(n3973), .A2(n2441), .B1(n2416), .B2(n3530), .ZN(n2746)
         );
  XNOR2_X1 U34770 ( .A(n2746), .B(n2782), .ZN(n3528) );
  OAI21_X1 U3478 ( .B1(n3453), .B2(n2748), .A(n2747), .ZN(n3525) );
  INV_X1 U34790 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3503) );
  AND2_X1 U3480 ( .A1(n2749), .A2(n3503), .ZN(n2750) );
  OR2_X1 U34810 ( .A1(n2750), .A2(n2759), .ZN(n3502) );
  AOI22_X1 U3482 ( .A1(n3424), .A2(REG0_REG_25__SCAN_IN), .B1(n2775), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n2752) );
  INV_X1 U34830 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3936) );
  OR2_X1 U3484 ( .A1(n2895), .A2(n3936), .ZN(n2751) );
  INV_X1 U34850 ( .A(n3926), .ZN(n3924) );
  NAND2_X1 U3486 ( .A1(n3924), .A2(n2416), .ZN(n2753) );
  NAND2_X1 U34870 ( .A1(n2754), .A2(n2753), .ZN(n2755) );
  XNOR2_X1 U3488 ( .A(n2755), .B(n2797), .ZN(n2758) );
  NOR2_X1 U34890 ( .A1(n3926), .A2(n2243), .ZN(n2756) );
  AOI21_X1 U3490 ( .B1(n3946), .B2(n2785), .A(n2756), .ZN(n2757) );
  NAND2_X1 U34910 ( .A1(n2758), .A2(n2757), .ZN(n3498) );
  NOR2_X1 U3492 ( .A1(n2758), .A2(n2757), .ZN(n3499) );
  NOR2_X1 U34930 ( .A1(n2759), .A2(REG3_REG_26__SCAN_IN), .ZN(n2760) );
  INV_X1 U3494 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U34950 ( .A1(n3424), .A2(REG0_REG_26__SCAN_IN), .ZN(n2762) );
  NAND2_X1 U3496 ( .A1(n2775), .A2(REG1_REG_26__SCAN_IN), .ZN(n2761) );
  OAI211_X1 U34970 ( .C1(n3911), .C2(n2895), .A(n2762), .B(n2761), .ZN(n2763)
         );
  INV_X1 U3498 ( .A(n2763), .ZN(n2764) );
  NAND2_X1 U34990 ( .A1(n3629), .A2(DATAI_26_), .ZN(n3905) );
  NAND2_X1 U3500 ( .A1(n3913), .A2(n2416), .ZN(n2765) );
  NAND2_X1 U35010 ( .A1(n2766), .A2(n2765), .ZN(n2767) );
  XNOR2_X1 U3502 ( .A(n2767), .B(n2797), .ZN(n2772) );
  INV_X1 U35030 ( .A(n2772), .ZN(n2770) );
  NOR2_X1 U3504 ( .A1(n3905), .A2(n2243), .ZN(n2768) );
  AOI21_X1 U35050 ( .B1(n3935), .B2(n2785), .A(n2768), .ZN(n2771) );
  INV_X1 U35060 ( .A(n2771), .ZN(n2769) );
  NAND2_X1 U35070 ( .A1(n2770), .A2(n2769), .ZN(n3589) );
  AND2_X1 U35080 ( .A1(n2772), .A2(n2771), .ZN(n3590) );
  NOR2_X1 U35090 ( .A1(n2773), .A2(REG3_REG_27__SCAN_IN), .ZN(n2774) );
  INV_X1 U35100 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3886) );
  NAND2_X1 U35110 ( .A1(n3424), .A2(REG0_REG_27__SCAN_IN), .ZN(n2777) );
  NAND2_X1 U35120 ( .A1(n2775), .A2(REG1_REG_27__SCAN_IN), .ZN(n2776) );
  OAI211_X1 U35130 ( .C1(n3886), .C2(n2895), .A(n2777), .B(n2776), .ZN(n2778)
         );
  INV_X1 U35140 ( .A(n2778), .ZN(n2779) );
  OAI21_X2 U35150 ( .B1(n3887), .B2(n2790), .A(n2779), .ZN(n3908) );
  NAND2_X1 U35160 ( .A1(n3908), .A2(n2682), .ZN(n2781) );
  NAND2_X1 U35170 ( .A1(n3629), .A2(DATAI_27_), .ZN(n3893) );
  NAND2_X1 U35180 ( .A1(n3883), .A2(n2416), .ZN(n2780) );
  NAND2_X1 U35190 ( .A1(n2781), .A2(n2780), .ZN(n2783) );
  XNOR2_X1 U35200 ( .A(n2783), .B(n2782), .ZN(n2828) );
  NOR2_X1 U35210 ( .A1(n3893), .A2(n2243), .ZN(n2784) );
  AOI21_X1 U35220 ( .B1(n3908), .B2(n2785), .A(n2784), .ZN(n2826) );
  XNOR2_X1 U35230 ( .A(n2828), .B(n2826), .ZN(n3446) );
  NAND2_X1 U35240 ( .A1(n2786), .A2(REG3_REG_28__SCAN_IN), .ZN(n3440) );
  INV_X1 U35250 ( .A(n2786), .ZN(n2788) );
  INV_X1 U35260 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U35270 ( .A1(n2788), .A2(n2787), .ZN(n2789) );
  NAND2_X1 U35280 ( .A1(n3440), .A2(n2789), .ZN(n3869) );
  INV_X1 U35290 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3879) );
  NAND2_X1 U35300 ( .A1(n3424), .A2(REG0_REG_28__SCAN_IN), .ZN(n2792) );
  NAND2_X1 U35310 ( .A1(n2775), .A2(REG1_REG_28__SCAN_IN), .ZN(n2791) );
  OAI211_X1 U35320 ( .C1(n3879), .C2(n2895), .A(n2792), .B(n2791), .ZN(n2793)
         );
  INV_X1 U35330 ( .A(n2793), .ZN(n2794) );
  OAI22_X1 U35340 ( .A1(n3394), .A2(n2243), .B1(n2796), .B2(n3876), .ZN(n2798)
         );
  XNOR2_X1 U35350 ( .A(n2798), .B(n2797), .ZN(n2801) );
  OAI22_X1 U35360 ( .A1(n3394), .A2(n2799), .B1(n2243), .B2(n3876), .ZN(n2800)
         );
  XNOR2_X1 U35370 ( .A(n2801), .B(n2800), .ZN(n2830) );
  INV_X1 U35380 ( .A(n2830), .ZN(n2824) );
  NAND2_X1 U35390 ( .A1(n2876), .A2(B_REG_SCAN_IN), .ZN(n2802) );
  MUX2_X1 U35400 ( .A(n2802), .B(B_REG_SCAN_IN), .S(n2198), .Z(n2803) );
  INV_X1 U35410 ( .A(n4360), .ZN(n2815) );
  NAND2_X1 U35420 ( .A1(n2815), .A2(n2804), .ZN(n2888) );
  INV_X1 U35430 ( .A(n3031), .ZN(n3056) );
  INV_X1 U35440 ( .A(n3000), .ZN(n2817) );
  NOR4_X1 U35450 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2808) );
  NOR4_X1 U35460 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2807) );
  NOR4_X1 U35470 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2806) );
  NOR4_X1 U35480 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2805) );
  NAND4_X1 U35490 ( .A1(n2808), .A2(n2807), .A3(n2806), .A4(n2805), .ZN(n2814)
         );
  NOR2_X1 U35500 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_9__SCAN_IN), .ZN(n2812)
         );
  NOR4_X1 U35510 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2811) );
  NOR4_X1 U35520 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2810) );
  NOR4_X1 U35530 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2809) );
  NAND4_X1 U35540 ( .A1(n2812), .A2(n2811), .A3(n2810), .A4(n2809), .ZN(n2813)
         );
  NOR2_X1 U35550 ( .A1(n2814), .A2(n2813), .ZN(n2998) );
  NAND2_X1 U35560 ( .A1(n2998), .A2(D_REG_1__SCAN_IN), .ZN(n2816) );
  NAND2_X1 U35570 ( .A1(n2815), .A2(n2876), .ZN(n2999) );
  INV_X1 U35580 ( .A(n2999), .ZN(n2890) );
  AOI21_X1 U35590 ( .B1(n2817), .B2(n2816), .A(n2890), .ZN(n3033) );
  OR2_X1 U35600 ( .A1(n2819), .A2(n2818), .ZN(n2820) );
  NAND2_X1 U35610 ( .A1(n2374), .A2(n3860), .ZN(n2833) );
  NAND2_X1 U35620 ( .A1(n2833), .A2(n3085), .ZN(n2822) );
  INV_X1 U35630 ( .A(n2988), .ZN(n2987) );
  NAND2_X1 U35640 ( .A1(n2822), .A2(n2987), .ZN(n2831) );
  OR2_X1 U35650 ( .A1(n3002), .A2(n2831), .ZN(n2823) );
  NAND2_X1 U35660 ( .A1(n2824), .A2(n3609), .ZN(n2825) );
  INV_X1 U35670 ( .A(n2826), .ZN(n2827) );
  NAND2_X1 U35680 ( .A1(n2828), .A2(n2827), .ZN(n2829) );
  NOR3_X1 U35690 ( .A1(n2830), .A2(n3577), .A3(n2829), .ZN(n2859) );
  INV_X1 U35700 ( .A(n2374), .ZN(n4361) );
  NAND2_X1 U35710 ( .A1(n2831), .A2(n4200), .ZN(n2832) );
  NAND2_X1 U35720 ( .A1(n2854), .A2(n2832), .ZN(n2835) );
  INV_X1 U35730 ( .A(n3001), .ZN(n2834) );
  NAND2_X1 U35740 ( .A1(n2835), .A2(n2834), .ZN(n2907) );
  NAND2_X1 U35750 ( .A1(n2864), .A2(n2922), .ZN(n2836) );
  OAI21_X1 U35760 ( .B1(n2907), .B2(n2836), .A(STATE_REG_SCAN_IN), .ZN(n2842)
         );
  INV_X1 U35770 ( .A(n2837), .ZN(n2838) );
  NAND2_X1 U35780 ( .A1(n2838), .A2(n4506), .ZN(n2839) );
  INV_X1 U35790 ( .A(n3755), .ZN(n2841) );
  NAND2_X1 U35800 ( .A1(n2854), .A2(n2841), .ZN(n2905) );
  OR2_X1 U35810 ( .A1(n2843), .A2(n2259), .ZN(n2844) );
  NOR2_X1 U3582 ( .A1(n3755), .A2(n4367), .ZN(n2845) );
  AND2_X2 U3583 ( .A1(n2852), .A2(n2845), .ZN(n3603) );
  AOI22_X1 U3584 ( .A1(n3908), .A2(n3603), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2857) );
  INV_X1 U3585 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4578) );
  NAND2_X1 U3586 ( .A1(n2467), .A2(REG2_REG_29__SCAN_IN), .ZN(n2847) );
  INV_X1 U3587 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4724) );
  OR2_X1 U3588 ( .A1(n2489), .A2(n4724), .ZN(n2846) );
  OAI211_X1 U3589 ( .C1(n2848), .C2(n4578), .A(n2847), .B(n2846), .ZN(n2849)
         );
  INV_X1 U3590 ( .A(n2849), .ZN(n2850) );
  NAND2_X1 U3591 ( .A1(n2050), .A2(n2850), .ZN(n3873) );
  INV_X1 U3592 ( .A(n4367), .ZN(n3799) );
  NOR2_X1 U3593 ( .A1(n3755), .A2(n3799), .ZN(n2851) );
  AND2_X2 U3594 ( .A1(n2852), .A2(n2851), .ZN(n3602) );
  OR2_X1 U3595 ( .A1(n3002), .A2(n4200), .ZN(n2853) );
  OR2_X1 U3596 ( .A1(n2854), .A2(n2853), .ZN(n2855) );
  NAND2_X1 U3597 ( .A1(n2374), .A2(n3850), .ZN(n3090) );
  AOI22_X1 U3598 ( .A1(n3873), .A2(n3602), .B1(n3868), .B2(n3604), .ZN(n2856)
         );
  OAI211_X1 U3599 ( .C1(n3607), .C2(n3869), .A(n2857), .B(n2856), .ZN(n2858)
         );
  AOI21_X1 U3600 ( .B1(n2860), .B2(n2047), .A(n2074), .ZN(n2861) );
  NAND2_X1 U3601 ( .A1(n2862), .A2(n2861), .ZN(U3217) );
  INV_X1 U3602 ( .A(n4506), .ZN(n2863) );
  MUX2_X1 U3603 ( .A(n2974), .B(n2497), .S(U3149), .Z(n2865) );
  INV_X1 U3604 ( .A(n2865), .ZN(U3347) );
  INV_X1 U3605 ( .A(DATAI_1_), .ZN(n2866) );
  MUX2_X1 U3606 ( .A(n3778), .B(n2866), .S(U3149), .Z(n2867) );
  INV_X1 U3607 ( .A(n2867), .ZN(U3351) );
  MUX2_X1 U3608 ( .A(n3828), .B(n2552), .S(U3149), .Z(n2868) );
  INV_X1 U3609 ( .A(n2868), .ZN(U3344) );
  INV_X1 U3610 ( .A(DATAI_21_), .ZN(n2870) );
  NAND2_X1 U3611 ( .A1(n3652), .A2(STATE_REG_SCAN_IN), .ZN(n2869) );
  OAI21_X1 U3612 ( .B1(STATE_REG_SCAN_IN), .B2(n2870), .A(n2869), .ZN(U3331)
         );
  INV_X1 U3613 ( .A(n3823), .ZN(n3855) );
  NAND2_X1 U3614 ( .A1(n3855), .A2(STATE_REG_SCAN_IN), .ZN(n2871) );
  OAI21_X1 U3615 ( .B1(STATE_REG_SCAN_IN), .B2(n2365), .A(n2871), .ZN(U3335)
         );
  INV_X1 U3616 ( .A(DATAI_22_), .ZN(n2873) );
  NAND2_X1 U3617 ( .A1(n3756), .A2(STATE_REG_SCAN_IN), .ZN(n2872) );
  OAI21_X1 U3618 ( .B1(STATE_REG_SCAN_IN), .B2(n2873), .A(n2872), .ZN(U3330)
         );
  INV_X1 U3619 ( .A(DATAI_19_), .ZN(n2874) );
  MUX2_X1 U3620 ( .A(n2874), .B(n3860), .S(STATE_REG_SCAN_IN), .Z(n2875) );
  INV_X1 U3621 ( .A(n2875), .ZN(U3333) );
  INV_X1 U3622 ( .A(DATAI_25_), .ZN(n2878) );
  NAND2_X1 U3623 ( .A1(n2197), .A2(STATE_REG_SCAN_IN), .ZN(n2877) );
  OAI21_X1 U3624 ( .B1(STATE_REG_SCAN_IN), .B2(n2878), .A(n2877), .ZN(U3327)
         );
  INV_X1 U3625 ( .A(DATAI_27_), .ZN(n2881) );
  XNOR2_X1 U3626 ( .A(n2879), .B(IR_REG_27__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U3627 ( .A1(n4377), .A2(STATE_REG_SCAN_IN), .ZN(n2880) );
  OAI21_X1 U3628 ( .B1(STATE_REG_SCAN_IN), .B2(n2881), .A(n2880), .ZN(U3325)
         );
  INV_X1 U3629 ( .A(DATAI_31_), .ZN(n2884) );
  OR4_X1 U3630 ( .A1(n2882), .A2(IR_REG_30__SCAN_IN), .A3(U3149), .A4(n2259), 
        .ZN(n2883) );
  OAI21_X1 U3631 ( .B1(STATE_REG_SCAN_IN), .B2(n2884), .A(n2883), .ZN(U3321)
         );
  INV_X1 U3632 ( .A(DATAI_30_), .ZN(n2887) );
  NAND2_X1 U3633 ( .A1(n2885), .A2(STATE_REG_SCAN_IN), .ZN(n2886) );
  OAI21_X1 U3634 ( .B1(STATE_REG_SCAN_IN), .B2(n2887), .A(n2886), .ZN(U3322)
         );
  INV_X1 U3635 ( .A(n3002), .ZN(n2904) );
  INV_X1 U3636 ( .A(D_REG_0__SCAN_IN), .ZN(n4738) );
  INV_X1 U3637 ( .A(n2888), .ZN(n2889) );
  AOI22_X1 U3638 ( .A1(n4505), .A2(n4738), .B1(n2889), .B2(n4506), .ZN(U3458)
         );
  INV_X1 U3639 ( .A(D_REG_1__SCAN_IN), .ZN(n2891) );
  AOI22_X1 U3640 ( .A1(n4505), .A2(n2891), .B1(n2890), .B2(n4506), .ZN(U3459)
         );
  INV_X1 U3641 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4577) );
  INV_X1 U3642 ( .A(REG2_REG_31__SCAN_IN), .ZN(n2894) );
  NAND2_X1 U3643 ( .A1(n2775), .A2(REG1_REG_31__SCAN_IN), .ZN(n2893) );
  NAND2_X1 U3644 ( .A1(n3424), .A2(REG0_REG_31__SCAN_IN), .ZN(n2892) );
  OAI211_X1 U3645 ( .C1(n2895), .C2(n2894), .A(n2893), .B(n2892), .ZN(n4191)
         );
  NAND2_X1 U3646 ( .A1(n4191), .A2(U4043), .ZN(n2896) );
  OAI21_X1 U3647 ( .B1(U4043), .B2(n4577), .A(n2896), .ZN(U3581) );
  INV_X1 U3648 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U3649 ( .A1(n2447), .A2(U4043), .ZN(n2897) );
  OAI21_X1 U3650 ( .B1(U4043), .B2(n4696), .A(n2897), .ZN(U3552) );
  INV_X1 U3651 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4713) );
  NAND2_X1 U3652 ( .A1(n3542), .A2(U4043), .ZN(n2898) );
  OAI21_X1 U3653 ( .B1(U4043), .B2(n4713), .A(n2898), .ZN(U3555) );
  INV_X1 U3654 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U3655 ( .A1(n3183), .A2(U4043), .ZN(n2899) );
  OAI21_X1 U3656 ( .B1(U4043), .B2(n4575), .A(n2899), .ZN(U3556) );
  INV_X1 U3657 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U3658 ( .A1(n3543), .A2(U4043), .ZN(n2900) );
  OAI21_X1 U3659 ( .B1(U4043), .B2(n4723), .A(n2900), .ZN(U3553) );
  INV_X1 U3660 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U3661 ( .A1(n3987), .A2(U4043), .ZN(n2901) );
  OAI21_X1 U3662 ( .B1(U4043), .B2(n4734), .A(n2901), .ZN(U3573) );
  INV_X1 U3663 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4728) );
  INV_X1 U3664 ( .A(n2984), .ZN(n2990) );
  NAND2_X1 U3665 ( .A1(n2984), .A2(U4043), .ZN(n2902) );
  OAI21_X1 U3666 ( .B1(U4043), .B2(n4728), .A(n2902), .ZN(U3550) );
  NAND2_X1 U3667 ( .A1(n2905), .A2(n2904), .ZN(n2906) );
  OR2_X1 U3668 ( .A1(n2907), .A2(n2906), .ZN(n3482) );
  INV_X1 U3669 ( .A(n3602), .ZN(n3568) );
  OAI22_X1 U3670 ( .A1(n3568), .A2(n3089), .B1(n3570), .B2(n3087), .ZN(n2908)
         );
  AOI21_X1 U3671 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3482), .A(n2908), .ZN(n2909)
         );
  OAI21_X1 U3672 ( .B1(n3577), .B2(n3800), .A(n2909), .ZN(U3229) );
  INV_X1 U3673 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2910) );
  XNOR2_X1 U3674 ( .A(n3778), .B(REG1_REG_1__SCAN_IN), .ZN(n3776) );
  NOR2_X1 U3675 ( .A1(n2316), .A2(n4558), .ZN(n3775) );
  NAND2_X1 U3676 ( .A1(n3776), .A2(n3775), .ZN(n3774) );
  NAND2_X1 U3677 ( .A1(n3777), .A2(REG1_REG_1__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U3678 ( .A1(n3774), .A2(n2911), .ZN(n3791) );
  NAND2_X1 U3679 ( .A1(n4365), .A2(REG1_REG_2__SCAN_IN), .ZN(n2912) );
  INV_X1 U3680 ( .A(n4364), .ZN(n2945) );
  XNOR2_X1 U3681 ( .A(n2913), .B(n2945), .ZN(n2939) );
  NAND2_X1 U3682 ( .A1(n2939), .A2(REG1_REG_3__SCAN_IN), .ZN(n2915) );
  NAND2_X1 U3683 ( .A1(n2913), .A2(n4364), .ZN(n2914) );
  NAND2_X1 U3684 ( .A1(n2915), .A2(n2914), .ZN(n2917) );
  INV_X1 U3685 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2916) );
  NAND2_X1 U3686 ( .A1(n2917), .A2(n4390), .ZN(n2918) );
  INV_X1 U3687 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2920) );
  MUX2_X1 U3688 ( .A(n2920), .B(REG1_REG_5__SCAN_IN), .S(n2974), .Z(n2919) );
  INV_X1 U3689 ( .A(n4363), .ZN(n2948) );
  XNOR2_X1 U3690 ( .A(n2946), .B(REG1_REG_6__SCAN_IN), .ZN(n2938) );
  NAND2_X1 U3691 ( .A1(n2988), .A2(n2922), .ZN(n2921) );
  AND2_X1 U3692 ( .A1(n3629), .A2(n2921), .ZN(n2931) );
  OR2_X1 U3693 ( .A1(n2922), .A2(U3149), .ZN(n3759) );
  NAND2_X1 U3694 ( .A1(n3002), .A2(n3759), .ZN(n2930) );
  NAND2_X1 U3695 ( .A1(n2931), .A2(n2930), .ZN(n4380) );
  INV_X1 U3696 ( .A(n2974), .ZN(n2929) );
  NAND2_X1 U3697 ( .A1(n3777), .A2(REG2_REG_1__SCAN_IN), .ZN(n2924) );
  INV_X1 U3698 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U3699 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3780) );
  AOI21_X1 U3700 ( .B1(n3778), .B2(n3779), .A(n3780), .ZN(n2923) );
  NAND2_X1 U3701 ( .A1(n2924), .A2(n2923), .ZN(n3783) );
  NAND2_X1 U3702 ( .A1(n3783), .A2(n2924), .ZN(n3789) );
  INV_X1 U3703 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3047) );
  AOI22_X1 U3704 ( .A1(n3789), .A2(n3788), .B1(n4365), .B2(REG2_REG_2__SCAN_IN), .ZN(n2925) );
  XOR2_X1 U3705 ( .A(n4364), .B(n2925), .Z(n2940) );
  INV_X1 U3706 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2926) );
  OAI22_X1 U3707 ( .A1(n2940), .A2(n2926), .B1(n2925), .B2(n2945), .ZN(n2927)
         );
  XNOR2_X1 U3708 ( .A(n2927), .B(n4390), .ZN(n4383) );
  INV_X1 U3709 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2928) );
  MUX2_X1 U3710 ( .A(REG2_REG_5__SCAN_IN), .B(n2928), .S(n2974), .Z(n2976) );
  XNOR2_X1 U3711 ( .A(n2950), .B(REG2_REG_6__SCAN_IN), .ZN(n2936) );
  INV_X1 U3712 ( .A(n4377), .ZN(n3798) );
  OR2_X1 U3713 ( .A1(n4367), .A2(n3798), .ZN(n3802) );
  INV_X1 U3714 ( .A(n2930), .ZN(n2932) );
  NOR2_X1 U3715 ( .A1(STATE_REG_SCAN_IN), .A2(n2933), .ZN(n3125) );
  AOI21_X1 U3716 ( .B1(n4457), .B2(ADDR_REG_6__SCAN_IN), .A(n3125), .ZN(n2934)
         );
  OAI21_X1 U3717 ( .B1(n2948), .B2(n4490), .A(n2934), .ZN(n2935) );
  AOI21_X1 U3718 ( .B1(n2936), .B2(n4487), .A(n2935), .ZN(n2937) );
  OAI21_X1 U3719 ( .B1(n2938), .B2(n4475), .A(n2937), .ZN(U3246) );
  NOR2_X1 U3720 ( .A1(n4457), .A2(U4043), .ZN(U3148) );
  XOR2_X1 U3721 ( .A(REG1_REG_3__SCAN_IN), .B(n2939), .Z(n2942) );
  XNOR2_X1 U3722 ( .A(n2940), .B(REG2_REG_3__SCAN_IN), .ZN(n2941) );
  AOI22_X1 U3723 ( .A1(n4471), .A2(n2942), .B1(n4487), .B2(n2941), .ZN(n2944)
         );
  AOI22_X1 U3724 ( .A1(n4457), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2943) );
  OAI211_X1 U3725 ( .C1(n2945), .C2(n4490), .A(n2944), .B(n2943), .ZN(U3243)
         );
  INV_X1 U3726 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4563) );
  XOR2_X1 U3727 ( .A(n4563), .B(n4362), .Z(n2947) );
  XNOR2_X1 U3728 ( .A(n2963), .B(n2947), .ZN(n2958) );
  OAI22_X1 U3729 ( .A1(n2950), .A2(n3168), .B1(n2949), .B2(n2948), .ZN(n2954)
         );
  MUX2_X1 U3730 ( .A(REG2_REG_7__SCAN_IN), .B(n2951), .S(n4362), .Z(n2953) );
  MUX2_X1 U3731 ( .A(n2951), .B(REG2_REG_7__SCAN_IN), .S(n4362), .Z(n2952) );
  OAI211_X1 U3732 ( .C1(n2954), .C2(n2953), .A(n4487), .B(n2959), .ZN(n2957)
         );
  AND2_X1 U3733 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3182) );
  INV_X1 U3734 ( .A(n4362), .ZN(n2960) );
  NOR2_X1 U3735 ( .A1(n4490), .A2(n2960), .ZN(n2955) );
  AOI211_X1 U3736 ( .C1(n4457), .C2(ADDR_REG_7__SCAN_IN), .A(n3182), .B(n2955), 
        .ZN(n2956) );
  OAI211_X1 U3737 ( .C1(n2958), .C2(n4475), .A(n2957), .B(n2956), .ZN(U3247)
         );
  XNOR2_X1 U3738 ( .A(n3826), .B(REG2_REG_8__SCAN_IN), .ZN(n2970) );
  AND2_X1 U3739 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3214) );
  NOR2_X1 U3740 ( .A1(n4490), .A2(n3828), .ZN(n2961) );
  AOI211_X1 U3741 ( .C1(n4457), .C2(ADDR_REG_8__SCAN_IN), .A(n3214), .B(n2961), 
        .ZN(n2969) );
  NAND2_X1 U3742 ( .A1(n4362), .A2(REG1_REG_7__SCAN_IN), .ZN(n2962) );
  OR2_X1 U3743 ( .A1(n4362), .A2(REG1_REG_7__SCAN_IN), .ZN(n2964) );
  NAND2_X1 U3744 ( .A1(n2965), .A2(n2964), .ZN(n3810) );
  INV_X1 U3745 ( .A(n2966), .ZN(n2967) );
  INV_X1 U3746 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3286) );
  OAI211_X1 U3747 ( .C1(n2967), .C2(REG1_REG_8__SCAN_IN), .A(n3809), .B(n4471), 
        .ZN(n2968) );
  OAI211_X1 U3748 ( .C1(n2970), .C2(n4443), .A(n2969), .B(n2968), .ZN(U3248)
         );
  MUX2_X1 U3749 ( .A(REG1_REG_5__SCAN_IN), .B(n2920), .S(n2974), .Z(n2972) );
  AOI211_X1 U3750 ( .C1(n2096), .C2(n2972), .A(n2971), .B(n4475), .ZN(n2980)
         );
  AND2_X1 U3751 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3065) );
  AOI21_X1 U3752 ( .B1(n4457), .B2(ADDR_REG_5__SCAN_IN), .A(n3065), .ZN(n2973)
         );
  OAI21_X1 U3753 ( .B1(n2974), .B2(n4490), .A(n2973), .ZN(n2979) );
  AOI211_X1 U3754 ( .C1(n2977), .C2(n2976), .A(n2975), .B(n4443), .ZN(n2978)
         );
  OR3_X1 U3755 ( .A1(n2980), .A2(n2979), .A3(n2978), .ZN(U3245) );
  INV_X1 U3756 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n2982) );
  NAND2_X1 U3757 ( .A1(n3908), .A2(U4043), .ZN(n2981) );
  OAI21_X1 U3758 ( .B1(U4043), .B2(n2982), .A(n2981), .ZN(U3577) );
  XNOR2_X1 U3759 ( .A(n3035), .B(n3756), .ZN(n2983) );
  NAND2_X1 U3760 ( .A1(n2986), .A2(n2985), .ZN(n3024) );
  OAI21_X1 U3761 ( .B1(n2985), .B2(n2986), .A(n3024), .ZN(n3095) );
  INV_X1 U3762 ( .A(n2447), .ZN(n3025) );
  INV_X1 U3763 ( .A(n4166), .ZN(n4139) );
  OAI22_X1 U3764 ( .A1(n3025), .A2(n4139), .B1(n4200), .B2(n2996), .ZN(n2994)
         );
  NAND2_X1 U3765 ( .A1(n2985), .A2(n3649), .ZN(n2992) );
  NAND2_X1 U3766 ( .A1(n4361), .A2(n3652), .ZN(n3749) );
  NAND2_X1 U3767 ( .A1(n3850), .A2(n3756), .ZN(n2991) );
  AOI21_X1 U3768 ( .B1(n3038), .B2(n2992), .A(n4147), .ZN(n2993) );
  AOI211_X1 U3769 ( .C1(n4143), .C2(n2984), .A(n2994), .B(n2993), .ZN(n2995)
         );
  OAI21_X1 U3770 ( .B1(n4175), .B2(n3095), .A(n2995), .ZN(n3094) );
  NAND2_X1 U3771 ( .A1(n3087), .A2(n2996), .ZN(n3044) );
  OAI21_X1 U3772 ( .B1(n2996), .B2(n3087), .A(n3044), .ZN(n3101) );
  OAI22_X1 U3773 ( .A1(n3095), .A2(n4531), .B1(n4530), .B2(n3101), .ZN(n2997)
         );
  NOR2_X1 U3774 ( .A1(n3094), .A2(n2997), .ZN(n4528) );
  OR2_X1 U3775 ( .A1(n3000), .A2(n2998), .ZN(n3005) );
  OAI21_X1 U3776 ( .B1(n3000), .B2(D_REG_1__SCAN_IN), .A(n2999), .ZN(n3004) );
  NOR2_X1 U3777 ( .A1(n3002), .A2(n3001), .ZN(n3032) );
  NAND4_X1 U3778 ( .A1(n3005), .A2(n3004), .A3(n3032), .A4(n3003), .ZN(n3057)
         );
  NAND2_X1 U3779 ( .A1(n4565), .A2(REG1_REG_1__SCAN_IN), .ZN(n3006) );
  OAI21_X1 U3780 ( .B1(n4528), .B2(n4565), .A(n3006), .ZN(U3519) );
  INV_X1 U3781 ( .A(n3008), .ZN(n3009) );
  AOI21_X1 U3782 ( .B1(n3007), .B2(n3010), .A(n3009), .ZN(n3014) );
  INV_X1 U3783 ( .A(n3043), .ZN(n3071) );
  AOI22_X1 U3784 ( .A1(n3602), .A2(n3543), .B1(n3603), .B2(n3773), .ZN(n3011)
         );
  OAI21_X1 U3785 ( .B1(n3570), .B2(n3071), .A(n3011), .ZN(n3012) );
  AOI21_X1 U3786 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3482), .A(n3012), .ZN(n3013)
         );
  OAI21_X1 U3787 ( .B1(n3014), .B2(n3577), .A(n3013), .ZN(U3234) );
  OAI21_X1 U3788 ( .B1(n3017), .B2(n3016), .A(n3015), .ZN(n3021) );
  MUX2_X1 U3789 ( .A(STATE_REG_SCAN_IN), .B(n3607), .S(n2456), .Z(n3019) );
  AOI22_X1 U3790 ( .A1(n3603), .A2(n2447), .B1(n3602), .B2(n3771), .ZN(n3018)
         );
  OAI211_X1 U3791 ( .C1(n3570), .C2(n3103), .A(n3019), .B(n3018), .ZN(n3020)
         );
  AOI21_X1 U3792 ( .B1(n3021), .B2(n3609), .A(n3020), .ZN(n3022) );
  INV_X1 U3793 ( .A(n3022), .ZN(U3215) );
  NAND2_X1 U3794 ( .A1(n3773), .A2(n3483), .ZN(n3023) );
  NAND2_X1 U3795 ( .A1(n3024), .A2(n3023), .ZN(n3028) );
  INV_X1 U3796 ( .A(n3028), .ZN(n3026) );
  NAND2_X1 U3797 ( .A1(n2447), .A2(n3071), .ZN(n3656) );
  NAND2_X1 U3798 ( .A1(n3028), .A2(n3027), .ZN(n3029) );
  AND2_X1 U3799 ( .A1(n3030), .A2(n3029), .ZN(n3051) );
  NAND3_X1 U3800 ( .A1(n3033), .A2(n3032), .A3(n3031), .ZN(n3034) );
  OR2_X1 U3801 ( .A1(n3035), .A2(n3860), .ZN(n3153) );
  INV_X1 U3802 ( .A(n3153), .ZN(n3036) );
  OAI22_X1 U3803 ( .A1(n3104), .A2(n4139), .B1(n3071), .B2(n4200), .ZN(n3041)
         );
  NAND3_X1 U3804 ( .A1(n3614), .A2(n3037), .A3(n3038), .ZN(n3039) );
  AOI21_X1 U3805 ( .B1(n3073), .B2(n3039), .A(n4147), .ZN(n3040) );
  AOI211_X1 U3806 ( .C1(n4143), .C2(n3773), .A(n3041), .B(n3040), .ZN(n3042)
         );
  OAI21_X1 U3807 ( .B1(n3051), .B2(n4175), .A(n3042), .ZN(n3052) );
  NAND2_X1 U3808 ( .A1(n3052), .A2(n4373), .ZN(n3050) );
  AND2_X1 U3809 ( .A1(n3044), .A2(n3043), .ZN(n3045) );
  NOR2_X1 U3810 ( .A1(n3079), .A2(n3045), .ZN(n3060) );
  OAI22_X1 U3811 ( .A1(n4183), .A2(n3047), .B1(n3046), .B2(n4180), .ZN(n3048)
         );
  AOI21_X1 U3812 ( .B1(n3060), .B2(n4498), .A(n3048), .ZN(n3049) );
  OAI211_X1 U3813 ( .C1(n3051), .C2(n4188), .A(n3050), .B(n3049), .ZN(U3288)
         );
  INV_X1 U3814 ( .A(n3051), .ZN(n3053) );
  AOI21_X1 U3815 ( .B1(n4540), .B2(n3053), .A(n3052), .ZN(n3062) );
  NOR2_X1 U3816 ( .A1(n4568), .A2(n2910), .ZN(n3054) );
  AOI21_X1 U3817 ( .B1(n3060), .B2(n4248), .A(n3054), .ZN(n3055) );
  OAI21_X1 U3818 ( .B1(n3062), .B2(n4565), .A(n3055), .ZN(U3520) );
  INV_X1 U3819 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3058) );
  NOR2_X1 U3820 ( .A1(n4756), .A2(n3058), .ZN(n3059) );
  AOI21_X1 U3821 ( .B1(n3060), .B2(n4330), .A(n3059), .ZN(n3061) );
  OAI21_X1 U3822 ( .B1(n3062), .B2(n4556), .A(n3061), .ZN(U3471) );
  XOR2_X1 U3823 ( .A(n3064), .B(n3063), .Z(n3069) );
  AOI21_X1 U3824 ( .B1(n3602), .B2(n3183), .A(n3065), .ZN(n3067) );
  AOI22_X1 U3825 ( .A1(n3604), .A2(n3191), .B1(n3603), .B2(n3771), .ZN(n3066)
         );
  OAI211_X1 U3826 ( .C1(n3607), .C2(n3205), .A(n3067), .B(n3066), .ZN(n3068)
         );
  AOI21_X1 U3827 ( .B1(n3069), .B2(n3609), .A(n3068), .ZN(n3070) );
  INV_X1 U3828 ( .A(n3070), .ZN(U3224) );
  NAND2_X1 U3829 ( .A1(n3025), .A2(n3071), .ZN(n3072) );
  NAND2_X1 U3830 ( .A1(n3104), .A2(n3102), .ZN(n3658) );
  NAND2_X1 U3831 ( .A1(n3543), .A2(n3103), .ZN(n3655) );
  XNOR2_X1 U3832 ( .A(n3142), .B(n3612), .ZN(n4532) );
  NAND2_X1 U3833 ( .A1(n3073), .A2(n3653), .ZN(n3074) );
  OAI21_X1 U3834 ( .B1(n3612), .B2(n3074), .A(n3110), .ZN(n3077) );
  AOI22_X1 U3835 ( .A1(n3771), .A2(n4166), .B1(n4192), .B2(n3102), .ZN(n3075)
         );
  OAI21_X1 U3836 ( .B1(n3025), .B2(n4169), .A(n3075), .ZN(n3076) );
  AOI21_X1 U3837 ( .B1(n3077), .B2(n4172), .A(n3076), .ZN(n3078) );
  OAI21_X1 U3838 ( .B1(n4532), .B2(n4175), .A(n3078), .ZN(n4534) );
  INV_X1 U3839 ( .A(n4534), .ZN(n3084) );
  INV_X1 U3840 ( .A(n4373), .ZN(n4368) );
  INV_X1 U3841 ( .A(n4532), .ZN(n3082) );
  NAND2_X1 U3842 ( .A1(n3079), .A2(n3103), .ZN(n3116) );
  OAI21_X1 U3843 ( .B1(n3079), .B2(n3103), .A(n3116), .ZN(n4529) );
  AOI22_X1 U3844 ( .A1(n4368), .A2(REG2_REG_3__SCAN_IN), .B1(n4496), .B2(n2456), .ZN(n3080) );
  OAI21_X1 U3845 ( .B1(n4151), .B2(n4529), .A(n3080), .ZN(n3081) );
  AOI21_X1 U3846 ( .B1(n3082), .B2(n4499), .A(n3081), .ZN(n3083) );
  OAI21_X1 U3847 ( .B1(n3084), .B2(n4368), .A(n3083), .ZN(U3287) );
  INV_X1 U3848 ( .A(n3085), .ZN(n3086) );
  NOR2_X1 U3849 ( .A1(n3087), .A2(n3086), .ZN(n4524) );
  INV_X1 U3850 ( .A(n4175), .ZN(n4494) );
  NAND2_X1 U3851 ( .A1(n2984), .A2(n3087), .ZN(n3651) );
  NAND2_X1 U3852 ( .A1(n3649), .A2(n3651), .ZN(n4525) );
  OAI21_X1 U3853 ( .B1(n4494), .B2(n4172), .A(n4525), .ZN(n3088) );
  OAI21_X1 U3854 ( .B1(n3089), .B2(n4139), .A(n3088), .ZN(n4523) );
  AOI21_X1 U3855 ( .B1(n4524), .B2(n3090), .A(n4523), .ZN(n3093) );
  AOI22_X1 U3856 ( .A1(n4368), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4496), .ZN(n3092) );
  NAND2_X1 U3857 ( .A1(n4525), .A2(n4499), .ZN(n3091) );
  OAI211_X1 U3858 ( .C1(n3093), .C2(n4368), .A(n3092), .B(n3091), .ZN(U3290)
         );
  NAND2_X1 U3859 ( .A1(n3094), .A2(n4373), .ZN(n3100) );
  INV_X1 U3860 ( .A(n3095), .ZN(n3098) );
  INV_X1 U3861 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3096) );
  OAI22_X1 U3862 ( .A1(n4183), .A2(n3779), .B1(n3096), .B2(n4180), .ZN(n3097)
         );
  AOI21_X1 U3863 ( .B1(n3098), .B2(n4499), .A(n3097), .ZN(n3099) );
  OAI211_X1 U3864 ( .C1(n3101), .C2(n4151), .A(n3100), .B(n3099), .ZN(U3289)
         );
  NAND2_X1 U3865 ( .A1(n3543), .A2(n3102), .ZN(n3140) );
  NAND2_X1 U3866 ( .A1(n3142), .A2(n3140), .ZN(n3105) );
  NAND2_X1 U3867 ( .A1(n3104), .A2(n3103), .ZN(n3144) );
  NAND2_X1 U3868 ( .A1(n3105), .A2(n3144), .ZN(n3107) );
  INV_X1 U3869 ( .A(n3771), .ZN(n3106) );
  INV_X1 U3870 ( .A(n3544), .ZN(n3117) );
  OR2_X1 U3871 ( .A1(n3107), .A2(n3616), .ZN(n3109) );
  NAND2_X1 U3872 ( .A1(n3107), .A2(n3616), .ZN(n3108) );
  NAND2_X1 U3873 ( .A1(n3109), .A2(n3108), .ZN(n4536) );
  XNOR2_X1 U3874 ( .A(n3132), .B(n3616), .ZN(n3114) );
  AOI22_X1 U3875 ( .A1(n3543), .A2(n4143), .B1(n3544), .B2(n4192), .ZN(n3112)
         );
  NAND2_X1 U3876 ( .A1(n3542), .A2(n4166), .ZN(n3111) );
  OAI211_X1 U3877 ( .C1(n4536), .C2(n4175), .A(n3112), .B(n3111), .ZN(n3113)
         );
  AOI21_X1 U3878 ( .B1(n3114), .B2(n4172), .A(n3113), .ZN(n3115) );
  INV_X1 U3879 ( .A(n3115), .ZN(n4538) );
  INV_X1 U3880 ( .A(n3116), .ZN(n3118) );
  OAI211_X1 U3881 ( .C1(n3118), .C2(n3117), .A(n4551), .B(n3190), .ZN(n4537)
         );
  OAI22_X1 U3882 ( .A1(n4537), .A2(n3850), .B1(n4180), .B2(n3545), .ZN(n3119)
         );
  OAI21_X1 U3883 ( .B1(n4538), .B2(n3119), .A(n4373), .ZN(n3121) );
  NAND2_X1 U3884 ( .A1(n4368), .A2(REG2_REG_4__SCAN_IN), .ZN(n3120) );
  OAI211_X1 U3885 ( .C1(n4536), .C2(n4188), .A(n3121), .B(n3120), .ZN(U3286)
         );
  NAND2_X1 U3886 ( .A1(n3174), .A2(n3122), .ZN(n3124) );
  NAND2_X1 U3887 ( .A1(n2062), .A2(n3175), .ZN(n3123) );
  XNOR2_X1 U3888 ( .A(n3124), .B(n3123), .ZN(n3129) );
  AOI21_X1 U3889 ( .B1(n3602), .B2(n3770), .A(n3125), .ZN(n3127) );
  AOI22_X1 U3890 ( .A1(n3604), .A2(n3159), .B1(n3603), .B2(n3542), .ZN(n3126)
         );
  OAI211_X1 U3891 ( .C1(n3607), .C2(n3167), .A(n3127), .B(n3126), .ZN(n3128)
         );
  AOI21_X1 U3892 ( .B1(n3129), .B2(n3609), .A(n3128), .ZN(n3130) );
  INV_X1 U3893 ( .A(n3130), .ZN(U3236) );
  INV_X1 U3894 ( .A(n3659), .ZN(n3131) );
  AND2_X1 U3895 ( .A1(n3542), .A2(n3197), .ZN(n3194) );
  INV_X1 U3896 ( .A(n3542), .ZN(n3161) );
  NAND2_X1 U3897 ( .A1(n3161), .A2(n3191), .ZN(n3679) );
  OAI21_X1 U3898 ( .B1(n3196), .B2(n3194), .A(n3679), .ZN(n3158) );
  NAND2_X1 U3899 ( .A1(n3183), .A2(n2274), .ZN(n3677) );
  NAND2_X1 U3900 ( .A1(n3158), .A2(n3677), .ZN(n3133) );
  NAND2_X1 U3901 ( .A1(n2275), .A2(n3159), .ZN(n3664) );
  NAND2_X1 U3902 ( .A1(n3133), .A2(n3664), .ZN(n3230) );
  INV_X1 U3903 ( .A(n3770), .ZN(n3250) );
  NAND2_X1 U3904 ( .A1(n3250), .A2(n3239), .ZN(n3228) );
  NAND2_X1 U3905 ( .A1(n3770), .A2(n3137), .ZN(n3667) );
  XNOR2_X1 U3906 ( .A(n3230), .B(n3665), .ZN(n3136) );
  AOI22_X1 U3907 ( .A1(n3769), .A2(n4166), .B1(n4192), .B2(n3239), .ZN(n3134)
         );
  OAI21_X1 U3908 ( .B1(n2275), .B2(n4169), .A(n3134), .ZN(n3135) );
  AOI21_X1 U3909 ( .B1(n3136), .B2(n4172), .A(n3135), .ZN(n4547) );
  NAND2_X1 U3910 ( .A1(n3166), .A2(n3137), .ZN(n3254) );
  OAI211_X1 U3911 ( .C1(n3166), .C2(n3137), .A(n4551), .B(n3254), .ZN(n4546)
         );
  INV_X1 U3912 ( .A(n4546), .ZN(n3139) );
  OAI22_X1 U3913 ( .A1(n4183), .A2(n2951), .B1(n3186), .B2(n4180), .ZN(n3138)
         );
  AOI21_X1 U3914 ( .B1(n3139), .B2(n4080), .A(n3138), .ZN(n3156) );
  NAND2_X1 U3915 ( .A1(n3771), .A2(n3544), .ZN(n3143) );
  AND2_X1 U3916 ( .A1(n3140), .A2(n3143), .ZN(n3141) );
  NAND2_X1 U3917 ( .A1(n3142), .A2(n3141), .ZN(n3193) );
  INV_X1 U3918 ( .A(n3143), .ZN(n3147) );
  NAND2_X1 U3919 ( .A1(n3659), .A2(n3661), .ZN(n3145) );
  AND2_X1 U3920 ( .A1(n3145), .A2(n3144), .ZN(n3146) );
  NAND2_X1 U3921 ( .A1(n3161), .A2(n3197), .ZN(n3148) );
  NAND3_X1 U3922 ( .A1(n3193), .A2(n3192), .A3(n3148), .ZN(n3150) );
  NAND2_X1 U3923 ( .A1(n3542), .A2(n3191), .ZN(n3149) );
  NAND2_X1 U3924 ( .A1(n3152), .A2(n3665), .ZN(n4543) );
  NAND2_X1 U3925 ( .A1(n4175), .A2(n3153), .ZN(n3154) );
  INV_X1 U3926 ( .A(n4133), .ZN(n4007) );
  NAND3_X1 U3927 ( .A1(n4544), .A2(n4543), .A3(n4007), .ZN(n3155) );
  OAI211_X1 U3928 ( .C1(n4547), .C2(n4368), .A(n3156), .B(n3155), .ZN(U3283)
         );
  NAND2_X1 U3929 ( .A1(n3664), .A2(n3677), .ZN(n3619) );
  XNOR2_X1 U3930 ( .A(n3157), .B(n3619), .ZN(n3220) );
  XOR2_X1 U3931 ( .A(n3619), .B(n3158), .Z(n3163) );
  AOI22_X1 U3932 ( .A1(n3770), .A2(n4166), .B1(n4192), .B2(n3159), .ZN(n3160)
         );
  OAI21_X1 U3933 ( .B1(n3161), .B2(n4169), .A(n3160), .ZN(n3162) );
  AOI21_X1 U3934 ( .B1(n3163), .B2(n4172), .A(n3162), .ZN(n3164) );
  OAI21_X1 U3935 ( .B1(n4175), .B2(n3220), .A(n3164), .ZN(n3221) );
  NAND2_X1 U3936 ( .A1(n3221), .A2(n4373), .ZN(n3172) );
  NOR2_X1 U3937 ( .A1(n3189), .A2(n2274), .ZN(n3165) );
  OR2_X1 U3938 ( .A1(n3166), .A2(n3165), .ZN(n3227) );
  INV_X1 U3939 ( .A(n3227), .ZN(n3170) );
  OAI22_X1 U3940 ( .A1(n4183), .A2(n3168), .B1(n3167), .B2(n4180), .ZN(n3169)
         );
  AOI21_X1 U3941 ( .B1(n3170), .B2(n4498), .A(n3169), .ZN(n3171) );
  OAI211_X1 U3942 ( .C1(n3220), .C2(n4188), .A(n3172), .B(n3171), .ZN(U3284)
         );
  AND2_X1 U3943 ( .A1(n3174), .A2(n3173), .ZN(n3178) );
  INV_X1 U3944 ( .A(n3178), .ZN(n3176) );
  NAND2_X1 U3945 ( .A1(n3176), .A2(n3175), .ZN(n3180) );
  NOR2_X1 U3946 ( .A1(n3178), .A2(n3177), .ZN(n3179) );
  AOI211_X1 U3947 ( .C1(n3181), .C2(n3180), .A(n3577), .B(n3179), .ZN(n3188)
         );
  AOI21_X1 U3948 ( .B1(n3602), .B2(n3769), .A(n3182), .ZN(n3185) );
  AOI22_X1 U3949 ( .A1(n3604), .A2(n3239), .B1(n3603), .B2(n3183), .ZN(n3184)
         );
  OAI211_X1 U3950 ( .C1(n3607), .C2(n3186), .A(n3185), .B(n3184), .ZN(n3187)
         );
  OR2_X1 U3951 ( .A1(n3188), .A2(n3187), .ZN(U3210) );
  AOI21_X1 U3952 ( .B1(n3191), .B2(n3190), .A(n3189), .ZN(n3206) );
  AND2_X1 U3953 ( .A1(n3193), .A2(n3192), .ZN(n3195) );
  INV_X1 U3954 ( .A(n3194), .ZN(n3662) );
  NAND2_X1 U3955 ( .A1(n3662), .A2(n3679), .ZN(n3628) );
  XNOR2_X1 U3956 ( .A(n3195), .B(n3628), .ZN(n3209) );
  INV_X1 U3957 ( .A(n4549), .ZN(n4245) );
  NOR2_X1 U3958 ( .A1(n3209), .A2(n4245), .ZN(n3201) );
  XOR2_X1 U3959 ( .A(n3628), .B(n3196), .Z(n3200) );
  OAI22_X1 U3960 ( .A1(n2275), .A2(n4139), .B1(n4200), .B2(n3197), .ZN(n3198)
         );
  AOI21_X1 U3961 ( .B1(n4143), .B2(n3771), .A(n3198), .ZN(n3199) );
  OAI21_X1 U3962 ( .B1(n3200), .B2(n4147), .A(n3199), .ZN(n3203) );
  AOI211_X1 U3963 ( .C1(n4551), .C2(n3206), .A(n3201), .B(n3203), .ZN(n4754)
         );
  OR2_X1 U3964 ( .A1(n4754), .A2(n4565), .ZN(n3202) );
  OAI21_X1 U3965 ( .B1(n4568), .B2(n2920), .A(n3202), .ZN(U3523) );
  INV_X1 U3966 ( .A(n3203), .ZN(n3204) );
  MUX2_X1 U3967 ( .A(n3204), .B(n2928), .S(n4368), .Z(n3208) );
  AOI22_X1 U3968 ( .A1(n3206), .A2(n4498), .B1(n2136), .B2(n4496), .ZN(n3207)
         );
  OAI211_X1 U3969 ( .C1(n4133), .C2(n3209), .A(n3208), .B(n3207), .ZN(U3285)
         );
  XNOR2_X1 U3970 ( .A(n3211), .B(n3210), .ZN(n3212) );
  XNOR2_X1 U3971 ( .A(n3213), .B(n3212), .ZN(n3218) );
  AOI21_X1 U3972 ( .B1(n3602), .B2(n3768), .A(n3214), .ZN(n3216) );
  AOI22_X1 U3973 ( .A1(n3604), .A2(n3248), .B1(n3603), .B2(n3770), .ZN(n3215)
         );
  OAI211_X1 U3974 ( .C1(n3607), .C2(n3258), .A(n3216), .B(n3215), .ZN(n3217)
         );
  AOI21_X1 U3975 ( .B1(n3218), .B2(n3609), .A(n3217), .ZN(n3219) );
  INV_X1 U3976 ( .A(n3219), .ZN(U3218) );
  INV_X1 U3977 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3223) );
  INV_X1 U3978 ( .A(n3220), .ZN(n3222) );
  AOI21_X1 U3979 ( .B1(n4540), .B2(n3222), .A(n3221), .ZN(n3225) );
  MUX2_X1 U3980 ( .A(n3223), .B(n3225), .S(n4756), .Z(n3224) );
  OAI21_X1 U3981 ( .B1(n3227), .B2(n4358), .A(n3224), .ZN(U3479) );
  INV_X1 U3982 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4570) );
  MUX2_X1 U3983 ( .A(n4570), .B(n3225), .S(n4568), .Z(n3226) );
  OAI21_X1 U3984 ( .B1(n3227), .B2(n4276), .A(n3226), .ZN(U3524) );
  INV_X1 U3985 ( .A(n3228), .ZN(n3229) );
  INV_X1 U3986 ( .A(n3769), .ZN(n3267) );
  NAND2_X1 U3987 ( .A1(n3267), .A2(n3248), .ZN(n3669) );
  NAND2_X1 U3988 ( .A1(n3769), .A2(n3256), .ZN(n3668) );
  INV_X1 U3989 ( .A(n3303), .ZN(n3304) );
  AND2_X1 U3990 ( .A1(n3768), .A2(n3304), .ZN(n3678) );
  INV_X1 U3991 ( .A(n3678), .ZN(n3231) );
  INV_X1 U3992 ( .A(n3768), .ZN(n3364) );
  NAND2_X1 U3993 ( .A1(n3364), .A2(n3303), .ZN(n3670) );
  NAND2_X1 U3994 ( .A1(n3231), .A2(n3670), .ZN(n3621) );
  XNOR2_X1 U3995 ( .A(n3299), .B(n3621), .ZN(n3235) );
  NAND2_X1 U3996 ( .A1(n3769), .A2(n4143), .ZN(n3233) );
  NAND2_X1 U3997 ( .A1(n3767), .A2(n4166), .ZN(n3232) );
  OAI211_X1 U3998 ( .C1(n4200), .C2(n3304), .A(n3233), .B(n3232), .ZN(n3234)
         );
  AOI21_X1 U3999 ( .B1(n3235), .B2(n4172), .A(n3234), .ZN(n4555) );
  AND2_X1 U4000 ( .A1(n3255), .A2(n3303), .ZN(n3236) );
  NOR2_X1 U4001 ( .A1(n3367), .A2(n3236), .ZN(n4552) );
  OAI22_X1 U4002 ( .A1(n4183), .A2(n3237), .B1(n3269), .B2(n4180), .ZN(n3238)
         );
  AOI21_X1 U4003 ( .B1(n4552), .B2(n4498), .A(n3238), .ZN(n3245) );
  NAND2_X1 U4004 ( .A1(n3770), .A2(n3239), .ZN(n3240) );
  NAND2_X1 U4005 ( .A1(n4544), .A2(n3240), .ZN(n3246) );
  NAND2_X1 U4006 ( .A1(n3267), .A2(n3256), .ZN(n3241) );
  NAND2_X1 U4007 ( .A1(n3769), .A2(n3248), .ZN(n3242) );
  INV_X1 U4008 ( .A(n3621), .ZN(n3243) );
  XNOR2_X1 U4009 ( .A(n3302), .B(n3243), .ZN(n4550) );
  NAND2_X1 U4010 ( .A1(n4550), .A2(n4007), .ZN(n3244) );
  OAI211_X1 U4011 ( .C1(n4555), .C2(n4368), .A(n3245), .B(n3244), .ZN(U3281)
         );
  NAND2_X1 U4012 ( .A1(n3669), .A2(n3668), .ZN(n3620) );
  XNOR2_X1 U4013 ( .A(n3246), .B(n3620), .ZN(n3283) );
  XNOR2_X1 U4014 ( .A(n3247), .B(n3620), .ZN(n3252) );
  AOI22_X1 U4015 ( .A1(n3768), .A2(n4166), .B1(n4192), .B2(n3248), .ZN(n3249)
         );
  OAI21_X1 U4016 ( .B1(n3250), .B2(n4169), .A(n3249), .ZN(n3251) );
  AOI21_X1 U4017 ( .B1(n3252), .B2(n4172), .A(n3251), .ZN(n3253) );
  OAI21_X1 U4018 ( .B1(n3283), .B2(n4175), .A(n3253), .ZN(n3284) );
  NAND2_X1 U4019 ( .A1(n3284), .A2(n4373), .ZN(n3262) );
  INV_X1 U4020 ( .A(n3254), .ZN(n3257) );
  OAI21_X1 U4021 ( .B1(n3257), .B2(n3256), .A(n3255), .ZN(n3291) );
  INV_X1 U4022 ( .A(n3291), .ZN(n3260) );
  OAI22_X1 U4023 ( .A1(n4183), .A2(n3829), .B1(n3258), .B2(n4180), .ZN(n3259)
         );
  AOI21_X1 U4024 ( .B1(n3260), .B2(n4498), .A(n3259), .ZN(n3261) );
  OAI211_X1 U4025 ( .C1(n3283), .C2(n4188), .A(n3262), .B(n3261), .ZN(U3282)
         );
  INV_X1 U4026 ( .A(n3263), .ZN(n3264) );
  AOI21_X1 U4027 ( .B1(n3266), .B2(n3265), .A(n3264), .ZN(n3272) );
  AND2_X1 U4028 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4396) );
  INV_X1 U4029 ( .A(n3603), .ZN(n3571) );
  OAI22_X1 U4030 ( .A1(n3267), .A2(n3571), .B1(n3570), .B2(n3304), .ZN(n3268)
         );
  AOI211_X1 U4031 ( .C1(n3602), .C2(n3767), .A(n4396), .B(n3268), .ZN(n3271)
         );
  INV_X1 U4032 ( .A(n3607), .ZN(n3574) );
  NAND2_X1 U4033 ( .A1(n3574), .A2(n2141), .ZN(n3270) );
  OAI211_X1 U4034 ( .C1(n3272), .C2(n3577), .A(n3271), .B(n3270), .ZN(U3228)
         );
  NAND2_X1 U4035 ( .A1(n3274), .A2(n3273), .ZN(n3275) );
  XNOR2_X1 U4036 ( .A(n3276), .B(n3275), .ZN(n3281) );
  INV_X1 U4037 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3277) );
  NOR2_X1 U4038 ( .A1(STATE_REG_SCAN_IN), .A2(n3277), .ZN(n4414) );
  AOI21_X1 U4039 ( .B1(n3602), .B2(n3765), .A(n4414), .ZN(n3279) );
  AOI22_X1 U4040 ( .A1(n3604), .A2(n3309), .B1(n3603), .B2(n3767), .ZN(n3278)
         );
  OAI211_X1 U4041 ( .C1(n3607), .C2(n3316), .A(n3279), .B(n3278), .ZN(n3280)
         );
  AOI21_X1 U4042 ( .B1(n3281), .B2(n3609), .A(n3280), .ZN(n3282) );
  INV_X1 U40430 ( .A(n3282), .ZN(U3233) );
  INV_X1 U4044 ( .A(n3283), .ZN(n3285) );
  AOI21_X1 U4045 ( .B1(n4540), .B2(n3285), .A(n3284), .ZN(n3288) );
  MUX2_X1 U4046 ( .A(n3286), .B(n3288), .S(n4568), .Z(n3287) );
  OAI21_X1 U4047 ( .B1(n3291), .B2(n4276), .A(n3287), .ZN(U3526) );
  INV_X1 U4048 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3289) );
  MUX2_X1 U4049 ( .A(n3289), .B(n3288), .S(n4756), .Z(n3290) );
  OAI21_X1 U4050 ( .B1(n3291), .B2(n4358), .A(n3290), .ZN(U3483) );
  XNOR2_X1 U4051 ( .A(n3347), .B(n3349), .ZN(n3293) );
  XNOR2_X1 U4052 ( .A(n3292), .B(n3293), .ZN(n3297) );
  AND2_X1 U4053 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4425) );
  AOI21_X1 U4054 ( .B1(n3602), .B2(n4142), .A(n4425), .ZN(n3295) );
  AOI22_X1 U4055 ( .A1(n3604), .A2(n3376), .B1(n3603), .B2(n3766), .ZN(n3294)
         );
  OAI211_X1 U4056 ( .C1(n3607), .C2(n3331), .A(n3295), .B(n3294), .ZN(n3296)
         );
  AOI21_X1 U4057 ( .B1(n3297), .B2(n3609), .A(n3296), .ZN(n3298) );
  INV_X1 U4058 ( .A(n3298), .ZN(U3221) );
  OR2_X1 U4059 ( .A1(n3299), .A2(n3678), .ZN(n3300) );
  NAND2_X1 U4060 ( .A1(n3300), .A2(n3670), .ZN(n3362) );
  NAND2_X1 U4061 ( .A1(n3767), .A2(n3315), .ZN(n3672) );
  NAND2_X1 U4062 ( .A1(n3362), .A2(n3672), .ZN(n3301) );
  INV_X1 U4063 ( .A(n3767), .ZN(n3307) );
  NAND2_X1 U4064 ( .A1(n3307), .A2(n3466), .ZN(n3682) );
  NAND2_X1 U4065 ( .A1(n3301), .A2(n3682), .ZN(n3399) );
  INV_X1 U4066 ( .A(n3766), .ZN(n3327) );
  NAND2_X1 U4067 ( .A1(n3327), .A2(n3309), .ZN(n3400) );
  NAND2_X1 U4068 ( .A1(n3766), .A2(n3326), .ZN(n3397) );
  XNOR2_X1 U4069 ( .A(n3399), .B(n3617), .ZN(n3313) );
  NAND2_X1 U4070 ( .A1(n3364), .A2(n3304), .ZN(n3305) );
  NAND2_X1 U4071 ( .A1(n3306), .A2(n3305), .ZN(n3361) );
  NOR2_X1 U4072 ( .A1(n3767), .A2(n3466), .ZN(n3308) );
  AOI21_X1 U4073 ( .B1(n3617), .B2(n3328), .A(n2083), .ZN(n3314) );
  AOI22_X1 U4074 ( .A1(n3765), .A2(n4166), .B1(n3309), .B2(n4192), .ZN(n3311)
         );
  NAND2_X1 U4075 ( .A1(n3767), .A2(n4143), .ZN(n3310) );
  OAI211_X1 U4076 ( .C1(n3314), .C2(n4175), .A(n3311), .B(n3310), .ZN(n3312)
         );
  AOI21_X1 U4077 ( .B1(n3313), .B2(n4172), .A(n3312), .ZN(n4271) );
  INV_X1 U4078 ( .A(n3314), .ZN(n4273) );
  OAI21_X1 U4079 ( .B1(n3368), .B2(n3326), .A(n3329), .ZN(n4359) );
  NOR2_X1 U4080 ( .A1(n4359), .A2(n4151), .ZN(n3319) );
  OAI22_X1 U4081 ( .A1(n4183), .A2(n3317), .B1(n3316), .B2(n4180), .ZN(n3318)
         );
  AOI211_X1 U4082 ( .C1(n4273), .C2(n4499), .A(n3319), .B(n3318), .ZN(n3320)
         );
  OAI21_X1 U4083 ( .B1(n4271), .B2(n4368), .A(n3320), .ZN(U3279) );
  INV_X1 U4084 ( .A(n3400), .ZN(n3321) );
  AOI21_X1 U4085 ( .B1(n3399), .B2(n3397), .A(n3321), .ZN(n4162) );
  INV_X1 U4086 ( .A(n3765), .ZN(n4170) );
  NAND2_X1 U4087 ( .A1(n4170), .A2(n3376), .ZN(n4161) );
  NAND2_X1 U4088 ( .A1(n3765), .A2(n3374), .ZN(n4159) );
  NAND2_X1 U4089 ( .A1(n4161), .A2(n4159), .ZN(n3627) );
  XNOR2_X1 U4090 ( .A(n4162), .B(n3627), .ZN(n3325) );
  NAND2_X1 U4091 ( .A1(n3766), .A2(n4143), .ZN(n3323) );
  NAND2_X1 U4092 ( .A1(n4142), .A2(n4166), .ZN(n3322) );
  OAI211_X1 U4093 ( .C1(n4200), .C2(n3374), .A(n3323), .B(n3322), .ZN(n3324)
         );
  AOI21_X1 U4094 ( .B1(n3325), .B2(n4172), .A(n3324), .ZN(n4268) );
  XNOR2_X1 U4095 ( .A(n3375), .B(n3627), .ZN(n4266) );
  NAND2_X1 U4096 ( .A1(n3329), .A2(n3376), .ZN(n3330) );
  NAND2_X1 U4097 ( .A1(n4176), .A2(n3330), .ZN(n4354) );
  NOR2_X1 U4098 ( .A1(n4354), .A2(n4151), .ZN(n3334) );
  OAI22_X1 U4099 ( .A1(n4183), .A2(n3332), .B1(n3331), .B2(n4180), .ZN(n3333)
         );
  AOI211_X1 U4100 ( .C1(n4266), .C2(n4007), .A(n3334), .B(n3333), .ZN(n3335)
         );
  OAI21_X1 U4101 ( .B1(n4368), .B2(n4268), .A(n3335), .ZN(U3278) );
  XNOR2_X1 U4102 ( .A(n3338), .B(n3337), .ZN(n3339) );
  XNOR2_X1 U4103 ( .A(n3336), .B(n3339), .ZN(n3344) );
  NAND2_X1 U4104 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4450) );
  INV_X1 U4105 ( .A(n4450), .ZN(n3340) );
  AOI21_X1 U4106 ( .B1(n3602), .B2(n3764), .A(n3340), .ZN(n3342) );
  AOI22_X1 U4107 ( .A1(n3604), .A2(n4148), .B1(n3603), .B2(n4142), .ZN(n3341)
         );
  OAI211_X1 U4108 ( .C1(n3607), .C2(n4152), .A(n3342), .B(n3341), .ZN(n3343)
         );
  AOI21_X1 U4109 ( .B1(n3344), .B2(n3609), .A(n3343), .ZN(n3345) );
  INV_X1 U4110 ( .A(n3345), .ZN(U3212) );
  INV_X1 U4111 ( .A(n3347), .ZN(n3346) );
  NOR2_X1 U4112 ( .A1(n3292), .A2(n3346), .ZN(n3350) );
  INV_X1 U4113 ( .A(n3292), .ZN(n3348) );
  OAI22_X1 U4114 ( .A1(n3350), .A2(n3349), .B1(n3348), .B2(n3347), .ZN(n3354)
         );
  NAND2_X1 U4115 ( .A1(n3352), .A2(n3351), .ZN(n3353) );
  XNOR2_X1 U4116 ( .A(n3354), .B(n3353), .ZN(n3359) );
  NOR2_X1 U4117 ( .A1(STATE_REG_SCAN_IN), .A2(n3355), .ZN(n4433) );
  AOI21_X1 U4118 ( .B1(n3602), .B2(n4167), .A(n4433), .ZN(n3357) );
  AOI22_X1 U4119 ( .A1(n3604), .A2(n4165), .B1(n3603), .B2(n3765), .ZN(n3356)
         );
  OAI211_X1 U4120 ( .C1(n3607), .C2(n4181), .A(n3357), .B(n3356), .ZN(n3358)
         );
  AOI21_X1 U4121 ( .B1(n3359), .B2(n3609), .A(n3358), .ZN(n3360) );
  INV_X1 U4122 ( .A(n3360), .ZN(U3231) );
  NAND2_X1 U4123 ( .A1(n3682), .A2(n3672), .ZN(n3626) );
  XOR2_X1 U4124 ( .A(n3626), .B(n3361), .Z(n4491) );
  XOR2_X1 U4125 ( .A(n3626), .B(n3362), .Z(n3366) );
  AOI22_X1 U4126 ( .A1(n3766), .A2(n4166), .B1(n4192), .B2(n3466), .ZN(n3363)
         );
  OAI21_X1 U4127 ( .B1(n3364), .B2(n4169), .A(n3363), .ZN(n3365) );
  AOI21_X1 U4128 ( .B1(n3366), .B2(n4172), .A(n3365), .ZN(n4492) );
  INV_X1 U4129 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4739) );
  MUX2_X1 U4130 ( .A(n4492), .B(n4739), .S(n4556), .Z(n3371) );
  INV_X1 U4131 ( .A(n3367), .ZN(n3369) );
  AOI21_X1 U4132 ( .B1(n3466), .B2(n3369), .A(n3368), .ZN(n4497) );
  NAND2_X1 U4133 ( .A1(n4497), .A2(n4330), .ZN(n3370) );
  OAI211_X1 U4134 ( .C1(n4491), .C2(n4341), .A(n3371), .B(n3370), .ZN(U3487)
         );
  INV_X1 U4135 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4405) );
  MUX2_X1 U4136 ( .A(n4492), .B(n4405), .S(n4565), .Z(n3373) );
  NAND2_X1 U4137 ( .A1(n4497), .A2(n4248), .ZN(n3372) );
  OAI211_X1 U4138 ( .C1(n4491), .C2(n4257), .A(n3373), .B(n3372), .ZN(U3528)
         );
  INV_X1 U4139 ( .A(n4142), .ZN(n3377) );
  AOI21_X1 U4140 ( .B1(n3377), .B2(n4178), .A(n4158), .ZN(n3378) );
  INV_X1 U4141 ( .A(n4167), .ZN(n4130) );
  NAND2_X1 U4142 ( .A1(n4130), .A2(n4148), .ZN(n3686) );
  INV_X1 U4143 ( .A(n4148), .ZN(n4138) );
  NAND2_X1 U4144 ( .A1(n4167), .A2(n4138), .ZN(n3674) );
  NAND2_X1 U4145 ( .A1(n3686), .A2(n3674), .ZN(n4136) );
  NAND2_X1 U4146 ( .A1(n3764), .A2(n4126), .ZN(n3379) );
  NAND2_X1 U4147 ( .A1(n4094), .A2(n4110), .ZN(n3730) );
  NAND2_X1 U4148 ( .A1(n4127), .A2(n3380), .ZN(n3694) );
  NAND2_X1 U4149 ( .A1(n3730), .A2(n3694), .ZN(n4100) );
  NAND2_X1 U4150 ( .A1(n4099), .A2(n3381), .ZN(n4083) );
  INV_X1 U4151 ( .A(n4111), .ZN(n4075) );
  NAND2_X1 U4152 ( .A1(n4075), .A2(n3411), .ZN(n3383) );
  INV_X1 U4153 ( .A(n4091), .ZN(n4056) );
  NAND2_X1 U4154 ( .A1(n4056), .A2(n4072), .ZN(n4048) );
  NAND2_X1 U4155 ( .A1(n4091), .A2(n4065), .ZN(n4049) );
  NAND2_X1 U4156 ( .A1(n4048), .A2(n4049), .ZN(n4071) );
  NAND2_X1 U4157 ( .A1(n4063), .A2(n4071), .ZN(n4062) );
  NOR2_X1 U4158 ( .A1(n4073), .A2(n4053), .ZN(n4018) );
  NAND2_X1 U4159 ( .A1(n4054), .A2(n3558), .ZN(n3634) );
  NAND2_X1 U4160 ( .A1(n4073), .A2(n4053), .ZN(n4019) );
  INV_X1 U4161 ( .A(n4054), .ZN(n3384) );
  NAND2_X1 U4162 ( .A1(n3384), .A2(n4035), .ZN(n3635) );
  NAND2_X1 U4163 ( .A1(n3763), .A2(n4009), .ZN(n3385) );
  INV_X1 U4164 ( .A(n3763), .ZN(n4021) );
  INV_X1 U4165 ( .A(n4002), .ZN(n3762) );
  NAND2_X1 U4166 ( .A1(n3762), .A2(n3569), .ZN(n3415) );
  NAND2_X1 U4167 ( .A1(n4002), .A2(n3990), .ZN(n3970) );
  NAND2_X1 U4168 ( .A1(n3415), .A2(n3970), .ZN(n3984) );
  NAND2_X1 U4169 ( .A1(n3983), .A2(n3984), .ZN(n3982) );
  NAND2_X1 U4170 ( .A1(n3944), .A2(n3975), .ZN(n3386) );
  NAND2_X1 U4171 ( .A1(n3973), .A2(n3530), .ZN(n3387) );
  INV_X1 U4172 ( .A(n3946), .ZN(n3906) );
  NAND2_X1 U4173 ( .A1(n3906), .A2(n3926), .ZN(n3388) );
  NAND2_X1 U4174 ( .A1(n3935), .A2(n3913), .ZN(n3389) );
  INV_X1 U4175 ( .A(n3935), .ZN(n3504) );
  NAND2_X1 U4176 ( .A1(n3504), .A2(n3905), .ZN(n3390) );
  NOR2_X1 U4177 ( .A1(n3908), .A2(n3883), .ZN(n3393) );
  NAND2_X1 U4178 ( .A1(n3908), .A2(n3883), .ZN(n3392) );
  NAND2_X1 U4179 ( .A1(n3895), .A2(n3876), .ZN(n3711) );
  NAND2_X1 U4180 ( .A1(n3394), .A2(n3868), .ZN(n3737) );
  NAND2_X1 U4181 ( .A1(n3711), .A2(n3737), .ZN(n3872) );
  AND2_X1 U4182 ( .A1(n3629), .A2(DATAI_29_), .ZN(n3713) );
  XNOR2_X1 U4183 ( .A(n3873), .B(n3713), .ZN(n3421) );
  NAND2_X1 U4184 ( .A1(n4142), .A2(n4178), .ZN(n3396) );
  NAND2_X1 U4185 ( .A1(n4159), .A2(n3396), .ZN(n3401) );
  INV_X1 U4186 ( .A(n3397), .ZN(n3398) );
  NOR2_X1 U4187 ( .A1(n3401), .A2(n3398), .ZN(n3673) );
  NAND2_X1 U4188 ( .A1(n3399), .A2(n3673), .ZN(n3405) );
  NAND2_X1 U4189 ( .A1(n3400), .A2(n4161), .ZN(n3404) );
  INV_X1 U4190 ( .A(n3401), .ZN(n3403) );
  NOR2_X1 U4191 ( .A1(n4142), .A2(n4178), .ZN(n3402) );
  AOI21_X1 U4192 ( .B1(n3404), .B2(n3403), .A(n3402), .ZN(n3687) );
  NAND2_X1 U4193 ( .A1(n3405), .A2(n3687), .ZN(n4134) );
  INV_X1 U4194 ( .A(n4136), .ZN(n3406) );
  NAND2_X1 U4195 ( .A1(n4140), .A2(n4126), .ZN(n3685) );
  NAND2_X1 U4196 ( .A1(n3764), .A2(n3433), .ZN(n3675) );
  NAND2_X1 U4197 ( .A1(n3685), .A2(n3675), .ZN(n4123) );
  INV_X1 U4198 ( .A(n4100), .ZN(n4108) );
  NAND2_X1 U4199 ( .A1(n4109), .A2(n4108), .ZN(n4107) );
  NAND2_X1 U4200 ( .A1(n4073), .A2(n4044), .ZN(n3407) );
  NAND2_X1 U4201 ( .A1(n4049), .A2(n3407), .ZN(n4025) );
  OAI22_X1 U4202 ( .A1(n4025), .A2(n4048), .B1(n4073), .B2(n4044), .ZN(n4026)
         );
  NAND2_X1 U4203 ( .A1(n4075), .A2(n4090), .ZN(n4023) );
  OAI22_X1 U4204 ( .A1(n4025), .A2(n4023), .B1(n4035), .B2(n4054), .ZN(n3408)
         );
  OR2_X1 U4205 ( .A1(n4026), .A2(n3408), .ZN(n3409) );
  NAND2_X1 U4206 ( .A1(n4054), .A2(n4035), .ZN(n3412) );
  NAND2_X1 U4207 ( .A1(n3409), .A2(n3412), .ZN(n3966) );
  OR2_X1 U4208 ( .A1(n3763), .A2(n3416), .ZN(n3968) );
  AND2_X1 U4209 ( .A1(n3968), .A2(n3970), .ZN(n3702) );
  INV_X1 U4210 ( .A(n3410), .ZN(n3732) );
  NAND2_X1 U4211 ( .A1(n4111), .A2(n3411), .ZN(n4022) );
  NAND2_X1 U4212 ( .A1(n4022), .A2(n3412), .ZN(n3413) );
  NOR2_X1 U4213 ( .A1(n4025), .A2(n3413), .ZN(n3964) );
  OR2_X1 U4214 ( .A1(n3732), .A2(n3964), .ZN(n3419) );
  NAND2_X1 U4215 ( .A1(n3987), .A2(n3975), .ZN(n3414) );
  NAND2_X1 U4216 ( .A1(n3415), .A2(n3414), .ZN(n3700) );
  AND2_X1 U4217 ( .A1(n3763), .A2(n3416), .ZN(n3698) );
  AND2_X1 U4218 ( .A1(n3970), .A2(n3698), .ZN(n3417) );
  NOR2_X1 U4219 ( .A1(n3700), .A2(n3417), .ZN(n3418) );
  OR2_X1 U4220 ( .A1(n3973), .A2(n3951), .ZN(n3632) );
  NAND2_X1 U4221 ( .A1(n3944), .A2(n3961), .ZN(n3940) );
  NAND2_X1 U4222 ( .A1(n3946), .A2(n3926), .ZN(n3641) );
  NAND2_X1 U4223 ( .A1(n3973), .A2(n3951), .ZN(n3928) );
  AND2_X1 U4224 ( .A1(n3641), .A2(n3928), .ZN(n3744) );
  NAND2_X1 U4225 ( .A1(n3929), .A2(n3744), .ZN(n3902) );
  OR2_X1 U4226 ( .A1(n3935), .A2(n3905), .ZN(n3640) );
  OR2_X1 U4227 ( .A1(n3946), .A2(n3926), .ZN(n3901) );
  AND2_X1 U4228 ( .A1(n3640), .A2(n3901), .ZN(n3739) );
  NAND2_X1 U4229 ( .A1(n3902), .A2(n3739), .ZN(n3420) );
  NAND2_X1 U4230 ( .A1(n3935), .A2(n3905), .ZN(n3706) );
  XNOR2_X1 U4231 ( .A(n3908), .B(n3893), .ZN(n3889) );
  OR2_X1 U4232 ( .A1(n3908), .A2(n3893), .ZN(n3736) );
  INV_X1 U4233 ( .A(n3737), .ZN(n3710) );
  INV_X1 U4234 ( .A(n3421), .ZN(n3646) );
  XNOR2_X1 U4235 ( .A(n3422), .B(n3646), .ZN(n3423) );
  NAND2_X1 U4236 ( .A1(n3423), .A2(n4172), .ZN(n3432) );
  INV_X1 U4237 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U4238 ( .A1(n2775), .A2(REG1_REG_30__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4239 ( .A1(n3424), .A2(REG0_REG_30__SCAN_IN), .ZN(n3425) );
  OAI211_X1 U4240 ( .C1(n2895), .C2(n3427), .A(n3426), .B(n3425), .ZN(n3761)
         );
  NAND2_X1 U4241 ( .A1(n4377), .A2(B_REG_SCAN_IN), .ZN(n3428) );
  AND2_X1 U4242 ( .A1(n4166), .A2(n3428), .ZN(n4190) );
  NAND2_X1 U4243 ( .A1(n3761), .A2(n4190), .ZN(n3429) );
  OAI21_X1 U4244 ( .B1(n3705), .B2(n4200), .A(n3429), .ZN(n3430) );
  AOI21_X1 U4245 ( .B1(n3895), .B2(n4143), .A(n3430), .ZN(n3431) );
  NAND2_X1 U4246 ( .A1(n4117), .A2(n3433), .ZN(n4118) );
  INV_X1 U4247 ( .A(n3866), .ZN(n3434) );
  NAND2_X1 U4248 ( .A1(n3434), .A2(n3713), .ZN(n3435) );
  OAI21_X1 U4249 ( .B1(n3445), .B2(n4257), .A(n3437), .ZN(U3547) );
  INV_X1 U4250 ( .A(n3438), .ZN(n3439) );
  AOI22_X1 U4251 ( .A1(n3439), .A2(n4498), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4368), .ZN(n3444) );
  NOR2_X1 U4252 ( .A1(n3440), .A2(n4180), .ZN(n3441) );
  OAI21_X1 U4253 ( .B1(n3442), .B2(n3441), .A(n4183), .ZN(n3443) );
  OAI211_X1 U4254 ( .C1(n3445), .C2(n4133), .A(n3444), .B(n3443), .ZN(U3354)
         );
  XNOR2_X1 U4255 ( .A(n3447), .B(n3446), .ZN(n3452) );
  NOR2_X1 U4256 ( .A1(n3887), .A2(n3607), .ZN(n3450) );
  AOI22_X1 U4257 ( .A1(n3935), .A2(n3603), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3448) );
  OAI21_X1 U4258 ( .B1(n3570), .B2(n3893), .A(n3448), .ZN(n3449) );
  AOI211_X1 U4259 ( .C1(n3602), .C2(n3895), .A(n3450), .B(n3449), .ZN(n3451)
         );
  OAI21_X1 U4260 ( .B1(n3452), .B2(n3577), .A(n3451), .ZN(U3211) );
  OAI21_X1 U4261 ( .B1(n3564), .B2(n3455), .A(n3454), .ZN(n3456) );
  NAND3_X1 U4262 ( .A1(n2238), .A2(n3609), .A3(n3456), .ZN(n3460) );
  AOI22_X1 U4263 ( .A1(n3973), .A2(n3602), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3459) );
  AOI22_X1 U4264 ( .A1(n3604), .A2(n3961), .B1(n3762), .B2(n3603), .ZN(n3458)
         );
  OR2_X1 U4265 ( .A1(n3607), .A2(n3962), .ZN(n3457) );
  NAND4_X1 U4266 ( .A1(n3460), .A2(n3459), .A3(n3458), .A4(n3457), .ZN(U3213)
         );
  AND2_X1 U4267 ( .A1(n3263), .A2(n3461), .ZN(n3464) );
  OAI211_X1 U4268 ( .C1(n3464), .C2(n3463), .A(n3609), .B(n3462), .ZN(n3470)
         );
  INV_X1 U4269 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3465) );
  NOR2_X1 U4270 ( .A1(STATE_REG_SCAN_IN), .A2(n3465), .ZN(n4406) );
  AOI21_X1 U4271 ( .B1(n3602), .B2(n3766), .A(n4406), .ZN(n3469) );
  AOI22_X1 U4272 ( .A1(n3604), .A2(n3466), .B1(n3603), .B2(n3768), .ZN(n3468)
         );
  OR2_X1 U4273 ( .A1(n3607), .A2(n4495), .ZN(n3467) );
  NAND4_X1 U4274 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(U3214)
         );
  XNOR2_X1 U4275 ( .A(n3472), .B(n3471), .ZN(n3477) );
  NAND2_X1 U4276 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3858) );
  INV_X1 U4277 ( .A(n3858), .ZN(n3473) );
  AOI21_X1 U4278 ( .B1(n3602), .B2(n4054), .A(n3473), .ZN(n3475) );
  AOI22_X1 U4279 ( .A1(n3604), .A2(n4053), .B1(n3603), .B2(n4091), .ZN(n3474)
         );
  OAI211_X1 U4280 ( .C1(n3607), .C2(n4047), .A(n3475), .B(n3474), .ZN(n3476)
         );
  AOI21_X1 U4281 ( .B1(n3477), .B2(n3609), .A(n3476), .ZN(n3478) );
  INV_X1 U4282 ( .A(n3478), .ZN(U3216) );
  XOR2_X1 U4283 ( .A(n3480), .B(n3479), .Z(n3481) );
  NAND2_X1 U4284 ( .A1(n3481), .A2(n3609), .ZN(n3487) );
  AOI22_X1 U4285 ( .A1(n3603), .A2(n2984), .B1(n3602), .B2(n2447), .ZN(n3486)
         );
  NAND2_X1 U4286 ( .A1(n3482), .A2(REG3_REG_1__SCAN_IN), .ZN(n3485) );
  NAND2_X1 U4287 ( .A1(n3604), .A2(n3483), .ZN(n3484) );
  NAND4_X1 U4288 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(U3219)
         );
  XNOR2_X1 U4289 ( .A(n3489), .B(n3488), .ZN(n3490) );
  XNOR2_X1 U4290 ( .A(n3491), .B(n3490), .ZN(n3496) );
  INV_X1 U4291 ( .A(n3492), .ZN(n4012) );
  AOI22_X1 U4292 ( .A1(n3762), .A2(n3602), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3494) );
  AOI22_X1 U4293 ( .A1(n3604), .A2(n4009), .B1(n3603), .B2(n4054), .ZN(n3493)
         );
  OAI211_X1 U4294 ( .C1(n3607), .C2(n4012), .A(n3494), .B(n3493), .ZN(n3495)
         );
  AOI21_X1 U4295 ( .B1(n3496), .B2(n3609), .A(n3495), .ZN(n3497) );
  INV_X1 U4296 ( .A(n3497), .ZN(U3220) );
  NOR2_X1 U4297 ( .A1(n3499), .A2(n2109), .ZN(n3500) );
  XNOR2_X1 U4298 ( .A(n3501), .B(n3500), .ZN(n3508) );
  INV_X1 U4299 ( .A(n3502), .ZN(n3925) );
  INV_X1 U4300 ( .A(n3973), .ZN(n3927) );
  OAI22_X1 U4301 ( .A1(n3927), .A2(n3571), .B1(n3570), .B2(n3926), .ZN(n3506)
         );
  OAI22_X1 U4302 ( .A1(n3504), .A2(n3568), .B1(STATE_REG_SCAN_IN), .B2(n3503), 
        .ZN(n3505) );
  AOI211_X1 U4303 ( .C1(n3925), .C2(n3574), .A(n3506), .B(n3505), .ZN(n3507)
         );
  OAI21_X1 U4304 ( .B1(n3508), .B2(n3577), .A(n3507), .ZN(U3222) );
  AOI21_X1 U4305 ( .B1(n3599), .B2(n3596), .A(n3598), .ZN(n3509) );
  XOR2_X1 U4306 ( .A(n3510), .B(n3509), .Z(n3514) );
  AND2_X1 U4307 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4464) );
  AOI21_X1 U4308 ( .B1(n3602), .B2(n4111), .A(n4464), .ZN(n3512) );
  AOI22_X1 U4309 ( .A1(n3604), .A2(n4110), .B1(n3603), .B2(n3764), .ZN(n3511)
         );
  OAI211_X1 U4310 ( .C1(n3607), .C2(n4104), .A(n3512), .B(n3511), .ZN(n3513)
         );
  AOI21_X1 U4311 ( .B1(n3514), .B2(n3609), .A(n3513), .ZN(n3515) );
  INV_X1 U4312 ( .A(n3515), .ZN(U3223) );
  XNOR2_X1 U4313 ( .A(n3517), .B(n3516), .ZN(n3518) );
  XNOR2_X1 U4314 ( .A(n3519), .B(n3518), .ZN(n3523) );
  NOR2_X1 U4315 ( .A1(STATE_REG_SCAN_IN), .A2(n4610), .ZN(n3822) );
  AOI21_X1 U4316 ( .B1(n3602), .B2(n4091), .A(n3822), .ZN(n3521) );
  AOI22_X1 U4317 ( .A1(n3604), .A2(n4090), .B1(n3603), .B2(n4127), .ZN(n3520)
         );
  OAI211_X1 U4318 ( .C1(n3607), .C2(n4085), .A(n3521), .B(n3520), .ZN(n3522)
         );
  AOI21_X1 U4319 ( .B1(n3523), .B2(n3609), .A(n3522), .ZN(n3524) );
  INV_X1 U4320 ( .A(n3524), .ZN(U3225) );
  INV_X1 U4321 ( .A(n3525), .ZN(n3526) );
  NOR2_X1 U4322 ( .A1(n3527), .A2(n3526), .ZN(n3529) );
  XNOR2_X1 U4323 ( .A(n3529), .B(n3528), .ZN(n3536) );
  NOR2_X1 U4324 ( .A1(n3607), .A2(n3949), .ZN(n3535) );
  NAND2_X1 U4325 ( .A1(n3946), .A2(n3602), .ZN(n3532) );
  AOI22_X1 U4326 ( .A1(n3604), .A2(n3530), .B1(n3603), .B2(n3987), .ZN(n3531)
         );
  OAI211_X1 U4327 ( .C1(STATE_REG_SCAN_IN), .C2(n3533), .A(n3532), .B(n3531), 
        .ZN(n3534) );
  AOI211_X1 U4328 ( .C1(n3536), .C2(n3609), .A(n3535), .B(n3534), .ZN(n3537)
         );
  INV_X1 U4329 ( .A(n3537), .ZN(U3226) );
  AND2_X1 U4330 ( .A1(n3015), .A2(n3538), .ZN(n3541) );
  OAI211_X1 U4331 ( .C1(n3541), .C2(n3540), .A(n3609), .B(n3539), .ZN(n3549)
         );
  AND2_X1 U4332 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4386) );
  AOI21_X1 U4333 ( .B1(n3602), .B2(n3542), .A(n4386), .ZN(n3548) );
  AOI22_X1 U4334 ( .A1(n3604), .A2(n3544), .B1(n3603), .B2(n3543), .ZN(n3547)
         );
  OR2_X1 U4335 ( .A1(n3607), .A2(n3545), .ZN(n3546) );
  NAND4_X1 U4336 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(U3227)
         );
  INV_X1 U4337 ( .A(n3550), .ZN(n3555) );
  AOI21_X1 U4338 ( .B1(n3554), .B2(n3552), .A(n3551), .ZN(n3553) );
  AOI21_X1 U4339 ( .B1(n3555), .B2(n3554), .A(n3553), .ZN(n3563) );
  NOR2_X1 U4340 ( .A1(n3556), .A2(STATE_REG_SCAN_IN), .ZN(n3557) );
  AOI21_X1 U4341 ( .B1(n3602), .B2(n3763), .A(n3557), .ZN(n3560) );
  AOI22_X1 U4342 ( .A1(n3604), .A2(n3558), .B1(n3603), .B2(n4073), .ZN(n3559)
         );
  OAI211_X1 U4343 ( .C1(n3607), .C2(n4037), .A(n3560), .B(n3559), .ZN(n3561)
         );
  INV_X1 U4344 ( .A(n3561), .ZN(n3562) );
  OAI21_X1 U4345 ( .B1(n3563), .B2(n3577), .A(n3562), .ZN(U3230) );
  AOI21_X1 U4346 ( .B1(n3566), .B2(n3565), .A(n3564), .ZN(n3578) );
  INV_X1 U4347 ( .A(n3991), .ZN(n3575) );
  INV_X1 U4348 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3567) );
  OAI22_X1 U4349 ( .A1(n3568), .A2(n3944), .B1(STATE_REG_SCAN_IN), .B2(n3567), 
        .ZN(n3573) );
  OAI22_X1 U4350 ( .A1(n4021), .A2(n3571), .B1(n3570), .B2(n3569), .ZN(n3572)
         );
  AOI211_X1 U4351 ( .C1(n3575), .C2(n3574), .A(n3573), .B(n3572), .ZN(n3576)
         );
  OAI21_X1 U4352 ( .B1(n3578), .B2(n3577), .A(n3576), .ZN(U3232) );
  INV_X1 U4353 ( .A(n3579), .ZN(n3581) );
  NOR2_X1 U4354 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  XNOR2_X1 U4355 ( .A(n3583), .B(n3582), .ZN(n3587) );
  AND2_X1 U4356 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4478) );
  AOI21_X1 U4357 ( .B1(n3602), .B2(n4073), .A(n4478), .ZN(n3585) );
  AOI22_X1 U4358 ( .A1(n3604), .A2(n4072), .B1(n3603), .B2(n4111), .ZN(n3584)
         );
  OAI211_X1 U4359 ( .C1(n3607), .C2(n4068), .A(n3585), .B(n3584), .ZN(n3586)
         );
  AOI21_X1 U4360 ( .B1(n3587), .B2(n3609), .A(n3586), .ZN(n3588) );
  INV_X1 U4361 ( .A(n3588), .ZN(U3235) );
  INV_X1 U4362 ( .A(n3589), .ZN(n3591) );
  NOR2_X1 U4363 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  AOI22_X1 U4364 ( .A1(n3908), .A2(n3602), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3594) );
  AOI22_X1 U4365 ( .A1(n3946), .A2(n3603), .B1(n3913), .B2(n3604), .ZN(n3593)
         );
  OAI211_X1 U4366 ( .C1(n3607), .C2(n3912), .A(n3594), .B(n3593), .ZN(n3595)
         );
  INV_X1 U4367 ( .A(n3596), .ZN(n3597) );
  NOR2_X1 U4368 ( .A1(n3598), .A2(n3597), .ZN(n3600) );
  XNOR2_X1 U4369 ( .A(n3600), .B(n3599), .ZN(n3610) );
  INV_X1 U4370 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3601) );
  NOR2_X1 U4371 ( .A1(STATE_REG_SCAN_IN), .A2(n3601), .ZN(n4456) );
  AOI21_X1 U4372 ( .B1(n3602), .B2(n4127), .A(n4456), .ZN(n3606) );
  AOI22_X1 U4373 ( .A1(n3604), .A2(n4126), .B1(n3603), .B2(n4167), .ZN(n3605)
         );
  OAI211_X1 U4374 ( .C1(n3607), .C2(n4120), .A(n3606), .B(n3605), .ZN(n3608)
         );
  AOI21_X1 U4375 ( .B1(n3610), .B2(n3609), .A(n3608), .ZN(n3611) );
  INV_X1 U4376 ( .A(n3611), .ZN(U3238) );
  INV_X1 U4377 ( .A(n3612), .ZN(n3613) );
  NOR4_X1 U4378 ( .A1(n3614), .A2(n3613), .A3(n4136), .A4(n4123), .ZN(n3625)
         );
  INV_X1 U4379 ( .A(n3698), .ZN(n3615) );
  INV_X1 U4380 ( .A(n4071), .ZN(n3618) );
  AND4_X1 U4381 ( .A1(n4005), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3624)
         );
  NOR4_X1 U4382 ( .A1(n2985), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3623)
         );
  NOR4_X1 U4383 ( .A1(n3151), .A2(n3984), .A3(n4525), .A4(n4100), .ZN(n3622)
         );
  NAND4_X1 U4384 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3639)
         );
  NAND2_X1 U4385 ( .A1(n4023), .A2(n4022), .ZN(n4087) );
  NOR4_X1 U4386 ( .A1(n4087), .A2(n3628), .A3(n3627), .A4(n3626), .ZN(n3637)
         );
  INV_X1 U4387 ( .A(n4191), .ZN(n3747) );
  NAND2_X1 U4388 ( .A1(n3629), .A2(DATAI_31_), .ZN(n4189) );
  INV_X1 U4389 ( .A(n4189), .ZN(n4193) );
  INV_X1 U4390 ( .A(n3761), .ZN(n3630) );
  AND2_X1 U4391 ( .A1(n3629), .A2(DATAI_30_), .ZN(n4197) );
  NOR2_X1 U4392 ( .A1(n3630), .A2(n4197), .ZN(n3748) );
  AOI21_X1 U4393 ( .B1(n3747), .B2(n4193), .A(n3748), .ZN(n3718) );
  INV_X1 U4394 ( .A(n4019), .ZN(n3631) );
  OR2_X1 U4395 ( .A1(n3631), .A2(n4018), .ZN(n4052) );
  INV_X1 U4396 ( .A(n4052), .ZN(n3633) );
  NAND2_X1 U4397 ( .A1(n3632), .A2(n3928), .ZN(n3942) );
  NOR2_X1 U4398 ( .A1(n3633), .A2(n3942), .ZN(n3636) );
  NAND2_X1 U4399 ( .A1(n3635), .A2(n3634), .ZN(n4028) );
  NAND4_X1 U4400 ( .A1(n3637), .A2(n3718), .A3(n3636), .A4(n4028), .ZN(n3638)
         );
  XNOR2_X1 U4401 ( .A(n4142), .B(n4178), .ZN(n4164) );
  NOR4_X1 U4402 ( .A1(n3889), .A2(n3639), .A3(n3638), .A4(n4164), .ZN(n3648)
         );
  NAND2_X1 U4403 ( .A1(n3706), .A2(n3640), .ZN(n3903) );
  INV_X1 U4404 ( .A(n3903), .ZN(n3644) );
  NAND2_X1 U4405 ( .A1(n3901), .A2(n3641), .ZN(n3931) );
  INV_X1 U4406 ( .A(n3931), .ZN(n3643) );
  XNOR2_X1 U4407 ( .A(n3987), .B(n3975), .ZN(n3958) );
  INV_X1 U4408 ( .A(n3958), .ZN(n3971) );
  NAND2_X1 U4409 ( .A1(n4191), .A2(n4189), .ZN(n3717) );
  INV_X1 U4410 ( .A(n4197), .ZN(n4201) );
  OR2_X1 U4411 ( .A1(n3761), .A2(n4201), .ZN(n3642) );
  AND2_X1 U4412 ( .A1(n3717), .A2(n3642), .ZN(n3740) );
  NAND4_X1 U4413 ( .A1(n3644), .A2(n3643), .A3(n3971), .A4(n3740), .ZN(n3645)
         );
  NOR3_X1 U4414 ( .A1(n3872), .A2(n3646), .A3(n3645), .ZN(n3647) );
  AOI21_X1 U4415 ( .B1(n3648), .B2(n3647), .A(n3652), .ZN(n3722) );
  OAI211_X1 U4416 ( .C1(n2150), .C2(n3652), .A(n3651), .B(n3650), .ZN(n3654)
         );
  NAND3_X1 U4417 ( .A1(n3654), .A2(n3653), .A3(n3037), .ZN(n3657) );
  NAND3_X1 U4418 ( .A1(n3657), .A2(n3656), .A3(n3655), .ZN(n3660) );
  NAND3_X1 U4419 ( .A1(n3660), .A2(n3659), .A3(n3658), .ZN(n3663) );
  NAND4_X1 U4420 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3677), .ZN(n3666)
         );
  AND3_X1 U4421 ( .A1(n3666), .A2(n3665), .A3(n3664), .ZN(n3671) );
  NAND2_X1 U4422 ( .A1(n3668), .A2(n3667), .ZN(n3680) );
  OAI211_X1 U4423 ( .C1(n3671), .C2(n3680), .A(n3670), .B(n3669), .ZN(n3693)
         );
  NAND2_X1 U4424 ( .A1(n3673), .A2(n3672), .ZN(n3689) );
  NAND2_X1 U4425 ( .A1(n3675), .A2(n3674), .ZN(n3676) );
  NOR3_X1 U4426 ( .A1(n3689), .A2(n3678), .A3(n3676), .ZN(n3692) );
  NAND2_X1 U4427 ( .A1(n3676), .A2(n3685), .ZN(n3727) );
  INV_X1 U4428 ( .A(n3677), .ZN(n3681) );
  NOR4_X1 U4429 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3684)
         );
  INV_X1 U4430 ( .A(n3682), .ZN(n3683) );
  NOR2_X1 U4431 ( .A1(n3684), .A2(n3683), .ZN(n3690) );
  NAND2_X1 U4432 ( .A1(n3686), .A2(n3685), .ZN(n3728) );
  INV_X1 U4433 ( .A(n3728), .ZN(n3688) );
  OAI211_X1 U4434 ( .C1(n3690), .C2(n3689), .A(n3688), .B(n3687), .ZN(n3691)
         );
  AOI22_X1 U4435 ( .A1(n3693), .A2(n3692), .B1(n3727), .B2(n3691), .ZN(n3695)
         );
  OAI21_X1 U4436 ( .B1(n3695), .B2(n2132), .A(n3730), .ZN(n3697) );
  INV_X1 U4437 ( .A(n3966), .ZN(n3696) );
  AOI21_X1 U4438 ( .B1(n3697), .B2(n3964), .A(n3696), .ZN(n3699) );
  OR2_X1 U4439 ( .A1(n3699), .A2(n3698), .ZN(n3701) );
  AOI21_X1 U4440 ( .B1(n3702), .B2(n3701), .A(n3700), .ZN(n3703) );
  OAI21_X1 U4441 ( .B1(n3703), .B2(n2128), .A(n3744), .ZN(n3708) );
  INV_X1 U4442 ( .A(n3908), .ZN(n3704) );
  NOR2_X1 U4443 ( .A1(n3704), .A2(n3883), .ZN(n3707) );
  NAND2_X1 U4444 ( .A1(n3873), .A2(n3705), .ZN(n3712) );
  NAND3_X1 U4445 ( .A1(n3712), .A2(n3711), .A3(n3706), .ZN(n3723) );
  AOI211_X1 U4446 ( .C1(n3739), .C2(n3708), .A(n3707), .B(n3723), .ZN(n3720)
         );
  INV_X1 U4447 ( .A(n3736), .ZN(n3709) );
  NOR2_X1 U4448 ( .A1(n3710), .A2(n3709), .ZN(n3716) );
  NAND2_X1 U4449 ( .A1(n3712), .A2(n3711), .ZN(n3715) );
  INV_X1 U4450 ( .A(n3873), .ZN(n3714) );
  NAND2_X1 U4451 ( .A1(n3714), .A2(n3713), .ZN(n3738) );
  OAI211_X1 U4452 ( .C1(n3716), .C2(n3715), .A(n3740), .B(n3738), .ZN(n3724)
         );
  INV_X1 U4453 ( .A(n3717), .ZN(n3719) );
  OAI22_X1 U4454 ( .A1(n3720), .A2(n3724), .B1(n3719), .B2(n3718), .ZN(n3721)
         );
  MUX2_X1 U4455 ( .A(n3722), .B(n3721), .S(n2374), .Z(n3753) );
  INV_X1 U4456 ( .A(n3889), .ZN(n3726) );
  INV_X1 U4457 ( .A(n3723), .ZN(n3725) );
  AOI21_X1 U4458 ( .B1(n3726), .B2(n3725), .A(n3724), .ZN(n3746) );
  OAI21_X1 U4459 ( .B1(n4134), .B2(n3728), .A(n3727), .ZN(n3729) );
  AOI21_X1 U4460 ( .B1(n3730), .B2(n3729), .A(n2132), .ZN(n3733) );
  OAI21_X1 U4461 ( .B1(n3733), .B2(n3732), .A(n3731), .ZN(n3735) );
  NAND2_X1 U4462 ( .A1(n3735), .A2(n3734), .ZN(n3743) );
  NAND4_X1 U4463 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3742)
         );
  INV_X1 U4464 ( .A(n3740), .ZN(n3741) );
  AOI211_X1 U4465 ( .C1(n3744), .C2(n3743), .A(n3742), .B(n3741), .ZN(n3745)
         );
  OAI22_X1 U4466 ( .A1(n3746), .A2(n3745), .B1(n4191), .B2(n4201), .ZN(n3751)
         );
  OAI21_X1 U4467 ( .B1(n3748), .B2(n3747), .A(n4193), .ZN(n3750) );
  AOI21_X1 U4468 ( .B1(n3751), .B2(n3750), .A(n3749), .ZN(n3752) );
  NOR2_X1 U4469 ( .A1(n3753), .A2(n3752), .ZN(n3754) );
  XNOR2_X1 U4470 ( .A(n3754), .B(n3850), .ZN(n3760) );
  NOR2_X1 U4471 ( .A1(n3755), .A2(n3802), .ZN(n3758) );
  OAI21_X1 U4472 ( .B1(n3759), .B2(n3756), .A(B_REG_SCAN_IN), .ZN(n3757) );
  OAI22_X1 U4473 ( .A1(n3760), .A2(n3759), .B1(n3758), .B2(n3757), .ZN(U3239)
         );
  MUX2_X1 U4474 ( .A(DATAO_REG_30__SCAN_IN), .B(n3761), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4475 ( .A(n3873), .B(DATAO_REG_29__SCAN_IN), .S(n3772), .Z(U3579)
         );
  MUX2_X1 U4476 ( .A(n3895), .B(DATAO_REG_28__SCAN_IN), .S(n3772), .Z(U3578)
         );
  MUX2_X1 U4477 ( .A(DATAO_REG_26__SCAN_IN), .B(n3935), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4478 ( .A(n3946), .B(DATAO_REG_25__SCAN_IN), .S(n3772), .Z(U3575)
         );
  MUX2_X1 U4479 ( .A(n3973), .B(DATAO_REG_24__SCAN_IN), .S(n3772), .Z(U3574)
         );
  MUX2_X1 U4480 ( .A(DATAO_REG_22__SCAN_IN), .B(n3762), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4481 ( .A(n3763), .B(DATAO_REG_21__SCAN_IN), .S(n3772), .Z(U3571)
         );
  MUX2_X1 U4482 ( .A(n4054), .B(DATAO_REG_20__SCAN_IN), .S(n3772), .Z(U3570)
         );
  MUX2_X1 U4483 ( .A(n4073), .B(DATAO_REG_19__SCAN_IN), .S(n3772), .Z(U3569)
         );
  MUX2_X1 U4484 ( .A(n4091), .B(DATAO_REG_18__SCAN_IN), .S(n3772), .Z(U3568)
         );
  MUX2_X1 U4485 ( .A(n4111), .B(DATAO_REG_17__SCAN_IN), .S(n3772), .Z(U3567)
         );
  MUX2_X1 U4486 ( .A(n4127), .B(DATAO_REG_16__SCAN_IN), .S(n3772), .Z(U3566)
         );
  MUX2_X1 U4487 ( .A(n3764), .B(DATAO_REG_15__SCAN_IN), .S(n3772), .Z(U3565)
         );
  MUX2_X1 U4488 ( .A(n4167), .B(DATAO_REG_14__SCAN_IN), .S(n3772), .Z(U3564)
         );
  MUX2_X1 U4489 ( .A(n4142), .B(DATAO_REG_13__SCAN_IN), .S(n3772), .Z(U3563)
         );
  MUX2_X1 U4490 ( .A(n3765), .B(DATAO_REG_12__SCAN_IN), .S(n3772), .Z(U3562)
         );
  MUX2_X1 U4491 ( .A(n3766), .B(DATAO_REG_11__SCAN_IN), .S(n3772), .Z(U3561)
         );
  MUX2_X1 U4492 ( .A(n3767), .B(DATAO_REG_10__SCAN_IN), .S(n3772), .Z(U3560)
         );
  MUX2_X1 U4493 ( .A(n3768), .B(DATAO_REG_9__SCAN_IN), .S(n3772), .Z(U3559) );
  MUX2_X1 U4494 ( .A(n3769), .B(DATAO_REG_8__SCAN_IN), .S(n3772), .Z(U3558) );
  MUX2_X1 U4495 ( .A(n3770), .B(DATAO_REG_7__SCAN_IN), .S(n3772), .Z(U3557) );
  MUX2_X1 U4496 ( .A(n3771), .B(DATAO_REG_4__SCAN_IN), .S(n3772), .Z(U3554) );
  MUX2_X1 U4497 ( .A(n3773), .B(DATAO_REG_1__SCAN_IN), .S(n3772), .Z(U3551) );
  AOI22_X1 U4498 ( .A1(n4457), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3787) );
  OAI211_X1 U4499 ( .C1(n3776), .C2(n3775), .A(n4471), .B(n3774), .ZN(n3786)
         );
  INV_X1 U4500 ( .A(n4490), .ZN(n4449) );
  NAND2_X1 U4501 ( .A1(n4449), .A2(n3777), .ZN(n3785) );
  MUX2_X1 U4502 ( .A(REG2_REG_1__SCAN_IN), .B(n3779), .S(n3778), .Z(n3781) );
  NAND2_X1 U4503 ( .A1(n3781), .A2(n3780), .ZN(n3782) );
  NAND3_X1 U4504 ( .A1(n4487), .A2(n3783), .A3(n3782), .ZN(n3784) );
  NAND4_X1 U4505 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(U3241)
         );
  XNOR2_X1 U4506 ( .A(n3789), .B(n3788), .ZN(n3790) );
  NOR2_X1 U4507 ( .A1(n4443), .A2(n3790), .ZN(n3797) );
  INV_X1 U4508 ( .A(n3791), .ZN(n3795) );
  MUX2_X1 U4509 ( .A(n2910), .B(REG1_REG_2__SCAN_IN), .S(n4365), .Z(n3794) );
  AOI211_X1 U4510 ( .C1(n3795), .C2(n3794), .A(n3793), .B(n4475), .ZN(n3796)
         );
  AOI211_X1 U4511 ( .C1(n4449), .C2(n4365), .A(n3797), .B(n3796), .ZN(n3808)
         );
  NAND3_X1 U4512 ( .A1(n3800), .A2(n3799), .A3(n3798), .ZN(n3806) );
  INV_X1 U4513 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3801) );
  AOI21_X1 U4514 ( .B1(n4377), .B2(n3801), .A(n4367), .ZN(n4376) );
  INV_X1 U4515 ( .A(n3802), .ZN(n3803) );
  NAND2_X1 U4516 ( .A1(n3803), .A2(REG2_REG_0__SCAN_IN), .ZN(n3804) );
  MUX2_X1 U4517 ( .A(n4376), .B(n3804), .S(IR_REG_0__SCAN_IN), .Z(n3805) );
  NAND3_X1 U4518 ( .A1(n3806), .A2(U4043), .A3(n3805), .ZN(n4391) );
  AOI22_X1 U4519 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4457), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3807) );
  NAND3_X1 U4520 ( .A1(n3808), .A2(n4391), .A3(n3807), .ZN(U3242) );
  XNOR2_X1 U4521 ( .A(n3823), .B(REG1_REG_17__SCAN_IN), .ZN(n3820) );
  INV_X1 U4522 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4566) );
  INV_X1 U4523 ( .A(n3825), .ZN(n4522) );
  AOI22_X1 U4524 ( .A1(n3825), .A2(n4566), .B1(REG1_REG_9__SCAN_IN), .B2(n4522), .ZN(n4394) );
  INV_X1 U4525 ( .A(n3830), .ZN(n4520) );
  NOR2_X1 U4526 ( .A1(n3812), .A2(n4520), .ZN(n3813) );
  INV_X1 U4527 ( .A(n3824), .ZN(n4518) );
  INV_X1 U4528 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4274) );
  AOI22_X1 U4529 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4518), .B1(n3824), .B2(
        n4274), .ZN(n4413) );
  NOR2_X1 U4530 ( .A1(n3814), .A2(n4516), .ZN(n3815) );
  INV_X1 U4531 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4423) );
  INV_X1 U4532 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4264) );
  AOI22_X1 U4533 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4514), .B1(n3837), .B2(
        n4264), .ZN(n4431) );
  INV_X1 U4534 ( .A(n4448), .ZN(n4513) );
  INV_X1 U4535 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4442) );
  XOR2_X1 U4536 ( .A(n4448), .B(n3816), .Z(n4441) );
  INV_X1 U4537 ( .A(n3839), .ZN(n4511) );
  INV_X1 U4538 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U4539 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4511), .B1(n3839), .B2(
        n4255), .ZN(n4454) );
  NAND2_X1 U4540 ( .A1(n3817), .A2(n4510), .ZN(n3818) );
  INV_X1 U4541 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4468) );
  OAI21_X1 U4542 ( .B1(n3820), .B2(n3819), .A(n3849), .ZN(n3821) );
  AOI22_X1 U4543 ( .A1(n3855), .A2(n4449), .B1(n4471), .B2(n3821), .ZN(n3847)
         );
  AOI21_X1 U4544 ( .B1(n4457), .B2(ADDR_REG_17__SCAN_IN), .A(n3822), .ZN(n3846) );
  XNOR2_X1 U4545 ( .A(n3823), .B(REG2_REG_17__SCAN_IN), .ZN(n3843) );
  NOR2_X1 U4546 ( .A1(n4182), .A2(n4514), .ZN(n4434) );
  NAND2_X1 U4547 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3824), .ZN(n3833) );
  AOI22_X1 U4548 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3824), .B1(n4518), .B2(
        n3317), .ZN(n4418) );
  AOI22_X1 U4549 ( .A1(n3825), .A2(REG2_REG_9__SCAN_IN), .B1(n3237), .B2(n4522), .ZN(n4400) );
  NAND2_X1 U4550 ( .A1(n4400), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U4551 ( .A1(n3830), .A2(n3831), .ZN(n3832) );
  NAND2_X1 U4552 ( .A1(n4418), .A2(n4417), .ZN(n4416) );
  NAND2_X1 U4553 ( .A1(n3834), .A2(n3835), .ZN(n3836) );
  NOR2_X1 U4554 ( .A1(n4153), .A2(n4445), .ZN(n4444) );
  AOI22_X1 U4555 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4511), .B1(n3839), .B2(
        n4121), .ZN(n4460) );
  NAND2_X1 U4556 ( .A1(n3840), .A2(n4510), .ZN(n3841) );
  NAND2_X1 U4557 ( .A1(n4466), .A2(n4105), .ZN(n4465) );
  OAI21_X1 U4558 ( .B1(n3843), .B2(n3842), .A(n3854), .ZN(n3844) );
  NAND2_X1 U4559 ( .A1(n4487), .A2(n3844), .ZN(n3845) );
  NAND3_X1 U4560 ( .A1(n3847), .A2(n3846), .A3(n3845), .ZN(U3257) );
  INV_X1 U4561 ( .A(n3856), .ZN(n4508) );
  INV_X1 U4562 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4563 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4508), .B1(n3856), .B2(
        n3848), .ZN(n4476) );
  XNOR2_X1 U4564 ( .A(n3850), .B(REG1_REG_19__SCAN_IN), .ZN(n3851) );
  XNOR2_X1 U4565 ( .A(n3852), .B(n3851), .ZN(n3864) );
  NAND2_X1 U4566 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3856), .ZN(n3853) );
  OAI21_X1 U4567 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3856), .A(n3853), .ZN(n4485) );
  MUX2_X1 U4568 ( .A(n4059), .B(REG2_REG_19__SCAN_IN), .S(n3860), .Z(n3857) );
  NAND2_X1 U4569 ( .A1(n4457), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3859) );
  OAI211_X1 U4570 ( .C1(n4490), .C2(n3860), .A(n3859), .B(n3858), .ZN(n3861)
         );
  AOI21_X1 U4571 ( .B1(n3862), .B2(n4487), .A(n3861), .ZN(n3863) );
  OAI21_X1 U4572 ( .B1(n3864), .B2(n4475), .A(n3863), .ZN(U3259) );
  XNOR2_X1 U4573 ( .A(n3865), .B(n3872), .ZN(n4287) );
  INV_X1 U4574 ( .A(n3885), .ZN(n3867) );
  AOI21_X1 U4575 ( .B1(n3868), .B2(n3867), .A(n3866), .ZN(n4285) );
  INV_X1 U4576 ( .A(n3869), .ZN(n3870) );
  AOI22_X1 U4577 ( .A1(n4285), .A2(n4498), .B1(n3870), .B2(n4496), .ZN(n3881)
         );
  XOR2_X1 U4578 ( .A(n3872), .B(n3871), .Z(n3878) );
  NAND2_X1 U4579 ( .A1(n3908), .A2(n4143), .ZN(n3875) );
  NAND2_X1 U4580 ( .A1(n3873), .A2(n4166), .ZN(n3874) );
  OAI211_X1 U4581 ( .C1(n3876), .C2(n4200), .A(n3875), .B(n3874), .ZN(n3877)
         );
  AOI21_X1 U4582 ( .B1(n3878), .B2(n4172), .A(n3877), .ZN(n4205) );
  MUX2_X1 U4583 ( .A(n3879), .B(n4205), .S(n4373), .Z(n3880) );
  OAI211_X1 U4584 ( .C1(n4287), .C2(n4133), .A(n3881), .B(n3880), .ZN(U3262)
         );
  XOR2_X1 U4585 ( .A(n3889), .B(n3882), .Z(n4291) );
  AND2_X1 U4586 ( .A1(n3915), .A2(n3883), .ZN(n3884) );
  NOR2_X1 U4587 ( .A1(n3885), .A2(n3884), .ZN(n4209) );
  OAI22_X1 U4588 ( .A1(n3887), .A2(n4180), .B1(n3886), .B2(n4373), .ZN(n3888)
         );
  AOI21_X1 U4589 ( .B1(n4209), .B2(n4498), .A(n3888), .ZN(n3899) );
  XNOR2_X1 U4590 ( .A(n3890), .B(n3889), .ZN(n3891) );
  NAND2_X1 U4591 ( .A1(n3891), .A2(n4172), .ZN(n3897) );
  NAND2_X1 U4592 ( .A1(n3935), .A2(n4143), .ZN(n3892) );
  OAI21_X1 U4593 ( .B1(n4200), .B2(n3893), .A(n3892), .ZN(n3894) );
  AOI21_X1 U4594 ( .B1(n3895), .B2(n4166), .A(n3894), .ZN(n3896) );
  NAND2_X1 U4595 ( .A1(n3897), .A2(n3896), .ZN(n4208) );
  NAND2_X1 U4596 ( .A1(n4208), .A2(n4373), .ZN(n3898) );
  OAI211_X1 U4597 ( .C1(n4291), .C2(n4133), .A(n3899), .B(n3898), .ZN(U3263)
         );
  XNOR2_X1 U4598 ( .A(n3900), .B(n3903), .ZN(n4213) );
  INV_X1 U4599 ( .A(n4213), .ZN(n3919) );
  NAND2_X1 U4600 ( .A1(n3902), .A2(n3901), .ZN(n3904) );
  XNOR2_X1 U4601 ( .A(n3904), .B(n3903), .ZN(n3910) );
  OAI22_X1 U4602 ( .A1(n3906), .A2(n4169), .B1(n3905), .B2(n4200), .ZN(n3907)
         );
  AOI21_X1 U4603 ( .B1(n4166), .B2(n3908), .A(n3907), .ZN(n3909) );
  OAI21_X1 U4604 ( .B1(n3910), .B2(n4147), .A(n3909), .ZN(n4212) );
  OAI22_X1 U4605 ( .A1(n3912), .A2(n4180), .B1(n3911), .B2(n4183), .ZN(n3917)
         );
  NAND2_X1 U4606 ( .A1(n3921), .A2(n3913), .ZN(n3914) );
  NAND2_X1 U4607 ( .A1(n3915), .A2(n3914), .ZN(n4295) );
  NOR2_X1 U4608 ( .A1(n4295), .A2(n4151), .ZN(n3916) );
  AOI211_X1 U4609 ( .C1(n4373), .C2(n4212), .A(n3917), .B(n3916), .ZN(n3918)
         );
  OAI21_X1 U4610 ( .B1(n3919), .B2(n4133), .A(n3918), .ZN(U3264) );
  XNOR2_X1 U4611 ( .A(n3920), .B(n3931), .ZN(n4300) );
  INV_X1 U4612 ( .A(n3953), .ZN(n3923) );
  INV_X1 U4613 ( .A(n3921), .ZN(n3922) );
  AOI21_X1 U4614 ( .B1(n3924), .B2(n3923), .A(n3922), .ZN(n4298) );
  AOI22_X1 U4615 ( .A1(n4298), .A2(n4498), .B1(n3925), .B2(n4496), .ZN(n3938)
         );
  OAI22_X1 U4616 ( .A1(n3927), .A2(n4169), .B1(n3926), .B2(n4200), .ZN(n3934)
         );
  NAND2_X1 U4617 ( .A1(n3929), .A2(n3928), .ZN(n3930) );
  XOR2_X1 U4618 ( .A(n3931), .B(n3930), .Z(n3932) );
  NOR2_X1 U4619 ( .A1(n3932), .A2(n4147), .ZN(n3933) );
  AOI211_X1 U4620 ( .C1(n4166), .C2(n3935), .A(n3934), .B(n3933), .ZN(n4216)
         );
  MUX2_X1 U4621 ( .A(n3936), .B(n4216), .S(n4183), .Z(n3937) );
  OAI211_X1 U4622 ( .C1(n4300), .C2(n4133), .A(n3938), .B(n3937), .ZN(U3265)
         );
  XNOR2_X1 U4623 ( .A(n3939), .B(n3942), .ZN(n4220) );
  INV_X1 U4624 ( .A(n4220), .ZN(n3957) );
  NAND2_X1 U4625 ( .A1(n3941), .A2(n3940), .ZN(n3943) );
  XNOR2_X1 U4626 ( .A(n3943), .B(n3942), .ZN(n3948) );
  OAI22_X1 U4627 ( .A1(n3944), .A2(n4169), .B1(n4200), .B2(n3951), .ZN(n3945)
         );
  AOI21_X1 U4628 ( .B1(n3946), .B2(n4166), .A(n3945), .ZN(n3947) );
  OAI21_X1 U4629 ( .B1(n3948), .B2(n4147), .A(n3947), .ZN(n4219) );
  OAI22_X1 U4630 ( .A1(n4183), .A2(n3950), .B1(n3949), .B2(n4180), .ZN(n3955)
         );
  NOR2_X1 U4631 ( .A1(n3960), .A2(n3951), .ZN(n3952) );
  NOR2_X1 U4632 ( .A1(n4304), .A2(n4151), .ZN(n3954) );
  AOI211_X1 U4633 ( .C1(n4373), .C2(n4219), .A(n3955), .B(n3954), .ZN(n3956)
         );
  OAI21_X1 U4634 ( .B1(n3957), .B2(n4133), .A(n3956), .ZN(U3266) );
  XNOR2_X1 U4635 ( .A(n3959), .B(n3958), .ZN(n4309) );
  INV_X1 U4636 ( .A(n3996), .ZN(n4227) );
  AOI21_X1 U4637 ( .B1(n3961), .B2(n4227), .A(n3960), .ZN(n4307) );
  INV_X1 U4638 ( .A(n3962), .ZN(n3963) );
  AOI22_X1 U4639 ( .A1(n4307), .A2(n4498), .B1(n3963), .B2(n4496), .ZN(n3981)
         );
  INV_X1 U4640 ( .A(n3964), .ZN(n3965) );
  OR2_X1 U4641 ( .A1(n4088), .A2(n3965), .ZN(n3967) );
  NAND2_X1 U4642 ( .A1(n3967), .A2(n3966), .ZN(n3999) );
  INV_X1 U4643 ( .A(n3968), .ZN(n3969) );
  AOI21_X1 U4644 ( .B1(n3999), .B2(n4005), .A(n3969), .ZN(n3985) );
  OAI21_X1 U4645 ( .B1(n3985), .B2(n3984), .A(n3970), .ZN(n3972) );
  XNOR2_X1 U4646 ( .A(n3972), .B(n3971), .ZN(n3978) );
  NOR2_X1 U4647 ( .A1(n4002), .A2(n4169), .ZN(n3977) );
  NAND2_X1 U4648 ( .A1(n3973), .A2(n4166), .ZN(n3974) );
  OAI21_X1 U4649 ( .B1(n4200), .B2(n3975), .A(n3974), .ZN(n3976) );
  AOI211_X1 U4650 ( .C1(n3978), .C2(n4172), .A(n3977), .B(n3976), .ZN(n4223)
         );
  MUX2_X1 U4651 ( .A(n3979), .B(n4223), .S(n4373), .Z(n3980) );
  OAI211_X1 U4652 ( .C1(n4309), .C2(n4133), .A(n3981), .B(n3980), .ZN(U3267)
         );
  OAI21_X1 U4653 ( .B1(n3983), .B2(n3984), .A(n3982), .ZN(n4313) );
  XNOR2_X1 U4654 ( .A(n3985), .B(n3984), .ZN(n3986) );
  NAND2_X1 U4655 ( .A1(n3986), .A2(n4172), .ZN(n3989) );
  AOI22_X1 U4656 ( .A1(n3987), .A2(n4166), .B1(n3990), .B2(n4192), .ZN(n3988)
         );
  OAI211_X1 U4657 ( .C1(n4021), .C2(n4169), .A(n3989), .B(n3988), .ZN(n4229)
         );
  NAND2_X1 U4658 ( .A1(n4011), .A2(n3990), .ZN(n4226) );
  NAND2_X1 U4659 ( .A1(n4226), .A2(n4498), .ZN(n3995) );
  OAI22_X1 U4660 ( .A1(n4183), .A2(n3992), .B1(n3991), .B2(n4180), .ZN(n3993)
         );
  INV_X1 U4661 ( .A(n3993), .ZN(n3994) );
  OAI21_X1 U4662 ( .B1(n3996), .B2(n3995), .A(n3994), .ZN(n3997) );
  AOI21_X1 U4663 ( .B1(n4229), .B2(n4183), .A(n3997), .ZN(n3998) );
  OAI21_X1 U4664 ( .B1(n4313), .B2(n4133), .A(n3998), .ZN(U3268) );
  XNOR2_X1 U4665 ( .A(n3999), .B(n4005), .ZN(n4004) );
  NAND2_X1 U4666 ( .A1(n4009), .A2(n4192), .ZN(n4001) );
  NAND2_X1 U4667 ( .A1(n4054), .A2(n4143), .ZN(n4000) );
  OAI211_X1 U4668 ( .C1(n4002), .C2(n4139), .A(n4001), .B(n4000), .ZN(n4003)
         );
  AOI21_X1 U4669 ( .B1(n4004), .B2(n4172), .A(n4003), .ZN(n4232) );
  XNOR2_X1 U4670 ( .A(n4006), .B(n4005), .ZN(n4317) );
  INV_X1 U4671 ( .A(n4317), .ZN(n4008) );
  NAND2_X1 U4672 ( .A1(n4008), .A2(n4007), .ZN(n4017) );
  NAND2_X1 U4673 ( .A1(n4034), .A2(n4009), .ZN(n4010) );
  NAND2_X1 U4674 ( .A1(n4011), .A2(n4010), .ZN(n4233) );
  INV_X1 U4675 ( .A(n4233), .ZN(n4015) );
  OAI22_X1 U4676 ( .A1(n4183), .A2(n4013), .B1(n4012), .B2(n4180), .ZN(n4014)
         );
  AOI21_X1 U4677 ( .B1(n4015), .B2(n4498), .A(n4014), .ZN(n4016) );
  OAI211_X1 U4678 ( .C1(n4368), .C2(n4232), .A(n4017), .B(n4016), .ZN(U3269)
         );
  AOI21_X1 U4679 ( .B1(n4043), .B2(n4019), .A(n4018), .ZN(n4020) );
  XOR2_X1 U4680 ( .A(n4028), .B(n4020), .Z(n4236) );
  OAI22_X1 U4681 ( .A1(n4021), .A2(n4139), .B1(n4200), .B2(n4035), .ZN(n4032)
         );
  INV_X1 U4682 ( .A(n4022), .ZN(n4024) );
  OAI21_X1 U4683 ( .B1(n4088), .B2(n4024), .A(n4023), .ZN(n4070) );
  INV_X1 U4684 ( .A(n4025), .ZN(n4027) );
  AOI21_X1 U4685 ( .B1(n4070), .B2(n4027), .A(n4026), .ZN(n4029) );
  XNOR2_X1 U4686 ( .A(n4029), .B(n4028), .ZN(n4030) );
  NOR2_X1 U4687 ( .A1(n4030), .A2(n4147), .ZN(n4031) );
  AOI211_X1 U4688 ( .C1(n4143), .C2(n4073), .A(n4032), .B(n4031), .ZN(n4033)
         );
  OAI21_X1 U4689 ( .B1(n4236), .B2(n4175), .A(n4033), .ZN(n4237) );
  NAND2_X1 U4690 ( .A1(n4237), .A2(n4373), .ZN(n4042) );
  INV_X1 U4691 ( .A(n4046), .ZN(n4036) );
  OAI21_X1 U4692 ( .B1(n4036), .B2(n4035), .A(n4034), .ZN(n4320) );
  INV_X1 U4693 ( .A(n4320), .ZN(n4040) );
  OAI22_X1 U4694 ( .A1(n4183), .A2(n4038), .B1(n4037), .B2(n4180), .ZN(n4039)
         );
  AOI21_X1 U4695 ( .B1(n4040), .B2(n4498), .A(n4039), .ZN(n4041) );
  OAI211_X1 U4696 ( .C1(n4236), .C2(n4188), .A(n4042), .B(n4041), .ZN(U3270)
         );
  XNOR2_X1 U4697 ( .A(n4043), .B(n4052), .ZN(n4326) );
  OR2_X1 U4698 ( .A1(n4066), .A2(n4044), .ZN(n4045) );
  AND2_X1 U4699 ( .A1(n4046), .A2(n4045), .ZN(n4324) );
  AOI22_X1 U4700 ( .A1(n4324), .A2(n4498), .B1(n2147), .B2(n4496), .ZN(n4061)
         );
  INV_X1 U4701 ( .A(n4048), .ZN(n4050) );
  OAI21_X1 U4702 ( .B1(n4070), .B2(n4050), .A(n4049), .ZN(n4051) );
  XOR2_X1 U4703 ( .A(n4052), .B(n4051), .Z(n4058) );
  AOI22_X1 U4704 ( .A1(n4054), .A2(n4166), .B1(n4192), .B2(n4053), .ZN(n4055)
         );
  OAI21_X1 U4705 ( .B1(n4056), .B2(n4169), .A(n4055), .ZN(n4057) );
  AOI21_X1 U4706 ( .B1(n4058), .B2(n4172), .A(n4057), .ZN(n4321) );
  MUX2_X1 U4707 ( .A(n4059), .B(n4321), .S(n4373), .Z(n4060) );
  OAI211_X1 U4708 ( .C1(n4326), .C2(n4133), .A(n4061), .B(n4060), .ZN(U3271)
         );
  OAI21_X1 U4709 ( .B1(n4063), .B2(n4071), .A(n4062), .ZN(n4064) );
  INV_X1 U4710 ( .A(n4064), .ZN(n4246) );
  OAI21_X1 U4711 ( .B1(n4084), .B2(n4065), .A(n4551), .ZN(n4067) );
  OR2_X1 U4712 ( .A1(n4067), .A2(n4066), .ZN(n4243) );
  INV_X1 U4713 ( .A(n4243), .ZN(n4081) );
  OAI22_X1 U4714 ( .A1(n4183), .A2(n4069), .B1(n4068), .B2(n4180), .ZN(n4079)
         );
  XOR2_X1 U4715 ( .A(n4071), .B(n4070), .Z(n4077) );
  AOI22_X1 U4716 ( .A1(n4073), .A2(n4166), .B1(n4072), .B2(n4192), .ZN(n4074)
         );
  OAI21_X1 U4717 ( .B1(n4075), .B2(n4169), .A(n4074), .ZN(n4076) );
  AOI21_X1 U4718 ( .B1(n4077), .B2(n4172), .A(n4076), .ZN(n4244) );
  NOR2_X1 U4719 ( .A1(n4244), .A2(n4368), .ZN(n4078) );
  AOI211_X1 U4720 ( .C1(n4081), .C2(n4080), .A(n4079), .B(n4078), .ZN(n4082)
         );
  OAI21_X1 U4721 ( .B1(n4246), .B2(n4133), .A(n4082), .ZN(U3272) );
  XNOR2_X1 U4722 ( .A(n4083), .B(n4087), .ZN(n4333) );
  AOI21_X1 U4723 ( .B1(n4090), .B2(n4103), .A(n4084), .ZN(n4331) );
  INV_X1 U4724 ( .A(n4085), .ZN(n4086) );
  AOI22_X1 U4725 ( .A1(n4331), .A2(n4498), .B1(n4086), .B2(n4496), .ZN(n4098)
         );
  XNOR2_X1 U4726 ( .A(n4088), .B(n4087), .ZN(n4089) );
  NAND2_X1 U4727 ( .A1(n4089), .A2(n4172), .ZN(n4093) );
  AOI22_X1 U4728 ( .A1(n4091), .A2(n4166), .B1(n4192), .B2(n4090), .ZN(n4092)
         );
  OAI211_X1 U4729 ( .C1(n4094), .C2(n4169), .A(n4093), .B(n4092), .ZN(n4328)
         );
  INV_X1 U4730 ( .A(n4328), .ZN(n4095) );
  MUX2_X1 U4731 ( .A(n4096), .B(n4095), .S(n4373), .Z(n4097) );
  OAI211_X1 U4732 ( .C1(n4333), .C2(n4133), .A(n4098), .B(n4097), .ZN(U3273)
         );
  OAI21_X1 U4733 ( .B1(n4101), .B2(n4100), .A(n4099), .ZN(n4337) );
  NAND2_X1 U4734 ( .A1(n4118), .A2(n4110), .ZN(n4102) );
  AND2_X1 U4735 ( .A1(n4103), .A2(n4102), .ZN(n4251) );
  OAI22_X1 U4736 ( .A1(n4183), .A2(n4105), .B1(n4104), .B2(n4180), .ZN(n4106)
         );
  AOI21_X1 U4737 ( .B1(n4251), .B2(n4498), .A(n4106), .ZN(n4115) );
  OAI211_X1 U4738 ( .C1(n4109), .C2(n4108), .A(n4107), .B(n4172), .ZN(n4113)
         );
  AOI22_X1 U4739 ( .A1(n4111), .A2(n4166), .B1(n4192), .B2(n4110), .ZN(n4112)
         );
  OAI211_X1 U4740 ( .C1(n4140), .C2(n4169), .A(n4113), .B(n4112), .ZN(n4250)
         );
  NAND2_X1 U4741 ( .A1(n4250), .A2(n4373), .ZN(n4114) );
  OAI211_X1 U4742 ( .C1(n4337), .C2(n4133), .A(n4115), .B(n4114), .ZN(U3274)
         );
  XOR2_X1 U4743 ( .A(n4123), .B(n4116), .Z(n4342) );
  INV_X1 U4744 ( .A(n4117), .ZN(n4150) );
  INV_X1 U4745 ( .A(n4118), .ZN(n4119) );
  AOI21_X1 U4746 ( .B1(n4126), .B2(n4150), .A(n4119), .ZN(n4254) );
  OAI22_X1 U4747 ( .A1(n4183), .A2(n4121), .B1(n4120), .B2(n4180), .ZN(n4122)
         );
  AOI21_X1 U4748 ( .B1(n4254), .B2(n4498), .A(n4122), .ZN(n4132) );
  INV_X1 U4749 ( .A(n4123), .ZN(n4125) );
  OAI211_X1 U4750 ( .C1(n2087), .C2(n4125), .A(n4172), .B(n4124), .ZN(n4129)
         );
  AOI22_X1 U4751 ( .A1(n4127), .A2(n4166), .B1(n4192), .B2(n4126), .ZN(n4128)
         );
  OAI211_X1 U4752 ( .C1(n4130), .C2(n4169), .A(n4129), .B(n4128), .ZN(n4253)
         );
  NAND2_X1 U4753 ( .A1(n4253), .A2(n4373), .ZN(n4131) );
  OAI211_X1 U4754 ( .C1(n4342), .C2(n4133), .A(n4132), .B(n4131), .ZN(U3275)
         );
  XNOR2_X1 U4755 ( .A(n4134), .B(n4136), .ZN(n4146) );
  OAI21_X1 U4756 ( .B1(n4137), .B2(n4136), .A(n4135), .ZN(n4259) );
  NAND2_X1 U4757 ( .A1(n4259), .A2(n4494), .ZN(n4145) );
  OAI22_X1 U4758 ( .A1(n4140), .A2(n4139), .B1(n4200), .B2(n4138), .ZN(n4141)
         );
  AOI21_X1 U4759 ( .B1(n4143), .B2(n4142), .A(n4141), .ZN(n4144) );
  OAI211_X1 U4760 ( .C1(n4147), .C2(n4146), .A(n4145), .B(n4144), .ZN(n4258)
         );
  INV_X1 U4761 ( .A(n4258), .ZN(n4157) );
  NAND2_X1 U4762 ( .A1(n4177), .A2(n4148), .ZN(n4149) );
  NAND2_X1 U4763 ( .A1(n4150), .A2(n4149), .ZN(n4346) );
  NOR2_X1 U4764 ( .A1(n4346), .A2(n4151), .ZN(n4155) );
  OAI22_X1 U4765 ( .A1(n4183), .A2(n4153), .B1(n4152), .B2(n4180), .ZN(n4154)
         );
  AOI211_X1 U4766 ( .C1(n4259), .C2(n4499), .A(n4155), .B(n4154), .ZN(n4156)
         );
  OAI21_X1 U4767 ( .B1(n4157), .B2(n4368), .A(n4156), .ZN(U3276) );
  XOR2_X1 U4768 ( .A(n4164), .B(n4158), .Z(n4261) );
  INV_X1 U4769 ( .A(n4159), .ZN(n4160) );
  AOI21_X1 U4770 ( .B1(n4162), .B2(n4161), .A(n4160), .ZN(n4163) );
  XOR2_X1 U4771 ( .A(n4164), .B(n4163), .Z(n4173) );
  AOI22_X1 U4772 ( .A1(n4167), .A2(n4166), .B1(n4192), .B2(n4165), .ZN(n4168)
         );
  OAI21_X1 U4773 ( .B1(n4170), .B2(n4169), .A(n4168), .ZN(n4171) );
  AOI21_X1 U4774 ( .B1(n4173), .B2(n4172), .A(n4171), .ZN(n4174) );
  OAI21_X1 U4775 ( .B1(n4261), .B2(n4175), .A(n4174), .ZN(n4262) );
  NAND2_X1 U4776 ( .A1(n4262), .A2(n4373), .ZN(n4187) );
  INV_X1 U4777 ( .A(n4176), .ZN(n4179) );
  OAI21_X1 U4778 ( .B1(n4179), .B2(n4178), .A(n4177), .ZN(n4350) );
  INV_X1 U4779 ( .A(n4350), .ZN(n4185) );
  OAI22_X1 U4780 ( .A1(n4183), .A2(n4182), .B1(n4181), .B2(n4180), .ZN(n4184)
         );
  AOI21_X1 U4781 ( .B1(n4185), .B2(n4498), .A(n4184), .ZN(n4186) );
  OAI211_X1 U4782 ( .C1(n4261), .C2(n4188), .A(n4187), .B(n4186), .ZN(U3277)
         );
  XOR2_X1 U4783 ( .A(n4189), .B(n4195), .Z(n4369) );
  INV_X1 U4784 ( .A(n4369), .ZN(n4279) );
  INV_X1 U4785 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4588) );
  AND2_X1 U4786 ( .A1(n4191), .A2(n4190), .ZN(n4198) );
  AOI21_X1 U4787 ( .B1(n4193), .B2(n4192), .A(n4198), .ZN(n4371) );
  MUX2_X1 U4788 ( .A(n4588), .B(n4371), .S(n4568), .Z(n4194) );
  OAI21_X1 U4789 ( .B1(n4279), .B2(n4276), .A(n4194), .ZN(U3549) );
  INV_X1 U4790 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4204) );
  AOI21_X1 U4791 ( .B1(n4197), .B2(n4196), .A(n4195), .ZN(n4374) );
  NAND2_X1 U4792 ( .A1(n4374), .A2(n4248), .ZN(n4203) );
  INV_X1 U4793 ( .A(n4198), .ZN(n4199) );
  OAI21_X1 U4794 ( .B1(n4201), .B2(n4200), .A(n4199), .ZN(n4372) );
  NAND2_X1 U4795 ( .A1(n4372), .A2(n4568), .ZN(n4202) );
  OAI211_X1 U4796 ( .C1(n4568), .C2(n4204), .A(n4203), .B(n4202), .ZN(U3548)
         );
  INV_X1 U4797 ( .A(n4205), .ZN(n4283) );
  MUX2_X1 U4798 ( .A(REG1_REG_28__SCAN_IN), .B(n4283), .S(n4568), .Z(n4206) );
  AOI21_X1 U4799 ( .B1(n4285), .B2(n4248), .A(n4206), .ZN(n4207) );
  OAI21_X1 U4800 ( .B1(n4287), .B2(n4257), .A(n4207), .ZN(U3546) );
  INV_X1 U4801 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4210) );
  AOI21_X1 U4802 ( .B1(n4209), .B2(n4551), .A(n4208), .ZN(n4288) );
  MUX2_X1 U4803 ( .A(n4210), .B(n4288), .S(n4568), .Z(n4211) );
  OAI21_X1 U4804 ( .B1(n4291), .B2(n4257), .A(n4211), .ZN(U3545) );
  INV_X1 U4805 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4214) );
  AOI21_X1 U4806 ( .B1(n4213), .B2(n4549), .A(n4212), .ZN(n4292) );
  OAI21_X1 U4807 ( .B1(n4276), .B2(n4295), .A(n4215), .ZN(U3544) );
  INV_X1 U4808 ( .A(n4216), .ZN(n4296) );
  MUX2_X1 U4809 ( .A(REG1_REG_25__SCAN_IN), .B(n4296), .S(n4568), .Z(n4217) );
  AOI21_X1 U4810 ( .B1(n4298), .B2(n4248), .A(n4217), .ZN(n4218) );
  OAI21_X1 U4811 ( .B1(n4300), .B2(n4257), .A(n4218), .ZN(U3543) );
  INV_X1 U4812 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4221) );
  AOI21_X1 U4813 ( .B1(n4220), .B2(n4549), .A(n4219), .ZN(n4301) );
  MUX2_X1 U4814 ( .A(n4221), .B(n4301), .S(n4568), .Z(n4222) );
  OAI21_X1 U4815 ( .B1(n4276), .B2(n4304), .A(n4222), .ZN(U3542) );
  INV_X1 U4816 ( .A(n4223), .ZN(n4305) );
  MUX2_X1 U4817 ( .A(REG1_REG_23__SCAN_IN), .B(n4305), .S(n4568), .Z(n4224) );
  AOI21_X1 U4818 ( .B1(n4307), .B2(n4248), .A(n4224), .ZN(n4225) );
  OAI21_X1 U4819 ( .B1(n4309), .B2(n4257), .A(n4225), .ZN(U3541) );
  INV_X1 U4820 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4230) );
  AND3_X1 U4821 ( .A1(n4227), .A2(n4551), .A3(n4226), .ZN(n4228) );
  NOR2_X1 U4822 ( .A1(n4229), .A2(n4228), .ZN(n4310) );
  MUX2_X1 U4823 ( .A(n4230), .B(n4310), .S(n4568), .Z(n4231) );
  OAI21_X1 U4824 ( .B1(n4313), .B2(n4257), .A(n4231), .ZN(U3540) );
  OAI21_X1 U4825 ( .B1(n4530), .B2(n4233), .A(n4232), .ZN(n4314) );
  MUX2_X1 U4826 ( .A(REG1_REG_21__SCAN_IN), .B(n4314), .S(n4568), .Z(n4234) );
  INV_X1 U4827 ( .A(n4234), .ZN(n4235) );
  OAI21_X1 U4828 ( .B1(n4317), .B2(n4257), .A(n4235), .ZN(U3539) );
  INV_X1 U4829 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4239) );
  INV_X1 U4830 ( .A(n4236), .ZN(n4238) );
  AOI21_X1 U4831 ( .B1(n4540), .B2(n4238), .A(n4237), .ZN(n4318) );
  MUX2_X1 U4832 ( .A(n4239), .B(n4318), .S(n4568), .Z(n4240) );
  OAI21_X1 U4833 ( .B1(n4276), .B2(n4320), .A(n4240), .ZN(U3538) );
  INV_X1 U4834 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4586) );
  MUX2_X1 U4835 ( .A(n4586), .B(n4321), .S(n4568), .Z(n4242) );
  NAND2_X1 U4836 ( .A1(n4324), .A2(n4248), .ZN(n4241) );
  OAI211_X1 U4837 ( .C1(n4326), .C2(n4257), .A(n4242), .B(n4241), .ZN(U3537)
         );
  OAI211_X1 U4838 ( .C1(n4246), .C2(n4245), .A(n4244), .B(n4243), .ZN(n4327)
         );
  MUX2_X1 U4839 ( .A(REG1_REG_18__SCAN_IN), .B(n4327), .S(n4568), .Z(U3536) );
  MUX2_X1 U4840 ( .A(REG1_REG_17__SCAN_IN), .B(n4328), .S(n4568), .Z(n4247) );
  AOI21_X1 U4841 ( .B1(n4331), .B2(n4248), .A(n4247), .ZN(n4249) );
  OAI21_X1 U4842 ( .B1(n4333), .B2(n4257), .A(n4249), .ZN(U3535) );
  AOI21_X1 U4843 ( .B1(n4551), .B2(n4251), .A(n4250), .ZN(n4334) );
  MUX2_X1 U4844 ( .A(n4468), .B(n4334), .S(n4568), .Z(n4252) );
  OAI21_X1 U4845 ( .B1(n4337), .B2(n4257), .A(n4252), .ZN(U3534) );
  AOI21_X1 U4846 ( .B1(n4551), .B2(n4254), .A(n4253), .ZN(n4338) );
  MUX2_X1 U4847 ( .A(n4255), .B(n4338), .S(n4568), .Z(n4256) );
  OAI21_X1 U4848 ( .B1(n4342), .B2(n4257), .A(n4256), .ZN(U3533) );
  AOI21_X1 U4849 ( .B1(n4540), .B2(n4259), .A(n4258), .ZN(n4343) );
  MUX2_X1 U4850 ( .A(n4442), .B(n4343), .S(n4568), .Z(n4260) );
  OAI21_X1 U4851 ( .B1(n4276), .B2(n4346), .A(n4260), .ZN(U3532) );
  INV_X1 U4852 ( .A(n4261), .ZN(n4263) );
  AOI21_X1 U4853 ( .B1(n4540), .B2(n4263), .A(n4262), .ZN(n4347) );
  MUX2_X1 U4854 ( .A(n4264), .B(n4347), .S(n4568), .Z(n4265) );
  OAI21_X1 U4855 ( .B1(n4276), .B2(n4350), .A(n4265), .ZN(U3531) );
  NAND2_X1 U4856 ( .A1(n4266), .A2(n4549), .ZN(n4267) );
  NAND2_X1 U4857 ( .A1(n4268), .A2(n4267), .ZN(n4351) );
  MUX2_X1 U4858 ( .A(REG1_REG_12__SCAN_IN), .B(n4351), .S(n4568), .Z(n4269) );
  INV_X1 U4859 ( .A(n4269), .ZN(n4270) );
  OAI21_X1 U4860 ( .B1(n4276), .B2(n4354), .A(n4270), .ZN(U3530) );
  INV_X1 U4861 ( .A(n4271), .ZN(n4272) );
  AOI21_X1 U4862 ( .B1(n4540), .B2(n4273), .A(n4272), .ZN(n4355) );
  MUX2_X1 U4863 ( .A(n4274), .B(n4355), .S(n4568), .Z(n4275) );
  OAI21_X1 U4864 ( .B1(n4276), .B2(n4359), .A(n4275), .ZN(U3529) );
  INV_X1 U4865 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4277) );
  MUX2_X1 U4866 ( .A(n4277), .B(n4371), .S(n4756), .Z(n4278) );
  OAI21_X1 U4867 ( .B1(n4279), .B2(n4358), .A(n4278), .ZN(U3517) );
  INV_X1 U4868 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U4869 ( .A1(n4374), .A2(n4330), .ZN(n4281) );
  NAND2_X1 U4870 ( .A1(n4372), .A2(n4756), .ZN(n4280) );
  OAI211_X1 U4871 ( .C1(n4756), .C2(n4282), .A(n4281), .B(n4280), .ZN(U3516)
         );
  MUX2_X1 U4872 ( .A(REG0_REG_28__SCAN_IN), .B(n4283), .S(n4756), .Z(n4284) );
  AOI21_X1 U4873 ( .B1(n4285), .B2(n4330), .A(n4284), .ZN(n4286) );
  OAI21_X1 U4874 ( .B1(n4287), .B2(n4341), .A(n4286), .ZN(U3514) );
  INV_X1 U4875 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4289) );
  MUX2_X1 U4876 ( .A(n4289), .B(n4288), .S(n4756), .Z(n4290) );
  OAI21_X1 U4877 ( .B1(n4291), .B2(n4341), .A(n4290), .ZN(U3513) );
  INV_X1 U4878 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4293) );
  OAI21_X1 U4879 ( .B1(n4295), .B2(n4358), .A(n4294), .ZN(U3512) );
  MUX2_X1 U4880 ( .A(REG0_REG_25__SCAN_IN), .B(n4296), .S(n4756), .Z(n4297) );
  AOI21_X1 U4881 ( .B1(n4298), .B2(n4330), .A(n4297), .ZN(n4299) );
  OAI21_X1 U4882 ( .B1(n4300), .B2(n4341), .A(n4299), .ZN(U3511) );
  INV_X1 U4883 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4302) );
  MUX2_X1 U4884 ( .A(n4302), .B(n4301), .S(n4756), .Z(n4303) );
  OAI21_X1 U4885 ( .B1(n4304), .B2(n4358), .A(n4303), .ZN(U3510) );
  MUX2_X1 U4886 ( .A(REG0_REG_23__SCAN_IN), .B(n4305), .S(n4756), .Z(n4306) );
  AOI21_X1 U4887 ( .B1(n4307), .B2(n4330), .A(n4306), .ZN(n4308) );
  OAI21_X1 U4888 ( .B1(n4309), .B2(n4341), .A(n4308), .ZN(U3509) );
  INV_X1 U4889 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4311) );
  MUX2_X1 U4890 ( .A(n4311), .B(n4310), .S(n4756), .Z(n4312) );
  OAI21_X1 U4891 ( .B1(n4313), .B2(n4341), .A(n4312), .ZN(U3508) );
  MUX2_X1 U4892 ( .A(REG0_REG_21__SCAN_IN), .B(n4314), .S(n4756), .Z(n4315) );
  INV_X1 U4893 ( .A(n4315), .ZN(n4316) );
  OAI21_X1 U4894 ( .B1(n4317), .B2(n4341), .A(n4316), .ZN(U3507) );
  INV_X1 U4895 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4571) );
  MUX2_X1 U4896 ( .A(n4571), .B(n4318), .S(n4756), .Z(n4319) );
  OAI21_X1 U4897 ( .B1(n4320), .B2(n4358), .A(n4319), .ZN(U3506) );
  INV_X1 U4898 ( .A(n4321), .ZN(n4322) );
  MUX2_X1 U4899 ( .A(REG0_REG_19__SCAN_IN), .B(n4322), .S(n4756), .Z(n4323) );
  AOI21_X1 U4900 ( .B1(n4324), .B2(n4330), .A(n4323), .ZN(n4325) );
  OAI21_X1 U4901 ( .B1(n4326), .B2(n4341), .A(n4325), .ZN(U3505) );
  MUX2_X1 U4902 ( .A(REG0_REG_18__SCAN_IN), .B(n4327), .S(n4756), .Z(U3503) );
  MUX2_X1 U4903 ( .A(REG0_REG_17__SCAN_IN), .B(n4328), .S(n4756), .Z(n4329) );
  AOI21_X1 U4904 ( .B1(n4331), .B2(n4330), .A(n4329), .ZN(n4332) );
  OAI21_X1 U4905 ( .B1(n4333), .B2(n4341), .A(n4332), .ZN(U3501) );
  INV_X1 U4906 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4335) );
  MUX2_X1 U4907 ( .A(n4335), .B(n4334), .S(n4756), .Z(n4336) );
  OAI21_X1 U4908 ( .B1(n4337), .B2(n4341), .A(n4336), .ZN(U3499) );
  INV_X1 U4909 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4339) );
  MUX2_X1 U4910 ( .A(n4339), .B(n4338), .S(n4756), .Z(n4340) );
  OAI21_X1 U4911 ( .B1(n4342), .B2(n4341), .A(n4340), .ZN(U3497) );
  INV_X1 U4912 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4344) );
  MUX2_X1 U4913 ( .A(n4344), .B(n4343), .S(n4756), .Z(n4345) );
  OAI21_X1 U4914 ( .B1(n4346), .B2(n4358), .A(n4345), .ZN(U3495) );
  INV_X1 U4915 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4348) );
  MUX2_X1 U4916 ( .A(n4348), .B(n4347), .S(n4756), .Z(n4349) );
  OAI21_X1 U4917 ( .B1(n4350), .B2(n4358), .A(n4349), .ZN(U3493) );
  MUX2_X1 U4918 ( .A(REG0_REG_12__SCAN_IN), .B(n4351), .S(n4756), .Z(n4352) );
  INV_X1 U4919 ( .A(n4352), .ZN(n4353) );
  OAI21_X1 U4920 ( .B1(n4354), .B2(n4358), .A(n4353), .ZN(U3491) );
  INV_X1 U4921 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4356) );
  MUX2_X1 U4922 ( .A(n4356), .B(n4355), .S(n4756), .Z(n4357) );
  OAI21_X1 U4923 ( .B1(n4359), .B2(n4358), .A(n4357), .ZN(U3489) );
  MUX2_X1 U4924 ( .A(DATAI_29_), .B(n2332), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4925 ( .A(n4360), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4926 ( .A(DATAI_24_), .B(n2198), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4927 ( .A(DATAI_20_), .B(n4361), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4928 ( .A(n4362), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4929 ( .A(n4363), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4930 ( .A(DATAI_4_), .B(n4390), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4931 ( .A(n4364), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4932 ( .A(n4365), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U4933 ( .A(DATAI_28_), .ZN(n4366) );
  AOI22_X1 U4934 ( .A1(STATE_REG_SCAN_IN), .A2(n4367), .B1(n4366), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4935 ( .A1(n4369), .A2(n4498), .B1(n4368), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4370) );
  OAI21_X1 U4936 ( .B1(n4368), .B2(n4371), .A(n4370), .ZN(U3260) );
  AOI22_X1 U4937 ( .A1(n4374), .A2(n4498), .B1(n4373), .B2(n4372), .ZN(n4375)
         );
  OAI21_X1 U4938 ( .B1(n3427), .B2(n4373), .A(n4375), .ZN(U3261) );
  OAI21_X1 U4939 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4377), .A(n4376), .ZN(n4378)
         );
  XOR2_X1 U4940 ( .A(n4378), .B(IR_REG_0__SCAN_IN), .Z(n4381) );
  AOI22_X1 U4941 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4457), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4379) );
  OAI21_X1 U4942 ( .B1(n4381), .B2(n4380), .A(n4379), .ZN(U3240) );
  XOR2_X1 U4943 ( .A(n4382), .B(REG1_REG_4__SCAN_IN), .Z(n4385) );
  XOR2_X1 U4944 ( .A(n4383), .B(REG2_REG_4__SCAN_IN), .Z(n4384) );
  OAI22_X1 U4945 ( .A1(n4385), .A2(n4475), .B1(n4443), .B2(n4384), .ZN(n4389)
         );
  AOI21_X1 U4946 ( .B1(n4457), .B2(ADDR_REG_4__SCAN_IN), .A(n4386), .ZN(n4387)
         );
  INV_X1 U4947 ( .A(n4387), .ZN(n4388) );
  AOI211_X1 U4948 ( .C1(n4390), .C2(n4449), .A(n4389), .B(n4388), .ZN(n4392)
         );
  NAND2_X1 U4949 ( .A1(n4392), .A2(n4391), .ZN(U3244) );
  AOI211_X1 U4950 ( .C1(n4395), .C2(n4394), .A(n4393), .B(n4475), .ZN(n4397)
         );
  AOI211_X1 U4951 ( .C1(n4457), .C2(ADDR_REG_9__SCAN_IN), .A(n4397), .B(n4396), 
        .ZN(n4402) );
  OAI211_X1 U4952 ( .C1(n4400), .C2(n4399), .A(n4487), .B(n4398), .ZN(n4401)
         );
  OAI211_X1 U4953 ( .C1(n4490), .C2(n4522), .A(n4402), .B(n4401), .ZN(U3249)
         );
  AOI211_X1 U4954 ( .C1(n4405), .C2(n4404), .A(n4403), .B(n4475), .ZN(n4407)
         );
  AOI211_X1 U4955 ( .C1(n4457), .C2(ADDR_REG_10__SCAN_IN), .A(n4407), .B(n4406), .ZN(n4411) );
  OAI211_X1 U4956 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4409), .A(n4487), .B(n4408), .ZN(n4410) );
  OAI211_X1 U4957 ( .C1(n4490), .C2(n4520), .A(n4411), .B(n4410), .ZN(U3250)
         );
  AOI211_X1 U4958 ( .C1(n2090), .C2(n4413), .A(n4412), .B(n4475), .ZN(n4415)
         );
  AOI211_X1 U4959 ( .C1(n4457), .C2(ADDR_REG_11__SCAN_IN), .A(n4415), .B(n4414), .ZN(n4420) );
  OAI211_X1 U4960 ( .C1(n4418), .C2(n4417), .A(n4487), .B(n4416), .ZN(n4419)
         );
  OAI211_X1 U4961 ( .C1(n4490), .C2(n4518), .A(n4420), .B(n4419), .ZN(U3251)
         );
  AOI211_X1 U4962 ( .C1(n4423), .C2(n4422), .A(n4421), .B(n4475), .ZN(n4424)
         );
  AOI211_X1 U4963 ( .C1(n4457), .C2(ADDR_REG_12__SCAN_IN), .A(n4425), .B(n4424), .ZN(n4429) );
  OAI211_X1 U4964 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4427), .A(n4487), .B(n4426), .ZN(n4428) );
  OAI211_X1 U4965 ( .C1(n4490), .C2(n4516), .A(n4429), .B(n4428), .ZN(U3252)
         );
  AOI211_X1 U4966 ( .C1(n2082), .C2(n4431), .A(n4430), .B(n4475), .ZN(n4432)
         );
  AOI211_X1 U4967 ( .C1(n4457), .C2(ADDR_REG_13__SCAN_IN), .A(n4433), .B(n4432), .ZN(n4439) );
  AOI21_X1 U4968 ( .B1(n4182), .B2(n4514), .A(n4434), .ZN(n4437) );
  AOI21_X1 U4969 ( .B1(n4437), .B2(n4436), .A(n4443), .ZN(n4435) );
  OAI21_X1 U4970 ( .B1(n4437), .B2(n4436), .A(n4435), .ZN(n4438) );
  OAI211_X1 U4971 ( .C1(n4490), .C2(n4514), .A(n4439), .B(n4438), .ZN(U3253)
         );
  NAND2_X1 U4972 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4457), .ZN(n4452) );
  AOI211_X1 U4973 ( .C1(n4442), .C2(n4441), .A(n4440), .B(n4475), .ZN(n4447)
         );
  AOI211_X1 U4974 ( .C1(n4153), .C2(n4445), .A(n4444), .B(n4443), .ZN(n4446)
         );
  AOI211_X1 U4975 ( .C1(n4449), .C2(n4448), .A(n4447), .B(n4446), .ZN(n4451)
         );
  NAND3_X1 U4976 ( .A1(n4452), .A2(n4451), .A3(n4450), .ZN(U3254) );
  AOI211_X1 U4977 ( .C1(n2078), .C2(n4454), .A(n4453), .B(n4475), .ZN(n4455)
         );
  AOI211_X1 U4978 ( .C1(n4457), .C2(ADDR_REG_15__SCAN_IN), .A(n4456), .B(n4455), .ZN(n4463) );
  AOI21_X1 U4979 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(n4461) );
  NAND2_X1 U4980 ( .A1(n4487), .A2(n4461), .ZN(n4462) );
  OAI211_X1 U4981 ( .C1(n4490), .C2(n4511), .A(n4463), .B(n4462), .ZN(U3255)
         );
  AOI21_X1 U4982 ( .B1(n4457), .B2(ADDR_REG_16__SCAN_IN), .A(n4464), .ZN(n4474) );
  OAI21_X1 U4983 ( .B1(n4466), .B2(n4105), .A(n4465), .ZN(n4472) );
  OAI21_X1 U4984 ( .B1(n4469), .B2(n4468), .A(n4467), .ZN(n4470) );
  AOI22_X1 U4985 ( .A1(n4487), .A2(n4472), .B1(n4471), .B2(n4470), .ZN(n4473)
         );
  OAI211_X1 U4986 ( .C1(n4510), .C2(n4490), .A(n4474), .B(n4473), .ZN(U3256)
         );
  NAND2_X1 U4987 ( .A1(n4457), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4480) );
  INV_X1 U4988 ( .A(n4478), .ZN(n4479) );
  NAND2_X1 U4989 ( .A1(n4480), .A2(n4479), .ZN(n4481) );
  AOI21_X1 U4990 ( .B1(n4485), .B2(n4484), .A(n4483), .ZN(n4486) );
  NAND2_X1 U4991 ( .A1(n4487), .A2(n4486), .ZN(n4488) );
  OAI211_X1 U4992 ( .C1(n4490), .C2(n4508), .A(n4489), .B(n4488), .ZN(U3258)
         );
  INV_X1 U4993 ( .A(n4491), .ZN(n4500) );
  INV_X1 U4994 ( .A(n4492), .ZN(n4493) );
  AOI21_X1 U4995 ( .B1(n4494), .B2(n4500), .A(n4493), .ZN(n4503) );
  AOI22_X1 U4996 ( .A1(n2140), .A2(n4496), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4368), .ZN(n4502) );
  AOI22_X1 U4997 ( .A1(n4500), .A2(n4499), .B1(n4498), .B2(n4497), .ZN(n4501)
         );
  OAI211_X1 U4998 ( .C1(n4368), .C2(n4503), .A(n4502), .B(n4501), .ZN(U3280)
         );
  AND2_X1 U4999 ( .A1(D_REG_31__SCAN_IN), .A2(n4505), .ZN(U3291) );
  AND2_X1 U5000 ( .A1(n4505), .A2(D_REG_30__SCAN_IN), .ZN(U3292) );
  AND2_X1 U5001 ( .A1(n4505), .A2(D_REG_29__SCAN_IN), .ZN(U3293) );
  AND2_X1 U5002 ( .A1(D_REG_28__SCAN_IN), .A2(n4505), .ZN(U3294) );
  INV_X1 U5003 ( .A(n4505), .ZN(n4504) );
  INV_X1 U5004 ( .A(D_REG_27__SCAN_IN), .ZN(n4700) );
  NOR2_X1 U5005 ( .A1(n4504), .A2(n4700), .ZN(U3295) );
  AND2_X1 U5006 ( .A1(D_REG_26__SCAN_IN), .A2(n4505), .ZN(U3296) );
  AND2_X1 U5007 ( .A1(D_REG_25__SCAN_IN), .A2(n4505), .ZN(U3297) );
  AND2_X1 U5008 ( .A1(D_REG_24__SCAN_IN), .A2(n4505), .ZN(U3298) );
  AND2_X1 U5009 ( .A1(n4505), .A2(D_REG_23__SCAN_IN), .ZN(U3299) );
  AND2_X1 U5010 ( .A1(D_REG_22__SCAN_IN), .A2(n4505), .ZN(U3300) );
  AND2_X1 U5011 ( .A1(D_REG_21__SCAN_IN), .A2(n4505), .ZN(U3301) );
  AND2_X1 U5012 ( .A1(D_REG_20__SCAN_IN), .A2(n4505), .ZN(U3302) );
  AND2_X1 U5013 ( .A1(D_REG_19__SCAN_IN), .A2(n4505), .ZN(U3303) );
  INV_X1 U5014 ( .A(D_REG_18__SCAN_IN), .ZN(n4721) );
  NOR2_X1 U5015 ( .A1(n4504), .A2(n4721), .ZN(U3304) );
  AND2_X1 U5016 ( .A1(D_REG_17__SCAN_IN), .A2(n4505), .ZN(U3305) );
  AND2_X1 U5017 ( .A1(D_REG_16__SCAN_IN), .A2(n4505), .ZN(U3306) );
  AND2_X1 U5018 ( .A1(D_REG_15__SCAN_IN), .A2(n4505), .ZN(U3307) );
  AND2_X1 U5019 ( .A1(D_REG_14__SCAN_IN), .A2(n4505), .ZN(U3308) );
  AND2_X1 U5020 ( .A1(D_REG_13__SCAN_IN), .A2(n4505), .ZN(U3309) );
  AND2_X1 U5021 ( .A1(D_REG_12__SCAN_IN), .A2(n4505), .ZN(U3310) );
  AND2_X1 U5022 ( .A1(D_REG_11__SCAN_IN), .A2(n4505), .ZN(U3311) );
  AND2_X1 U5023 ( .A1(n4505), .A2(D_REG_10__SCAN_IN), .ZN(U3312) );
  INV_X1 U5024 ( .A(D_REG_9__SCAN_IN), .ZN(n4574) );
  NOR2_X1 U5025 ( .A1(n4504), .A2(n4574), .ZN(U3313) );
  AND2_X1 U5026 ( .A1(D_REG_8__SCAN_IN), .A2(n4505), .ZN(U3314) );
  AND2_X1 U5027 ( .A1(D_REG_7__SCAN_IN), .A2(n4505), .ZN(U3315) );
  AND2_X1 U5028 ( .A1(n4505), .A2(D_REG_6__SCAN_IN), .ZN(U3316) );
  AND2_X1 U5029 ( .A1(D_REG_5__SCAN_IN), .A2(n4505), .ZN(U3317) );
  AND2_X1 U5030 ( .A1(D_REG_4__SCAN_IN), .A2(n4505), .ZN(U3318) );
  AND2_X1 U5031 ( .A1(D_REG_3__SCAN_IN), .A2(n4505), .ZN(U3319) );
  AND2_X1 U5032 ( .A1(D_REG_2__SCAN_IN), .A2(n4505), .ZN(U3320) );
  INV_X1 U5033 ( .A(DATAI_23_), .ZN(n4507) );
  AOI21_X1 U5034 ( .B1(U3149), .B2(n4507), .A(n4506), .ZN(U3329) );
  INV_X1 U5035 ( .A(DATAI_18_), .ZN(n4701) );
  AOI22_X1 U5036 ( .A1(STATE_REG_SCAN_IN), .A2(n4508), .B1(n4701), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5037 ( .A(DATAI_16_), .ZN(n4509) );
  AOI22_X1 U5038 ( .A1(STATE_REG_SCAN_IN), .A2(n4510), .B1(n4509), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5039 ( .A(DATAI_15_), .ZN(n4594) );
  AOI22_X1 U5040 ( .A1(STATE_REG_SCAN_IN), .A2(n4511), .B1(n4594), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5041 ( .A(DATAI_14_), .ZN(n4512) );
  AOI22_X1 U5042 ( .A1(STATE_REG_SCAN_IN), .A2(n4513), .B1(n4512), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5043 ( .A1(STATE_REG_SCAN_IN), .A2(n4514), .B1(n2628), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5044 ( .A1(STATE_REG_SCAN_IN), .A2(n4516), .B1(n4515), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5045 ( .A(DATAI_11_), .ZN(n4517) );
  AOI22_X1 U5046 ( .A1(STATE_REG_SCAN_IN), .A2(n4518), .B1(n4517), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5047 ( .A(DATAI_10_), .ZN(n4519) );
  AOI22_X1 U5048 ( .A1(STATE_REG_SCAN_IN), .A2(n4520), .B1(n4519), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5049 ( .A(DATAI_9_), .ZN(n4521) );
  AOI22_X1 U5050 ( .A1(STATE_REG_SCAN_IN), .A2(n4522), .B1(n4521), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5051 ( .A1(STATE_REG_SCAN_IN), .A2(n2316), .B1(n2201), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5052 ( .C1(n4540), .C2(n4525), .A(n4524), .B(n4523), .ZN(n4559)
         );
  INV_X1 U5053 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5054 ( .A1(n4756), .A2(n4559), .B1(n4526), .B2(n4556), .ZN(U3467)
         );
  INV_X1 U5055 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5056 ( .A1(n4756), .A2(n4528), .B1(n4527), .B2(n4556), .ZN(U3469)
         );
  OAI22_X1 U5057 ( .A1(n4532), .A2(n4531), .B1(n4530), .B2(n4529), .ZN(n4533)
         );
  NOR2_X1 U5058 ( .A1(n4534), .A2(n4533), .ZN(n4561) );
  INV_X1 U5059 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5060 ( .A1(n4756), .A2(n4561), .B1(n4535), .B2(n4556), .ZN(U3473)
         );
  INV_X1 U5061 ( .A(n4536), .ZN(n4541) );
  INV_X1 U5062 ( .A(n4537), .ZN(n4539) );
  AOI211_X1 U5063 ( .C1(n4541), .C2(n4540), .A(n4539), .B(n4538), .ZN(n4562)
         );
  INV_X1 U5064 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5065 ( .A1(n4756), .A2(n4562), .B1(n4542), .B2(n4556), .ZN(U3475)
         );
  NAND3_X1 U5066 ( .A1(n4544), .A2(n4543), .A3(n4549), .ZN(n4545) );
  AND3_X1 U5067 ( .A1(n4547), .A2(n4546), .A3(n4545), .ZN(n4564) );
  INV_X1 U5068 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4548) );
  AOI22_X1 U5069 ( .A1(n4756), .A2(n4564), .B1(n4548), .B2(n4556), .ZN(U3481)
         );
  NAND2_X1 U5070 ( .A1(n4550), .A2(n4549), .ZN(n4554) );
  NAND2_X1 U5071 ( .A1(n4552), .A2(n4551), .ZN(n4553) );
  INV_X1 U5072 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U5073 ( .A1(n4756), .A2(n4567), .B1(n4557), .B2(n4556), .ZN(U3485)
         );
  AOI22_X1 U5074 ( .A1(n4568), .A2(n4559), .B1(n4558), .B2(n4565), .ZN(U3518)
         );
  INV_X1 U5075 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5076 ( .A1(n4568), .A2(n4561), .B1(n4560), .B2(n4565), .ZN(U3521)
         );
  AOI22_X1 U5077 ( .A1(n4568), .A2(n4562), .B1(n2916), .B2(n4565), .ZN(U3522)
         );
  AOI22_X1 U5078 ( .A1(n4568), .A2(n4564), .B1(n4563), .B2(n4565), .ZN(U3525)
         );
  AOI22_X1 U5079 ( .A1(n4568), .A2(n4567), .B1(n4566), .B2(n4565), .ZN(U3527)
         );
  AOI22_X1 U5080 ( .A1(n4571), .A2(keyinput99), .B1(keyinput112), .B2(n4570), 
        .ZN(n4569) );
  OAI221_X1 U5081 ( .B1(n4571), .B2(keyinput99), .C1(n4570), .C2(keyinput112), 
        .A(n4569), .ZN(n4582) );
  INV_X1 U5082 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5083 ( .A1(n4182), .A2(keyinput122), .B1(keyinput121), .B2(n4697), 
        .ZN(n4572) );
  OAI221_X1 U5084 ( .B1(n4182), .B2(keyinput122), .C1(n4697), .C2(keyinput121), 
        .A(n4572), .ZN(n4581) );
  AOI22_X1 U5085 ( .A1(n4575), .A2(keyinput91), .B1(n4574), .B2(keyinput116), 
        .ZN(n4573) );
  OAI221_X1 U5086 ( .B1(n4575), .B2(keyinput91), .C1(n4574), .C2(keyinput116), 
        .A(n4573), .ZN(n4580) );
  AOI22_X1 U5087 ( .A1(n4578), .A2(keyinput114), .B1(keyinput88), .B2(n4577), 
        .ZN(n4576) );
  OAI221_X1 U5088 ( .B1(n4578), .B2(keyinput114), .C1(n4577), .C2(keyinput88), 
        .A(n4576), .ZN(n4579) );
  NOR4_X1 U5089 ( .A1(n4582), .A2(n4581), .A3(n4580), .A4(n4579), .ZN(n4620)
         );
  AOI22_X1 U5090 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput95), .B1(
        IR_REG_26__SCAN_IN), .B2(keyinput87), .ZN(n4583) );
  OAI221_X1 U5091 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput95), .C1(
        IR_REG_26__SCAN_IN), .C2(keyinput87), .A(n4583), .ZN(n4592) );
  AOI22_X1 U5092 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput69), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput74), .ZN(n4584) );
  OAI221_X1 U5093 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput69), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput74), .A(n4584), .ZN(n4591) );
  AOI22_X1 U5094 ( .A1(n4586), .A2(keyinput110), .B1(keyinput100), .B2(n4069), 
        .ZN(n4585) );
  OAI221_X1 U5095 ( .B1(n4586), .B2(keyinput110), .C1(n4069), .C2(keyinput100), 
        .A(n4585), .ZN(n4590) );
  AOI22_X1 U5096 ( .A1(n4724), .A2(keyinput106), .B1(keyinput77), .B2(n4588), 
        .ZN(n4587) );
  OAI221_X1 U5097 ( .B1(n4724), .B2(keyinput106), .C1(n4588), .C2(keyinput77), 
        .A(n4587), .ZN(n4589) );
  NOR4_X1 U5098 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), .ZN(n4619)
         );
  AOI22_X1 U5099 ( .A1(n4594), .A2(keyinput71), .B1(n4721), .B2(keyinput82), 
        .ZN(n4593) );
  OAI221_X1 U5100 ( .B1(n4594), .B2(keyinput71), .C1(n4721), .C2(keyinput82), 
        .A(n4593), .ZN(n4605) );
  XNOR2_X1 U5101 ( .A(n4595), .B(keyinput97), .ZN(n4598) );
  XNOR2_X1 U5102 ( .A(n4596), .B(keyinput98), .ZN(n4597) );
  NOR2_X1 U5103 ( .A1(n4598), .A2(n4597), .ZN(n4602) );
  XNOR2_X1 U5104 ( .A(keyinput68), .B(DATAI_18_), .ZN(n4601) );
  XNOR2_X1 U5105 ( .A(IR_REG_22__SCAN_IN), .B(keyinput65), .ZN(n4600) );
  XNOR2_X1 U5106 ( .A(IR_REG_5__SCAN_IN), .B(keyinput67), .ZN(n4599) );
  NAND4_X1 U5107 ( .A1(n4602), .A2(n4601), .A3(n4600), .A4(n4599), .ZN(n4604)
         );
  XNOR2_X1 U5108 ( .A(n4700), .B(keyinput109), .ZN(n4603) );
  NOR3_X1 U5109 ( .A1(n4605), .A2(n4604), .A3(n4603), .ZN(n4618) );
  INV_X1 U5110 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4607) );
  AOI22_X1 U5111 ( .A1(n4607), .A2(keyinput103), .B1(n2548), .B2(keyinput90), 
        .ZN(n4606) );
  OAI221_X1 U5112 ( .B1(n4607), .B2(keyinput103), .C1(n2548), .C2(keyinput90), 
        .A(n4606), .ZN(n4616) );
  AOI22_X1 U5113 ( .A1(n2327), .A2(keyinput84), .B1(keyinput102), .B2(n4723), 
        .ZN(n4608) );
  OAI221_X1 U5114 ( .B1(n2327), .B2(keyinput84), .C1(n4723), .C2(keyinput102), 
        .A(n4608), .ZN(n4615) );
  AOI22_X1 U5115 ( .A1(n4728), .A2(keyinput83), .B1(n4610), .B2(keyinput70), 
        .ZN(n4609) );
  OAI221_X1 U5116 ( .B1(n4728), .B2(keyinput83), .C1(n4610), .C2(keyinput70), 
        .A(n4609), .ZN(n4614) );
  XOR2_X1 U5117 ( .A(n2317), .B(keyinput81), .Z(n4612) );
  XNOR2_X1 U5118 ( .A(IR_REG_9__SCAN_IN), .B(keyinput72), .ZN(n4611) );
  NAND2_X1 U5119 ( .A1(n4612), .A2(n4611), .ZN(n4613) );
  NOR4_X1 U5120 ( .A1(n4616), .A2(n4615), .A3(n4614), .A4(n4613), .ZN(n4617)
         );
  AND4_X1 U5121 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4753)
         );
  OAI22_X1 U5122 ( .A1(REG3_REG_18__SCAN_IN), .A2(keyinput85), .B1(
        ADDR_REG_7__SCAN_IN), .B2(keyinput75), .ZN(n4621) );
  AOI221_X1 U5123 ( .B1(REG3_REG_18__SCAN_IN), .B2(keyinput85), .C1(keyinput75), .C2(ADDR_REG_7__SCAN_IN), .A(n4621), .ZN(n4628) );
  OAI22_X1 U5124 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput124), .B1(keyinput126), 
        .B2(DATAO_REG_23__SCAN_IN), .ZN(n4622) );
  AOI221_X1 U5125 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput124), .C1(
        DATAO_REG_23__SCAN_IN), .C2(keyinput126), .A(n4622), .ZN(n4627) );
  OAI22_X1 U5126 ( .A1(REG2_REG_21__SCAN_IN), .A2(keyinput96), .B1(
        DATAO_REG_5__SCAN_IN), .B2(keyinput73), .ZN(n4623) );
  AOI221_X1 U5127 ( .B1(REG2_REG_21__SCAN_IN), .B2(keyinput96), .C1(keyinput73), .C2(DATAO_REG_5__SCAN_IN), .A(n4623), .ZN(n4626) );
  OAI22_X1 U5128 ( .A1(REG2_REG_30__SCAN_IN), .A2(keyinput86), .B1(keyinput64), 
        .B2(ADDR_REG_12__SCAN_IN), .ZN(n4624) );
  AOI221_X1 U5129 ( .B1(REG2_REG_30__SCAN_IN), .B2(keyinput86), .C1(
        ADDR_REG_12__SCAN_IN), .C2(keyinput64), .A(n4624), .ZN(n4625) );
  NAND4_X1 U5130 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4656)
         );
  OAI22_X1 U5131 ( .A1(REG0_REG_10__SCAN_IN), .A2(keyinput123), .B1(
        keyinput105), .B2(REG2_REG_0__SCAN_IN), .ZN(n4629) );
  AOI221_X1 U5132 ( .B1(REG0_REG_10__SCAN_IN), .B2(keyinput123), .C1(
        REG2_REG_0__SCAN_IN), .C2(keyinput105), .A(n4629), .ZN(n4636) );
  OAI22_X1 U5133 ( .A1(REG1_REG_26__SCAN_IN), .A2(keyinput115), .B1(
        REG2_REG_2__SCAN_IN), .B2(keyinput92), .ZN(n4630) );
  AOI221_X1 U5134 ( .B1(REG1_REG_26__SCAN_IN), .B2(keyinput115), .C1(
        keyinput92), .C2(REG2_REG_2__SCAN_IN), .A(n4630), .ZN(n4635) );
  OAI22_X1 U5135 ( .A1(REG1_REG_1__SCAN_IN), .A2(keyinput94), .B1(
        DATAO_REG_27__SCAN_IN), .B2(keyinput78), .ZN(n4631) );
  AOI221_X1 U5136 ( .B1(REG1_REG_1__SCAN_IN), .B2(keyinput94), .C1(keyinput78), 
        .C2(DATAO_REG_27__SCAN_IN), .A(n4631), .ZN(n4634) );
  OAI22_X1 U5137 ( .A1(REG0_REG_5__SCAN_IN), .A2(keyinput113), .B1(
        REG1_REG_4__SCAN_IN), .B2(keyinput127), .ZN(n4632) );
  AOI221_X1 U5138 ( .B1(REG0_REG_5__SCAN_IN), .B2(keyinput113), .C1(
        keyinput127), .C2(REG1_REG_4__SCAN_IN), .A(n4632), .ZN(n4633) );
  NAND4_X1 U5139 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4655)
         );
  OAI22_X1 U5140 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput119), .B1(keyinput108), 
        .B2(D_REG_6__SCAN_IN), .ZN(n4637) );
  AOI221_X1 U5141 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput119), .C1(
        D_REG_6__SCAN_IN), .C2(keyinput108), .A(n4637), .ZN(n4644) );
  OAI22_X1 U5142 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput89), .B1(keyinput79), 
        .B2(DATAI_14_), .ZN(n4638) );
  AOI221_X1 U5143 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput89), .C1(DATAI_14_), 
        .C2(keyinput79), .A(n4638), .ZN(n4643) );
  OAI22_X1 U5144 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput111), .B1(keyinput118), 
        .B2(D_REG_23__SCAN_IN), .ZN(n4639) );
  AOI221_X1 U5145 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput111), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput118), .A(n4639), .ZN(n4642) );
  OAI22_X1 U5146 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput107), .B1(keyinput125), 
        .B2(D_REG_30__SCAN_IN), .ZN(n4640) );
  AOI221_X1 U5147 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput107), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput125), .A(n4640), .ZN(n4641) );
  NAND4_X1 U5148 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4654)
         );
  OAI22_X1 U5149 ( .A1(DATAI_20_), .A2(keyinput120), .B1(keyinput93), .B2(
        DATAI_6_), .ZN(n4645) );
  AOI221_X1 U5150 ( .B1(DATAI_20_), .B2(keyinput120), .C1(DATAI_6_), .C2(
        keyinput93), .A(n4645), .ZN(n4652) );
  OAI22_X1 U5151 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput101), .B1(
        keyinput117), .B2(DATAO_REG_2__SCAN_IN), .ZN(n4646) );
  AOI221_X1 U5152 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput101), .C1(
        DATAO_REG_2__SCAN_IN), .C2(keyinput117), .A(n4646), .ZN(n4651) );
  OAI22_X1 U5153 ( .A1(DATAI_8_), .A2(keyinput66), .B1(keyinput104), .B2(
        DATAI_7_), .ZN(n4647) );
  AOI221_X1 U5154 ( .B1(DATAI_8_), .B2(keyinput66), .C1(DATAI_7_), .C2(
        keyinput104), .A(n4647), .ZN(n4650) );
  OAI22_X1 U5155 ( .A1(DATAI_28_), .A2(keyinput76), .B1(keyinput80), .B2(
        DATAI_24_), .ZN(n4648) );
  AOI221_X1 U5156 ( .B1(DATAI_28_), .B2(keyinput76), .C1(DATAI_24_), .C2(
        keyinput80), .A(n4648), .ZN(n4649) );
  NAND4_X1 U5157 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4653)
         );
  NOR4_X1 U5158 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4752)
         );
  AOI22_X1 U5159 ( .A1(DATAI_14_), .A2(keyinput15), .B1(IR_REG_26__SCAN_IN), 
        .B2(keyinput23), .ZN(n4657) );
  OAI221_X1 U5160 ( .B1(DATAI_14_), .B2(keyinput15), .C1(IR_REG_26__SCAN_IN), 
        .C2(keyinput23), .A(n4657), .ZN(n4664) );
  AOI22_X1 U5161 ( .A1(ADDR_REG_7__SCAN_IN), .A2(keyinput11), .B1(DATAI_15_), 
        .B2(keyinput7), .ZN(n4658) );
  OAI221_X1 U5162 ( .B1(ADDR_REG_7__SCAN_IN), .B2(keyinput11), .C1(DATAI_15_), 
        .C2(keyinput7), .A(n4658), .ZN(n4663) );
  AOI22_X1 U5163 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput27), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput3), .ZN(n4659) );
  OAI221_X1 U5164 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput27), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput3), .A(n4659), .ZN(n4662) );
  AOI22_X1 U5165 ( .A1(REG1_REG_6__SCAN_IN), .A2(keyinput48), .B1(
        REG2_REG_21__SCAN_IN), .B2(keyinput32), .ZN(n4660) );
  OAI221_X1 U5166 ( .B1(REG1_REG_6__SCAN_IN), .B2(keyinput48), .C1(
        REG2_REG_21__SCAN_IN), .C2(keyinput32), .A(n4660), .ZN(n4661) );
  NOR4_X1 U5167 ( .A1(n4664), .A2(n4663), .A3(n4662), .A4(n4661), .ZN(n4692)
         );
  AOI22_X1 U5168 ( .A1(DATAI_7_), .A2(keyinput40), .B1(D_REG_29__SCAN_IN), 
        .B2(keyinput43), .ZN(n4665) );
  OAI221_X1 U5169 ( .B1(DATAI_7_), .B2(keyinput40), .C1(D_REG_29__SCAN_IN), 
        .C2(keyinput43), .A(n4665), .ZN(n4672) );
  AOI22_X1 U5170 ( .A1(REG0_REG_20__SCAN_IN), .A2(keyinput35), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput60), .ZN(n4666) );
  OAI221_X1 U5171 ( .B1(REG0_REG_20__SCAN_IN), .B2(keyinput35), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput60), .A(n4666), .ZN(n4671) );
  AOI22_X1 U5172 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput39), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput52), .ZN(n4667) );
  OAI221_X1 U5173 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput39), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput52), .A(n4667), .ZN(n4670) );
  AOI22_X1 U5174 ( .A1(REG0_REG_29__SCAN_IN), .A2(keyinput50), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput54), .ZN(n4668) );
  OAI221_X1 U5175 ( .B1(REG0_REG_29__SCAN_IN), .B2(keyinput50), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput54), .A(n4668), .ZN(n4669) );
  NOR4_X1 U5176 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(n4691)
         );
  AOI22_X1 U5177 ( .A1(REG1_REG_19__SCAN_IN), .A2(keyinput46), .B1(
        IR_REG_28__SCAN_IN), .B2(keyinput34), .ZN(n4673) );
  OAI221_X1 U5178 ( .B1(REG1_REG_19__SCAN_IN), .B2(keyinput46), .C1(
        IR_REG_28__SCAN_IN), .C2(keyinput34), .A(n4673), .ZN(n4680) );
  AOI22_X1 U5179 ( .A1(DATAO_REG_27__SCAN_IN), .A2(keyinput14), .B1(
        REG1_REG_1__SCAN_IN), .B2(keyinput30), .ZN(n4674) );
  OAI221_X1 U5180 ( .B1(DATAO_REG_27__SCAN_IN), .B2(keyinput14), .C1(
        REG1_REG_1__SCAN_IN), .C2(keyinput30), .A(n4674), .ZN(n4679) );
  AOI22_X1 U5181 ( .A1(DATAI_8_), .A2(keyinput2), .B1(REG3_REG_17__SCAN_IN), 
        .B2(keyinput6), .ZN(n4675) );
  OAI221_X1 U5182 ( .B1(DATAI_8_), .B2(keyinput2), .C1(REG3_REG_17__SCAN_IN), 
        .C2(keyinput6), .A(n4675), .ZN(n4678) );
  AOI22_X1 U5183 ( .A1(DATAI_24_), .A2(keyinput16), .B1(REG3_REG_28__SCAN_IN), 
        .B2(keyinput37), .ZN(n4676) );
  OAI221_X1 U5184 ( .B1(DATAI_24_), .B2(keyinput16), .C1(REG3_REG_28__SCAN_IN), 
        .C2(keyinput37), .A(n4676), .ZN(n4677) );
  NOR4_X1 U5185 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4690)
         );
  AOI22_X1 U5186 ( .A1(DATAI_28_), .A2(keyinput12), .B1(REG3_REG_18__SCAN_IN), 
        .B2(keyinput21), .ZN(n4681) );
  OAI221_X1 U5187 ( .B1(DATAI_28_), .B2(keyinput12), .C1(REG3_REG_18__SCAN_IN), 
        .C2(keyinput21), .A(n4681), .ZN(n4688) );
  AOI22_X1 U5188 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput25), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput61), .ZN(n4682) );
  OAI221_X1 U5189 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput25), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput61), .A(n4682), .ZN(n4687) );
  AOI22_X1 U5190 ( .A1(REG0_REG_5__SCAN_IN), .A2(keyinput49), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput44), .ZN(n4683) );
  OAI221_X1 U5191 ( .B1(REG0_REG_5__SCAN_IN), .B2(keyinput49), .C1(
        D_REG_6__SCAN_IN), .C2(keyinput44), .A(n4683), .ZN(n4686) );
  AOI22_X1 U5192 ( .A1(REG2_REG_0__SCAN_IN), .A2(keyinput41), .B1(
        IR_REG_29__SCAN_IN), .B2(keyinput20), .ZN(n4684) );
  OAI221_X1 U5193 ( .B1(REG2_REG_0__SCAN_IN), .B2(keyinput41), .C1(
        IR_REG_29__SCAN_IN), .C2(keyinput20), .A(n4684), .ZN(n4685) );
  NOR4_X1 U5194 ( .A1(n4688), .A2(n4687), .A3(n4686), .A4(n4685), .ZN(n4689)
         );
  NAND4_X1 U5195 ( .A1(n4692), .A2(n4691), .A3(n4690), .A4(n4689), .ZN(n4751)
         );
  INV_X1 U5196 ( .A(DATAI_20_), .ZN(n4694) );
  AOI22_X1 U5197 ( .A1(n4069), .A2(keyinput36), .B1(n4694), .B2(keyinput56), 
        .ZN(n4693) );
  OAI221_X1 U5198 ( .B1(n4069), .B2(keyinput36), .C1(n4694), .C2(keyinput56), 
        .A(n4693), .ZN(n4707) );
  AOI22_X1 U5199 ( .A1(n4697), .A2(keyinput57), .B1(keyinput53), .B2(n4696), 
        .ZN(n4695) );
  OAI221_X1 U5200 ( .B1(n4697), .B2(keyinput57), .C1(n4696), .C2(keyinput53), 
        .A(n4695), .ZN(n4706) );
  INV_X1 U5201 ( .A(DATAI_6_), .ZN(n4699) );
  AOI22_X1 U5202 ( .A1(n4700), .A2(keyinput45), .B1(keyinput29), .B2(n4699), 
        .ZN(n4698) );
  OAI221_X1 U5203 ( .B1(n4700), .B2(keyinput45), .C1(n4699), .C2(keyinput29), 
        .A(n4698), .ZN(n4705) );
  XOR2_X1 U5204 ( .A(n4701), .B(keyinput4), .Z(n4703) );
  XNOR2_X1 U5205 ( .A(REG2_REG_2__SCAN_IN), .B(keyinput28), .ZN(n4702) );
  NAND2_X1 U5206 ( .A1(n4703), .A2(n4702), .ZN(n4704) );
  NOR4_X1 U5207 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n4749)
         );
  AOI22_X1 U5208 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput24), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput17), .ZN(n4708) );
  OAI221_X1 U5209 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput24), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput17), .A(n4708), .ZN(n4711) );
  AOI22_X1 U5210 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput8), .B1(
        IR_REG_14__SCAN_IN), .B2(keyinput33), .ZN(n4709) );
  OAI221_X1 U5211 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput8), .C1(
        IR_REG_14__SCAN_IN), .C2(keyinput33), .A(n4709), .ZN(n4710) );
  NOR2_X1 U5212 ( .A1(n4711), .A2(n4710), .ZN(n4719) );
  INV_X1 U5213 ( .A(keyinput9), .ZN(n4712) );
  XNOR2_X1 U5214 ( .A(n4713), .B(n4712), .ZN(n4718) );
  XNOR2_X1 U5215 ( .A(IR_REG_12__SCAN_IN), .B(keyinput5), .ZN(n4717) );
  AOI22_X1 U5216 ( .A1(REG1_REG_31__SCAN_IN), .A2(keyinput13), .B1(
        IR_REG_22__SCAN_IN), .B2(keyinput1), .ZN(n4714) );
  OAI221_X1 U5217 ( .B1(REG1_REG_31__SCAN_IN), .B2(keyinput13), .C1(
        IR_REG_22__SCAN_IN), .C2(keyinput1), .A(n4714), .ZN(n4715) );
  INV_X1 U5218 ( .A(n4715), .ZN(n4716) );
  AND4_X1 U5219 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4748)
         );
  AOI22_X1 U5220 ( .A1(n2548), .A2(keyinput26), .B1(keyinput18), .B2(n4721), 
        .ZN(n4720) );
  OAI221_X1 U5221 ( .B1(n2548), .B2(keyinput26), .C1(n4721), .C2(keyinput18), 
        .A(n4720), .ZN(n4732) );
  AOI22_X1 U5222 ( .A1(n4724), .A2(keyinput42), .B1(keyinput38), .B2(n4723), 
        .ZN(n4722) );
  OAI221_X1 U5223 ( .B1(n4724), .B2(keyinput42), .C1(n4723), .C2(keyinput38), 
        .A(n4722), .ZN(n4731) );
  XOR2_X1 U5224 ( .A(n3427), .B(keyinput22), .Z(n4727) );
  XNOR2_X1 U5225 ( .A(IR_REG_27__SCAN_IN), .B(keyinput31), .ZN(n4726) );
  XNOR2_X1 U5226 ( .A(IR_REG_31__SCAN_IN), .B(keyinput10), .ZN(n4725) );
  NAND3_X1 U5227 ( .A1(n4727), .A2(n4726), .A3(n4725), .ZN(n4730) );
  XNOR2_X1 U5228 ( .A(n4728), .B(keyinput19), .ZN(n4729) );
  NOR4_X1 U5229 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n4729), .ZN(n4747)
         );
  INV_X1 U5230 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4735) );
  AOI22_X1 U5231 ( .A1(n4735), .A2(keyinput0), .B1(n4734), .B2(keyinput62), 
        .ZN(n4733) );
  OAI221_X1 U5232 ( .B1(n4735), .B2(keyinput0), .C1(n4734), .C2(keyinput62), 
        .A(n4733), .ZN(n4745) );
  AOI22_X1 U5233 ( .A1(n2916), .A2(keyinput63), .B1(n4182), .B2(keyinput58), 
        .ZN(n4736) );
  OAI221_X1 U5234 ( .B1(n2916), .B2(keyinput63), .C1(n4182), .C2(keyinput58), 
        .A(n4736), .ZN(n4744) );
  AOI22_X1 U5235 ( .A1(n4739), .A2(keyinput59), .B1(n4738), .B2(keyinput55), 
        .ZN(n4737) );
  OAI221_X1 U5236 ( .B1(n4739), .B2(keyinput59), .C1(n4738), .C2(keyinput55), 
        .A(n4737), .ZN(n4743) );
  XNOR2_X1 U5237 ( .A(REG1_REG_26__SCAN_IN), .B(keyinput51), .ZN(n4741) );
  XNOR2_X1 U5238 ( .A(IR_REG_11__SCAN_IN), .B(keyinput47), .ZN(n4740) );
  NAND2_X1 U5239 ( .A1(n4741), .A2(n4740), .ZN(n4742) );
  NOR4_X1 U5240 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4746)
         );
  NAND4_X1 U5241 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n4750)
         );
  AOI211_X1 U5242 ( .C1(n4753), .C2(n4752), .A(n4751), .B(n4750), .ZN(n4758)
         );
  NAND2_X1 U5243 ( .A1(n4754), .A2(n4756), .ZN(n4755) );
  OAI21_X1 U5244 ( .B1(REG0_REG_5__SCAN_IN), .B2(n4756), .A(n4755), .ZN(n4757)
         );
  XNOR2_X1 U5245 ( .A(n4758), .B(n4757), .ZN(U3477) );
endmodule

