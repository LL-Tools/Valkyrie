

module b21_C_AntiSAT_k_128_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137;

  INV_X2 U4820 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OR2_X1 U4821 ( .A1(n9223), .A2(n9354), .ZN(n9209) );
  BUF_X1 U4822 ( .A(n5097), .Z(n5675) );
  NAND2_X1 U4823 ( .A1(n5140), .A2(n5139), .ZN(n9704) );
  OAI211_X1 U4824 ( .C1(n5856), .C2(n6095), .A(n5810), .B(n5809), .ZN(n7965)
         );
  OAI211_X2 U4825 ( .C1(n5290), .C2(n6088), .A(n5048), .B(n5047), .ZN(n9676)
         );
  INV_X1 U4826 ( .A(n5622), .ZN(n5051) );
  INV_X1 U4827 ( .A(n7956), .ZN(n7790) );
  INV_X1 U4828 ( .A(n7082), .ZN(n5800) );
  AND2_X1 U4831 ( .A1(n4941), .A2(n6495), .ZN(n4940) );
  INV_X2 U4832 ( .A(n5096), .ZN(n4935) );
  NAND2_X1 U4833 ( .A1(n6147), .A2(n5590), .ZN(n4939) );
  AND4_X1 U4834 ( .A1(n5729), .A2(n5728), .A3(n5727), .A4(n5726), .ZN(n5733)
         );
  CLKBUF_X1 U4835 ( .A(n8165), .Z(n4315) );
  OAI21_X1 U4836 ( .B1(n6075), .B2(n6060), .A(n8485), .ZN(n8165) );
  INV_X2 U4837 ( .A(n9763), .ZN(n8467) );
  INV_X1 U4839 ( .A(n7953), .ZN(n7829) );
  CLKBUF_X2 U4840 ( .A(n4940), .Z(n5549) );
  INV_X1 U4841 ( .A(n4940), .ZN(n5672) );
  INV_X1 U4842 ( .A(n4939), .ZN(n5040) );
  INV_X1 U4843 ( .A(n6263), .ZN(n7515) );
  OAI21_X1 U4844 ( .B1(n8404), .B2(n4736), .A(n4354), .ZN(n8351) );
  NAND2_X1 U4845 ( .A1(n8719), .A2(n8715), .ZN(n8659) );
  CLKBUF_X2 U4846 ( .A(n5030), .Z(n5683) );
  NOR2_X1 U4847 ( .A1(n9321), .A2(n9676), .ZN(n9608) );
  INV_X1 U4848 ( .A(n6672), .ZN(n9683) );
  INV_X1 U4849 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4880) );
  OAI21_X1 U4850 ( .B1(n5263), .B2(n4898), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4903) );
  NAND2_X1 U4851 ( .A1(n4787), .A2(n5072), .ZN(n5090) );
  NAND2_X1 U4852 ( .A1(n5245), .A2(n5244), .ZN(n9400) );
  NAND2_X1 U4853 ( .A1(n5185), .A2(n5184), .ZN(n7426) );
  INV_X1 U4854 ( .A(n4914), .ZN(n7775) );
  XNOR2_X1 U4855 ( .A(n5090), .B(n5088), .ZN(n6098) );
  BUF_X1 U4856 ( .A(n4925), .Z(n7118) );
  INV_X2 U4857 ( .A(n7995), .ZN(n7593) );
  NAND2_X1 U4858 ( .A1(n5503), .A2(n5504), .ZN(n8652) );
  OAI21_X2 U4859 ( .B1(n7123), .B2(n7120), .A(n7121), .ZN(n5258) );
  OAI21_X2 U4860 ( .B1(n5788), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5787) );
  NAND2_X2 U4861 ( .A1(n7137), .A2(n7134), .ZN(n7123) );
  OAI21_X2 U4862 ( .B1(n8659), .B2(n4657), .A(n4654), .ZN(n8671) );
  AOI21_X2 U4863 ( .B1(n8700), .B2(n8701), .A(n5481), .ZN(n5503) );
  XNOR2_X2 U4864 ( .A(n4963), .B(n4916), .ZN(n4962) );
  XNOR2_X2 U4865 ( .A(n4517), .B(n4516), .ZN(n9072) );
  NAND2_X1 U4866 ( .A1(n4748), .A2(n4362), .ZN(n7467) );
  BUF_X2 U4867 ( .A(n5049), .Z(n5552) );
  INV_X1 U4868 ( .A(n6513), .ZN(n6313) );
  INV_X2 U4869 ( .A(n8170), .ZN(n9820) );
  INV_X2 U4870 ( .A(n5067), .ZN(n8733) );
  NAND2_X2 U4871 ( .A1(n6502), .A2(n8999), .ZN(n5580) );
  BUF_X2 U4872 ( .A(n5026), .Z(n8093) );
  AND2_X2 U4873 ( .A1(n5767), .A2(n5766), .ZN(n5816) );
  AND4_X1 U4874 ( .A1(n5731), .A2(n5730), .A3(n5898), .A4(n5839), .ZN(n5732)
         );
  AND2_X1 U4875 ( .A1(n4425), .A2(n4424), .ZN(n7964) );
  NOR2_X1 U4876 ( .A1(n4669), .A2(n4482), .ZN(n4481) );
  NAND2_X1 U4877 ( .A1(n5388), .A2(n5387), .ZN(n8715) );
  AOI22_X1 U4878 ( .A1(n4848), .A2(n4318), .B1(n9272), .B2(n4329), .ZN(n9222)
         );
  AOI21_X1 U4879 ( .B1(n9286), .B2(n8075), .A(n8074), .ZN(n9272) );
  NAND2_X1 U4880 ( .A1(n8073), .A2(n8072), .ZN(n9286) );
  OR2_X1 U4881 ( .A1(n7644), .A2(n8896), .ZN(n8073) );
  AND2_X1 U4882 ( .A1(n7391), .A2(n4610), .ZN(n9287) );
  NOR2_X1 U4883 ( .A1(n8045), .A2(n8602), .ZN(n8488) );
  AND2_X1 U4884 ( .A1(n7862), .A2(n7859), .ZN(n7799) );
  AND2_X1 U4885 ( .A1(n7854), .A2(n7858), .ZN(n7853) );
  XNOR2_X1 U4886 ( .A(n5179), .B(n4860), .ZN(n6184) );
  NAND2_X1 U4887 ( .A1(n5122), .A2(n5121), .ZN(n7096) );
  NAND2_X2 U4888 ( .A1(n6745), .A2(n8485), .ZN(n9763) );
  NAND2_X1 U4889 ( .A1(n5093), .A2(n5092), .ZN(n5112) );
  INV_X2 U4890 ( .A(n9646), .ZN(n9648) );
  CLKBUF_X1 U4891 ( .A(n6559), .Z(n9666) );
  NAND2_X1 U4892 ( .A1(n5039), .A2(n5038), .ZN(n5070) );
  OAI211_X1 U4893 ( .C1(n5290), .C2(n6091), .A(n5000), .B(n4999), .ZN(n6513)
         );
  NAND2_X2 U4894 ( .A1(n7290), .A2(n4933), .ZN(n5049) );
  NAND2_X1 U4895 ( .A1(n5007), .A2(n5006), .ZN(n5036) );
  AND4_X1 U4896 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n6790)
         );
  AND2_X2 U4897 ( .A1(n6132), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND4_X1 U4898 ( .A1(n4948), .A2(n4947), .A3(n4946), .A4(n4945), .ZN(n6488)
         );
  INV_X1 U4899 ( .A(n8080), .ZN(n5290) );
  AND4_X1 U4900 ( .A1(n4987), .A2(n4986), .A3(n4985), .A4(n4984), .ZN(n6620)
         );
  NAND4_X2 U4901 ( .A1(n4888), .A2(n4887), .A3(n4886), .A4(n4885), .ZN(n6489)
         );
  AND4_X1 U4902 ( .A1(n5804), .A2(n5803), .A3(n5802), .A4(n5801), .ZN(n6412)
         );
  AND2_X1 U4903 ( .A1(n4939), .A2(n7775), .ZN(n8080) );
  NAND2_X1 U4904 ( .A1(n4993), .A2(n4992), .ZN(n5003) );
  NAND2_X1 U4905 ( .A1(n4941), .A2(n4933), .ZN(n5096) );
  OR2_X2 U4906 ( .A1(n6052), .A2(n7956), .ZN(n9881) );
  CLKBUF_X1 U4907 ( .A(n4941), .Z(n5723) );
  NAND2_X2 U4908 ( .A1(n8014), .A2(n7953), .ZN(n6052) );
  AND2_X2 U4909 ( .A1(n5765), .A2(n5766), .ZN(n7764) );
  AND2_X1 U4910 ( .A1(n9423), .A2(n4884), .ZN(n5026) );
  AND2_X1 U4911 ( .A1(n9426), .A2(n9423), .ZN(n5030) );
  XNOR2_X1 U4912 ( .A(n4893), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5554) );
  AND2_X1 U4913 ( .A1(n4883), .A2(n4884), .ZN(n5025) );
  INV_X1 U4914 ( .A(n4884), .ZN(n9426) );
  XNOR2_X1 U4915 ( .A(n4931), .B(n5573), .ZN(n5579) );
  NAND2_X2 U4916 ( .A1(n4902), .A2(n4923), .ZN(n4926) );
  XNOR2_X1 U4917 ( .A(n4877), .B(n4876), .ZN(n4883) );
  NAND2_X1 U4918 ( .A1(n4892), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4893) );
  OAI211_X1 U4919 ( .C1(n4882), .C2(n4875), .A(n4879), .B(n4881), .ZN(n4884)
         );
  NAND2_X1 U4920 ( .A1(n5776), .A2(n5778), .ZN(n6280) );
  NAND2_X1 U4921 ( .A1(n4786), .A2(n5764), .ZN(n8642) );
  NAND2_X1 U4922 ( .A1(n4909), .A2(n4908), .ZN(n4911) );
  OAI21_X1 U4923 ( .B1(n5393), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4994), .ZN(
        n5004) );
  XNOR2_X1 U4924 ( .A(n4891), .B(n4653), .ZN(n7318) );
  NAND2_X1 U4925 ( .A1(n5760), .A2(n5757), .ZN(n5782) );
  INV_X1 U4926 ( .A(n6541), .ZN(n6542) );
  CLKBUF_X1 U4927 ( .A(n4895), .Z(n5263) );
  NAND2_X1 U4928 ( .A1(n4817), .A2(n4815), .ZN(n4965) );
  AND4_X1 U4929 ( .A1(n4458), .A2(n4457), .A3(n4865), .A4(n4864), .ZN(n4866)
         );
  NOR3_X1 U4930 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_26__SCAN_IN), .ZN(n4874) );
  INV_X1 U4931 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4896) );
  NOR2_X1 U4932 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4454) );
  NOR2_X1 U4933 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4453) );
  INV_X1 U4934 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5264) );
  NOR2_X1 U4935 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4456) );
  NOR2_X1 U4936 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4455) );
  INV_X1 U4937 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5572) );
  NOR2_X1 U4938 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4457) );
  NOR2_X1 U4939 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4458) );
  INV_X1 U4940 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5573) );
  INV_X2 U4941 ( .A(n6492), .ZN(n4970) );
  AND3_X2 U4942 ( .A1(n4969), .A2(n4968), .A3(n4967), .ZN(n6492) );
  NAND2_X2 U4943 ( .A1(n4911), .A2(n4910), .ZN(n5590) );
  OAI22_X2 U4944 ( .A1(n6436), .A2(n4648), .B1(n4647), .B2(n6437), .ZN(n6516)
         );
  NAND2_X1 U4945 ( .A1(n5061), .A2(n5060), .ZN(n6436) );
  AOI21_X2 U4946 ( .B1(n8649), .B2(n8682), .A(n8681), .ZN(n8685) );
  XNOR2_X2 U4947 ( .A(n4906), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U4948 ( .A1(n5260), .A2(n5259), .ZN(n4814) );
  OR2_X1 U4949 ( .A1(n9333), .A2(n9173), .ZN(n8987) );
  OR2_X2 U4950 ( .A1(n4926), .A2(n9032), .ZN(n4933) );
  NAND2_X1 U4951 ( .A1(n4418), .A2(n7656), .ZN(n7758) );
  NAND2_X1 U4952 ( .A1(n7653), .A2(n7652), .ZN(n4418) );
  NAND2_X1 U4953 ( .A1(n5510), .A2(n5509), .ZN(n5537) );
  NAND2_X1 U4954 ( .A1(n4814), .A2(n5261), .ZN(n5282) );
  NAND2_X1 U4955 ( .A1(n7827), .A2(n7947), .ZN(n4524) );
  NAND2_X1 U4956 ( .A1(n4546), .A2(n7874), .ZN(n4545) );
  NAND2_X1 U4957 ( .A1(n4558), .A2(n8384), .ZN(n4557) );
  INV_X1 U4958 ( .A(n5341), .ZN(n4583) );
  INV_X1 U4959 ( .A(n5180), .ZN(n4800) );
  NAND2_X1 U4960 ( .A1(n5159), .A2(n4862), .ZN(n5161) );
  OAI21_X1 U4961 ( .B1(n4686), .B2(n4573), .A(n4580), .ZN(n4572) );
  AOI21_X1 U4962 ( .B1(n4762), .B2(n8308), .A(n4764), .ZN(n4760) );
  INV_X1 U4963 ( .A(n5767), .ZN(n5765) );
  OR2_X1 U4964 ( .A1(n8533), .A2(n8007), .ZN(n7940) );
  OR2_X1 U4965 ( .A1(n8582), .A2(n7676), .ZN(n7910) );
  OR2_X1 U4966 ( .A1(n8602), .A2(n8497), .ZN(n7895) );
  OR2_X1 U4967 ( .A1(n8607), .A2(n7535), .ZN(n7889) );
  NAND2_X1 U4968 ( .A1(n8507), .A2(n9831), .ZN(n9743) );
  OAI21_X1 U4969 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n6038), .A(n9800), .ZN(n6410)
         );
  AND2_X1 U4970 ( .A1(n6048), .A2(n9766), .ZN(n6739) );
  INV_X1 U4971 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5757) );
  NOR2_X1 U4972 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4682) );
  OR2_X1 U4973 ( .A1(n5929), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5931) );
  OR2_X1 U4974 ( .A1(n4507), .A2(n6160), .ZN(n4506) );
  INV_X1 U4975 ( .A(n6157), .ZN(n4507) );
  INV_X1 U4976 ( .A(n9563), .ZN(n4508) );
  AOI21_X1 U4977 ( .B1(n4790), .B2(n8982), .A(n8089), .ZN(n4789) );
  INV_X1 U4978 ( .A(n4483), .ZN(n9187) );
  OR2_X1 U4979 ( .A1(n7399), .A2(n7398), .ZN(n7403) );
  NAND2_X1 U4980 ( .A1(n4894), .A2(n5554), .ZN(n4941) );
  NOR2_X1 U4981 ( .A1(n7479), .A2(n7318), .ZN(n4894) );
  OAI21_X1 U4982 ( .B1(n5484), .B2(n5483), .A(n5482), .ZN(n5508) );
  NAND2_X1 U4983 ( .A1(n8024), .A2(n7980), .ZN(n7981) );
  NAND2_X1 U4984 ( .A1(n6263), .A2(n7775), .ZN(n5869) );
  AND2_X1 U4985 ( .A1(n7732), .A2(n7731), .ZN(n8143) );
  CLKBUF_X1 U4986 ( .A(n7082), .Z(n7742) );
  INV_X1 U4987 ( .A(n5816), .ZN(n7763) );
  NAND2_X1 U4988 ( .A1(n5767), .A2(n8642), .ZN(n7082) );
  AND2_X1 U4989 ( .A1(n7940), .A2(n7941), .ZN(n8053) );
  OR2_X1 U4990 ( .A1(n8543), .A2(n8340), .ZN(n8042) );
  AOI21_X1 U4991 ( .B1(n8408), .B2(n4739), .A(n4330), .ZN(n4737) );
  NAND2_X1 U4992 ( .A1(n4745), .A2(n8038), .ZN(n4744) );
  NAND2_X1 U4993 ( .A1(n4742), .A2(n4746), .ZN(n4741) );
  INV_X1 U4994 ( .A(n8404), .ZN(n4742) );
  AND2_X1 U4995 ( .A1(n7919), .A2(n7918), .ZN(n8379) );
  INV_X1 U4996 ( .A(n4732), .ZN(n4731) );
  OR2_X1 U4997 ( .A1(n8612), .A2(n7451), .ZN(n7883) );
  AOI21_X1 U4998 ( .B1(n6987), .B2(n7800), .A(n4775), .ZN(n4863) );
  INV_X1 U4999 ( .A(n7872), .ZN(n4775) );
  NOR2_X2 U5000 ( .A1(n6539), .A2(n4480), .ZN(n5760) );
  NAND2_X1 U5001 ( .A1(n9632), .A2(n4940), .ZN(n4975) );
  AND4_X1 U5002 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(n8079)
         );
  NAND2_X1 U5004 ( .A1(n6661), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4501) );
  NOR2_X1 U5005 ( .A1(n4353), .A2(n4845), .ZN(n4844) );
  INV_X1 U5006 ( .A(n4335), .ZN(n4845) );
  AND2_X1 U5007 ( .A1(n9264), .A2(n9280), .ZN(n4850) );
  NAND2_X1 U5008 ( .A1(n9317), .A2(n4829), .ZN(n9606) );
  AND2_X1 U5009 ( .A1(n6680), .A2(n6679), .ZN(n4829) );
  XNOR2_X1 U5010 ( .A(n9632), .B(n6492), .ZN(n6526) );
  NOR2_X1 U5011 ( .A1(n6488), .A2(n9637), .ZN(n9629) );
  INV_X1 U5012 ( .A(n9616), .ZN(n9631) );
  NAND2_X1 U5013 ( .A1(n8082), .A2(n8081), .ZN(n9327) );
  NAND2_X1 U5014 ( .A1(n5665), .A2(n5664), .ZN(n9333) );
  AND2_X1 U5015 ( .A1(n6249), .A2(n5583), .ZN(n9677) );
  OR2_X1 U5016 ( .A1(n6251), .A2(n9032), .ZN(n9706) );
  NAND2_X1 U5017 ( .A1(n7118), .A2(n4926), .ZN(n6251) );
  INV_X1 U5018 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4876) );
  NAND2_X1 U5019 ( .A1(n4879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U5020 ( .A1(n4416), .A2(n5535), .ZN(n5611) );
  OR2_X1 U5021 ( .A1(n5537), .A2(n5536), .ZN(n4416) );
  XNOR2_X1 U5022 ( .A(n4903), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U5023 ( .A1(n4584), .A2(n4590), .ZN(n5340) );
  NAND2_X1 U5024 ( .A1(n5282), .A2(n4592), .ZN(n4584) );
  AOI21_X1 U5025 ( .B1(n8102), .B2(n9313), .A(n4861), .ZN(n9330) );
  NAND2_X1 U5026 ( .A1(n4530), .A2(n4520), .ZN(n4519) );
  NAND2_X1 U5027 ( .A1(n7834), .A2(n7833), .ZN(n4530) );
  AND2_X1 U5028 ( .A1(n4524), .A2(n4525), .ZN(n4520) );
  NAND2_X1 U5029 ( .A1(n4548), .A2(n7939), .ZN(n4547) );
  NAND2_X1 U5030 ( .A1(n4545), .A2(n7947), .ZN(n4544) );
  NAND2_X1 U5031 ( .A1(n4550), .A2(n4549), .ZN(n4548) );
  OAI211_X1 U5032 ( .C1(n7916), .C2(n7947), .A(n4556), .B(n4553), .ZN(n7921)
         );
  AND2_X1 U5033 ( .A1(n8379), .A2(n4554), .ZN(n4553) );
  NAND2_X1 U5034 ( .A1(n4557), .A2(n7947), .ZN(n4556) );
  OAI21_X1 U5035 ( .B1(n4538), .B2(n4537), .A(n4536), .ZN(n7933) );
  AND2_X1 U5036 ( .A1(n7929), .A2(n7947), .ZN(n4537) );
  NOR2_X1 U5037 ( .A1(n8323), .A2(n7932), .ZN(n4536) );
  AOI21_X1 U5038 ( .B1(n4542), .B2(n4540), .A(n4539), .ZN(n4538) );
  OAI21_X1 U5039 ( .B1(n7887), .B2(n4770), .A(n7894), .ZN(n4769) );
  INV_X1 U5040 ( .A(n7889), .ZN(n4770) );
  INV_X1 U5041 ( .A(n7895), .ZN(n4767) );
  INV_X1 U5042 ( .A(n4585), .ZN(n4405) );
  NAND2_X1 U5043 ( .A1(n4585), .A2(n4404), .ZN(n4403) );
  AOI21_X1 U5044 ( .B1(n4585), .B2(n4588), .A(n4583), .ZN(n4582) );
  INV_X1 U5045 ( .A(n5261), .ZN(n4404) );
  INV_X1 U5046 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4818) );
  NAND2_X1 U5047 ( .A1(n6705), .A2(n5868), .ZN(n8106) );
  NOR2_X1 U5048 ( .A1(n7974), .A2(n4573), .ZN(n4576) );
  INV_X1 U5049 ( .A(n4690), .ZN(n4575) );
  INV_X1 U5050 ( .A(n7974), .ZN(n4571) );
  NAND2_X1 U5051 ( .A1(n4689), .A2(n7307), .ZN(n4695) );
  NOR2_X1 U5052 ( .A1(n7593), .A2(n4596), .ZN(n4598) );
  XNOR2_X1 U5053 ( .A(n8178), .B(n7593), .ZN(n5922) );
  OR2_X1 U5054 ( .A1(n7781), .A2(n7780), .ZN(n7946) );
  AND2_X1 U5055 ( .A1(n7790), .A2(n8499), .ZN(n6061) );
  INV_X1 U5056 ( .A(n7922), .ZN(n4782) );
  OAI21_X1 U5057 ( .B1(n8039), .B2(n4782), .A(n7926), .ZN(n4781) );
  OAI21_X1 U5058 ( .B1(n4756), .B2(n4475), .A(n7682), .ZN(n4474) );
  NOR2_X1 U5059 ( .A1(n8397), .A2(n4680), .ZN(n4679) );
  INV_X1 U5060 ( .A(n4681), .ZN(n4680) );
  INV_X1 U5061 ( .A(n4757), .ZN(n4754) );
  OR2_X1 U5062 ( .A1(n8599), .A2(n7673), .ZN(n7824) );
  NOR2_X1 U5063 ( .A1(n8492), .A2(n4733), .ZN(n4732) );
  INV_X1 U5064 ( .A(n8025), .ZN(n4733) );
  NOR2_X1 U5065 ( .A1(n7881), .A2(n7148), .ZN(n4677) );
  INV_X1 U5066 ( .A(n6961), .ZN(n4716) );
  INV_X1 U5067 ( .A(n6983), .ZN(n4719) );
  NAND2_X1 U5068 ( .A1(n4715), .A2(n7853), .ZN(n4714) );
  NAND2_X1 U5069 ( .A1(n6965), .A2(n6970), .ZN(n4720) );
  AND2_X1 U5070 ( .A1(n7853), .A2(n7851), .ZN(n4771) );
  NAND2_X1 U5071 ( .A1(n6862), .A2(n4773), .ZN(n4772) );
  NOR2_X1 U5072 ( .A1(n6863), .A2(n4774), .ZN(n4773) );
  INV_X1 U5073 ( .A(n7848), .ZN(n4774) );
  AND2_X1 U5074 ( .A1(n7851), .A2(n7850), .ZN(n7847) );
  NAND2_X1 U5075 ( .A1(n7836), .A2(n6836), .ZN(n7831) );
  NAND2_X1 U5076 ( .A1(n6691), .A2(n9820), .ZN(n7839) );
  INV_X1 U5077 ( .A(n8507), .ZN(n6860) );
  NOR2_X1 U5078 ( .A1(n6539), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6541) );
  NOR2_X1 U5079 ( .A1(n5931), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5967) );
  INV_X1 U5080 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5870) );
  INV_X1 U5081 ( .A(n5439), .ZN(n4655) );
  INV_X1 U5082 ( .A(n5723), .ZN(n4942) );
  NAND2_X1 U5083 ( .A1(n4664), .A2(n4663), .ZN(n4662) );
  INV_X1 U5084 ( .A(n8661), .ZN(n4663) );
  INV_X1 U5085 ( .A(n8660), .ZN(n4664) );
  NOR2_X1 U5086 ( .A1(n9200), .A2(n4843), .ZN(n4842) );
  NOR2_X1 U5087 ( .A1(n4844), .A2(n4320), .ZN(n4843) );
  OR2_X1 U5088 ( .A1(n9364), .A2(n8676), .ZN(n8973) );
  AND2_X1 U5089 ( .A1(n9285), .A2(n9294), .ZN(n4794) );
  AND2_X1 U5090 ( .A1(n4613), .A2(n4614), .ZN(n4612) );
  NOR2_X1 U5091 ( .A1(n7623), .A2(n9395), .ZN(n4614) );
  NOR2_X1 U5092 ( .A1(n8938), .A2(n4437), .ZN(n4436) );
  INV_X1 U5093 ( .A(n8934), .ZN(n4437) );
  AOI21_X1 U5094 ( .B1(n7419), .B2(n7327), .A(n4357), .ZN(n7330) );
  NOR2_X1 U5095 ( .A1(n5079), .A2(n5078), .ZN(n5104) );
  XNOR2_X1 U5096 ( .A(n4643), .B(n6489), .ZN(n8874) );
  NAND2_X1 U5097 ( .A1(n4447), .A2(n4446), .ZN(n9615) );
  NAND2_X1 U5098 ( .A1(n4361), .A2(n8945), .ZN(n4446) );
  OAI21_X1 U5099 ( .B1(n7758), .B2(n7661), .A(n7660), .ZN(n7774) );
  NAND2_X1 U5100 ( .A1(n5661), .A2(n5660), .ZN(n7653) );
  NAND2_X1 U5101 ( .A1(n4417), .A2(n5632), .ZN(n5659) );
  NAND2_X1 U5102 ( .A1(n4410), .A2(n4407), .ZN(n4417) );
  AOI21_X1 U5103 ( .B1(n4412), .B2(n4409), .A(n4408), .ZN(n4407) );
  OR2_X1 U5104 ( .A1(n5537), .A2(n4411), .ZN(n4410) );
  NOR2_X1 U5105 ( .A1(n5610), .A2(n4415), .ZN(n4414) );
  INV_X1 U5106 ( .A(n5535), .ZN(n4415) );
  AOI21_X1 U5107 ( .B1(n4414), .B2(n5536), .A(n4413), .ZN(n4412) );
  INV_X1 U5108 ( .A(n5609), .ZN(n4413) );
  AND2_X1 U5109 ( .A1(n5509), .A2(n5490), .ZN(n5507) );
  OAI21_X1 U5110 ( .B1(n5459), .B2(n4423), .A(n5462), .ZN(n5484) );
  INV_X1 U5111 ( .A(n5460), .ZN(n4423) );
  OAI21_X1 U5112 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n5441) );
  AND2_X1 U5113 ( .A1(n5442), .A2(n5420), .ZN(n5440) );
  NOR2_X1 U5114 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4927) );
  NAND2_X1 U5115 ( .A1(n4402), .A2(n4400), .ZN(n5416) );
  AOI21_X1 U5116 ( .B1(n4317), .B2(n4344), .A(n4401), .ZN(n4400) );
  NAND2_X1 U5117 ( .A1(n4814), .A2(n4348), .ZN(n4402) );
  INV_X1 U5118 ( .A(n4792), .ZN(n4401) );
  OAI21_X1 U5119 ( .B1(n4814), .B2(n4405), .A(n4317), .ZN(n5369) );
  NAND2_X1 U5120 ( .A1(n4873), .A2(n4857), .ZN(n5343) );
  AND2_X1 U5121 ( .A1(n4797), .A2(n4802), .ZN(n4795) );
  INV_X1 U5122 ( .A(n5232), .ZN(n4802) );
  NAND2_X1 U5123 ( .A1(n5112), .A2(n5111), .ZN(n4421) );
  AOI21_X1 U5124 ( .B1(n4703), .B2(n4701), .A(n4700), .ZN(n4699) );
  INV_X1 U5125 ( .A(n7987), .ZN(n4700) );
  INV_X1 U5126 ( .A(n4707), .ZN(n4701) );
  NAND2_X1 U5127 ( .A1(n7586), .A2(n7587), .ZN(n4580) );
  NAND2_X1 U5128 ( .A1(n8158), .A2(n8157), .ZN(n4565) );
  NAND2_X1 U5129 ( .A1(n6921), .A2(n6920), .ZN(n7062) );
  NAND2_X1 U5130 ( .A1(n8132), .A2(n8131), .ZN(n4569) );
  NOR2_X1 U5131 ( .A1(n7984), .A2(n4564), .ZN(n4563) );
  INV_X1 U5132 ( .A(n8131), .ZN(n4564) );
  NAND2_X1 U5133 ( .A1(n6637), .A2(n5961), .ZN(n6645) );
  INV_X1 U5134 ( .A(n7985), .ZN(n5895) );
  OR2_X1 U5135 ( .A1(n7311), .A2(n6117), .ZN(n7522) );
  AND2_X1 U5136 ( .A1(n4687), .A2(n4693), .ZN(n4686) );
  AOI21_X1 U5137 ( .B1(n4390), .B2(n4854), .A(n4694), .ZN(n4693) );
  NAND2_X1 U5138 ( .A1(n4689), .A2(n4688), .ZN(n4687) );
  INV_X1 U5139 ( .A(n7553), .ZN(n4694) );
  NAND2_X1 U5140 ( .A1(n4691), .A2(n4390), .ZN(n4690) );
  INV_X1 U5141 ( .A(n4695), .ZN(n4691) );
  OR2_X1 U5142 ( .A1(n6078), .A2(n9765), .ZN(n6075) );
  AND2_X1 U5143 ( .A1(n8140), .A2(n8139), .ZN(n4705) );
  NOR2_X1 U5144 ( .A1(n8292), .A2(n8294), .ZN(n7949) );
  NAND2_X1 U5145 ( .A1(n4759), .A2(n4758), .ZN(n7783) );
  AOI21_X1 U5146 ( .B1(n4760), .B2(n4761), .A(n4319), .ZN(n4758) );
  AND2_X1 U5147 ( .A1(n7946), .A2(n7943), .ZN(n7818) );
  AND3_X1 U5148 ( .A1(n7526), .A2(n7525), .A3(n7524), .ZN(n7676) );
  OR2_X1 U5149 ( .A1(n6326), .A2(n6325), .ZN(n4626) );
  NAND2_X1 U5150 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  NAND2_X1 U5151 ( .A1(n6271), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4625) );
  AND2_X1 U5152 ( .A1(n4624), .A2(n4623), .ZN(n6336) );
  INV_X1 U5153 ( .A(n6337), .ZN(n4623) );
  NOR2_X1 U5154 ( .A1(n6600), .A2(n4382), .ZN(n6604) );
  NOR2_X1 U5155 ( .A1(n7026), .A2(n4634), .ZN(n7028) );
  AND2_X1 U5156 ( .A1(n7027), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4634) );
  NOR2_X1 U5157 ( .A1(n8252), .A2(n8251), .ZN(n8263) );
  NOR2_X1 U5158 ( .A1(n8263), .A2(n4627), .ZN(n8274) );
  AND2_X1 U5159 ( .A1(n8264), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5160 ( .A1(n4459), .A2(n7931), .ZN(n8318) );
  OR2_X1 U5161 ( .A1(n8554), .A2(n8339), .ZN(n8040) );
  NAND2_X1 U5162 ( .A1(n7708), .A2(n8039), .ZN(n8374) );
  INV_X1 U5163 ( .A(n4744), .ZN(n4740) );
  INV_X1 U5164 ( .A(n4725), .ZN(n4724) );
  AND2_X1 U5165 ( .A1(n7910), .A2(n8452), .ZN(n4757) );
  OR2_X1 U5166 ( .A1(n8588), .A2(n8476), .ZN(n8031) );
  AND2_X1 U5167 ( .A1(n7910), .A2(n7911), .ZN(n8437) );
  AND2_X1 U5168 ( .A1(n7901), .A2(n8432), .ZN(n8452) );
  OR2_X1 U5169 ( .A1(n8471), .A2(n8472), .ZN(n8473) );
  AND2_X1 U5170 ( .A1(n7824), .A2(n7822), .ZN(n8492) );
  NAND2_X1 U5171 ( .A1(n8026), .A2(n4732), .ZN(n8482) );
  NAND2_X1 U5172 ( .A1(n7539), .A2(n7788), .ZN(n8026) );
  AND4_X1 U5173 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(n7535)
         );
  NAND2_X1 U5174 ( .A1(n7145), .A2(n4339), .ZN(n7455) );
  NOR2_X1 U5175 ( .A1(n7879), .A2(n4750), .ZN(n4749) );
  OR2_X1 U5176 ( .A1(n5992), .A2(n5991), .ZN(n6010) );
  NAND2_X1 U5177 ( .A1(n7004), .A2(n7867), .ZN(n4776) );
  NAND2_X1 U5178 ( .A1(n6962), .A2(n6961), .ZN(n7040) );
  AND4_X1 U5179 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n7042)
         );
  AND2_X1 U5180 ( .A1(n7846), .A2(n7848), .ZN(n8516) );
  NAND2_X1 U5181 ( .A1(n6782), .A2(n6787), .ZN(n6851) );
  NAND2_X1 U5182 ( .A1(n4460), .A2(n7834), .ZN(n6859) );
  INV_X1 U5183 ( .A(n8506), .ZN(n8498) );
  OR2_X1 U5184 ( .A1(n9881), .A2(n8499), .ZN(n6407) );
  AND2_X1 U5185 ( .A1(n6076), .A2(n6269), .ZN(n8506) );
  NAND2_X1 U5186 ( .A1(n7957), .A2(n7786), .ZN(n8511) );
  NAND2_X1 U5187 ( .A1(n8533), .A2(n9836), .ZN(n4670) );
  NAND2_X1 U5188 ( .A1(n7723), .A2(n7722), .ZN(n8549) );
  NAND2_X1 U5189 ( .A1(n7438), .A2(n7437), .ZN(n8592) );
  INV_X1 U5190 ( .A(n8178), .ZN(n9835) );
  AND2_X1 U5191 ( .A1(n5903), .A2(n5902), .ZN(n9831) );
  NOR2_X1 U5192 ( .A1(n7533), .A2(n6037), .ZN(n9766) );
  AND2_X1 U5193 ( .A1(n7484), .A2(n6036), .ZN(n6037) );
  NAND2_X1 U5194 ( .A1(n4479), .A2(n5744), .ZN(n5745) );
  INV_X1 U5195 ( .A(n5760), .ZN(n5752) );
  INV_X1 U5196 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U5197 ( .A1(n5736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5755) );
  INV_X1 U5198 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U5199 ( .A(n5793), .B(P2_IR_REG_20__SCAN_IN), .ZN(n7956) );
  NOR2_X1 U5200 ( .A1(n5897), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5908) );
  OR2_X1 U5201 ( .A1(n5859), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5897) );
  OAI21_X1 U5202 ( .B1(n5821), .B2(n4631), .A(n4629), .ZN(n4628) );
  NAND2_X1 U5203 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4631) );
  NAND2_X1 U5204 ( .A1(n5838), .A2(n4630), .ZN(n4629) );
  OR2_X1 U5205 ( .A1(n5169), .A2(n6298), .ZN(n5187) );
  XNOR2_X1 U5206 ( .A(n4934), .B(n5049), .ZN(n4957) );
  NAND2_X1 U5207 ( .A1(n4643), .A2(n4935), .ZN(n4641) );
  XNOR2_X1 U5208 ( .A(n5050), .B(n5552), .ZN(n6456) );
  OAI22_X1 U5209 ( .A1(n6619), .A2(n5672), .B1(n6670), .B2(n5096), .ZN(n5050)
         );
  NOR2_X1 U5210 ( .A1(n5701), .A2(n5702), .ZN(n5627) );
  NOR2_X1 U5211 ( .A1(n5588), .A2(n6212), .ZN(n5603) );
  AND2_X1 U5212 ( .A1(n9327), .A2(n8860), .ZN(n9023) );
  AND4_X1 U5213 ( .A1(n5066), .A2(n5065), .A3(n5064), .A4(n5063), .ZN(n6681)
         );
  NAND2_X1 U5214 ( .A1(n9087), .A2(n4380), .ZN(n9550) );
  OR2_X1 U5215 ( .A1(n4508), .A2(n4506), .ZN(n4505) );
  AOI21_X1 U5216 ( .B1(n4508), .B2(n4333), .A(n4381), .ZN(n6293) );
  AND2_X1 U5217 ( .A1(n4506), .A2(n4333), .ZN(n4504) );
  NAND2_X1 U5218 ( .A1(n4496), .A2(n4495), .ZN(n6903) );
  AOI21_X1 U5219 ( .B1(n4503), .B2(n4334), .A(n4391), .ZN(n4495) );
  NAND2_X1 U5220 ( .A1(n4500), .A2(n4498), .ZN(n4502) );
  NOR2_X1 U5221 ( .A1(n9112), .A2(n4393), .ZN(n9116) );
  OR2_X1 U5222 ( .A1(n9116), .A2(n9115), .ZN(n4514) );
  NOR2_X1 U5223 ( .A1(n9485), .A2(n4616), .ZN(n4615) );
  INV_X1 U5224 ( .A(n4617), .ZN(n4616) );
  NAND2_X1 U5225 ( .A1(n4452), .A2(n8835), .ZN(n4483) );
  INV_X1 U5226 ( .A(n9201), .ZN(n4452) );
  AND4_X1 U5227 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n9214)
         );
  OR2_X1 U5228 ( .A1(n9358), .A2(n9246), .ZN(n8077) );
  AND2_X1 U5229 ( .A1(n8973), .A2(n8828), .ZN(n9244) );
  NAND2_X1 U5230 ( .A1(n9272), .A2(n8076), .ZN(n4849) );
  AND2_X1 U5231 ( .A1(n4849), .A2(n4323), .ZN(n9256) );
  NOR2_X1 U5232 ( .A1(n4494), .A2(n8811), .ZN(n4444) );
  NAND2_X1 U5233 ( .A1(n9295), .A2(n4794), .ZN(n4445) );
  OR2_X1 U5234 ( .A1(n7634), .A2(n8921), .ZN(n9295) );
  INV_X1 U5235 ( .A(n4435), .ZN(n4434) );
  OAI21_X1 U5236 ( .B1(n4436), .B2(n8801), .A(n7410), .ZN(n4435) );
  NAND2_X1 U5237 ( .A1(n7386), .A2(n4436), .ZN(n4433) );
  AND2_X1 U5238 ( .A1(n4834), .A2(n4372), .ZN(n4833) );
  NAND2_X1 U5239 ( .A1(n5268), .A2(n5267), .ZN(n7395) );
  OR2_X1 U5240 ( .A1(n7293), .A2(n7323), .ZN(n7415) );
  NOR2_X2 U5241 ( .A1(n7415), .A2(n9400), .ZN(n7414) );
  NAND2_X1 U5242 ( .A1(n9615), .A2(n8949), .ZN(n4493) );
  AND2_X1 U5243 ( .A1(n8945), .A2(n8948), .ZN(n9318) );
  AND3_X1 U5244 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5062) );
  NOR2_X1 U5245 ( .A1(n4608), .A2(n4970), .ZN(n6528) );
  INV_X1 U5246 ( .A(n8874), .ZN(n6496) );
  NAND3_X2 U5247 ( .A1(n4932), .A2(n5580), .A3(n5579), .ZN(n7290) );
  NAND2_X1 U5248 ( .A1(n7118), .A2(n4933), .ZN(n4932) );
  NAND2_X1 U5249 ( .A1(n5618), .A2(n5617), .ZN(n9343) );
  NAND2_X1 U5250 ( .A1(n5512), .A2(n5511), .ZN(n9354) );
  INV_X1 U5251 ( .A(n9677), .ZN(n9705) );
  XNOR2_X1 U5252 ( .A(n5577), .B(n5576), .ZN(n7229) );
  INV_X1 U5253 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5576) );
  AND2_X1 U5254 ( .A1(n4880), .A2(n4904), .ZN(n4650) );
  XNOR2_X1 U5255 ( .A(n5484), .B(n5483), .ZN(n7678) );
  XNOR2_X1 U5256 ( .A(n5416), .B(n5415), .ZN(n7514) );
  AND2_X1 U5257 ( .A1(n5086), .A2(n4866), .ZN(n5214) );
  NAND2_X1 U5258 ( .A1(n4796), .A2(n4797), .ZN(n5233) );
  XNOR2_X1 U5259 ( .A(n4998), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9083) );
  INV_X1 U5260 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4516) );
  NOR2_X1 U5261 ( .A1(n9515), .A2(n4880), .ZN(n4517) );
  XNOR2_X1 U5262 ( .A(n7981), .B(n7982), .ZN(n8132) );
  AND4_X1 U5263 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n6849)
         );
  NAND2_X1 U5264 ( .A1(n7069), .A2(n7068), .ZN(n8602) );
  AND4_X1 U5265 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n7451)
         );
  AND4_X1 U5266 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n6985)
         );
  NAND2_X1 U5267 ( .A1(n4706), .A2(n4703), .ZN(n4708) );
  NAND2_X1 U5268 ( .A1(n8197), .A2(n8198), .ZN(n4605) );
  NAND2_X1 U5269 ( .A1(n4706), .A2(n4702), .ZN(n8197) );
  INV_X1 U5270 ( .A(n4705), .ZN(n4702) );
  INV_X1 U5271 ( .A(n8206), .ZN(n4602) );
  XNOR2_X1 U5272 ( .A(n4712), .B(n8053), .ZN(n8535) );
  NAND2_X1 U5273 ( .A1(n8307), .A2(n8043), .ZN(n4712) );
  OR2_X1 U5274 ( .A1(n8298), .A2(n4672), .ZN(n4671) );
  NOR2_X1 U5275 ( .A1(n4674), .A2(n4673), .ZN(n4672) );
  NAND2_X1 U5276 ( .A1(n8436), .A2(n8034), .ZN(n8420) );
  INV_X1 U5277 ( .A(n8400), .ZN(n8521) );
  AND2_X1 U5278 ( .A1(n4368), .A2(n5759), .ZN(n4784) );
  INV_X1 U5279 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4785) );
  AND4_X1 U5280 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n7225)
         );
  NAND2_X1 U5281 ( .A1(n5543), .A2(n5542), .ZN(n9348) );
  OAI21_X1 U5282 ( .B1(n5703), .B2(n5702), .A(n5701), .ZN(n5705) );
  AND4_X1 U5283 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n7492)
         );
  INV_X1 U5284 ( .A(n9214), .ZN(n9189) );
  INV_X1 U5285 ( .A(n6681), .ZN(n9311) );
  NAND2_X1 U5286 ( .A1(n5030), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U5287 ( .A1(n5026), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U5288 ( .A1(n5030), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4947) );
  NOR2_X1 U5289 ( .A1(n9536), .A2(n9535), .ZN(n9534) );
  AOI21_X1 U5290 ( .B1(n7117), .B2(n6575), .A(n6574), .ZN(n9596) );
  XNOR2_X1 U5291 ( .A(n7353), .B(n7359), .ZN(n7208) );
  AND2_X1 U5292 ( .A1(n9162), .A2(n9161), .ZN(n9336) );
  AOI22_X1 U5293 ( .A1(n9160), .A2(n9631), .B1(n9633), .B2(n9190), .ZN(n9161)
         );
  NAND2_X1 U5294 ( .A1(n9159), .A2(n9313), .ZN(n9162) );
  AND2_X1 U5295 ( .A1(n4489), .A2(n4488), .ZN(n9341) );
  AOI21_X1 U5296 ( .B1(n9203), .B2(n9633), .A(n9177), .ZN(n4488) );
  NAND2_X1 U5297 ( .A1(n4491), .A2(n4490), .ZN(n4489) );
  INV_X1 U5298 ( .A(n9343), .ZN(n9185) );
  NAND2_X1 U5299 ( .A1(n5445), .A2(n5444), .ZN(n9264) );
  AND2_X1 U5300 ( .A1(n9317), .A2(n6679), .ZN(n9607) );
  NAND2_X1 U5301 ( .A1(n9646), .A2(n6482), .ZN(n9623) );
  XNOR2_X1 U5302 ( .A(n6496), .B(n9628), .ZN(n9653) );
  AND2_X1 U5303 ( .A1(n9646), .A2(n6483), .ZN(n9612) );
  NAND2_X1 U5304 ( .A1(n8905), .A2(n4828), .ZN(n4822) );
  OR2_X1 U5305 ( .A1(n9149), .A2(n4825), .ZN(n4824) );
  AND2_X1 U5306 ( .A1(n9330), .A2(n9329), .ZN(n9331) );
  NAND2_X1 U5307 ( .A1(n7828), .A2(n7947), .ZN(n4525) );
  OAI21_X1 U5308 ( .B1(n7845), .B2(n4521), .A(n4518), .ZN(n4528) );
  INV_X1 U5309 ( .A(n4524), .ZN(n4521) );
  AND2_X1 U5310 ( .A1(n4519), .A2(n4529), .ZN(n4518) );
  OAI21_X1 U5311 ( .B1(n7845), .B2(n4523), .A(n4522), .ZN(n4526) );
  OR2_X1 U5312 ( .A1(n7844), .A2(n4527), .ZN(n4523) );
  AOI21_X1 U5313 ( .B1(n4331), .B2(n7846), .A(n7947), .ZN(n4522) );
  OR2_X1 U5314 ( .A1(n7881), .A2(n7882), .ZN(n4549) );
  NAND2_X1 U5315 ( .A1(n4543), .A2(n7885), .ZN(n7888) );
  NAND2_X1 U5316 ( .A1(n4555), .A2(n7939), .ZN(n4554) );
  INV_X1 U5317 ( .A(n7917), .ZN(n4555) );
  NAND2_X1 U5318 ( .A1(n7925), .A2(n4346), .ZN(n4542) );
  AND2_X1 U5319 ( .A1(n7931), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U5320 ( .A1(n4779), .A2(n7939), .ZN(n4541) );
  INV_X1 U5321 ( .A(n7930), .ZN(n4539) );
  INV_X1 U5322 ( .A(n4590), .ZN(n4588) );
  AOI21_X1 U5323 ( .B1(n4590), .B2(n4587), .A(n4586), .ZN(n4585) );
  INV_X1 U5324 ( .A(n5339), .ZN(n4586) );
  INV_X1 U5325 ( .A(n4592), .ZN(n4587) );
  AND2_X1 U5326 ( .A1(n8053), .A2(n7934), .ZN(n4762) );
  NOR2_X1 U5327 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5727) );
  NOR2_X1 U5328 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5726) );
  NOR2_X1 U5329 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5728) );
  NOR2_X1 U5330 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5731) );
  INV_X1 U5331 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5839) );
  INV_X1 U5332 ( .A(n4412), .ZN(n4411) );
  INV_X1 U5333 ( .A(n4414), .ZN(n4409) );
  INV_X1 U5334 ( .A(n5630), .ZN(n4408) );
  AOI21_X1 U5335 ( .B1(n5390), .B2(n4793), .A(n4383), .ZN(n4792) );
  INV_X1 U5336 ( .A(n5367), .ZN(n4793) );
  INV_X1 U5337 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5342) );
  INV_X1 U5338 ( .A(SI_16_), .ZN(n5315) );
  INV_X1 U5339 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5262) );
  AND2_X1 U5340 ( .A1(n7440), .A2(n4390), .ZN(n4688) );
  OR2_X1 U5341 ( .A1(n8140), .A2(n8139), .ZN(n4707) );
  AOI21_X1 U5342 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n7955) );
  INV_X1 U5343 ( .A(n4762), .ZN(n4761) );
  OR2_X1 U5344 ( .A1(n8549), .A2(n8143), .ZN(n7931) );
  OR2_X1 U5345 ( .A1(n8571), .A2(n8038), .ZN(n8384) );
  NOR2_X1 U5346 ( .A1(n8571), .A2(n8576), .ZN(n4681) );
  OAI21_X1 U5347 ( .B1(n8033), .B2(n4726), .A(n8035), .ZN(n4725) );
  NAND2_X1 U5348 ( .A1(n4732), .A2(n7892), .ZN(n4730) );
  OR2_X1 U5349 ( .A1(n6026), .A2(n7247), .ZN(n6066) );
  INV_X1 U5350 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5952) );
  OR2_X1 U5351 ( .A1(n5953), .A2(n5952), .ZN(n5975) );
  NAND2_X1 U5352 ( .A1(n6860), .A2(n9831), .ZN(n4729) );
  AND2_X1 U5353 ( .A1(n9754), .A2(n9743), .ZN(n7843) );
  NAND2_X1 U5354 ( .A1(n7790), .A2(n7829), .ZN(n6742) );
  AND2_X1 U5355 ( .A1(n4763), .A2(n7934), .ZN(n8052) );
  AOI21_X1 U5356 ( .B1(n4768), .B2(n4770), .A(n4767), .ZN(n4766) );
  INV_X1 U5357 ( .A(n4769), .ZN(n4768) );
  AND2_X1 U5358 ( .A1(n5759), .A2(n5750), .ZN(n4751) );
  NAND2_X1 U5359 ( .A1(n5748), .A2(n4751), .ZN(n5779) );
  AND3_X1 U5360 ( .A1(n5741), .A2(n5742), .A3(n5743), .ZN(n4479) );
  AND3_X1 U5361 ( .A1(n5794), .A2(n5740), .A3(n5739), .ZN(n5744) );
  OR3_X1 U5362 ( .A1(n6005), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n6023) );
  INV_X1 U5363 ( .A(n5049), .ZN(n5097) );
  INV_X1 U5364 ( .A(n5628), .ZN(n4646) );
  OR2_X1 U5365 ( .A1(n5628), .A2(n5530), .ZN(n4644) );
  OR2_X1 U5366 ( .A1(n9339), .A2(n8079), .ZN(n8984) );
  AND2_X1 U5367 ( .A1(n8852), .A2(n8740), .ZN(n9029) );
  INV_X1 U5368 ( .A(SI_21_), .ZN(n10054) );
  INV_X1 U5369 ( .A(n6663), .ZN(n4497) );
  INV_X1 U5370 ( .A(n6584), .ZN(n4499) );
  NOR2_X1 U5371 ( .A1(n9327), .A2(n4618), .ZN(n4617) );
  INV_X1 U5372 ( .A(n4619), .ZN(n4618) );
  NOR2_X1 U5373 ( .A1(n9333), .A2(n9339), .ZN(n4619) );
  NAND2_X1 U5374 ( .A1(n4483), .A2(n8983), .ZN(n4791) );
  AND2_X1 U5375 ( .A1(n8984), .A2(n8917), .ZN(n8901) );
  NAND2_X1 U5376 ( .A1(n4813), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5377 ( .A1(n8829), .A2(n9231), .ZN(n4812) );
  NOR2_X1 U5378 ( .A1(n4850), .A2(n4847), .ZN(n4846) );
  INV_X1 U5379 ( .A(n8076), .ZN(n4847) );
  INV_X1 U5380 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5322) );
  AND2_X1 U5381 ( .A1(n7408), .A2(n4366), .ZN(n4835) );
  INV_X1 U5382 ( .A(n7401), .ZN(n4836) );
  NAND2_X1 U5383 ( .A1(n7268), .A2(n7272), .ZN(n7293) );
  INV_X1 U5384 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6298) );
  AND2_X1 U5385 ( .A1(n6877), .A2(n8762), .ZN(n4492) );
  INV_X1 U5386 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5141) );
  OR2_X1 U5387 ( .A1(n5142), .A2(n5141), .ZN(n5169) );
  NOR2_X1 U5388 ( .A1(n6884), .A2(n7096), .ZN(n4607) );
  NAND2_X1 U5389 ( .A1(n4493), .A2(n4492), .ZN(n6879) );
  INV_X1 U5390 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5078) );
  NOR2_X1 U5391 ( .A1(n8873), .A2(n4449), .ZN(n4448) );
  INV_X1 U5392 ( .A(n9003), .ZN(n4449) );
  NAND2_X1 U5393 ( .A1(n6487), .A2(n9637), .ZN(n4608) );
  AND2_X1 U5394 ( .A1(n8949), .A2(n8762), .ZN(n9614) );
  NAND2_X1 U5395 ( .A1(n9310), .A2(n6675), .ZN(n9307) );
  INV_X1 U5396 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5571) );
  AND2_X1 U5397 ( .A1(n5660), .A2(n5637), .ZN(n5658) );
  INV_X1 U5398 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5399 ( .A1(n5443), .A2(n5442), .ZN(n5459) );
  NOR2_X1 U5400 ( .A1(n5313), .A2(n4593), .ZN(n4592) );
  INV_X1 U5401 ( .A(n5285), .ZN(n4593) );
  AOI21_X1 U5402 ( .B1(n4592), .B2(n5281), .A(n4591), .ZN(n4590) );
  INV_X1 U5403 ( .A(n5312), .ZN(n4591) );
  AND2_X1 U5404 ( .A1(n5261), .A2(n5240), .ZN(n5259) );
  AOI21_X1 U5405 ( .B1(n4798), .B2(n4799), .A(n4359), .ZN(n4797) );
  INV_X1 U5406 ( .A(n4860), .ZN(n4798) );
  NAND2_X1 U5407 ( .A1(n5161), .A2(n4600), .ZN(n4796) );
  AND2_X1 U5408 ( .A1(n4799), .A2(n5160), .ZN(n4600) );
  NAND2_X1 U5409 ( .A1(n4422), .A2(n5127), .ZN(n5159) );
  NAND2_X1 U5410 ( .A1(n4421), .A2(n4419), .ZN(n4422) );
  NOR2_X1 U5411 ( .A1(n5128), .A2(n4420), .ZN(n4419) );
  INV_X1 U5412 ( .A(n5114), .ZN(n4420) );
  INV_X1 U5413 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4816) );
  OR2_X1 U5414 ( .A1(n5924), .A2(n8182), .ZN(n8108) );
  NAND2_X1 U5415 ( .A1(n5920), .A2(n5919), .ZN(n6550) );
  CLKBUF_X1 U5416 ( .A(n8106), .Z(n8149) );
  OR2_X1 U5417 ( .A1(n7973), .A2(n7972), .ZN(n4579) );
  NAND2_X1 U5418 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  BUF_X1 U5419 ( .A(n5895), .Z(n7994) );
  NAND2_X1 U5420 ( .A1(n6645), .A2(n4683), .ZN(n6757) );
  AND2_X1 U5421 ( .A1(n5985), .A2(n5965), .ZN(n4683) );
  OAI21_X1 U5422 ( .B1(n4692), .B2(n4695), .A(n4685), .ZN(n7513) );
  OR2_X1 U5423 ( .A1(n7441), .A2(n7442), .ZN(n4685) );
  NAND2_X1 U5424 ( .A1(n4595), .A2(n4594), .ZN(n7439) );
  NAND2_X1 U5425 ( .A1(n4599), .A2(n4598), .ZN(n4595) );
  NOR2_X1 U5426 ( .A1(n7995), .A2(n5856), .ZN(n4597) );
  AND2_X1 U5427 ( .A1(n5911), .A2(n5910), .ZN(n8178) );
  NAND2_X1 U5428 ( .A1(n7062), .A2(n4327), .ZN(n7179) );
  INV_X1 U5429 ( .A(n4355), .ZN(n4684) );
  INV_X1 U5430 ( .A(n8053), .ZN(n8044) );
  NAND2_X1 U5431 ( .A1(n4534), .A2(n7790), .ZN(n4533) );
  NAND2_X1 U5432 ( .A1(n7955), .A2(n7957), .ZN(n4534) );
  AND2_X1 U5433 ( .A1(n7770), .A2(n7769), .ZN(n8007) );
  AND2_X1 U5434 ( .A1(n7757), .A2(n7756), .ZN(n8126) );
  AND2_X1 U5435 ( .A1(n7745), .A2(n7744), .ZN(n8201) );
  OR2_X1 U5436 ( .A1(n8327), .A2(n7763), .ZN(n7745) );
  AND4_X1 U5437 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n8497)
         );
  XNOR2_X1 U5438 ( .A(n6372), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6368) );
  NOR2_X1 U5439 ( .A1(n6336), .A2(n4622), .ZN(n6277) );
  NOR2_X1 U5440 ( .A1(n6349), .A2(n6272), .ZN(n4622) );
  NOR2_X1 U5441 ( .A1(n6466), .A2(n4632), .ZN(n6469) );
  AND2_X1 U5442 ( .A1(n6472), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4632) );
  NOR2_X1 U5443 ( .A1(n6469), .A2(n6468), .ZN(n6600) );
  NOR2_X1 U5444 ( .A1(n6604), .A2(n6603), .ZN(n6765) );
  NOR2_X1 U5445 ( .A1(n7028), .A2(n7029), .ZN(n7165) );
  NOR2_X1 U5446 ( .A1(n7165), .A2(n4633), .ZN(n7169) );
  AND2_X1 U5447 ( .A1(n7166), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U5448 ( .A1(n7169), .A2(n7168), .ZN(n7251) );
  NAND2_X1 U5449 ( .A1(n7253), .A2(n7254), .ZN(n7375) );
  NAND2_X1 U5450 ( .A1(n7375), .A2(n4621), .ZN(n7377) );
  OR2_X1 U5451 ( .A1(n7376), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5452 ( .A1(n7377), .A2(n7378), .ZN(n7576) );
  NAND2_X1 U5453 ( .A1(n7576), .A2(n4620), .ZN(n8223) );
  OR2_X1 U5454 ( .A1(n7577), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5455 ( .A1(n8249), .A2(n4392), .ZN(n8252) );
  AND2_X1 U5456 ( .A1(n7669), .A2(n7668), .ZN(n8299) );
  OR2_X1 U5457 ( .A1(n7751), .A2(n7750), .ZN(n8048) );
  NAND2_X1 U5458 ( .A1(n4777), .A2(n4778), .ZN(n8338) );
  AOI21_X1 U5459 ( .B1(n4780), .B2(n4782), .A(n4779), .ZN(n4778) );
  INV_X1 U5460 ( .A(n4781), .ZN(n4780) );
  NAND2_X1 U5461 ( .A1(n4737), .A2(n8370), .ZN(n4736) );
  OAI21_X1 U5462 ( .B1(n4472), .B2(n4470), .A(n4468), .ZN(n8371) );
  AOI21_X1 U5463 ( .B1(n4474), .B2(n7696), .A(n4465), .ZN(n4468) );
  INV_X1 U5464 ( .A(n7918), .ZN(n4465) );
  AND2_X1 U5465 ( .A1(n7720), .A2(n7719), .ZN(n8372) );
  NAND2_X1 U5466 ( .A1(n8439), .A2(n4324), .ZN(n8365) );
  NAND2_X1 U5467 ( .A1(n8439), .A2(n4679), .ZN(n8393) );
  NAND2_X1 U5468 ( .A1(n4467), .A2(n4466), .ZN(n8387) );
  AND2_X1 U5469 ( .A1(n7694), .A2(n7693), .ZN(n8413) );
  NAND2_X1 U5470 ( .A1(n8439), .A2(n8426), .ZN(n8421) );
  AND2_X1 U5471 ( .A1(n8444), .A2(n8456), .ZN(n8439) );
  NAND2_X1 U5472 ( .A1(n8451), .A2(n8452), .ZN(n8450) );
  OR2_X1 U5473 ( .A1(n8489), .A2(n8592), .ZN(n8464) );
  NAND2_X1 U5474 ( .A1(n6115), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U5475 ( .A1(n7534), .A2(n7889), .ZN(n7672) );
  AND2_X1 U5476 ( .A1(n7456), .A2(n7874), .ZN(n4783) );
  NAND2_X1 U5477 ( .A1(n7457), .A2(n7887), .ZN(n7534) );
  NAND2_X1 U5478 ( .A1(n6992), .A2(n4326), .ZN(n8045) );
  NAND2_X1 U5479 ( .A1(n6992), .A2(n4677), .ZN(n7471) );
  NAND2_X1 U5480 ( .A1(n6992), .A2(n4321), .ZN(n7469) );
  AND2_X1 U5481 ( .A1(n6992), .A2(n9880), .ZN(n7155) );
  NAND2_X1 U5482 ( .A1(n4713), .A2(n4350), .ZN(n6986) );
  NAND2_X1 U5483 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  NOR2_X1 U5484 ( .A1(n7013), .A2(n6980), .ZN(n6992) );
  INV_X1 U5485 ( .A(n4720), .ZN(n6982) );
  NAND2_X1 U5486 ( .A1(n4722), .A2(n4721), .ZN(n6965) );
  INV_X1 U5487 ( .A(n6964), .ZN(n4721) );
  INV_X1 U5488 ( .A(n6999), .ZN(n4722) );
  INV_X1 U5489 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5991) );
  INV_X1 U5490 ( .A(n7858), .ZN(n4464) );
  INV_X1 U5491 ( .A(n6856), .ZN(n4717) );
  NAND2_X1 U5492 ( .A1(n4772), .A2(n4771), .ZN(n6969) );
  AND2_X1 U5493 ( .A1(n4772), .A2(n7851), .ZN(n6865) );
  AND4_X1 U5494 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n7005)
         );
  AND4_X1 U5495 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n8179)
         );
  NAND2_X1 U5496 ( .A1(n5873), .A2(n5872), .ZN(n6854) );
  NOR2_X1 U5497 ( .A1(n6949), .A2(n6854), .ZN(n6950) );
  NAND2_X1 U5498 ( .A1(n6859), .A2(n7826), .ZN(n9755) );
  OR2_X1 U5499 ( .A1(n9817), .A2(n6692), .ZN(n6784) );
  NOR2_X1 U5500 ( .A1(n6784), .A2(n6783), .ZN(n9746) );
  AND4_X1 U5501 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n6696)
         );
  NAND2_X1 U5502 ( .A1(n6420), .A2(n6421), .ZN(n6748) );
  NAND2_X1 U5503 ( .A1(n7749), .A2(n7748), .ZN(n8537) );
  NAND2_X1 U5504 ( .A1(n7735), .A2(n7734), .ZN(n8543) );
  NAND2_X1 U5505 ( .A1(n9820), .A2(n6840), .ZN(n9817) );
  INV_X1 U5506 ( .A(n9881), .ZN(n9837) );
  INV_X1 U5507 ( .A(n9836), .ZN(n9879) );
  INV_X1 U5508 ( .A(n6737), .ZN(n6432) );
  AND2_X1 U5509 ( .A1(n6411), .A2(n6410), .ZN(n6433) );
  AND2_X1 U5510 ( .A1(n5758), .A2(n5757), .ZN(n5759) );
  INV_X1 U5511 ( .A(n6280), .ZN(n6269) );
  INV_X1 U5512 ( .A(n5779), .ZN(n5781) );
  INV_X1 U5513 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5734) );
  INV_X1 U5514 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U5515 ( .A1(n5791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U5516 ( .A1(n6541), .A2(n10083), .ZN(n6652) );
  AND2_X1 U5517 ( .A1(n5987), .A2(n5970), .ZN(n7027) );
  AND2_X1 U5518 ( .A1(n5933), .A2(n5932), .ZN(n6601) );
  CLKBUF_X1 U5519 ( .A(n5806), .Z(n5821) );
  NOR2_X1 U5520 ( .A1(n5640), .A2(n5717), .ZN(n5667) );
  INV_X1 U5521 ( .A(n5425), .ZN(n5423) );
  AOI21_X1 U5522 ( .B1(n4658), .B2(n4656), .A(n4655), .ZN(n4654) );
  INV_X1 U5523 ( .A(n4658), .ZN(n4657) );
  INV_X1 U5524 ( .A(n4662), .ZN(n4656) );
  INV_X1 U5525 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8675) );
  NOR2_X1 U5526 ( .A1(n5599), .A2(n5544), .ZN(n5593) );
  NOR2_X1 U5527 ( .A1(n4341), .A2(n4639), .ZN(n4637) );
  NAND2_X1 U5528 ( .A1(n5337), .A2(n5336), .ZN(n7497) );
  NOR2_X1 U5529 ( .A1(n5323), .A2(n5322), .ZN(n5349) );
  NAND2_X1 U5530 ( .A1(n5506), .A2(n5505), .ZN(n8682) );
  AND2_X1 U5531 ( .A1(n5493), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U5532 ( .A1(n6591), .A2(n6592), .ZN(n4667) );
  NAND2_X1 U5533 ( .A1(n6590), .A2(n4668), .ZN(n4666) );
  OR2_X1 U5534 ( .A1(n6591), .A2(n6592), .ZN(n4668) );
  AND2_X1 U5535 ( .A1(n4944), .A2(n4943), .ZN(n4950) );
  AOI21_X1 U5536 ( .B1(n6509), .B2(n4935), .A(n4951), .ZN(n4952) );
  NAND2_X1 U5537 ( .A1(n6207), .A2(n6209), .ZN(n6208) );
  NAND2_X1 U5538 ( .A1(n8660), .A2(n8661), .ZN(n4661) );
  NOR2_X1 U5539 ( .A1(n8691), .A2(n4659), .ZN(n4658) );
  INV_X1 U5540 ( .A(n4661), .ZN(n4659) );
  NAND2_X1 U5541 ( .A1(n8663), .A2(n4662), .ZN(n4660) );
  NAND2_X1 U5542 ( .A1(n5402), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5425) );
  INV_X1 U5543 ( .A(n5403), .ZN(n5402) );
  NAND2_X1 U5544 ( .A1(n5423), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5446) );
  AND2_X1 U5545 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5469), .ZN(n5493) );
  NOR2_X1 U5546 ( .A1(n5446), .A2(n8675), .ZN(n5469) );
  INV_X1 U5547 ( .A(n5580), .ZN(n6504) );
  NAND2_X1 U5548 ( .A1(n5385), .A2(n5386), .ZN(n8714) );
  NAND2_X1 U5549 ( .A1(n5374), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5403) );
  AND2_X1 U5550 ( .A1(n5349), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5374) );
  INV_X1 U5551 ( .A(n6454), .ZN(n5056) );
  AND2_X1 U5552 ( .A1(n5579), .A2(n8912), .ZN(n9033) );
  AND4_X1 U5553 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n8860)
         );
  NOR2_X1 U5554 ( .A1(n9550), .A2(n9551), .ZN(n9549) );
  NOR2_X1 U5555 ( .A1(n6171), .A2(n6170), .ZN(n6169) );
  NOR2_X1 U5556 ( .A1(n6143), .A2(n9559), .ZN(n6146) );
  INV_X1 U5557 ( .A(n4505), .ZN(n6195) );
  NOR2_X1 U5558 ( .A1(n6286), .A2(n6285), .ZN(n9572) );
  NAND2_X1 U5559 ( .A1(n6657), .A2(n4397), .ZN(n6658) );
  NAND2_X1 U5560 ( .A1(n4399), .A2(n4398), .ZN(n4397) );
  NAND2_X1 U5561 ( .A1(n6658), .A2(n6659), .ZN(n6900) );
  XNOR2_X1 U5562 ( .A(n4512), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U5563 ( .A1(n4514), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U5564 ( .A1(n9126), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5565 ( .A1(n4788), .A2(n4325), .ZN(n9157) );
  AND4_X1 U5566 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n9173)
         );
  NOR2_X1 U5567 ( .A1(n8091), .A2(n9174), .ZN(n4490) );
  AND2_X1 U5568 ( .A1(n4791), .A2(n4790), .ZN(n9174) );
  NAND2_X1 U5569 ( .A1(n9175), .A2(n9176), .ZN(n4491) );
  NAND2_X1 U5570 ( .A1(n4791), .A2(n8914), .ZN(n9175) );
  NAND2_X1 U5571 ( .A1(n4841), .A2(n4840), .ZN(n9180) );
  AOI21_X1 U5572 ( .B1(n4842), .B2(n4320), .A(n4356), .ZN(n4840) );
  NAND2_X1 U5573 ( .A1(n4484), .A2(n4808), .ZN(n9201) );
  NAND2_X1 U5574 ( .A1(n4811), .A2(n4351), .ZN(n4808) );
  NAND2_X1 U5575 ( .A1(n9232), .A2(n4485), .ZN(n4484) );
  AND2_X1 U5576 ( .A1(n4351), .A2(n8829), .ZN(n4485) );
  NAND2_X1 U5577 ( .A1(n9232), .A2(n8829), .ZN(n4809) );
  INV_X1 U5578 ( .A(n4811), .ZN(n4810) );
  NOR2_X1 U5579 ( .A1(n9230), .A2(n8087), .ZN(n9216) );
  NOR2_X1 U5580 ( .A1(n9232), .A2(n9231), .ZN(n9230) );
  OR2_X1 U5581 ( .A1(n9264), .A2(n8703), .ZN(n9240) );
  OAI21_X1 U5582 ( .B1(n9295), .B2(n4442), .A(n4438), .ZN(n9258) );
  AOI21_X1 U5583 ( .B1(n4441), .B2(n4440), .A(n4439), .ZN(n4438) );
  INV_X1 U5584 ( .A(n8872), .ZN(n4439) );
  INV_X1 U5585 ( .A(n4794), .ZN(n4440) );
  NAND2_X1 U5586 ( .A1(n9258), .A2(n9259), .ZN(n9257) );
  NAND2_X1 U5587 ( .A1(n8815), .A2(n8966), .ZN(n9296) );
  NOR2_X1 U5588 ( .A1(n9386), .A2(n4611), .ZN(n4610) );
  INV_X1 U5589 ( .A(n4612), .ZN(n4611) );
  AOI21_X1 U5590 ( .B1(n4434), .B2(n8801), .A(n4432), .ZN(n4431) );
  NAND2_X1 U5591 ( .A1(n7391), .A2(n4614), .ZN(n7626) );
  AND2_X1 U5592 ( .A1(n8747), .A2(n8085), .ZN(n8895) );
  NOR2_X1 U5593 ( .A1(n8775), .A2(n8771), .ZN(n4450) );
  AND2_X1 U5594 ( .A1(n8933), .A2(n8959), .ZN(n8890) );
  AND2_X1 U5595 ( .A1(n5218), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5246) );
  NOR2_X1 U5596 ( .A1(n5187), .A2(n5186), .ZN(n5218) );
  AOI21_X1 U5597 ( .B1(n8887), .B2(n7263), .A(n4328), .ZN(n4839) );
  AND2_X1 U5598 ( .A1(n8776), .A2(n8791), .ZN(n8888) );
  NAND2_X1 U5599 ( .A1(n7260), .A2(n8768), .ZN(n7283) );
  NOR2_X1 U5600 ( .A1(n7220), .A2(n7262), .ZN(n7268) );
  NAND2_X1 U5601 ( .A1(n4429), .A2(n8767), .ZN(n7259) );
  OAI21_X1 U5602 ( .B1(n4493), .B2(n4428), .A(n4426), .ZN(n4429) );
  INV_X1 U5603 ( .A(n4427), .ZN(n4426) );
  OAI21_X1 U5604 ( .B1(n4492), .B2(n4428), .A(n8927), .ZN(n4427) );
  NAND2_X1 U5605 ( .A1(n4607), .A2(n4606), .ZN(n7220) );
  INV_X1 U5606 ( .A(n4607), .ZN(n7218) );
  NAND2_X1 U5607 ( .A1(n6313), .A2(n6528), .ZN(n6631) );
  OAI211_X1 U5608 ( .C1(n5290), .C2(n6089), .A(n5012), .B(n5011), .ZN(n6559)
         );
  NAND2_X1 U5609 ( .A1(n6622), .A2(n4448), .ZN(n9308) );
  INV_X1 U5610 ( .A(n6615), .ZN(n8876) );
  AND4_X1 U5611 ( .A1(n5017), .A2(n5016), .A3(n5015), .A4(n5014), .ZN(n6676)
         );
  INV_X1 U5612 ( .A(n4608), .ZN(n9639) );
  NAND2_X1 U5613 ( .A1(n8870), .A2(n4826), .ZN(n4825) );
  INV_X1 U5614 ( .A(n4828), .ZN(n4826) );
  AND2_X1 U5615 ( .A1(n9333), .A2(n9052), .ZN(n4828) );
  NAND2_X1 U5616 ( .A1(n5492), .A2(n5491), .ZN(n9358) );
  NAND2_X1 U5617 ( .A1(n5401), .A2(n5400), .ZN(n9381) );
  INV_X1 U5618 ( .A(n7395), .ZN(n9493) );
  INV_X1 U5619 ( .A(n9706), .ZN(n9667) );
  NAND2_X1 U5620 ( .A1(n8733), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4969) );
  INV_X1 U5621 ( .A(n7111), .ZN(n6480) );
  AND3_X1 U5622 ( .A1(n4873), .A2(n4370), .A3(n4872), .ZN(n4878) );
  XNOR2_X1 U5623 ( .A(n7774), .B(n7773), .ZN(n8737) );
  XNOR2_X1 U5624 ( .A(n7758), .B(n7760), .ZN(n8640) );
  XNOR2_X1 U5625 ( .A(n7653), .B(n7652), .ZN(n8643) );
  NAND2_X1 U5626 ( .A1(n4406), .A2(n4412), .ZN(n5631) );
  NAND2_X1 U5627 ( .A1(n5537), .A2(n4414), .ZN(n4406) );
  NAND2_X1 U5628 ( .A1(n4652), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U5629 ( .A1(n4905), .A2(n4889), .ZN(n4892) );
  XNOR2_X1 U5630 ( .A(n4924), .B(n5570), .ZN(n4925) );
  NAND2_X1 U5631 ( .A1(n4923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U5632 ( .A1(n4930), .A2(n4929), .ZN(n5575) );
  OAI21_X1 U5633 ( .B1(n5369), .B2(n5368), .A(n5367), .ZN(n5391) );
  INV_X1 U5634 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U5635 ( .A1(n4589), .A2(n5285), .ZN(n5314) );
  INV_X1 U5636 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U5637 ( .A1(n4801), .A2(n5180), .ZN(n5209) );
  NAND2_X1 U5638 ( .A1(n5179), .A2(n4860), .ZN(n4801) );
  INV_X1 U5639 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U5640 ( .A1(n4421), .A2(n5114), .ZN(n5129) );
  AND2_X1 U5641 ( .A1(n4635), .A2(n4995), .ZN(n5041) );
  NOR2_X1 U5642 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4635) );
  AND2_X1 U5643 ( .A1(n5926), .A2(n5886), .ZN(n8111) );
  OR2_X1 U5644 ( .A1(n6553), .A2(n5885), .ZN(n5886) );
  INV_X1 U5645 ( .A(n4708), .ZN(n8195) );
  NAND2_X1 U5646 ( .A1(n4698), .A2(n4696), .ZN(n8124) );
  AOI21_X1 U5647 ( .B1(n4699), .B2(n4704), .A(n4697), .ZN(n4696) );
  INV_X1 U5648 ( .A(n8120), .ZN(n4697) );
  NAND2_X1 U5649 ( .A1(n6645), .A2(n5965), .ZN(n6759) );
  AND4_X1 U5650 ( .A1(n5770), .A2(n5768), .A3(n5771), .A4(n5769), .ZN(n8064)
         );
  AND2_X1 U5651 ( .A1(n8065), .A2(n5798), .ZN(n7968) );
  NAND2_X1 U5652 ( .A1(n4690), .A2(n4686), .ZN(n4577) );
  NAND2_X1 U5653 ( .A1(n4692), .A2(n4686), .ZN(n4578) );
  AND4_X1 U5654 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n7006)
         );
  NOR2_X1 U5655 ( .A1(n6075), .A2(n6074), .ZN(n8152) );
  NAND2_X1 U5656 ( .A1(n4562), .A2(n4559), .ZN(n8158) );
  AND2_X1 U5657 ( .A1(n4561), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U5658 ( .A1(n4566), .A2(n4569), .ZN(n4562) );
  OR2_X1 U5660 ( .A1(n5850), .A2(n5799), .ZN(n5804) );
  OR2_X1 U5661 ( .A1(n6846), .A2(n5895), .ZN(n8065) );
  OAI21_X1 U5662 ( .B1(n4692), .B2(n4690), .A(n4686), .ZN(n7589) );
  NAND2_X1 U5663 ( .A1(n7557), .A2(n7556), .ZN(n8582) );
  INV_X1 U5664 ( .A(n8205), .ZN(n8162) );
  OR2_X1 U5665 ( .A1(n8196), .A2(n7994), .ZN(n8189) );
  OAI21_X1 U5666 ( .B1(n5869), .B2(n6094), .A(n4476), .ZN(n8170) );
  INV_X1 U5667 ( .A(n4477), .ZN(n4476) );
  OAI22_X1 U5668 ( .A1(n5856), .A2(n6093), .B1(n4478), .B2(n6263), .ZN(n4477)
         );
  NAND2_X1 U5669 ( .A1(n5828), .A2(n5827), .ZN(n8173) );
  AND2_X1 U5670 ( .A1(n8152), .A2(n8508), .ZN(n8168) );
  AND4_X1 U5671 ( .A1(n7087), .A2(n7086), .A3(n7085), .A4(n7084), .ZN(n7673)
         );
  INV_X1 U5672 ( .A(n8168), .ZN(n8202) );
  AND2_X1 U5673 ( .A1(n8067), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8205) );
  NAND2_X1 U5674 ( .A1(n4531), .A2(n4535), .ZN(n4425) );
  NAND2_X1 U5675 ( .A1(n4533), .A2(n4532), .ZN(n4531) );
  INV_X1 U5676 ( .A(n7958), .ZN(n4535) );
  NAND2_X1 U5677 ( .A1(n7954), .A2(n7953), .ZN(n4532) );
  OR2_X1 U5678 ( .A1(n7785), .A2(n4394), .ZN(n4424) );
  AOI21_X1 U5679 ( .B1(n7783), .B2(n7818), .A(n7949), .ZN(n7784) );
  INV_X1 U5680 ( .A(n8014), .ZN(n7960) );
  INV_X1 U5681 ( .A(n8126), .ZN(n8319) );
  INV_X1 U5682 ( .A(n8143), .ZN(n8320) );
  INV_X1 U5683 ( .A(n8372), .ZN(n8339) );
  NAND2_X1 U5684 ( .A1(n5894), .A2(n4551), .ZN(n8507) );
  NOR2_X1 U5685 ( .A1(n4552), .A2(n4343), .ZN(n4551) );
  NAND2_X1 U5686 ( .A1(n5892), .A2(n5893), .ZN(n4552) );
  INV_X2 U5687 ( .A(P2_U3966), .ZN(n8222) );
  INV_X1 U5688 ( .A(n8064), .ZN(n6418) );
  INV_X1 U5689 ( .A(n4626), .ZN(n6324) );
  INV_X1 U5690 ( .A(n4624), .ZN(n6338) );
  INV_X1 U5691 ( .A(n8291), .ZN(n9738) );
  NAND2_X1 U5692 ( .A1(n9733), .A2(n6269), .ZN(n8282) );
  NAND2_X1 U5693 ( .A1(n8274), .A2(n8275), .ZN(n8278) );
  AND2_X1 U5694 ( .A1(n6281), .A2(n6280), .ZN(n8285) );
  INV_X1 U5695 ( .A(n8299), .ZN(n8528) );
  NAND2_X1 U5696 ( .A1(n8374), .A2(n7922), .ZN(n8356) );
  NAND2_X1 U5697 ( .A1(n7711), .A2(n7710), .ZN(n8554) );
  NAND2_X1 U5698 ( .A1(n4734), .A2(n4737), .ZN(n8364) );
  NAND2_X1 U5699 ( .A1(n8404), .A2(n4739), .ZN(n4734) );
  NAND2_X1 U5700 ( .A1(n4741), .A2(n4739), .ZN(n8382) );
  NAND2_X1 U5701 ( .A1(n4741), .A2(n4744), .ZN(n8380) );
  NAND2_X1 U5702 ( .A1(n4752), .A2(n4756), .ZN(n8427) );
  NAND2_X1 U5703 ( .A1(n8451), .A2(n4757), .ZN(n4752) );
  NAND2_X1 U5704 ( .A1(n4727), .A2(n8033), .ZN(n8436) );
  NAND2_X1 U5705 ( .A1(n7517), .A2(n7516), .ZN(n8588) );
  NAND2_X1 U5706 ( .A1(n4599), .A2(n7305), .ZN(n8599) );
  NAND2_X1 U5707 ( .A1(n8026), .A2(n8025), .ZN(n8484) );
  NAND2_X1 U5708 ( .A1(n7455), .A2(n7874), .ZN(n7474) );
  AND2_X1 U5709 ( .A1(n7145), .A2(n7876), .ZN(n7146) );
  NAND2_X1 U5710 ( .A1(n6862), .A2(n7848), .ZN(n6953) );
  INV_X1 U5711 ( .A(n6852), .ZN(n8517) );
  INV_X1 U5712 ( .A(n8485), .ZN(n9751) );
  INV_X1 U5713 ( .A(n8499), .ZN(n9753) );
  NAND2_X1 U5714 ( .A1(n6851), .A2(n6850), .ZN(n9745) );
  OR2_X1 U5715 ( .A1(n6745), .A2(n7985), .ZN(n8400) );
  OR2_X1 U5716 ( .A1(n9765), .A2(n6407), .ZN(n8485) );
  OR2_X1 U5717 ( .A1(n6263), .A2(n6391), .ZN(n5809) );
  AND2_X1 U5718 ( .A1(n7775), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4709) );
  INV_X1 U5719 ( .A(n8504), .ZN(n8518) );
  INV_X1 U5720 ( .A(n8469), .ZN(n8514) );
  AND2_X2 U5721 ( .A1(n6433), .A2(n6737), .ZN(n9906) );
  NAND2_X1 U5722 ( .A1(n4322), .A2(n4481), .ZN(n8619) );
  NOR2_X1 U5723 ( .A1(n4671), .A2(n9881), .ZN(n4482) );
  OAI21_X1 U5724 ( .B1(n8535), .B2(n9871), .A(n4670), .ZN(n4669) );
  NAND2_X1 U5725 ( .A1(n4786), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5762) );
  MUX2_X1 U5726 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5763), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5764) );
  NAND2_X1 U5727 ( .A1(n5784), .A2(n5785), .ZN(n8056) );
  NOR2_X1 U5728 ( .A1(n5781), .A2(n5780), .ZN(n5785) );
  OR2_X1 U5729 ( .A1(n5783), .A2(n5758), .ZN(n5784) );
  NOR2_X1 U5730 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5780) );
  NAND2_X1 U5731 ( .A1(n5747), .A2(n5782), .ZN(n7533) );
  INV_X1 U5732 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7482) );
  INV_X1 U5733 ( .A(n5748), .ZN(n5749) );
  XNOR2_X1 U5734 ( .A(n5738), .B(n5739), .ZN(n7321) );
  NAND2_X1 U5735 ( .A1(n5737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5738) );
  INV_X1 U5736 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8017) );
  XNOR2_X1 U5737 ( .A(n5787), .B(n5786), .ZN(n8014) );
  XNOR2_X1 U5738 ( .A(n5790), .B(n5789), .ZN(n7953) );
  INV_X1 U5739 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U5740 ( .A1(n5788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5790) );
  INV_X1 U5741 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6898) );
  INV_X1 U5742 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9961) );
  INV_X1 U5743 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6573) );
  INV_X1 U5744 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6451) );
  INV_X1 U5745 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6323) );
  INV_X1 U5746 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6309) );
  INV_X1 U5747 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6231) );
  INV_X1 U5748 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6187) );
  INV_X1 U5749 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6131) );
  AND2_X1 U5750 ( .A1(n5901), .A2(n5900), .ZN(n6355) );
  AND2_X1 U5751 ( .A1(n7775), .A2(P2_U3152), .ZN(n8644) );
  NOR2_X1 U5752 ( .A1(n5723), .A2(n5722), .ZN(n6132) );
  INV_X1 U5753 ( .A(n6438), .ZN(n4647) );
  CLKBUF_X1 U5754 ( .A(n8659), .Z(n8663) );
  NAND2_X1 U5755 ( .A1(n5714), .A2(n5657), .ZN(n5680) );
  OR2_X1 U5756 ( .A1(n5067), .A2(n4918), .ZN(n4920) );
  AND4_X1 U5757 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n7261)
         );
  NAND2_X1 U5758 ( .A1(n4666), .A2(n4667), .ZN(n6728) );
  NAND2_X1 U5759 ( .A1(n4660), .A2(n4661), .ZN(n8690) );
  NAND2_X1 U5760 ( .A1(n5422), .A2(n5421), .ZN(n9375) );
  NAND2_X1 U5761 ( .A1(n5468), .A2(n5467), .ZN(n9364) );
  INV_X1 U5762 ( .A(n8723), .ZN(n8664) );
  OR2_X1 U5763 ( .A1(n5589), .A2(n6210), .ZN(n8726) );
  AND4_X1 U5764 ( .A1(n5084), .A2(n5083), .A3(n5082), .A4(n5081), .ZN(n9617)
         );
  NAND2_X1 U5765 ( .A1(n5603), .A2(n5592), .ZN(n8706) );
  INV_X1 U5766 ( .A(n4639), .ZN(n4636) );
  INV_X1 U5767 ( .A(n8730), .ZN(n8709) );
  INV_X1 U5768 ( .A(n9203), .ZN(n10115) );
  NAND2_X1 U5769 ( .A1(n5033), .A2(n5032), .ZN(n9064) );
  XNOR2_X1 U5770 ( .A(n9072), .B(n4515), .ZN(n9071) );
  OAI21_X1 U5771 ( .B1(n9534), .B2(n9084), .A(n6150), .ZN(n9087) );
  AND2_X1 U5772 ( .A1(n4505), .A2(n4333), .ZN(n6199) );
  OR2_X1 U5773 ( .A1(n6576), .A2(n9592), .ZN(n9594) );
  NAND2_X1 U5774 ( .A1(n4500), .A2(n4503), .ZN(n9599) );
  AND2_X1 U5775 ( .A1(n4502), .A2(n4501), .ZN(n6664) );
  XNOR2_X1 U5776 ( .A(n7358), .B(n7359), .ZN(n7211) );
  NOR2_X1 U5777 ( .A1(n7208), .A2(n7207), .ZN(n7354) );
  NAND2_X1 U5778 ( .A1(n4511), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5779 ( .A1(n7355), .A2(n4511), .ZN(n4509) );
  INV_X1 U5780 ( .A(n7357), .ZN(n4511) );
  AOI21_X1 U5781 ( .B1(n9100), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9099), .ZN(
        n9102) );
  INV_X1 U5782 ( .A(n4514), .ZN(n9124) );
  INV_X1 U5783 ( .A(n9573), .ZN(n9593) );
  AND2_X1 U5784 ( .A1(n9585), .A2(n5590), .ZN(n9578) );
  INV_X1 U5785 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9135) );
  INV_X1 U5786 ( .A(n8857), .ZN(n9465) );
  XNOR2_X1 U5787 ( .A(n4451), .B(n8904), .ZN(n9191) );
  NAND2_X1 U5788 ( .A1(n4483), .A2(n9186), .ZN(n4451) );
  AOI21_X1 U5789 ( .B1(n8078), .B2(n4844), .A(n4320), .ZN(n9195) );
  NOR2_X1 U5790 ( .A1(n9256), .A2(n4850), .ZN(n9238) );
  NAND2_X1 U5791 ( .A1(n4445), .A2(n4444), .ZN(n9277) );
  NAND2_X1 U5792 ( .A1(n4433), .A2(n8924), .ZN(n7387) );
  OAI21_X1 U5793 ( .B1(n7386), .B2(n8801), .A(n4434), .ZN(n7628) );
  NAND2_X1 U5794 ( .A1(n5321), .A2(n5320), .ZN(n7623) );
  NAND2_X1 U5795 ( .A1(n7386), .A2(n8934), .ZN(n7491) );
  NAND2_X1 U5796 ( .A1(n4837), .A2(n7408), .ZN(n7486) );
  NAND2_X1 U5797 ( .A1(n7402), .A2(n7401), .ZN(n4837) );
  NAND2_X1 U5798 ( .A1(n5217), .A2(n5216), .ZN(n7323) );
  NAND2_X1 U5799 ( .A1(n7264), .A2(n7263), .ZN(n7276) );
  NAND2_X1 U5800 ( .A1(n4493), .A2(n8762), .ZN(n6876) );
  INV_X1 U5801 ( .A(n9318), .ZN(n4830) );
  XNOR2_X1 U5802 ( .A(n9629), .B(n6496), .ZN(n9636) );
  INV_X1 U5803 ( .A(n9641), .ZN(n9314) );
  INV_X1 U5804 ( .A(n9623), .ZN(n9316) );
  AOI211_X1 U5805 ( .C1(n9677), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9503)
         );
  NAND2_X1 U5806 ( .A1(n4807), .A2(n9710), .ZN(n4806) );
  INV_X1 U5807 ( .A(n9332), .ZN(n4807) );
  OR2_X1 U5808 ( .A1(n9368), .A2(n9696), .ZN(n9374) );
  OAI22_X1 U5809 ( .A1(n6241), .A2(P1_D_REG_0__SCAN_IN), .B1(n5554), .B2(n5557), .ZN(n7112) );
  NAND2_X1 U5810 ( .A1(n5723), .A2(n5578), .ZN(n6212) );
  INV_X1 U5811 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7480) );
  OAI21_X1 U5812 ( .B1(n4889), .B2(n4905), .A(n4892), .ZN(n7479) );
  INV_X1 U5813 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10071) );
  INV_X1 U5814 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7119) );
  INV_X1 U5815 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6935) );
  INV_X1 U5816 ( .A(n9032), .ZN(n8912) );
  AND2_X1 U5817 ( .A1(n5346), .A2(n5370), .ZN(n9113) );
  INV_X1 U5818 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6453) );
  AND2_X1 U5819 ( .A1(n5266), .A2(n5291), .ZN(n7210) );
  INV_X1 U5820 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6233) );
  INV_X1 U5821 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6185) );
  INV_X1 U5822 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6129) );
  NOR2_X1 U5823 ( .A1(n9458), .A2(n10127), .ZN(n9934) );
  AOI21_X1 U5824 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9932), .ZN(n9931) );
  NOR2_X1 U5825 ( .A1(n9931), .A2(n9930), .ZN(n9929) );
  AOI21_X1 U5826 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9929), .ZN(n9928) );
  OAI21_X1 U5827 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9926), .ZN(n9924) );
  INV_X1 U5828 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4912) );
  NAND2_X1 U5829 ( .A1(n4604), .A2(n4601), .ZN(P2_U3242) );
  NOR2_X1 U5830 ( .A1(n4603), .A2(n4602), .ZN(n4601) );
  NOR2_X1 U5831 ( .A1(n8336), .A2(n8207), .ZN(n4603) );
  AOI211_X1 U5832 ( .C1(n8534), .C2(n8521), .A(n8061), .B(n8060), .ZN(n8062)
         );
  INV_X1 U5833 ( .A(n4671), .ZN(n8534) );
  NAND2_X1 U5834 ( .A1(n4711), .A2(n4710), .ZN(P2_U3517) );
  NAND2_X1 U5835 ( .A1(n9887), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5836 ( .A1(n8619), .A2(n9888), .ZN(n4711) );
  NAND2_X1 U5837 ( .A1(n6162), .A2(n4939), .ZN(n5725) );
  OAI21_X1 U5838 ( .B1(n9185), .B2(n8730), .A(n5708), .ZN(n5709) );
  AOI211_X1 U5839 ( .C1(n9328), .C2(n9612), .A(n8104), .B(n8103), .ZN(n8105)
         );
  NOR2_X1 U5840 ( .A1(n9336), .A2(n9648), .ZN(n9163) );
  INV_X1 U5841 ( .A(n4486), .ZN(n9179) );
  OAI21_X1 U5842 ( .B1(n9341), .B2(n9648), .A(n4487), .ZN(n4486) );
  AOI21_X1 U5843 ( .B1(n9338), .B2(n9322), .A(n9178), .ZN(n4487) );
  NAND2_X1 U5844 ( .A1(n9726), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4827) );
  OR2_X1 U5845 ( .A1(n9696), .A2(n9726), .ZN(n4821) );
  NAND2_X1 U5846 ( .A1(n4804), .A2(n4803), .ZN(P1_U3520) );
  NAND2_X1 U5847 ( .A1(n9712), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4803) );
  NAND2_X1 U5848 ( .A1(n4805), .A2(n9714), .ZN(n4804) );
  NAND2_X1 U5849 ( .A1(n9331), .A2(n4806), .ZN(n4805) );
  AND2_X1 U5850 ( .A1(n4582), .A2(n4403), .ZN(n4317) );
  OR2_X1 U5851 ( .A1(n9239), .A2(n8676), .ZN(n4318) );
  INV_X1 U5852 ( .A(n7846), .ZN(n4527) );
  AND2_X1 U5853 ( .A1(n7787), .A2(n7771), .ZN(n4319) );
  NOR2_X1 U5854 ( .A1(n9354), .A2(n9202), .ZN(n4320) );
  OR2_X1 U5855 ( .A1(n9358), .A2(n8705), .ZN(n8829) );
  AND2_X1 U5856 ( .A1(n4677), .A2(n4676), .ZN(n4321) );
  NAND2_X1 U5857 ( .A1(n4360), .A2(n7910), .ZN(n4756) );
  NAND2_X1 U5858 ( .A1(n6619), .A2(n9676), .ZN(n8945) );
  AND2_X1 U5859 ( .A1(n8059), .A2(n8058), .ZN(n4322) );
  AND2_X1 U5860 ( .A1(n9254), .A2(n4376), .ZN(n4323) );
  NAND2_X1 U5861 ( .A1(n8310), .A2(n8047), .ZN(n8311) );
  INV_X1 U5862 ( .A(n8311), .ZN(n4674) );
  AND2_X1 U5863 ( .A1(n4679), .A2(n4678), .ZN(n4324) );
  AND2_X1 U5864 ( .A1(n4789), .A2(n9158), .ZN(n4325) );
  AND2_X1 U5865 ( .A1(n4321), .A2(n4675), .ZN(n4326) );
  AND2_X1 U5866 ( .A1(n4684), .A2(n7061), .ZN(n4327) );
  AND2_X1 U5867 ( .A1(n7426), .A2(n9059), .ZN(n4328) );
  AND2_X1 U5868 ( .A1(n4318), .A2(n4846), .ZN(n4329) );
  NOR2_X1 U5869 ( .A1(n8563), .A2(n8413), .ZN(n4330) );
  INV_X1 U5870 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10083) );
  INV_X1 U5871 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4867) );
  AND2_X1 U5872 ( .A1(n7843), .A2(n7842), .ZN(n4331) );
  OAI21_X1 U5873 ( .B1(n8451), .B2(n4755), .A(n4753), .ZN(n8407) );
  NOR2_X1 U5874 ( .A1(n5368), .A2(n5389), .ZN(n4332) );
  OR2_X1 U5875 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6194), .ZN(n4333) );
  INV_X1 U5876 ( .A(n8955), .ZN(n4428) );
  OR2_X1 U5877 ( .A1(n6582), .A2(n9591), .ZN(n4500) );
  AND2_X1 U5878 ( .A1(n4389), .A2(n9591), .ZN(n4334) );
  INV_X1 U5879 ( .A(n4474), .ZN(n4473) );
  OR2_X1 U5880 ( .A1(n9228), .A2(n8705), .ZN(n4335) );
  INV_X1 U5881 ( .A(n5025), .ZN(n8097) );
  INV_X1 U5882 ( .A(n7588), .ZN(n4573) );
  INV_X1 U5883 ( .A(n7441), .ZN(n4689) );
  OR2_X1 U5884 ( .A1(n6947), .A2(n7847), .ZN(n4336) );
  NAND2_X1 U5885 ( .A1(n7881), .A2(n8213), .ZN(n4337) );
  AND2_X1 U5886 ( .A1(n8439), .A2(n4681), .ZN(n4338) );
  INV_X1 U5887 ( .A(n4643), .ZN(n6487) );
  NAND2_X1 U5888 ( .A1(n4642), .A2(n4920), .ZN(n4643) );
  AND2_X1 U5889 ( .A1(n7879), .A2(n7876), .ZN(n4339) );
  XNOR2_X1 U5890 ( .A(n5762), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5767) );
  OR2_X1 U5891 ( .A1(n9395), .A2(n9055), .ZN(n4340) );
  INV_X1 U5892 ( .A(n9064), .ZN(n6619) );
  NAND2_X1 U5893 ( .A1(n8078), .A2(n4335), .ZN(n9208) );
  AND2_X1 U5894 ( .A1(n8384), .A2(n7917), .ZN(n8408) );
  INV_X1 U5895 ( .A(n8408), .ZN(n4746) );
  INV_X1 U5896 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4653) );
  AND2_X1 U5897 ( .A1(n7344), .A2(n5308), .ZN(n4341) );
  OR2_X1 U5898 ( .A1(n6412), .A2(n7965), .ZN(n6419) );
  AND2_X1 U5899 ( .A1(n4567), .A2(n4565), .ZN(n4342) );
  NOR2_X1 U5900 ( .A1(n9176), .A2(n8915), .ZN(n4790) );
  NAND2_X1 U5901 ( .A1(n9381), .A2(n8692), .ZN(n8966) );
  OR2_X1 U5902 ( .A1(n8537), .A2(n8126), .ZN(n7934) );
  NAND2_X1 U5903 ( .A1(n6025), .A2(n6024), .ZN(n7881) );
  NAND2_X1 U5904 ( .A1(n5373), .A2(n5372), .ZN(n9386) );
  NAND2_X1 U5905 ( .A1(n7592), .A2(n7591), .ZN(n8576) );
  NAND2_X1 U5906 ( .A1(n7685), .A2(n7684), .ZN(n8397) );
  NOR2_X1 U5907 ( .A1(n7742), .A2(n5890), .ZN(n4343) );
  AND2_X1 U5908 ( .A1(n4405), .A2(n4332), .ZN(n4344) );
  OR2_X1 U5909 ( .A1(n9364), .A2(n9260), .ZN(n4345) );
  AND2_X1 U5910 ( .A1(n7926), .A2(n7924), .ZN(n4346) );
  INV_X1 U5911 ( .A(n9339), .ZN(n9172) );
  NAND2_X1 U5912 ( .A1(n5639), .A2(n5638), .ZN(n9339) );
  AND2_X1 U5913 ( .A1(n4660), .A2(n4658), .ZN(n4347) );
  AND2_X1 U5914 ( .A1(n4317), .A2(n4332), .ZN(n4348) );
  OR2_X1 U5915 ( .A1(n9348), .A2(n9214), .ZN(n9186) );
  AND2_X1 U5916 ( .A1(n8987), .A2(n8918), .ZN(n9158) );
  AND2_X1 U5917 ( .A1(n4810), .A2(n4809), .ZN(n4349) );
  AND2_X1 U5918 ( .A1(n4714), .A2(n4718), .ZN(n4350) );
  NAND2_X1 U5919 ( .A1(n8919), .A2(n8978), .ZN(n4351) );
  INV_X1 U5920 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5761) );
  OR2_X1 U5921 ( .A1(n8554), .A2(n8372), .ZN(n7927) );
  INV_X1 U5922 ( .A(n7927), .ZN(n4779) );
  AND2_X1 U5923 ( .A1(n4788), .A2(n4789), .ZN(n4352) );
  AND2_X1 U5924 ( .A1(n9354), .A2(n9202), .ZN(n4353) );
  AND2_X1 U5925 ( .A1(n4735), .A2(n4743), .ZN(n4354) );
  XOR2_X1 U5926 ( .A(n8607), .B(n7995), .Z(n4355) );
  NOR2_X1 U5927 ( .A1(n8989), .A2(n9023), .ZN(n8870) );
  NOR2_X1 U5928 ( .A1(n9348), .A2(n9189), .ZN(n4356) );
  INV_X1 U5929 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5740) );
  AND2_X1 U5930 ( .A1(n8890), .A2(n8795), .ZN(n4357) );
  NAND2_X1 U5931 ( .A1(n4569), .A2(n4568), .ZN(n4358) );
  OAI21_X1 U5932 ( .B1(n4323), .B2(n4850), .A(n4345), .ZN(n4848) );
  INV_X1 U5933 ( .A(n8419), .ZN(n7677) );
  AND2_X1 U5934 ( .A1(n5207), .A2(SI_11_), .ZN(n4359) );
  INV_X1 U5935 ( .A(n4442), .ZN(n4441) );
  NAND2_X1 U5936 ( .A1(n4444), .A2(n4443), .ZN(n4442) );
  OR2_X1 U5937 ( .A1(n8033), .A2(n7907), .ZN(n4360) );
  OAI21_X1 U5938 ( .B1(n8299), .B2(n7771), .A(n7941), .ZN(n4764) );
  NAND2_X1 U5939 ( .A1(n9307), .A2(n8948), .ZN(n4361) );
  NAND2_X1 U5940 ( .A1(n4473), .A2(n4471), .ZN(n8383) );
  AND2_X1 U5941 ( .A1(n7886), .A2(n4337), .ZN(n4362) );
  AND2_X1 U5942 ( .A1(n8926), .A2(n8768), .ZN(n8887) );
  AOI21_X1 U5943 ( .B1(n4756), .B2(n4754), .A(n8419), .ZN(n4753) );
  AND2_X1 U5944 ( .A1(n6850), .A2(n4729), .ZN(n4363) );
  AND2_X1 U5945 ( .A1(n4904), .A2(n4653), .ZN(n4364) );
  OR2_X1 U5946 ( .A1(n6860), .A2(n9831), .ZN(n4365) );
  NOR2_X1 U5947 ( .A1(n5208), .A2(n4800), .ZN(n4799) );
  AND2_X1 U5948 ( .A1(n4340), .A2(n7279), .ZN(n4366) );
  AND2_X1 U5949 ( .A1(n5627), .A2(n4644), .ZN(n4367) );
  NOR2_X1 U5950 ( .A1(n6984), .A2(n4716), .ZN(n4715) );
  AND2_X1 U5951 ( .A1(n5761), .A2(n4785), .ZN(n4368) );
  AND2_X1 U5952 ( .A1(n4751), .A2(n5761), .ZN(n4369) );
  AND2_X1 U5953 ( .A1(n4852), .A2(n4851), .ZN(n4370) );
  AND2_X1 U5954 ( .A1(n4730), .A2(n8028), .ZN(n4371) );
  INV_X1 U5955 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4630) );
  OR2_X1 U5956 ( .A1(n7490), .A2(n7409), .ZN(n4372) );
  INV_X1 U5957 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5750) );
  AND2_X1 U5958 ( .A1(n4874), .A2(n4653), .ZN(n4852) );
  INV_X1 U5959 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4851) );
  OR2_X1 U5960 ( .A1(n9137), .A2(n9136), .ZN(P1_U3260) );
  AOI21_X1 U5961 ( .B1(n8732), .B2(n5928), .A(n4853), .ZN(n8292) );
  INV_X1 U5962 ( .A(n7305), .ZN(n4596) );
  AND2_X1 U5963 ( .A1(n7391), .A2(n4612), .ZN(n4374) );
  NAND2_X1 U5964 ( .A1(n7280), .A2(n7279), .ZN(n7402) );
  AND2_X1 U5965 ( .A1(n7391), .A2(n7490), .ZN(n4375) );
  OR2_X1 U5966 ( .A1(n9375), .A2(n9301), .ZN(n4376) );
  NOR2_X1 U5967 ( .A1(n7513), .A2(n4854), .ZN(n7554) );
  AND2_X1 U5968 ( .A1(n4638), .A2(n4636), .ZN(n7342) );
  AND3_X1 U5969 ( .A1(n5693), .A2(n8683), .A3(n5692), .ZN(n4377) );
  OR2_X1 U5970 ( .A1(n9172), .A2(n8730), .ZN(n4378) );
  INV_X1 U5971 ( .A(n8920), .ZN(n4432) );
  NAND2_X1 U5972 ( .A1(n7762), .A2(n7761), .ZN(n8533) );
  INV_X1 U5973 ( .A(n8533), .ZN(n4673) );
  INV_X1 U5974 ( .A(n4739), .ZN(n4738) );
  NOR2_X1 U5975 ( .A1(n8379), .A2(n4740), .ZN(n4739) );
  NOR2_X1 U5976 ( .A1(n7354), .A2(n7355), .ZN(n4379) );
  INV_X1 U5977 ( .A(n8871), .ZN(n4443) );
  INV_X1 U5978 ( .A(n4704), .ZN(n4703) );
  OR2_X1 U5979 ( .A1(n8198), .A2(n4705), .ZN(n4704) );
  OR2_X1 U5980 ( .A1(n9081), .A2(n6151), .ZN(n4380) );
  INV_X1 U5981 ( .A(n9485), .ZN(n9144) );
  NAND2_X1 U5982 ( .A1(n8739), .A2(n8738), .ZN(n9485) );
  OR2_X1 U5983 ( .A1(n4504), .A2(n6198), .ZN(n4381) );
  NOR2_X1 U5984 ( .A1(n9288), .A2(n9375), .ZN(n9263) );
  INV_X1 U5985 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9515) );
  AND2_X1 U5986 ( .A1(n6601), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4382) );
  INV_X1 U5987 ( .A(n8086), .ZN(n4494) );
  OR2_X1 U5988 ( .A1(n7102), .A2(n8887), .ZN(n7264) );
  AND2_X1 U5989 ( .A1(n5392), .A2(SI_18_), .ZN(n4383) );
  INV_X1 U5990 ( .A(n4756), .ZN(n4755) );
  AND2_X1 U5991 ( .A1(n4581), .A2(n4580), .ZN(n4384) );
  INV_X1 U5992 ( .A(n8034), .ZN(n4726) );
  AND2_X1 U5993 ( .A1(n4747), .A2(n4337), .ZN(n4385) );
  AND2_X1 U5994 ( .A1(n4849), .A2(n4376), .ZN(n4386) );
  AND2_X1 U5995 ( .A1(n4445), .A2(n8086), .ZN(n4387) );
  AND2_X1 U5996 ( .A1(n7593), .A2(n4596), .ZN(n4388) );
  INV_X1 U5997 ( .A(n5067), .ZN(n5399) );
  NAND2_X2 U5998 ( .A1(n8014), .A2(n7816), .ZN(n7947) );
  NAND2_X1 U5999 ( .A1(n7065), .A2(n7064), .ZN(n8607) );
  INV_X1 U6000 ( .A(n8607), .ZN(n4675) );
  NAND2_X1 U6001 ( .A1(n6054), .A2(n6053), .ZN(n8196) );
  NAND2_X1 U6002 ( .A1(n5348), .A2(n5347), .ZN(n9391) );
  INV_X1 U6003 ( .A(n9391), .ZN(n4613) );
  NAND2_X1 U6004 ( .A1(n6879), .A2(n8955), .ZN(n7103) );
  NAND2_X1 U6005 ( .A1(n7680), .A2(n7679), .ZN(n8571) );
  INV_X1 U6006 ( .A(n8571), .ZN(n4745) );
  NAND2_X1 U6007 ( .A1(n6969), .A2(n7858), .ZN(n7041) );
  NAND2_X1 U6008 ( .A1(n4776), .A2(n7866), .ZN(n6987) );
  AND2_X1 U6009 ( .A1(n4497), .A2(n4499), .ZN(n4389) );
  NAND2_X1 U6010 ( .A1(n6918), .A2(n6917), .ZN(n8612) );
  INV_X1 U6011 ( .A(n8612), .ZN(n4676) );
  OR2_X1 U6012 ( .A1(n7519), .A2(n7518), .ZN(n4390) );
  NAND2_X1 U6013 ( .A1(n7699), .A2(n7698), .ZN(n8558) );
  INV_X1 U6014 ( .A(n8558), .ZN(n4678) );
  NAND2_X1 U6015 ( .A1(n4717), .A2(n6864), .ZN(n6962) );
  NOR2_X1 U6016 ( .A1(n6663), .A2(n4501), .ZN(n4391) );
  INV_X1 U6017 ( .A(n6696), .ZN(n6691) );
  AND2_X2 U6018 ( .A1(n6433), .A2(n6432), .ZN(n9888) );
  NAND2_X1 U6019 ( .A1(n4831), .A2(n4830), .ZN(n9317) );
  AND2_X2 U6020 ( .A1(n7114), .A2(n7113), .ZN(n9729) );
  INV_X1 U6021 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n4398) );
  INV_X1 U6022 ( .A(n4925), .ZN(n6502) );
  INV_X1 U6023 ( .A(n9704), .ZN(n4606) );
  AND2_X1 U6024 ( .A1(n4950), .A2(n4949), .ZN(n6207) );
  OR2_X1 U6025 ( .A1(n8250), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4392) );
  AND2_X1 U6026 ( .A1(n9113), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4393) );
  AND2_X1 U6027 ( .A1(n7985), .A2(n7786), .ZN(n4394) );
  AND2_X1 U6028 ( .A1(n4939), .A2(P1_STATE_REG_SCAN_IN), .ZN(n4395) );
  INV_X1 U6029 ( .A(n6661), .ZN(n4399) );
  NOR2_X1 U6030 ( .A1(n5822), .A2(n4628), .ZN(n6372) );
  INV_X1 U6031 ( .A(n6372), .ZN(n4478) );
  INV_X1 U6032 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U6033 ( .A1(n4914), .A2(n4913), .ZN(n5774) );
  NAND2_X1 U6034 ( .A1(n4396), .A2(n4964), .ZN(n4989) );
  NAND2_X1 U6035 ( .A1(n4962), .A2(n4961), .ZN(n4396) );
  INV_X1 U6036 ( .A(n5680), .ZN(n5716) );
  NAND2_X1 U6037 ( .A1(n4645), .A2(n4367), .ZN(n5714) );
  NAND2_X1 U6038 ( .A1(n6938), .A2(n5200), .ZN(n6939) );
  NAND2_X1 U6039 ( .A1(n4638), .A2(n4637), .ZN(n5311) );
  NAND2_X1 U6040 ( .A1(n7386), .A2(n4434), .ZN(n4430) );
  NAND2_X1 U6041 ( .A1(n4431), .A2(n4430), .ZN(n7634) );
  NAND3_X1 U6042 ( .A1(n6622), .A2(n4448), .A3(n8945), .ZN(n4447) );
  NAND2_X1 U6043 ( .A1(n6622), .A2(n9003), .ZN(n6623) );
  NAND2_X1 U6044 ( .A1(n7260), .A2(n4450), .ZN(n7419) );
  INV_X2 U6045 ( .A(n4895), .ZN(n4873) );
  NAND3_X1 U6046 ( .A1(n4866), .A2(n5086), .A3(n4453), .ZN(n4895) );
  AND3_X2 U6047 ( .A1(n4456), .A2(n4455), .A3(n4454), .ZN(n5086) );
  NAND2_X1 U6048 ( .A1(n8318), .A2(n7808), .ZN(n7746) );
  NAND2_X1 U6049 ( .A1(n8338), .A2(n7810), .ZN(n4459) );
  NAND2_X1 U6050 ( .A1(n6748), .A2(n7838), .ZN(n4460) );
  INV_X1 U6051 ( .A(n4771), .ZN(n4462) );
  OAI211_X1 U6052 ( .C1(n4772), .C2(n4464), .A(n4461), .B(n7799), .ZN(n4463)
         );
  NAND2_X1 U6053 ( .A1(n4462), .A2(n7858), .ZN(n4461) );
  NAND2_X1 U6054 ( .A1(n4463), .A2(n7859), .ZN(n7004) );
  INV_X1 U6055 ( .A(n4753), .ZN(n4475) );
  AOI21_X1 U6056 ( .B1(n4473), .B2(n4475), .A(n4469), .ZN(n4466) );
  NAND2_X1 U6057 ( .A1(n4472), .A2(n4473), .ZN(n4467) );
  INV_X1 U6058 ( .A(n7696), .ZN(n4469) );
  NAND2_X1 U6059 ( .A1(n4753), .A2(n7696), .ZN(n4470) );
  NAND2_X1 U6060 ( .A1(n8451), .A2(n4753), .ZN(n4471) );
  INV_X1 U6061 ( .A(n8451), .ZN(n4472) );
  NAND2_X2 U6062 ( .A1(n6263), .A2(n4914), .ZN(n5856) );
  NAND2_X2 U6063 ( .A1(n8056), .A2(n6280), .ZN(n6263) );
  NAND3_X1 U6064 ( .A1(n4479), .A2(n5744), .A3(n5750), .ZN(n4480) );
  NAND3_X2 U6065 ( .A1(n5733), .A2(n5732), .A3(n5822), .ZN(n6539) );
  NAND2_X1 U6066 ( .A1(n4863), .A2(n6988), .ZN(n7145) );
  NAND2_X1 U6067 ( .A1(n7455), .A2(n4783), .ZN(n7458) );
  NOR2_X2 U6068 ( .A1(n4871), .A2(n4870), .ZN(n4872) );
  NAND3_X1 U6069 ( .A1(n6582), .A2(n4389), .A3(n4503), .ZN(n4496) );
  AND2_X1 U6070 ( .A1(n4503), .A2(n4499), .ZN(n4498) );
  OR2_X1 U6071 ( .A1(n9601), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4503) );
  INV_X1 U6072 ( .A(n4502), .ZN(n6660) );
  NAND2_X1 U6073 ( .A1(n9563), .A2(n6157), .ZN(n6161) );
  OAI21_X1 U6074 ( .B1(n7208), .B2(n4510), .A(n4509), .ZN(n9095) );
  AOI21_X1 U6075 ( .B1(n4528), .B2(n4526), .A(n7849), .ZN(n7856) );
  AND2_X1 U6076 ( .A1(n7841), .A2(n7846), .ZN(n4529) );
  NAND3_X1 U6077 ( .A1(n4547), .A2(n4544), .A3(n7456), .ZN(n4543) );
  NAND3_X1 U6078 ( .A1(n7873), .A2(n7879), .A3(n7876), .ZN(n4546) );
  NAND3_X1 U6079 ( .A1(n7880), .A2(n7879), .A3(n7878), .ZN(n4550) );
  NAND2_X1 U6080 ( .A1(n5748), .A2(n4369), .ZN(n5776) );
  NAND2_X1 U6081 ( .A1(n5776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5763) );
  NAND3_X1 U6082 ( .A1(n7905), .A2(n7917), .A3(n8409), .ZN(n4558) );
  OR2_X1 U6083 ( .A1(n4568), .A2(n7984), .ZN(n4560) );
  NAND2_X1 U6084 ( .A1(n8132), .A2(n4563), .ZN(n4561) );
  NAND3_X1 U6085 ( .A1(n4567), .A2(n4707), .A3(n4565), .ZN(n4706) );
  AND2_X1 U6086 ( .A1(n4568), .A2(n7984), .ZN(n4566) );
  NAND2_X1 U6087 ( .A1(n4358), .A2(n7984), .ZN(n4567) );
  NAND2_X1 U6088 ( .A1(n7983), .A2(n7982), .ZN(n4568) );
  NAND3_X1 U6089 ( .A1(n4574), .A2(n4579), .A3(n4570), .ZN(n7979) );
  NAND3_X1 U6090 ( .A1(n7308), .A2(n4576), .A3(n4575), .ZN(n4574) );
  NAND3_X1 U6091 ( .A1(n4578), .A2(n4577), .A3(n7588), .ZN(n4581) );
  XNOR2_X1 U6092 ( .A(n7979), .B(n7975), .ZN(n8018) );
  OR2_X1 U6093 ( .A1(n5282), .A2(n5281), .ZN(n4589) );
  AOI21_X1 U6094 ( .B1(n7304), .B2(n4597), .A(n4388), .ZN(n4594) );
  NAND2_X1 U6095 ( .A1(n7304), .A2(n5928), .ZN(n4599) );
  NOR2_X1 U6096 ( .A1(n7439), .A2(n7306), .ZN(n7440) );
  NAND2_X1 U6097 ( .A1(n5161), .A2(n5160), .ZN(n5179) );
  NAND2_X1 U6098 ( .A1(n4796), .A2(n4795), .ZN(n5235) );
  NAND3_X1 U6099 ( .A1(n4605), .A2(n4708), .A3(n8185), .ZN(n4604) );
  NAND3_X1 U6100 ( .A1(n4873), .A2(n4852), .A3(n4872), .ZN(n4609) );
  NAND2_X1 U6101 ( .A1(n4609), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U6102 ( .A1(n4873), .A2(n4872), .ZN(n4890) );
  AND2_X1 U6103 ( .A1(n9181), .A2(n4617), .ZN(n9143) );
  NAND2_X1 U6104 ( .A1(n9181), .A2(n4615), .ZN(n9142) );
  NAND2_X1 U6105 ( .A1(n9181), .A2(n4619), .ZN(n9152) );
  NAND2_X1 U6106 ( .A1(n9181), .A2(n9172), .ZN(n9167) );
  NOR2_X2 U6107 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5806) );
  NAND3_X1 U6108 ( .A1(n5258), .A2(n4640), .A3(n5257), .ZN(n4638) );
  NAND2_X1 U6109 ( .A1(n5258), .A2(n5257), .ZN(n7233) );
  NOR2_X1 U6110 ( .A1(n7234), .A2(n7235), .ZN(n4639) );
  NAND2_X1 U6111 ( .A1(n7234), .A2(n7235), .ZN(n4640) );
  NAND2_X1 U6112 ( .A1(n4922), .A2(n4641), .ZN(n4934) );
  AND2_X1 U6113 ( .A1(n4921), .A2(n4919), .ZN(n4642) );
  NOR2_X1 U6114 ( .A1(n8685), .A2(n5531), .ZN(n5629) );
  NAND2_X1 U6115 ( .A1(n8685), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U6116 ( .A1(n6516), .A2(n6517), .ZN(n5103) );
  NOR2_X1 U6117 ( .A1(n5077), .A2(n6438), .ZN(n4648) );
  AND2_X1 U6118 ( .A1(n4872), .A2(n4653), .ZN(n4649) );
  AND2_X1 U6119 ( .A1(n4364), .A2(n4872), .ZN(n4651) );
  NAND2_X1 U6120 ( .A1(n4873), .A2(n4649), .ZN(n4652) );
  AOI21_X1 U6121 ( .B1(n4873), .B2(n4651), .A(n4650), .ZN(n4906) );
  MUX2_X1 U6122 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9433), .S(n4939), .Z(n6509) );
  NAND2_X1 U6123 ( .A1(n4666), .A2(n4665), .ZN(n6726) );
  AND2_X1 U6124 ( .A1(n5157), .A2(n4667), .ZN(n4665) );
  OAI22_X1 U6125 ( .A1(n6620), .A2(n5672), .B1(n6313), .B2(n5096), .ZN(n5001)
         );
  NAND2_X1 U6126 ( .A1(n6819), .A2(n6820), .ZN(n6938) );
  NAND2_X1 U6127 ( .A1(n8671), .A2(n8672), .ZN(n8670) );
  NAND2_X1 U6128 ( .A1(n7132), .A2(n7133), .ZN(n7137) );
  NAND2_X1 U6129 ( .A1(n6726), .A2(n5158), .ZN(n6819) );
  NAND2_X1 U6130 ( .A1(n7611), .A2(n7614), .ZN(n5385) );
  NOR2_X2 U6131 ( .A1(n7965), .A2(n9804), .ZN(n6840) );
  NAND2_X1 U6132 ( .A1(n6541), .A2(n4682), .ZN(n5791) );
  INV_X1 U6133 ( .A(n5791), .ZN(n5735) );
  NAND2_X1 U6134 ( .A1(n7062), .A2(n7061), .ZN(n7066) );
  INV_X1 U6135 ( .A(n7308), .ZN(n4692) );
  NAND2_X1 U6136 ( .A1(n7308), .A2(n7307), .ZN(n7443) );
  NAND2_X1 U6137 ( .A1(n4342), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U6138 ( .A1(n6263), .A2(n4709), .ZN(n5810) );
  NAND2_X1 U6139 ( .A1(n4715), .A2(n6856), .ZN(n4713) );
  INV_X1 U6140 ( .A(n8438), .ZN(n4727) );
  NAND2_X1 U6141 ( .A1(n4723), .A2(n4724), .ZN(n8037) );
  NAND2_X1 U6142 ( .A1(n8438), .A2(n8034), .ZN(n4723) );
  NAND2_X1 U6143 ( .A1(n6851), .A2(n4363), .ZN(n4728) );
  NAND2_X1 U6144 ( .A1(n4728), .A2(n4365), .ZN(n6852) );
  OAI21_X1 U6145 ( .B1(n7539), .B2(n4731), .A(n4371), .ZN(n8030) );
  NAND3_X1 U6146 ( .A1(n4737), .A2(n4738), .A3(n8370), .ZN(n4735) );
  OR2_X1 U6147 ( .A1(n8558), .A2(n8390), .ZN(n4743) );
  NAND2_X1 U6148 ( .A1(n7150), .A2(n4749), .ZN(n4748) );
  CLKBUF_X1 U6149 ( .A(n4748), .Z(n4747) );
  NAND2_X1 U6150 ( .A1(n7150), .A2(n7149), .ZN(n7151) );
  INV_X1 U6151 ( .A(n7149), .ZN(n4750) );
  NOR2_X2 U6152 ( .A1(n6539), .A2(n5745), .ZN(n5748) );
  NAND2_X1 U6153 ( .A1(n8304), .A2(n4760), .ZN(n4759) );
  NAND2_X1 U6154 ( .A1(n8304), .A2(n7811), .ZN(n4763) );
  NAND2_X1 U6155 ( .A1(n4763), .A2(n4762), .ZN(n8051) );
  NAND2_X1 U6156 ( .A1(n7457), .A2(n4768), .ZN(n4765) );
  NAND2_X1 U6157 ( .A1(n4765), .A2(n4766), .ZN(n8493) );
  NAND2_X1 U6158 ( .A1(n7708), .A2(n4780), .ZN(n4777) );
  NAND2_X1 U6159 ( .A1(n8064), .A2(n9804), .ZN(n6836) );
  NAND2_X1 U6160 ( .A1(n5760), .A2(n4784), .ZN(n4786) );
  NAND2_X1 U6161 ( .A1(n5090), .A2(n5089), .ZN(n5093) );
  NAND2_X1 U6162 ( .A1(n5070), .A2(n5069), .ZN(n4787) );
  NAND2_X1 U6163 ( .A1(n9187), .A2(n4790), .ZN(n4788) );
  INV_X1 U6164 ( .A(n9215), .ZN(n4813) );
  NAND3_X1 U6165 ( .A1(n4816), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4815) );
  NAND3_X1 U6166 ( .A1(n4912), .A2(n9135), .A3(n4818), .ZN(n4817) );
  AOI22_X1 U6167 ( .A1(n9632), .A2(n5622), .B1(n4940), .B2(n4970), .ZN(n4979)
         );
  NAND4_X2 U6168 ( .A1(n4973), .A2(n4971), .A3(n4972), .A4(n4974), .ZN(n9632)
         );
  INV_X1 U6169 ( .A(n9331), .ZN(n4819) );
  NAND2_X1 U6170 ( .A1(n4819), .A2(n9729), .ZN(n4820) );
  OAI211_X1 U6171 ( .C1(n9332), .C2(n4821), .A(n4820), .B(n4827), .ZN(P1_U3552) );
  NAND2_X1 U6172 ( .A1(n9149), .A2(n8905), .ZN(n4823) );
  NAND3_X1 U6173 ( .A1(n4824), .A2(n4823), .A3(n4822), .ZN(n9332) );
  INV_X1 U6174 ( .A(n9319), .ZN(n4831) );
  NAND2_X1 U6175 ( .A1(n7280), .A2(n4835), .ZN(n4832) );
  NAND2_X1 U6176 ( .A1(n4832), .A2(n4833), .ZN(n7622) );
  NAND3_X1 U6177 ( .A1(n4836), .A2(n7408), .A3(n4340), .ZN(n4834) );
  NAND2_X1 U6178 ( .A1(n4838), .A2(n4839), .ZN(n7278) );
  NAND2_X1 U6179 ( .A1(n7102), .A2(n7263), .ZN(n4838) );
  NAND2_X1 U6180 ( .A1(n8078), .A2(n4842), .ZN(n4841) );
  NAND3_X1 U6181 ( .A1(n5086), .A2(n4866), .A3(n4867), .ZN(n5241) );
  AND2_X1 U6182 ( .A1(n8382), .A2(n8381), .ZN(n8568) );
  AOI21_X1 U6183 ( .B1(n5716), .B2(n5698), .A(n5697), .ZN(n5699) );
  NAND2_X1 U6184 ( .A1(n4939), .A2(n4914), .ZN(n5067) );
  NAND2_X2 U6185 ( .A1(n5765), .A2(n8642), .ZN(n5850) );
  INV_X1 U6186 ( .A(n5385), .ZN(n5388) );
  NAND2_X1 U6187 ( .A1(n6488), .A2(n5622), .ZN(n4949) );
  INV_X1 U6188 ( .A(n6412), .ZN(n6829) );
  OAI21_X1 U6189 ( .B1(n5716), .B2(n5715), .A(n8683), .ZN(n5721) );
  NAND2_X1 U6190 ( .A1(n7278), .A2(n7277), .ZN(n7281) );
  AND2_X1 U6191 ( .A1(n5629), .A2(n5628), .ZN(n5582) );
  AOI21_X1 U6192 ( .B1(n5714), .B2(n5656), .A(n5651), .ZN(n5715) );
  NAND2_X1 U6193 ( .A1(n6208), .A2(n4955), .ZN(n6223) );
  INV_X1 U6194 ( .A(n8683), .ZN(n8716) );
  AND2_X1 U6195 ( .A1(n5603), .A2(n5581), .ZN(n8683) );
  AND2_X1 U6196 ( .A1(n7747), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n4853) );
  AND2_X1 U6197 ( .A1(n7512), .A2(n7511), .ZN(n4854) );
  OR2_X1 U6198 ( .A1(n8100), .A2(n8099), .ZN(n4855) );
  AND2_X1 U6199 ( .A1(n5794), .A2(n5734), .ZN(n4856) );
  AND2_X1 U6200 ( .A1(n5264), .A2(n5292), .ZN(n4857) );
  AND2_X1 U6201 ( .A1(n5024), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4858) );
  AND2_X1 U6202 ( .A1(n6504), .A2(n9512), .ZN(n9633) );
  NOR2_X1 U6203 ( .A1(n5374), .A2(n5350), .ZN(n4859) );
  INV_X1 U6204 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5394) );
  AND2_X1 U6205 ( .A1(n5180), .A2(n5165), .ZN(n4860) );
  NAND2_X1 U6206 ( .A1(n8101), .A2(n4855), .ZN(n4861) );
  NAND2_X1 U6207 ( .A1(n6503), .A2(n8868), .ZN(n9313) );
  AND2_X1 U6208 ( .A1(n5160), .A2(n5133), .ZN(n4862) );
  AND2_X1 U6209 ( .A1(n7605), .A2(n7604), .ZN(n8038) );
  INV_X1 U6210 ( .A(n8038), .ZN(n7976) );
  INV_X1 U6211 ( .A(n5579), .ZN(n5398) );
  INV_X1 U6212 ( .A(n8775), .ZN(n7284) );
  INV_X1 U6213 ( .A(n8310), .ZN(n8325) );
  INV_X1 U6214 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5758) );
  NOR4_X1 U6215 ( .A1(n7814), .A2(n7813), .A3(n8044), .A4(n7812), .ZN(n7815)
         );
  INV_X1 U6216 ( .A(n7071), .ZN(n6114) );
  INV_X1 U6217 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6218 ( .A1(n4942), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6219 ( .A1(n4970), .A2(n4935), .ZN(n4976) );
  INV_X1 U6220 ( .A(n8880), .ZN(n6877) );
  NAND2_X1 U6221 ( .A1(n4851), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4908) );
  INV_X1 U6222 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4864) );
  AND2_X1 U6223 ( .A1(n7953), .A2(n8499), .ZN(n5796) );
  INV_X1 U6224 ( .A(n7522), .ZN(n7521) );
  OR2_X1 U6225 ( .A1(n7598), .A2(n7597), .ZN(n7688) );
  INV_X1 U6226 ( .A(n7802), .ZN(n6988) );
  INV_X1 U6227 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9970) );
  INV_X1 U6228 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5297) );
  INV_X1 U6229 ( .A(n8888), .ZN(n7279) );
  INV_X1 U6230 ( .A(n8945), .ZN(n6671) );
  INV_X1 U6231 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4875) );
  OR2_X1 U6232 ( .A1(n4880), .A2(n5571), .ZN(n4899) );
  INV_X1 U6233 ( .A(SI_19_), .ZN(n9958) );
  INV_X1 U6234 ( .A(SI_15_), .ZN(n5286) );
  NOR2_X1 U6235 ( .A1(n5925), .A2(n8107), .ZN(n5919) );
  INV_X1 U6236 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6065) );
  OR2_X1 U6237 ( .A1(n7700), .A2(n8161), .ZN(n7714) );
  NAND2_X1 U6238 ( .A1(n7521), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7598) );
  INV_X1 U6239 ( .A(n8642), .ZN(n5766) );
  AND2_X1 U6240 ( .A1(n6267), .A2(n6266), .ZN(n6274) );
  INV_X1 U6241 ( .A(n8537), .ZN(n8047) );
  OR2_X1 U6242 ( .A1(n8549), .A2(n8320), .ZN(n8041) );
  INV_X1 U6243 ( .A(n8437), .ZN(n8033) );
  INV_X1 U6244 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5898) );
  AND2_X1 U6245 ( .A1(n5655), .A2(n5654), .ZN(n5712) );
  INV_X1 U6246 ( .A(n7499), .ZN(n5336) );
  AND2_X1 U6247 ( .A1(n5246), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5269) );
  INV_X1 U6248 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5186) );
  OR2_X1 U6249 ( .A1(n5298), .A2(n5297), .ZN(n5323) );
  NAND2_X1 U6250 ( .A1(n9263), .A2(n9370), .ZN(n9265) );
  INV_X1 U6251 ( .A(n9614), .ZN(n6680) );
  NAND2_X1 U6252 ( .A1(n4875), .A2(n4880), .ZN(n4881) );
  NAND2_X1 U6253 ( .A1(n4903), .A2(n4899), .ZN(n4900) );
  INV_X1 U6254 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5344) );
  OR2_X1 U6255 ( .A1(n5119), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6256 ( .A1(n5393), .A2(n6084), .ZN(n4994) );
  OR2_X1 U6257 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  INV_X1 U6258 ( .A(n6061), .ZN(n6074) );
  AND2_X1 U6259 ( .A1(n7301), .A2(n7300), .ZN(n7302) );
  NAND2_X1 U6260 ( .A1(n6720), .A2(n6019), .ZN(n6811) );
  INV_X1 U6261 ( .A(n8171), .ZN(n5827) );
  OR2_X1 U6262 ( .A1(n7724), .A2(n8199), .ZN(n7738) );
  OR2_X1 U6263 ( .A1(n6066), .A2(n6065), .ZN(n7071) );
  OR2_X1 U6264 ( .A1(n8313), .A2(n7763), .ZN(n7757) );
  INV_X1 U6265 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7247) );
  INV_X1 U6266 ( .A(n9734), .ZN(n9731) );
  NAND2_X1 U6267 ( .A1(n7960), .A2(n7829), .ZN(n6264) );
  OR2_X1 U6268 ( .A1(n8537), .A2(n8319), .ZN(n8043) );
  OR2_X1 U6269 ( .A1(n7040), .A2(n7799), .ZN(n7038) );
  AOI22_X1 U6270 ( .A1(n8319), .A2(n8506), .B1(n8293), .B2(n8208), .ZN(n8058)
         );
  AND2_X1 U6271 ( .A1(n9805), .A2(n6074), .ZN(n9836) );
  OR2_X1 U6272 ( .A1(n6269), .A2(n6264), .ZN(n8496) );
  INV_X4 U6273 ( .A(n4914), .ZN(n5393) );
  NAND2_X1 U6274 ( .A1(n5269), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5298) );
  NOR2_X1 U6275 ( .A1(n5713), .A2(n5712), .ZN(n5657) );
  INV_X1 U6276 ( .A(n9202), .ZN(n9229) );
  NAND2_X1 U6277 ( .A1(n5515), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5544) );
  INV_X1 U6278 ( .A(n9246), .ZN(n8705) );
  INV_X1 U6279 ( .A(n4926), .ZN(n8999) );
  AND4_X1 U6280 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n8703)
         );
  AND2_X1 U6281 ( .A1(n6162), .A2(n7550), .ZN(n9585) );
  AND2_X1 U6282 ( .A1(n8809), .A2(n9297), .ZN(n8896) );
  OR2_X1 U6283 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  OR2_X1 U6284 ( .A1(n6212), .A2(n6211), .ZN(n7111) );
  INV_X1 U6285 ( .A(n8893), .ZN(n7410) );
  NAND2_X1 U6286 ( .A1(n6504), .A2(n5590), .ZN(n9616) );
  INV_X1 U6287 ( .A(n6889), .ZN(n9692) );
  OAI21_X1 U6288 ( .B1(n7774), .B2(n7773), .A(n7772), .ZN(n7779) );
  AND2_X1 U6289 ( .A1(n5632), .A2(n5616), .ZN(n5630) );
  AND2_X1 U6290 ( .A1(n5341), .A2(n5318), .ZN(n5339) );
  OR3_X1 U6291 ( .A1(n7321), .A2(n7533), .A3(n7484), .ZN(n6261) );
  INV_X1 U6292 ( .A(n6075), .ZN(n6054) );
  AND2_X1 U6293 ( .A1(n7738), .A2(n7725), .ZN(n8345) );
  INV_X1 U6294 ( .A(n8196), .ZN(n8185) );
  INV_X1 U6295 ( .A(n7764), .ZN(n7728) );
  INV_X1 U6296 ( .A(n8282), .ZN(n9735) );
  AND2_X1 U6297 ( .A1(n6275), .A2(n8056), .ZN(n9734) );
  INV_X1 U6298 ( .A(n8039), .ZN(n8370) );
  INV_X1 U6299 ( .A(n7537), .ZN(n7887) );
  INV_X1 U6300 ( .A(n8496), .ZN(n8508) );
  AND2_X1 U6301 ( .A1(n9798), .A2(n6050), .ZN(n6737) );
  AND2_X1 U6302 ( .A1(n8532), .A2(n9849), .ZN(n9871) );
  INV_X1 U6303 ( .A(n9871), .ZN(n9885) );
  NAND2_X1 U6304 ( .A1(n6261), .A2(n9797), .ZN(n9765) );
  INV_X1 U6305 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5786) );
  INV_X1 U6306 ( .A(n4957), .ZN(n6226) );
  INV_X1 U6307 ( .A(n8703), .ZN(n9280) );
  AND4_X1 U6308 ( .A1(n5379), .A2(n5378), .A3(n5377), .A4(n5376), .ZN(n7633)
         );
  AND4_X1 U6309 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n7322)
         );
  AND2_X1 U6310 ( .A1(n9585), .A2(n9512), .ZN(n9598) );
  INV_X1 U6311 ( .A(n9578), .ZN(n9587) );
  INV_X1 U6312 ( .A(n9598), .ZN(n9553) );
  INV_X1 U6313 ( .A(n5602), .ZN(n6482) );
  INV_X1 U6314 ( .A(n8901), .ZN(n9176) );
  AND2_X1 U6315 ( .A1(n9186), .A2(n8835), .ZN(n9200) );
  INV_X1 U6316 ( .A(n9296), .ZN(n9285) );
  OR2_X1 U6317 ( .A1(n5604), .A2(n9706), .ZN(n9641) );
  AND2_X1 U6318 ( .A1(n7290), .A2(n9671), .ZN(n9696) );
  INV_X1 U6319 ( .A(n9696), .ZN(n9710) );
  INV_X1 U6320 ( .A(n6246), .ZN(n7114) );
  OR2_X1 U6321 ( .A1(n5568), .A2(n5556), .ZN(n6241) );
  AND2_X1 U6322 ( .A1(n5046), .A2(n5045), .ZN(n6178) );
  AND2_X1 U6323 ( .A1(n6124), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9797) );
  INV_X1 U6324 ( .A(n8397), .ZN(n8563) );
  INV_X1 U6325 ( .A(n4315), .ZN(n8207) );
  INV_X1 U6326 ( .A(n8201), .ZN(n8340) );
  INV_X1 U6327 ( .A(n7676), .ZN(n8454) );
  INV_X1 U6328 ( .A(n6985), .ZN(n8214) );
  INV_X1 U6329 ( .A(n8285), .ZN(n9730) );
  NAND2_X1 U6330 ( .A1(n9763), .A2(n9749), .ZN(n8469) );
  NAND2_X1 U6331 ( .A1(n9763), .A2(n9762), .ZN(n8504) );
  INV_X1 U6332 ( .A(n9906), .ZN(n9904) );
  AND2_X1 U6333 ( .A1(n9878), .A2(n9877), .ZN(n9903) );
  INV_X1 U6334 ( .A(n9888), .ZN(n9887) );
  NOR2_X1 U6335 ( .A1(n9766), .A2(n9765), .ZN(n9780) );
  CLKBUF_X1 U6336 ( .A(n9780), .Z(n9802) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7319) );
  INV_X1 U6338 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10103) );
  CLKBUF_X1 U6339 ( .A(n8647), .Z(n8016) );
  INV_X1 U6340 ( .A(n9358), .ZN(n9228) );
  OAI21_X1 U6341 ( .B1(n5582), .B2(n5703), .A(n8683), .ZN(n5608) );
  AND2_X1 U6342 ( .A1(n5605), .A2(n9641), .ZN(n8730) );
  INV_X1 U6343 ( .A(n8079), .ZN(n9190) );
  INV_X1 U6344 ( .A(n7633), .ZN(n9300) );
  INV_X1 U6345 ( .A(n7225), .ZN(n9062) );
  OR2_X1 U6346 ( .A1(n9521), .A2(n9036), .ZN(n9573) );
  OR2_X1 U6347 ( .A1(P1_U3083), .A2(n6132), .ZN(n9584) );
  OR2_X1 U6348 ( .A1(n9256), .A2(n9255), .ZN(n9368) );
  NAND2_X1 U6349 ( .A1(n9646), .A2(n6684), .ZN(n9306) );
  NAND2_X1 U6350 ( .A1(n6685), .A2(n9641), .ZN(n9646) );
  INV_X1 U6351 ( .A(n9729), .ZN(n9726) );
  INV_X1 U6352 ( .A(n9714), .ZN(n9712) );
  AND2_X2 U6353 ( .A1(n6247), .A2(n7114), .ZN(n9714) );
  NAND2_X1 U6354 ( .A1(n9038), .A2(n6241), .ZN(n9650) );
  INV_X1 U6355 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10072) );
  INV_X1 U6356 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6188) );
  NOR2_X1 U6357 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  AND2_X1 U6358 ( .A1(n5756), .A2(n9797), .ZN(P2_U3966) );
  INV_X2 U6359 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U6360 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4869) );
  NOR2_X1 U6361 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4868) );
  NAND4_X1 U6362 ( .A1(n4869), .A2(n4868), .A3(n5572), .A4(n9970), .ZN(n4871)
         );
  NAND4_X1 U6363 ( .A1(n5344), .A2(n5264), .A3(n5573), .A4(n4896), .ZN(n4870)
         );
  NAND2_X1 U6364 ( .A1(n4878), .A2(n4875), .ZN(n4879) );
  INV_X1 U6365 ( .A(n4878), .ZN(n4910) );
  NAND2_X1 U6366 ( .A1(n4910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U6367 ( .A1(n5025), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4888) );
  INV_X1 U6368 ( .A(n4883), .ZN(n9423) );
  NAND2_X1 U6369 ( .A1(n5030), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4887) );
  AND2_X2 U6370 ( .A1(n9426), .A2(n4883), .ZN(n5024) );
  NAND2_X1 U6371 ( .A1(n5024), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U6372 ( .A1(n5026), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4885) );
  INV_X1 U6373 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6374 ( .A1(n4890), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4891) );
  NOR2_X1 U6375 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4897) );
  NAND4_X1 U6376 ( .A1(n4927), .A2(n4897), .A3(n4896), .A4(n5292), .ZN(n4898)
         );
  NAND2_X1 U6377 ( .A1(n4900), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4902) );
  INV_X1 U6378 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6379 ( .A1(n4901), .A2(n5572), .ZN(n4923) );
  INV_X1 U6380 ( .A(n4933), .ZN(n6495) );
  NAND2_X1 U6381 ( .A1(n6489), .A2(n4940), .ZN(n4922) );
  OAI21_X1 U6382 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U6383 ( .A1(n4907), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4909) );
  INV_X2 U6384 ( .A(n4965), .ZN(n4914) );
  AND2_X1 U6385 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4913) );
  NAND3_X1 U6386 ( .A1(n4965), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4915) );
  NAND2_X1 U6387 ( .A1(n5774), .A2(n4915), .ZN(n4963) );
  INV_X1 U6388 ( .A(SI_1_), .ZN(n4916) );
  MUX2_X1 U6389 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4965), .Z(n4961) );
  XNOR2_X1 U6390 ( .A(n4962), .B(n4961), .ZN(n6095) );
  INV_X1 U6391 ( .A(n6095), .ZN(n4917) );
  NAND2_X1 U6392 ( .A1(n8080), .A2(n4917), .ZN(n4921) );
  INV_X1 U6393 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U6394 ( .A1(n5040), .A2(n9072), .ZN(n4919) );
  INV_X1 U6395 ( .A(n5343), .ZN(n4930) );
  INV_X1 U6396 ( .A(n4927), .ZN(n4928) );
  NOR2_X1 U6397 ( .A1(n4928), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U6398 ( .A1(n5575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4931) );
  AND2_X4 U6399 ( .A1(n4935), .A2(n6251), .ZN(n5622) );
  NAND2_X1 U6400 ( .A1(n6489), .A2(n5622), .ZN(n4937) );
  OR2_X1 U6401 ( .A1(n6487), .A2(n5672), .ZN(n4936) );
  NAND2_X1 U6402 ( .A1(n4937), .A2(n4936), .ZN(n4958) );
  NAND2_X1 U6403 ( .A1(n4957), .A2(n4958), .ZN(n4956) );
  NAND2_X1 U6404 ( .A1(n7775), .A2(SI_0_), .ZN(n4938) );
  XNOR2_X1 U6405 ( .A(n4938), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U6406 ( .A1(n6509), .A2(n4940), .ZN(n4944) );
  NAND2_X1 U6407 ( .A1(n5026), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U6408 ( .A1(n5025), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U6409 ( .A1(n5024), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U6410 ( .A1(n6488), .A2(n4940), .ZN(n4953) );
  INV_X1 U6411 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9510) );
  NOR2_X1 U6412 ( .A1(n5723), .A2(n9510), .ZN(n4951) );
  NAND2_X1 U6413 ( .A1(n4953), .A2(n4952), .ZN(n6209) );
  INV_X1 U6414 ( .A(n6209), .ZN(n4954) );
  NAND2_X1 U6415 ( .A1(n4954), .A2(n5049), .ZN(n4955) );
  NAND2_X1 U6416 ( .A1(n4956), .A2(n6223), .ZN(n4960) );
  INV_X1 U6417 ( .A(n4958), .ZN(n6224) );
  NAND2_X1 U6418 ( .A1(n6226), .A2(n6224), .ZN(n4959) );
  NAND2_X1 U6419 ( .A1(n4960), .A2(n4959), .ZN(n6235) );
  NOR2_X1 U6420 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5042) );
  OR2_X1 U6421 ( .A1(n5042), .A2(n4880), .ZN(n4996) );
  INV_X1 U6422 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4995) );
  XNOR2_X1 U6423 ( .A(n4996), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U6424 ( .A1(n5040), .A2(n9529), .ZN(n4968) );
  NAND2_X1 U6425 ( .A1(n4963), .A2(SI_1_), .ZN(n4964) );
  INV_X1 U6426 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6094) );
  INV_X1 U6427 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6083) );
  MUX2_X1 U6428 ( .A(n6094), .B(n6083), .S(n4965), .Z(n4990) );
  XNOR2_X1 U6429 ( .A(n4990), .B(SI_2_), .ZN(n4988) );
  XNOR2_X1 U6430 ( .A(n4989), .B(n4988), .ZN(n6093) );
  INV_X1 U6431 ( .A(n6093), .ZN(n4966) );
  NAND2_X1 U6432 ( .A1(n8080), .A2(n4966), .ZN(n4967) );
  NAND2_X1 U6433 ( .A1(n5024), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6434 ( .A1(n5025), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6435 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  XNOR2_X1 U6436 ( .A(n4977), .B(n5049), .ZN(n4978) );
  XNOR2_X1 U6437 ( .A(n4978), .B(n4979), .ZN(n6234) );
  NAND2_X1 U6438 ( .A1(n6235), .A2(n6234), .ZN(n4982) );
  INV_X1 U6439 ( .A(n4978), .ZN(n4980) );
  NAND2_X1 U6440 ( .A1(n4980), .A2(n4979), .ZN(n4981) );
  NAND2_X1 U6441 ( .A1(n4982), .A2(n4981), .ZN(n6310) );
  NAND2_X1 U6442 ( .A1(n5024), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U6443 ( .A1(n5025), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4986) );
  INV_X1 U6444 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U6445 ( .A1(n5030), .A2(n4983), .ZN(n4985) );
  NAND2_X1 U6446 ( .A1(n5026), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6447 ( .A1(n4989), .A2(n4988), .ZN(n4993) );
  INV_X1 U6448 ( .A(n4990), .ZN(n4991) );
  NAND2_X1 U6449 ( .A1(n4991), .A2(SI_2_), .ZN(n4992) );
  INV_X1 U6450 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6092) );
  INV_X1 U6451 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U6452 ( .A(n5004), .B(SI_3_), .ZN(n5002) );
  XNOR2_X1 U6453 ( .A(n5003), .B(n5002), .ZN(n6091) );
  OR2_X1 U6454 ( .A1(n5067), .A2(n6084), .ZN(n5000) );
  NAND2_X1 U6455 ( .A1(n4996), .A2(n4995), .ZN(n4997) );
  NAND2_X1 U6456 ( .A1(n4997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6457 ( .A1(n5040), .A2(n9083), .ZN(n4999) );
  XNOR2_X1 U6458 ( .A(n5001), .B(n5097), .ZN(n5021) );
  OAI22_X1 U6459 ( .A1(n6620), .A2(n5051), .B1(n6313), .B2(n5672), .ZN(n5019)
         );
  XNOR2_X1 U6460 ( .A(n5021), .B(n5019), .ZN(n6311) );
  NAND2_X1 U6461 ( .A1(n6310), .A2(n6311), .ZN(n6562) );
  NAND2_X1 U6462 ( .A1(n5003), .A2(n5002), .ZN(n5007) );
  INV_X1 U6463 ( .A(n5004), .ZN(n5005) );
  NAND2_X1 U6464 ( .A1(n5005), .A2(SI_3_), .ZN(n5006) );
  MUX2_X1 U6465 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5393), .Z(n5037) );
  XNOR2_X1 U6466 ( .A(n5037), .B(SI_4_), .ZN(n5034) );
  XNOR2_X1 U6467 ( .A(n5036), .B(n5034), .ZN(n5857) );
  INV_X1 U6468 ( .A(n5857), .ZN(n6089) );
  NAND2_X1 U6469 ( .A1(n8733), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5012) );
  NOR2_X1 U6470 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5008) );
  NAND2_X1 U6471 ( .A1(n5042), .A2(n5008), .ZN(n5009) );
  NAND2_X1 U6472 ( .A1(n5009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5010) );
  XNOR2_X1 U6473 ( .A(n5010), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U6474 ( .A1(n4316), .A2(n9541), .ZN(n5011) );
  INV_X1 U6475 ( .A(n6559), .ZN(n6675) );
  NAND2_X1 U6476 ( .A1(n5024), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5017) );
  INV_X1 U6477 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5013) );
  XNOR2_X1 U6478 ( .A(n5013), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U6479 ( .A1(n5030), .A2(n6632), .ZN(n5016) );
  NAND2_X1 U6480 ( .A1(n5025), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U6481 ( .A1(n5026), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5014) );
  OAI22_X1 U6482 ( .A1(n6675), .A2(n5096), .B1(n6676), .B2(n5672), .ZN(n5018)
         );
  XNOR2_X1 U6483 ( .A(n5018), .B(n5049), .ZN(n5055) );
  OAI22_X1 U6484 ( .A1(n6676), .A2(n5051), .B1(n6675), .B2(n5672), .ZN(n5054)
         );
  XNOR2_X1 U6485 ( .A(n5055), .B(n5054), .ZN(n6561) );
  INV_X1 U6486 ( .A(n5019), .ZN(n5020) );
  NAND2_X1 U6487 ( .A1(n5021), .A2(n5020), .ZN(n6563) );
  INV_X1 U6488 ( .A(n6563), .ZN(n5022) );
  NOR2_X1 U6489 ( .A1(n6561), .A2(n5022), .ZN(n5023) );
  NAND2_X1 U6490 ( .A1(n6562), .A2(n5023), .ZN(n6564) );
  INV_X4 U6491 ( .A(n8097), .ZN(n6217) );
  NAND2_X1 U6492 ( .A1(n6217), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6493 ( .A1(n5026), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6494 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  NOR2_X1 U6495 ( .A1(n4858), .A2(n5029), .ZN(n5033) );
  AOI21_X1 U6496 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U6497 ( .A1(n5031), .A2(n5062), .ZN(n9315) );
  NAND2_X1 U6498 ( .A1(n5683), .A2(n9315), .ZN(n5032) );
  INV_X1 U6499 ( .A(n5034), .ZN(n5035) );
  NAND2_X1 U6500 ( .A1(n5036), .A2(n5035), .ZN(n5039) );
  NAND2_X1 U6501 ( .A1(n5037), .A2(SI_4_), .ZN(n5038) );
  MUX2_X1 U6502 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5393), .Z(n5071) );
  XNOR2_X1 U6503 ( .A(n5071), .B(SI_5_), .ZN(n5068) );
  XNOR2_X1 U6504 ( .A(n5070), .B(n5068), .ZN(n5896) );
  INV_X1 U6505 ( .A(n5896), .ZN(n6088) );
  NAND2_X1 U6506 ( .A1(n8733), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6507 ( .A1(n5042), .A2(n5041), .ZN(n5043) );
  NAND2_X1 U6508 ( .A1(n5043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5044) );
  MUX2_X1 U6509 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5044), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5046) );
  INV_X1 U6510 ( .A(n5086), .ZN(n5045) );
  NAND2_X1 U6511 ( .A1(n4316), .A2(n6178), .ZN(n5047) );
  INV_X1 U6512 ( .A(n9676), .ZN(n6670) );
  OR2_X1 U6513 ( .A1(n6619), .A2(n5051), .ZN(n5053) );
  NAND2_X1 U6514 ( .A1(n9676), .A2(n5549), .ZN(n5052) );
  NAND2_X1 U6515 ( .A1(n5053), .A2(n5052), .ZN(n5058) );
  NAND2_X1 U6516 ( .A1(n5055), .A2(n5054), .ZN(n6454) );
  AOI21_X1 U6517 ( .B1(n6456), .B2(n5058), .A(n5056), .ZN(n5057) );
  NAND2_X1 U6518 ( .A1(n6564), .A2(n5057), .ZN(n5061) );
  INV_X1 U6519 ( .A(n6456), .ZN(n5059) );
  INV_X1 U6520 ( .A(n5058), .ZN(n6455) );
  NAND2_X1 U6521 ( .A1(n5059), .A2(n6455), .ZN(n5060) );
  NAND2_X1 U6522 ( .A1(n5024), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6523 ( .A1(n5062), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5079) );
  OAI21_X1 U6524 ( .B1(n5062), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5079), .ZN(
        n9622) );
  INV_X1 U6525 ( .A(n9622), .ZN(n6441) );
  NAND2_X1 U6526 ( .A1(n5683), .A2(n6441), .ZN(n5065) );
  NAND2_X1 U6527 ( .A1(n6217), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6528 ( .A1(n8093), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5063) );
  INV_X1 U6529 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6102) );
  INV_X1 U6530 ( .A(n5068), .ZN(n5069) );
  NAND2_X1 U6531 ( .A1(n5071), .A2(SI_5_), .ZN(n5072) );
  MUX2_X1 U6532 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5393), .Z(n5091) );
  XNOR2_X1 U6533 ( .A(n5091), .B(SI_6_), .ZN(n5088) );
  NAND2_X1 U6534 ( .A1(n8080), .A2(n6098), .ZN(n5075) );
  OR2_X1 U6535 ( .A1(n5086), .A2(n4880), .ZN(n5073) );
  XNOR2_X1 U6536 ( .A(n5073), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U6537 ( .A1(n4316), .A2(n9558), .ZN(n5074) );
  OAI211_X1 U6538 ( .C1(n5067), .C2(n6102), .A(n5075), .B(n5074), .ZN(n6672)
         );
  OAI22_X1 U6539 ( .A1(n6681), .A2(n5672), .B1(n9683), .B2(n5096), .ZN(n5076)
         );
  XNOR2_X1 U6540 ( .A(n5076), .B(n5675), .ZN(n6437) );
  OAI22_X1 U6541 ( .A1(n6681), .A2(n5051), .B1(n9683), .B2(n5672), .ZN(n6438)
         );
  INV_X1 U6542 ( .A(n6437), .ZN(n5077) );
  NAND2_X1 U6543 ( .A1(n5024), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5084) );
  AND2_X1 U6544 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  NOR2_X1 U6545 ( .A1(n5104), .A2(n5080), .ZN(n6686) );
  NAND2_X1 U6546 ( .A1(n5683), .A2(n6686), .ZN(n5083) );
  NAND2_X1 U6547 ( .A1(n6217), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6548 ( .A1(n8093), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5081) );
  INV_X1 U6549 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6550 ( .A1(n5086), .A2(n5085), .ZN(n5119) );
  NAND2_X1 U6551 ( .A1(n5119), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U6552 ( .A(n5087), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6194) );
  AOI22_X1 U6553 ( .A1(n5399), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4316), .B2(
        n6194), .ZN(n5095) );
  INV_X1 U6554 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6555 ( .A1(n5091), .A2(SI_6_), .ZN(n5092) );
  MUX2_X1 U6556 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5393), .Z(n5113) );
  XNOR2_X1 U6557 ( .A(n5113), .B(SI_7_), .ZN(n5110) );
  XNOR2_X1 U6558 ( .A(n5112), .B(n5110), .ZN(n6103) );
  INV_X2 U6559 ( .A(n5290), .ZN(n8736) );
  NAND2_X1 U6560 ( .A1(n6103), .A2(n8736), .ZN(n5094) );
  NAND2_X1 U6561 ( .A1(n5095), .A2(n5094), .ZN(n6889) );
  OAI22_X1 U6562 ( .A1(n9617), .A2(n5672), .B1(n9692), .B2(n5096), .ZN(n5098)
         );
  XNOR2_X1 U6563 ( .A(n5098), .B(n5675), .ZN(n5099) );
  OAI22_X1 U6564 ( .A1(n9617), .A2(n5051), .B1(n9692), .B2(n5672), .ZN(n5100)
         );
  XNOR2_X1 U6565 ( .A(n5099), .B(n5100), .ZN(n6517) );
  INV_X1 U6566 ( .A(n5099), .ZN(n5101) );
  NAND2_X1 U6567 ( .A1(n5101), .A2(n5100), .ZN(n5102) );
  NAND2_X1 U6568 ( .A1(n5103), .A2(n5102), .ZN(n6590) );
  NAND2_X1 U6569 ( .A1(n5024), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6570 ( .A1(n5104), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5142) );
  OR2_X1 U6571 ( .A1(n5104), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5105) );
  AND2_X1 U6572 ( .A1(n5142), .A2(n5105), .ZN(n6886) );
  NAND2_X1 U6573 ( .A1(n5683), .A2(n6886), .ZN(n5108) );
  NAND2_X1 U6574 ( .A1(n6217), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6575 ( .A1(n8093), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5106) );
  OR2_X1 U6576 ( .A1(n7225), .A2(n5051), .ZN(n5124) );
  INV_X1 U6577 ( .A(n5110), .ZN(n5111) );
  NAND2_X1 U6578 ( .A1(n5113), .A2(SI_7_), .ZN(n5114) );
  INV_X1 U6579 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6108) );
  INV_X1 U6580 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6110) );
  MUX2_X1 U6581 ( .A(n6108), .B(n6110), .S(n5393), .Z(n5116) );
  INV_X1 U6582 ( .A(SI_8_), .ZN(n5115) );
  NAND2_X1 U6583 ( .A1(n5116), .A2(n5115), .ZN(n5127) );
  INV_X1 U6584 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U6585 ( .A1(n5117), .A2(SI_8_), .ZN(n5118) );
  NAND2_X1 U6586 ( .A1(n5127), .A2(n5118), .ZN(n5128) );
  XNOR2_X1 U6587 ( .A(n5129), .B(n5128), .ZN(n6107) );
  NAND2_X1 U6588 ( .A1(n6107), .A2(n8736), .ZN(n5122) );
  NAND2_X1 U6589 ( .A1(n5134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5120) );
  XNOR2_X1 U6590 ( .A(n5120), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6292) );
  AOI22_X1 U6591 ( .A1(n5399), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4316), .B2(
        n6292), .ZN(n5121) );
  NAND2_X1 U6592 ( .A1(n7096), .A2(n5549), .ZN(n5123) );
  NAND2_X1 U6593 ( .A1(n5124), .A2(n5123), .ZN(n6592) );
  NAND2_X1 U6594 ( .A1(n7096), .A2(n5666), .ZN(n5125) );
  OAI21_X1 U6595 ( .B1(n7225), .B2(n5672), .A(n5125), .ZN(n5126) );
  XNOR2_X1 U6596 ( .A(n5126), .B(n5552), .ZN(n6591) );
  MUX2_X1 U6597 ( .A(n6131), .B(n6129), .S(n5393), .Z(n5131) );
  INV_X1 U6598 ( .A(SI_9_), .ZN(n5130) );
  NAND2_X1 U6599 ( .A1(n5131), .A2(n5130), .ZN(n5160) );
  INV_X1 U6600 ( .A(n5131), .ZN(n5132) );
  NAND2_X1 U6601 ( .A1(n5132), .A2(SI_9_), .ZN(n5133) );
  XNOR2_X1 U6602 ( .A(n5159), .B(n4862), .ZN(n6128) );
  NAND2_X1 U6603 ( .A1(n6128), .A2(n8736), .ZN(n5140) );
  NOR2_X1 U6604 ( .A1(n5134), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6605 ( .A1(n5137), .A2(n4880), .ZN(n5135) );
  MUX2_X1 U6606 ( .A(n5135), .B(P1_IR_REG_31__SCAN_IN), .S(n5136), .Z(n5138)
         );
  NAND2_X1 U6607 ( .A1(n5137), .A2(n5136), .ZN(n5182) );
  NAND2_X1 U6608 ( .A1(n5138), .A2(n5182), .ZN(n6289) );
  INV_X1 U6609 ( .A(n6289), .ZN(n9577) );
  AOI22_X1 U6610 ( .A1(n5399), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4316), .B2(
        n9577), .ZN(n5139) );
  NAND2_X1 U6611 ( .A1(n9704), .A2(n5666), .ZN(n5149) );
  NAND2_X1 U6612 ( .A1(n5024), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6613 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  AND2_X1 U6614 ( .A1(n5169), .A2(n5143), .ZN(n7221) );
  NAND2_X1 U6615 ( .A1(n5683), .A2(n7221), .ZN(n5146) );
  NAND2_X1 U6616 ( .A1(n6217), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6617 ( .A1(n8093), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5144) );
  NAND4_X1 U6618 ( .A1(n5147), .A2(n5146), .A3(n5145), .A4(n5144), .ZN(n9061)
         );
  NAND2_X1 U6619 ( .A1(n9061), .A2(n5549), .ZN(n5148) );
  NAND2_X1 U6620 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  XNOR2_X1 U6621 ( .A(n5150), .B(n5675), .ZN(n5152) );
  AND2_X1 U6622 ( .A1(n9061), .A2(n5622), .ZN(n5151) );
  AOI21_X1 U6623 ( .B1(n9704), .B2(n5549), .A(n5151), .ZN(n5153) );
  NAND2_X1 U6624 ( .A1(n5152), .A2(n5153), .ZN(n5158) );
  INV_X1 U6625 ( .A(n5152), .ZN(n5155) );
  INV_X1 U6626 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6627 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  NAND2_X1 U6628 ( .A1(n5158), .A2(n5156), .ZN(n6729) );
  INV_X1 U6629 ( .A(n6729), .ZN(n5157) );
  MUX2_X1 U6630 ( .A(n6187), .B(n6185), .S(n5393), .Z(n5163) );
  INV_X1 U6631 ( .A(SI_10_), .ZN(n5162) );
  NAND2_X1 U6632 ( .A1(n5163), .A2(n5162), .ZN(n5180) );
  INV_X1 U6633 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6634 ( .A1(n5164), .A2(SI_10_), .ZN(n5165) );
  NAND2_X1 U6635 ( .A1(n6184), .A2(n8736), .ZN(n5168) );
  NAND2_X1 U6636 ( .A1(n5182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6637 ( .A(n5166), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U6638 ( .A1(n5399), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4316), .B2(
        n6578), .ZN(n5167) );
  NAND2_X2 U6639 ( .A1(n5168), .A2(n5167), .ZN(n7262) );
  NAND2_X1 U6640 ( .A1(n7262), .A2(n5666), .ZN(n5176) );
  NAND2_X1 U6641 ( .A1(n5024), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6642 ( .A1(n5169), .A2(n6298), .ZN(n5170) );
  AND2_X1 U6643 ( .A1(n5187), .A2(n5170), .ZN(n7192) );
  NAND2_X1 U6644 ( .A1(n5683), .A2(n7192), .ZN(n5173) );
  NAND2_X1 U6645 ( .A1(n6217), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6646 ( .A1(n8093), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5171) );
  OR2_X1 U6647 ( .A1(n7261), .A2(n5672), .ZN(n5175) );
  NAND2_X1 U6648 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  XNOR2_X1 U6649 ( .A(n5177), .B(n5552), .ZN(n5197) );
  NOR2_X1 U6650 ( .A1(n7261), .A2(n5051), .ZN(n5178) );
  AOI21_X1 U6651 ( .B1(n7262), .B2(n5549), .A(n5178), .ZN(n5198) );
  XNOR2_X1 U6652 ( .A(n5197), .B(n5198), .ZN(n6820) );
  INV_X1 U6653 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5181) );
  MUX2_X1 U6654 ( .A(n5181), .B(n6188), .S(n5393), .Z(n5206) );
  XNOR2_X1 U6655 ( .A(n5206), .B(SI_11_), .ZN(n5205) );
  XNOR2_X1 U6656 ( .A(n5209), .B(n5205), .ZN(n6182) );
  NAND2_X1 U6657 ( .A1(n6182), .A2(n8736), .ZN(n5185) );
  OAI21_X1 U6658 ( .B1(n5182), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5183) );
  XNOR2_X1 U6659 ( .A(n5183), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9591) );
  AOI22_X1 U6660 ( .A1(n5399), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4316), .B2(
        n9591), .ZN(n5184) );
  NAND2_X1 U6661 ( .A1(n7426), .A2(n5666), .ZN(n5194) );
  NAND2_X1 U6662 ( .A1(n8092), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5192) );
  AND2_X1 U6663 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NOR2_X1 U6664 ( .A1(n5218), .A2(n5188), .ZN(n7270) );
  NAND2_X1 U6665 ( .A1(n5683), .A2(n7270), .ZN(n5191) );
  NAND2_X1 U6666 ( .A1(n6217), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6667 ( .A1(n8093), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5189) );
  NAND4_X1 U6668 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n9059)
         );
  NAND2_X1 U6669 ( .A1(n9059), .A2(n5549), .ZN(n5193) );
  NAND2_X1 U6670 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  XNOR2_X1 U6671 ( .A(n5195), .B(n5552), .ZN(n5203) );
  AND2_X1 U6672 ( .A1(n9059), .A2(n5622), .ZN(n5196) );
  AOI21_X1 U6673 ( .B1(n7426), .B2(n5549), .A(n5196), .ZN(n5201) );
  XNOR2_X1 U6674 ( .A(n5203), .B(n5201), .ZN(n6940) );
  INV_X1 U6675 ( .A(n5197), .ZN(n5199) );
  NAND2_X1 U6676 ( .A1(n5199), .A2(n5198), .ZN(n6937) );
  AND2_X1 U6677 ( .A1(n6940), .A2(n6937), .ZN(n5200) );
  INV_X1 U6678 ( .A(n5201), .ZN(n5202) );
  NAND2_X1 U6679 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  NAND2_X1 U6680 ( .A1(n6939), .A2(n5204), .ZN(n7132) );
  INV_X1 U6681 ( .A(n5205), .ZN(n5208) );
  INV_X1 U6682 ( .A(n5206), .ZN(n5207) );
  MUX2_X1 U6683 ( .A(n6231), .B(n6233), .S(n5393), .Z(n5211) );
  INV_X1 U6684 ( .A(SI_12_), .ZN(n5210) );
  NAND2_X1 U6685 ( .A1(n5211), .A2(n5210), .ZN(n5234) );
  INV_X1 U6686 ( .A(n5211), .ZN(n5212) );
  NAND2_X1 U6687 ( .A1(n5212), .A2(SI_12_), .ZN(n5213) );
  NAND2_X1 U6688 ( .A1(n5234), .A2(n5213), .ZN(n5232) );
  XNOR2_X1 U6689 ( .A(n5233), .B(n5232), .ZN(n6230) );
  NAND2_X1 U6690 ( .A1(n6230), .A2(n8736), .ZN(n5217) );
  OR2_X1 U6691 ( .A1(n5214), .A2(n4880), .ZN(n5215) );
  XNOR2_X1 U6692 ( .A(n5215), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6661) );
  AOI22_X1 U6693 ( .A1(n5399), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4316), .B2(
        n6661), .ZN(n5216) );
  NAND2_X1 U6694 ( .A1(n7323), .A2(n5666), .ZN(n5225) );
  NAND2_X1 U6695 ( .A1(n8092), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5223) );
  NOR2_X1 U6696 ( .A1(n5218), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5219) );
  OR2_X1 U6697 ( .A1(n5246), .A2(n5219), .ZN(n7291) );
  INV_X1 U6698 ( .A(n7291), .ZN(n7142) );
  NAND2_X1 U6699 ( .A1(n5683), .A2(n7142), .ZN(n5222) );
  NAND2_X1 U6700 ( .A1(n6217), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6701 ( .A1(n8093), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6702 ( .A1(n7322), .A2(n5672), .ZN(n5224) );
  NAND2_X1 U6703 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  XNOR2_X1 U6704 ( .A(n5226), .B(n5675), .ZN(n5228) );
  NOR2_X1 U6705 ( .A1(n7322), .A2(n5051), .ZN(n5227) );
  AOI21_X1 U6706 ( .B1(n7323), .B2(n5549), .A(n5227), .ZN(n5229) );
  NAND2_X1 U6707 ( .A1(n5228), .A2(n5229), .ZN(n7133) );
  INV_X1 U6708 ( .A(n5228), .ZN(n5231) );
  INV_X1 U6709 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6710 ( .A1(n5231), .A2(n5230), .ZN(n7134) );
  NAND2_X1 U6711 ( .A1(n5235), .A2(n5234), .ZN(n5260) );
  INV_X1 U6712 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5236) );
  MUX2_X1 U6713 ( .A(n6309), .B(n5236), .S(n5393), .Z(n5238) );
  INV_X1 U6714 ( .A(SI_13_), .ZN(n5237) );
  NAND2_X1 U6715 ( .A1(n5238), .A2(n5237), .ZN(n5261) );
  INV_X1 U6716 ( .A(n5238), .ZN(n5239) );
  NAND2_X1 U6717 ( .A1(n5239), .A2(SI_13_), .ZN(n5240) );
  XNOR2_X1 U6718 ( .A(n5260), .B(n5259), .ZN(n6306) );
  NAND2_X1 U6719 ( .A1(n6306), .A2(n8736), .ZN(n5245) );
  NAND2_X1 U6720 ( .A1(n5241), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5242) );
  MUX2_X1 U6721 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5242), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5243) );
  AND2_X1 U6722 ( .A1(n5263), .A2(n5243), .ZN(n6904) );
  AOI22_X1 U6723 ( .A1(n5399), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4316), .B2(
        n6904), .ZN(n5244) );
  NAND2_X1 U6724 ( .A1(n9400), .A2(n5666), .ZN(n5253) );
  NAND2_X1 U6725 ( .A1(n8092), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5251) );
  NOR2_X1 U6726 ( .A1(n5246), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6727 ( .A1(n5269), .A2(n5247), .ZN(n7127) );
  INV_X1 U6728 ( .A(n7127), .ZN(n7416) );
  NAND2_X1 U6729 ( .A1(n5683), .A2(n7416), .ZN(n5250) );
  NAND2_X1 U6730 ( .A1(n8093), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6731 ( .A1(n6217), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5248) );
  NAND4_X1 U6732 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n9057)
         );
  NAND2_X1 U6733 ( .A1(n9057), .A2(n5549), .ZN(n5252) );
  NAND2_X1 U6734 ( .A1(n5253), .A2(n5252), .ZN(n5254) );
  XNOR2_X1 U6735 ( .A(n5254), .B(n5552), .ZN(n7120) );
  NAND2_X1 U6736 ( .A1(n9400), .A2(n5549), .ZN(n5256) );
  NAND2_X1 U6737 ( .A1(n9057), .A2(n5622), .ZN(n5255) );
  NAND2_X1 U6738 ( .A1(n5256), .A2(n5255), .ZN(n7121) );
  NAND2_X1 U6739 ( .A1(n7123), .A2(n7120), .ZN(n5257) );
  MUX2_X1 U6740 ( .A(n6323), .B(n5262), .S(n5393), .Z(n5283) );
  XNOR2_X1 U6741 ( .A(n5283), .B(SI_14_), .ZN(n5280) );
  XNOR2_X1 U6742 ( .A(n5282), .B(n5280), .ZN(n6916) );
  NAND2_X1 U6743 ( .A1(n6916), .A2(n8736), .ZN(n5268) );
  NAND2_X1 U6744 ( .A1(n5263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5265) );
  OR2_X1 U6745 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6746 ( .A1(n5265), .A2(n5264), .ZN(n5291) );
  AOI22_X1 U6747 ( .A1(n5399), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4316), .B2(
        n7210), .ZN(n5267) );
  NAND2_X1 U6748 ( .A1(n7395), .A2(n5549), .ZN(n5276) );
  NAND2_X1 U6749 ( .A1(n8092), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6750 ( .A1(n5269), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5270) );
  AND2_X1 U6751 ( .A1(n5270), .A2(n5298), .ZN(n7336) );
  NAND2_X1 U6752 ( .A1(n5683), .A2(n7336), .ZN(n5273) );
  NAND2_X1 U6753 ( .A1(n6217), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6754 ( .A1(n8093), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5271) );
  NAND4_X1 U6755 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n9056)
         );
  NAND2_X1 U6756 ( .A1(n9056), .A2(n5622), .ZN(n5275) );
  NAND2_X1 U6757 ( .A1(n5276), .A2(n5275), .ZN(n7235) );
  NAND2_X1 U6758 ( .A1(n7395), .A2(n5666), .ZN(n5278) );
  NAND2_X1 U6759 ( .A1(n9056), .A2(n5549), .ZN(n5277) );
  NAND2_X1 U6760 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  XNOR2_X1 U6761 ( .A(n5279), .B(n5552), .ZN(n7234) );
  INV_X1 U6762 ( .A(n5280), .ZN(n5281) );
  INV_X1 U6763 ( .A(n5283), .ZN(n5284) );
  NAND2_X1 U6764 ( .A1(n5284), .A2(SI_14_), .ZN(n5285) );
  MUX2_X1 U6765 ( .A(n6451), .B(n6453), .S(n5393), .Z(n5287) );
  NAND2_X1 U6766 ( .A1(n5287), .A2(n5286), .ZN(n5312) );
  INV_X1 U6767 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U6768 ( .A1(n5288), .A2(SI_15_), .ZN(n5289) );
  NAND2_X1 U6769 ( .A1(n5312), .A2(n5289), .ZN(n5313) );
  XNOR2_X1 U6770 ( .A(n5314), .B(n5313), .ZN(n7063) );
  NAND2_X1 U6771 ( .A1(n7063), .A2(n8736), .ZN(n5296) );
  NAND2_X1 U6772 ( .A1(n5291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5293) );
  XNOR2_X1 U6773 ( .A(n5293), .B(n5292), .ZN(n7359) );
  INV_X1 U6774 ( .A(n7359), .ZN(n5294) );
  AOI22_X1 U6775 ( .A1(n8733), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4316), .B2(
        n5294), .ZN(n5295) );
  NAND2_X2 U6776 ( .A1(n5296), .A2(n5295), .ZN(n9395) );
  NAND2_X1 U6777 ( .A1(n9395), .A2(n5666), .ZN(n5305) );
  NAND2_X1 U6778 ( .A1(n8092), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6779 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  AND2_X1 U6780 ( .A1(n5323), .A2(n5299), .ZN(n7488) );
  NAND2_X1 U6781 ( .A1(n5683), .A2(n7488), .ZN(n5302) );
  NAND2_X1 U6782 ( .A1(n6217), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6783 ( .A1(n8093), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5300) );
  NAND4_X1 U6784 ( .A1(n5303), .A2(n5302), .A3(n5301), .A4(n5300), .ZN(n9055)
         );
  NAND2_X1 U6785 ( .A1(n9055), .A2(n5549), .ZN(n5304) );
  NAND2_X1 U6786 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  XNOR2_X1 U6787 ( .A(n5306), .B(n5675), .ZN(n7344) );
  AND2_X1 U6788 ( .A1(n9055), .A2(n5622), .ZN(n5307) );
  AOI21_X1 U6789 ( .B1(n9395), .B2(n5549), .A(n5307), .ZN(n5308) );
  INV_X1 U6790 ( .A(n7344), .ZN(n5309) );
  INV_X1 U6791 ( .A(n5308), .ZN(n7343) );
  NAND2_X1 U6792 ( .A1(n5309), .A2(n7343), .ZN(n5310) );
  NAND2_X1 U6793 ( .A1(n5311), .A2(n5310), .ZN(n7500) );
  INV_X1 U6794 ( .A(n7500), .ZN(n5337) );
  MUX2_X1 U6795 ( .A(n10103), .B(n10072), .S(n5393), .Z(n5316) );
  NAND2_X1 U6796 ( .A1(n5316), .A2(n5315), .ZN(n5341) );
  INV_X1 U6797 ( .A(n5316), .ZN(n5317) );
  NAND2_X1 U6798 ( .A1(n5317), .A2(SI_16_), .ZN(n5318) );
  XNOR2_X1 U6799 ( .A(n5340), .B(n5339), .ZN(n7067) );
  NAND2_X1 U6800 ( .A1(n7067), .A2(n8736), .ZN(n5321) );
  NAND2_X1 U6801 ( .A1(n5343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5319) );
  XNOR2_X1 U6802 ( .A(n5319), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9100) );
  AOI22_X1 U6803 ( .A1(n5399), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4316), .B2(
        n9100), .ZN(n5320) );
  NAND2_X1 U6804 ( .A1(n7623), .A2(n5666), .ZN(n5330) );
  NAND2_X1 U6805 ( .A1(n8092), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5328) );
  AND2_X1 U6806 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  NOR2_X1 U6807 ( .A1(n5349), .A2(n5324), .ZN(n7503) );
  NAND2_X1 U6808 ( .A1(n5683), .A2(n7503), .ZN(n5327) );
  NAND2_X1 U6809 ( .A1(n6217), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6810 ( .A1(n8093), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5325) );
  OR2_X1 U6811 ( .A1(n7492), .A2(n5672), .ZN(n5329) );
  NAND2_X1 U6812 ( .A1(n5330), .A2(n5329), .ZN(n5331) );
  XNOR2_X1 U6813 ( .A(n5331), .B(n5675), .ZN(n5334) );
  NOR2_X1 U6814 ( .A1(n7492), .A2(n5051), .ZN(n5332) );
  AOI21_X1 U6815 ( .B1(n7623), .B2(n5549), .A(n5332), .ZN(n5333) );
  NAND2_X1 U6816 ( .A1(n5334), .A2(n5333), .ZN(n5338) );
  OR2_X1 U6817 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  NAND2_X1 U6818 ( .A1(n5338), .A2(n5335), .ZN(n7499) );
  NAND2_X1 U6819 ( .A1(n7497), .A2(n5338), .ZN(n7612) );
  MUX2_X1 U6820 ( .A(n6573), .B(n5342), .S(n5393), .Z(n5365) );
  XNOR2_X1 U6821 ( .A(n5365), .B(SI_17_), .ZN(n5364) );
  XNOR2_X1 U6822 ( .A(n5369), .B(n5364), .ZN(n7304) );
  NAND2_X1 U6823 ( .A1(n7304), .A2(n8736), .ZN(n5348) );
  OAI21_X1 U6824 ( .B1(n5343), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5345) );
  OR2_X1 U6825 ( .A1(n5345), .A2(n5344), .ZN(n5346) );
  NAND2_X1 U6826 ( .A1(n5345), .A2(n5344), .ZN(n5370) );
  AOI22_X1 U6827 ( .A1(n5399), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4316), .B2(
        n9113), .ZN(n5347) );
  NAND2_X1 U6828 ( .A1(n9391), .A2(n5666), .ZN(n5356) );
  NAND2_X1 U6829 ( .A1(n8092), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5354) );
  NOR2_X1 U6830 ( .A1(n5349), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6831 ( .A1(n5683), .A2(n4859), .ZN(n5353) );
  NAND2_X1 U6832 ( .A1(n6217), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6833 ( .A1(n8093), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5351) );
  NAND4_X1 U6834 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n9053)
         );
  NAND2_X1 U6835 ( .A1(n9053), .A2(n5549), .ZN(n5355) );
  NAND2_X1 U6836 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  XNOR2_X1 U6837 ( .A(n5357), .B(n5552), .ZN(n5360) );
  NAND2_X1 U6838 ( .A1(n9391), .A2(n5549), .ZN(n5359) );
  NAND2_X1 U6839 ( .A1(n9053), .A2(n5622), .ZN(n5358) );
  NAND2_X1 U6840 ( .A1(n5359), .A2(n5358), .ZN(n5361) );
  NAND2_X1 U6841 ( .A1(n5360), .A2(n5361), .ZN(n7613) );
  NAND2_X1 U6842 ( .A1(n7612), .A2(n7613), .ZN(n7611) );
  INV_X1 U6843 ( .A(n5360), .ZN(n5363) );
  INV_X1 U6844 ( .A(n5361), .ZN(n5362) );
  NAND2_X1 U6845 ( .A1(n5363), .A2(n5362), .ZN(n7614) );
  INV_X1 U6846 ( .A(n5364), .ZN(n5368) );
  INV_X1 U6847 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U6848 ( .A1(n5366), .A2(SI_17_), .ZN(n5367) );
  MUX2_X1 U6849 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5393), .Z(n5392) );
  XNOR2_X1 U6850 ( .A(n5392), .B(SI_18_), .ZN(n5389) );
  XNOR2_X1 U6851 ( .A(n5391), .B(n5389), .ZN(n7436) );
  NAND2_X1 U6852 ( .A1(n7436), .A2(n8736), .ZN(n5373) );
  NAND2_X1 U6853 ( .A1(n5370), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U6854 ( .A(n5371), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9126) );
  AOI22_X1 U6855 ( .A1(n5399), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4316), .B2(
        n9126), .ZN(n5372) );
  NAND2_X1 U6856 ( .A1(n9386), .A2(n5666), .ZN(n5381) );
  OR2_X1 U6857 ( .A1(n5374), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5375) );
  AND2_X1 U6858 ( .A1(n5375), .A2(n5403), .ZN(n8727) );
  NAND2_X1 U6859 ( .A1(n8727), .A2(n5683), .ZN(n5379) );
  NAND2_X1 U6860 ( .A1(n8092), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6861 ( .A1(n8093), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6862 ( .A1(n6217), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5376) );
  OR2_X1 U6863 ( .A1(n7633), .A2(n5672), .ZN(n5380) );
  NAND2_X1 U6864 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  XNOR2_X1 U6865 ( .A(n5382), .B(n5675), .ZN(n5386) );
  NAND2_X1 U6866 ( .A1(n9386), .A2(n5549), .ZN(n5384) );
  OR2_X1 U6867 ( .A1(n7633), .A2(n5051), .ZN(n5383) );
  NAND2_X1 U6868 ( .A1(n5384), .A2(n5383), .ZN(n8713) );
  NAND2_X1 U6869 ( .A1(n8714), .A2(n8713), .ZN(n8719) );
  INV_X1 U6870 ( .A(n5386), .ZN(n5387) );
  INV_X1 U6871 ( .A(n5389), .ZN(n5390) );
  MUX2_X1 U6872 ( .A(n9961), .B(n5394), .S(n5393), .Z(n5395) );
  NAND2_X1 U6873 ( .A1(n5395), .A2(n9958), .ZN(n5414) );
  INV_X1 U6874 ( .A(n5395), .ZN(n5396) );
  NAND2_X1 U6875 ( .A1(n5396), .A2(SI_19_), .ZN(n5397) );
  NAND2_X1 U6876 ( .A1(n5414), .A2(n5397), .ZN(n5415) );
  NAND2_X1 U6877 ( .A1(n7514), .A2(n8736), .ZN(n5401) );
  AOI22_X1 U6878 ( .A1(n5399), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4316), .B2(
        n5398), .ZN(n5400) );
  NAND2_X1 U6879 ( .A1(n9381), .A2(n5666), .ZN(n5410) );
  NAND2_X1 U6880 ( .A1(n8092), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5408) );
  INV_X1 U6881 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5404) );
  AOI21_X1 U6882 ( .B1(n5404), .B2(n5403), .A(n5423), .ZN(n9291) );
  NAND2_X1 U6883 ( .A1(n5683), .A2(n9291), .ZN(n5407) );
  NAND2_X1 U6884 ( .A1(n6217), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6885 ( .A1(n8093), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5405) );
  NAND4_X1 U6886 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n9279)
         );
  NAND2_X1 U6887 ( .A1(n9279), .A2(n5549), .ZN(n5409) );
  NAND2_X1 U6888 ( .A1(n5410), .A2(n5409), .ZN(n5411) );
  XNOR2_X1 U6889 ( .A(n5411), .B(n5552), .ZN(n8660) );
  NAND2_X1 U6890 ( .A1(n9381), .A2(n5549), .ZN(n5413) );
  NAND2_X1 U6891 ( .A1(n9279), .A2(n5622), .ZN(n5412) );
  NAND2_X1 U6892 ( .A1(n5413), .A2(n5412), .ZN(n8661) );
  MUX2_X1 U6893 ( .A(n6898), .B(n6935), .S(n7775), .Z(n5418) );
  INV_X1 U6894 ( .A(SI_20_), .ZN(n5417) );
  NAND2_X1 U6895 ( .A1(n5418), .A2(n5417), .ZN(n5442) );
  INV_X1 U6896 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U6897 ( .A1(n5419), .A2(SI_20_), .ZN(n5420) );
  XNOR2_X1 U6898 ( .A(n5441), .B(n5440), .ZN(n7555) );
  NAND2_X1 U6899 ( .A1(n7555), .A2(n8736), .ZN(n5422) );
  NAND2_X1 U6900 ( .A1(n8733), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6901 ( .A1(n9375), .A2(n5666), .ZN(n5431) );
  NAND2_X1 U6902 ( .A1(n8092), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5429) );
  INV_X1 U6903 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8693) );
  INV_X1 U6904 ( .A(n5446), .ZN(n5424) );
  AOI21_X1 U6905 ( .B1(n8693), .B2(n5425), .A(n5424), .ZN(n9274) );
  NAND2_X1 U6906 ( .A1(n5683), .A2(n9274), .ZN(n5428) );
  NAND2_X1 U6907 ( .A1(n8093), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6908 ( .A1(n6217), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5426) );
  NAND4_X1 U6909 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n9301)
         );
  NAND2_X1 U6910 ( .A1(n9301), .A2(n5549), .ZN(n5430) );
  NAND2_X1 U6911 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  XNOR2_X1 U6912 ( .A(n5432), .B(n5675), .ZN(n5434) );
  AND2_X1 U6913 ( .A1(n9301), .A2(n5622), .ZN(n5433) );
  AOI21_X1 U6914 ( .B1(n9375), .B2(n5549), .A(n5433), .ZN(n5435) );
  NAND2_X1 U6915 ( .A1(n5434), .A2(n5435), .ZN(n5439) );
  INV_X1 U6916 ( .A(n5434), .ZN(n5437) );
  INV_X1 U6917 ( .A(n5435), .ZN(n5436) );
  NAND2_X1 U6918 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  NAND2_X1 U6919 ( .A1(n5439), .A2(n5438), .ZN(n8691) );
  NAND2_X1 U6920 ( .A1(n5441), .A2(n5440), .ZN(n5443) );
  MUX2_X1 U6921 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7775), .Z(n5461) );
  XNOR2_X1 U6922 ( .A(n5461), .B(n10054), .ZN(n5460) );
  XNOR2_X1 U6923 ( .A(n5459), .B(n5460), .ZN(n7590) );
  NAND2_X1 U6924 ( .A1(n7590), .A2(n8736), .ZN(n5445) );
  NAND2_X1 U6925 ( .A1(n8733), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6926 ( .A1(n9264), .A2(n5666), .ZN(n5452) );
  NAND2_X1 U6927 ( .A1(n6217), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6928 ( .A1(n8092), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5449) );
  AOI21_X1 U6929 ( .B1(n5446), .B2(n8675), .A(n5469), .ZN(n9267) );
  NAND2_X1 U6930 ( .A1(n5683), .A2(n9267), .ZN(n5448) );
  NAND2_X1 U6931 ( .A1(n8093), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6932 ( .A1(n9280), .A2(n5549), .ZN(n5451) );
  NAND2_X1 U6933 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  XNOR2_X1 U6934 ( .A(n5453), .B(n5552), .ZN(n5455) );
  NOR2_X1 U6935 ( .A1(n8703), .A2(n5051), .ZN(n5454) );
  AOI21_X1 U6936 ( .B1(n9264), .B2(n5549), .A(n5454), .ZN(n5456) );
  XNOR2_X1 U6937 ( .A(n5455), .B(n5456), .ZN(n8672) );
  INV_X1 U6938 ( .A(n5455), .ZN(n5457) );
  NAND2_X1 U6939 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U6940 ( .A1(n8670), .A2(n5458), .ZN(n5480) );
  NAND2_X1 U6941 ( .A1(n5461), .A2(SI_21_), .ZN(n5462) );
  MUX2_X1 U6942 ( .A(n8017), .B(n7119), .S(n7775), .Z(n5464) );
  INV_X1 U6943 ( .A(SI_22_), .ZN(n5463) );
  NAND2_X1 U6944 ( .A1(n5464), .A2(n5463), .ZN(n5482) );
  INV_X1 U6945 ( .A(n5464), .ZN(n5465) );
  NAND2_X1 U6946 ( .A1(n5465), .A2(SI_22_), .ZN(n5466) );
  NAND2_X1 U6947 ( .A1(n5482), .A2(n5466), .ZN(n5483) );
  NAND2_X1 U6948 ( .A1(n7678), .A2(n8736), .ZN(n5468) );
  NAND2_X1 U6949 ( .A1(n8733), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U6950 ( .A1(n8092), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5474) );
  NOR2_X1 U6951 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5469), .ZN(n5470) );
  NOR2_X1 U6952 ( .A1(n5493), .A2(n5470), .ZN(n9249) );
  NAND2_X1 U6953 ( .A1(n5683), .A2(n9249), .ZN(n5473) );
  NAND2_X1 U6954 ( .A1(n6217), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6955 ( .A1(n8093), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5471) );
  NAND4_X1 U6956 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n9260)
         );
  AND2_X1 U6957 ( .A1(n9260), .A2(n5622), .ZN(n5475) );
  AOI21_X1 U6958 ( .B1(n9364), .B2(n5549), .A(n5475), .ZN(n5479) );
  OR2_X2 U6959 ( .A1(n5480), .A2(n5479), .ZN(n8700) );
  NAND2_X1 U6960 ( .A1(n9364), .A2(n5666), .ZN(n5477) );
  NAND2_X1 U6961 ( .A1(n9260), .A2(n5549), .ZN(n5476) );
  NAND2_X1 U6962 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  XNOR2_X1 U6963 ( .A(n5478), .B(n5675), .ZN(n8701) );
  NAND2_X1 U6964 ( .A1(n5480), .A2(n5479), .ZN(n8699) );
  INV_X1 U6965 ( .A(n8699), .ZN(n5481) );
  INV_X1 U6966 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5486) );
  INV_X1 U6967 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5485) );
  MUX2_X1 U6968 ( .A(n5486), .B(n5485), .S(n7775), .Z(n5488) );
  INV_X1 U6969 ( .A(SI_23_), .ZN(n5487) );
  NAND2_X1 U6970 ( .A1(n5488), .A2(n5487), .ZN(n5509) );
  INV_X1 U6971 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U6972 ( .A1(n5489), .A2(SI_23_), .ZN(n5490) );
  XNOR2_X1 U6973 ( .A(n5508), .B(n5507), .ZN(n7683) );
  NAND2_X1 U6974 ( .A1(n7683), .A2(n8736), .ZN(n5492) );
  NAND2_X1 U6975 ( .A1(n5399), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6976 ( .A1(n9358), .A2(n5666), .ZN(n5500) );
  NAND2_X1 U6977 ( .A1(n8092), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5498) );
  NOR2_X1 U6978 ( .A1(n5493), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5494) );
  NOR2_X1 U6979 ( .A1(n5515), .A2(n5494), .ZN(n9226) );
  NAND2_X1 U6980 ( .A1(n5683), .A2(n9226), .ZN(n5497) );
  NAND2_X1 U6981 ( .A1(n6217), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6982 ( .A1(n8093), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5495) );
  NAND4_X1 U6983 ( .A1(n5498), .A2(n5497), .A3(n5496), .A4(n5495), .ZN(n9246)
         );
  NAND2_X1 U6984 ( .A1(n9246), .A2(n5549), .ZN(n5499) );
  NAND2_X1 U6985 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  XNOR2_X1 U6986 ( .A(n5501), .B(n5552), .ZN(n5504) );
  AND2_X1 U6987 ( .A1(n9246), .A2(n5622), .ZN(n5502) );
  AOI21_X1 U6988 ( .B1(n9358), .B2(n5549), .A(n5502), .ZN(n8651) );
  NAND2_X1 U6989 ( .A1(n8652), .A2(n8651), .ZN(n8649) );
  INV_X1 U6990 ( .A(n5503), .ZN(n5506) );
  INV_X1 U6991 ( .A(n5504), .ZN(n5505) );
  NAND2_X1 U6992 ( .A1(n5508), .A2(n5507), .ZN(n5510) );
  MUX2_X1 U6993 ( .A(n7319), .B(n10071), .S(n7775), .Z(n5533) );
  XNOR2_X1 U6994 ( .A(n5533), .B(SI_24_), .ZN(n5532) );
  XNOR2_X1 U6995 ( .A(n5537), .B(n5532), .ZN(n7697) );
  NAND2_X1 U6996 ( .A1(n7697), .A2(n8736), .ZN(n5512) );
  NAND2_X1 U6997 ( .A1(n8733), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U6998 ( .A1(n9354), .A2(n5666), .ZN(n5522) );
  NAND2_X1 U6999 ( .A1(n8092), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5520) );
  INV_X1 U7000 ( .A(n5515), .ZN(n5514) );
  INV_X1 U7001 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7002 ( .A1(n5514), .A2(n5513), .ZN(n5516) );
  AND2_X1 U7003 ( .A1(n5516), .A2(n5544), .ZN(n9211) );
  NAND2_X1 U7004 ( .A1(n5683), .A2(n9211), .ZN(n5519) );
  NAND2_X1 U7005 ( .A1(n8093), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7006 ( .A1(n6217), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5517) );
  NAND4_X1 U7007 ( .A1(n5520), .A2(n5519), .A3(n5518), .A4(n5517), .ZN(n9202)
         );
  NAND2_X1 U7008 ( .A1(n9202), .A2(n5549), .ZN(n5521) );
  NAND2_X1 U7009 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  XNOR2_X1 U7010 ( .A(n5523), .B(n5675), .ZN(n5525) );
  AND2_X1 U7011 ( .A1(n9202), .A2(n5622), .ZN(n5524) );
  AOI21_X1 U7012 ( .B1(n9354), .B2(n5549), .A(n5524), .ZN(n5526) );
  NAND2_X1 U7013 ( .A1(n5525), .A2(n5526), .ZN(n5530) );
  INV_X1 U7014 ( .A(n5525), .ZN(n5528) );
  INV_X1 U7015 ( .A(n5526), .ZN(n5527) );
  NAND2_X1 U7016 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  NAND2_X1 U7017 ( .A1(n5530), .A2(n5529), .ZN(n8681) );
  INV_X1 U7018 ( .A(n5530), .ZN(n5531) );
  INV_X1 U7019 ( .A(n5532), .ZN(n5536) );
  INV_X1 U7020 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7021 ( .A1(n5534), .A2(SI_24_), .ZN(n5535) );
  MUX2_X1 U7022 ( .A(n7482), .B(n7480), .S(n7775), .Z(n5539) );
  INV_X1 U7023 ( .A(SI_25_), .ZN(n5538) );
  NAND2_X1 U7024 ( .A1(n5539), .A2(n5538), .ZN(n5609) );
  INV_X1 U7025 ( .A(n5539), .ZN(n5540) );
  NAND2_X1 U7026 ( .A1(n5540), .A2(SI_25_), .ZN(n5541) );
  NAND2_X1 U7027 ( .A1(n5609), .A2(n5541), .ZN(n5610) );
  XNOR2_X1 U7028 ( .A(n5611), .B(n5610), .ZN(n7709) );
  NAND2_X1 U7029 ( .A1(n7709), .A2(n8736), .ZN(n5543) );
  NAND2_X1 U7030 ( .A1(n8733), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7031 ( .A1(n8092), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7032 ( .A1(n6217), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5547) );
  INV_X1 U7033 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5599) );
  AOI21_X1 U7034 ( .B1(n5544), .B2(n5599), .A(n5593), .ZN(n9197) );
  NAND2_X1 U7035 ( .A1(n5683), .A2(n9197), .ZN(n5546) );
  NAND2_X1 U7036 ( .A1(n8093), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5545) );
  AOI22_X1 U7037 ( .A1(n9348), .A2(n5549), .B1(n5622), .B2(n9189), .ZN(n5624)
         );
  NAND2_X1 U7038 ( .A1(n9348), .A2(n5666), .ZN(n5551) );
  NAND2_X1 U7039 ( .A1(n9189), .A2(n5549), .ZN(n5550) );
  NAND2_X1 U7040 ( .A1(n5551), .A2(n5550), .ZN(n5553) );
  XNOR2_X1 U7041 ( .A(n5553), .B(n5552), .ZN(n5626) );
  XOR2_X1 U7042 ( .A(n5624), .B(n5626), .Z(n5628) );
  NOR2_X1 U7043 ( .A1(n5629), .A2(n5628), .ZN(n5703) );
  INV_X1 U7044 ( .A(n5554), .ZN(n5568) );
  NAND3_X1 U7045 ( .A1(n7479), .A2(P1_B_REG_SCAN_IN), .A3(n7318), .ZN(n5555)
         );
  OAI21_X1 U7046 ( .B1(P1_B_REG_SCAN_IN), .B2(n7318), .A(n5555), .ZN(n5556) );
  INV_X1 U7047 ( .A(n7318), .ZN(n5557) );
  NOR4_X1 U7048 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5561) );
  NOR4_X1 U7049 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5560) );
  NOR4_X1 U7050 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5559) );
  NOR4_X1 U7051 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5558) );
  AND4_X1 U7052 ( .A1(n5561), .A2(n5560), .A3(n5559), .A4(n5558), .ZN(n5567)
         );
  NOR2_X1 U7053 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n5565) );
  NOR4_X1 U7054 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5564) );
  NOR4_X1 U7055 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5563) );
  NOR4_X1 U7056 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5562) );
  AND4_X1 U7057 ( .A1(n5565), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n5566)
         );
  NAND2_X1 U7058 ( .A1(n5567), .A2(n5566), .ZN(n6242) );
  INV_X1 U7059 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6112) );
  NOR2_X1 U7060 ( .A1(n6242), .A2(n6112), .ZN(n5569) );
  NAND2_X1 U7061 ( .A1(n5568), .A2(n7479), .ZN(n6240) );
  OAI21_X1 U7062 ( .B1(n6241), .B2(n5569), .A(n6240), .ZN(n6479) );
  OR2_X1 U7063 ( .A1(n7112), .A2(n6479), .ZN(n5588) );
  NAND4_X1 U7064 ( .A1(n5573), .A2(n5572), .A3(n5571), .A4(n5570), .ZN(n5574)
         );
  OAI21_X1 U7065 ( .B1(n5575), .B2(n5574), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5577) );
  AND2_X1 U7066 ( .A1(n7229), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5578) );
  INV_X1 U7067 ( .A(n6251), .ZN(n6249) );
  INV_X1 U7068 ( .A(n9033), .ZN(n5583) );
  NOR2_X1 U7069 ( .A1(n9677), .A2(n6504), .ZN(n5581) );
  NAND2_X1 U7070 ( .A1(n5588), .A2(n9705), .ZN(n6213) );
  NAND2_X1 U7071 ( .A1(n6213), .A2(n5580), .ZN(n5584) );
  OR2_X1 U7072 ( .A1(n5580), .A2(n5583), .ZN(n6248) );
  NAND2_X1 U7073 ( .A1(n5584), .A2(n6248), .ZN(n5586) );
  AND2_X1 U7074 ( .A1(n5723), .A2(n7229), .ZN(n5585) );
  AOI21_X1 U7075 ( .B1(n5586), .B2(n5585), .A(P1_U3084), .ZN(n5589) );
  OR2_X1 U7076 ( .A1(n6251), .A2(n8912), .ZN(n5602) );
  AOI21_X1 U7077 ( .B1(n5602), .B2(n6248), .A(n6212), .ZN(n5587) );
  AND2_X1 U7078 ( .A1(n5588), .A2(n5587), .ZN(n6210) );
  NOR2_X1 U7079 ( .A1(n6248), .A2(n5590), .ZN(n5591) );
  NAND2_X1 U7080 ( .A1(n5603), .A2(n5591), .ZN(n8723) );
  NOR2_X1 U7081 ( .A1(n8723), .A2(n9229), .ZN(n5601) );
  INV_X1 U7082 ( .A(n5590), .ZN(n9512) );
  NOR2_X1 U7083 ( .A1(n6248), .A2(n9512), .ZN(n5592) );
  NAND2_X1 U7084 ( .A1(n8092), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7085 ( .A1(n5593), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5640) );
  OAI21_X1 U7086 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5593), .A(n5640), .ZN(
        n5594) );
  INV_X1 U7087 ( .A(n5594), .ZN(n9183) );
  NAND2_X1 U7088 ( .A1(n5683), .A2(n9183), .ZN(n5597) );
  NAND2_X1 U7089 ( .A1(n6217), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7090 ( .A1(n8093), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5595) );
  NAND4_X1 U7091 ( .A1(n5598), .A2(n5597), .A3(n5596), .A4(n5595), .ZN(n9203)
         );
  OAI22_X1 U7092 ( .A1(n8706), .A2(n10115), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5599), .ZN(n5600) );
  AOI211_X1 U7093 ( .C1(n9197), .C2(n8726), .A(n5601), .B(n5600), .ZN(n5607)
         );
  NAND2_X1 U7094 ( .A1(n5603), .A2(n6482), .ZN(n5605) );
  OR2_X1 U7095 ( .A1(n6212), .A2(n5579), .ZN(n5604) );
  NAND2_X1 U7096 ( .A1(n9348), .A2(n8709), .ZN(n5606) );
  NAND3_X1 U7097 ( .A1(n5608), .A2(n5607), .A3(n5606), .ZN(P1_U3223) );
  INV_X1 U7098 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10116) );
  INV_X1 U7099 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5612) );
  MUX2_X1 U7100 ( .A(n10116), .B(n5612), .S(n7775), .Z(n5614) );
  INV_X1 U7101 ( .A(SI_26_), .ZN(n5613) );
  NAND2_X1 U7102 ( .A1(n5614), .A2(n5613), .ZN(n5632) );
  INV_X1 U7103 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7104 ( .A1(n5615), .A2(SI_26_), .ZN(n5616) );
  XNOR2_X1 U7105 ( .A(n5631), .B(n5630), .ZN(n7721) );
  NAND2_X1 U7106 ( .A1(n7721), .A2(n8736), .ZN(n5618) );
  NAND2_X1 U7107 ( .A1(n5399), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7108 ( .A1(n9343), .A2(n5666), .ZN(n5620) );
  NAND2_X1 U7109 ( .A1(n9203), .A2(n5549), .ZN(n5619) );
  NAND2_X1 U7110 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  XNOR2_X1 U7111 ( .A(n5621), .B(n5675), .ZN(n5652) );
  AND2_X1 U7112 ( .A1(n9203), .A2(n5622), .ZN(n5623) );
  AOI21_X1 U7113 ( .B1(n9343), .B2(n5549), .A(n5623), .ZN(n5653) );
  XNOR2_X1 U7114 ( .A(n5652), .B(n5653), .ZN(n5701) );
  INV_X1 U7115 ( .A(n5624), .ZN(n5625) );
  NOR2_X1 U7116 ( .A1(n5626), .A2(n5625), .ZN(n5702) );
  INV_X1 U7117 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7569) );
  INV_X1 U7118 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5633) );
  MUX2_X1 U7119 ( .A(n7569), .B(n5633), .S(n7775), .Z(n5635) );
  INV_X1 U7120 ( .A(SI_27_), .ZN(n5634) );
  NAND2_X1 U7121 ( .A1(n5635), .A2(n5634), .ZN(n5660) );
  INV_X1 U7122 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7123 ( .A1(n5636), .A2(SI_27_), .ZN(n5637) );
  XNOR2_X1 U7124 ( .A(n5659), .B(n5658), .ZN(n7733) );
  NAND2_X1 U7125 ( .A1(n7733), .A2(n8736), .ZN(n5639) );
  NAND2_X1 U7126 ( .A1(n5399), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7127 ( .A1(n9339), .A2(n5666), .ZN(n5646) );
  NAND2_X1 U7128 ( .A1(n6217), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7129 ( .A1(n8092), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5643) );
  INV_X1 U7130 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5717) );
  AOI21_X1 U7131 ( .B1(n5717), .B2(n5640), .A(n5667), .ZN(n9170) );
  NAND2_X1 U7132 ( .A1(n5683), .A2(n9170), .ZN(n5642) );
  NAND2_X1 U7133 ( .A1(n8093), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7134 ( .A1(n9190), .A2(n5549), .ZN(n5645) );
  NAND2_X1 U7135 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  XNOR2_X1 U7136 ( .A(n5647), .B(n5675), .ZN(n5650) );
  NOR2_X1 U7137 ( .A1(n8079), .A2(n5051), .ZN(n5648) );
  AOI21_X1 U7138 ( .B1(n9339), .B2(n5549), .A(n5648), .ZN(n5649) );
  NAND2_X1 U7139 ( .A1(n5650), .A2(n5649), .ZN(n5692) );
  OAI21_X1 U7140 ( .B1(n5650), .B2(n5649), .A(n5692), .ZN(n5713) );
  INV_X1 U7141 ( .A(n5713), .ZN(n5651) );
  INV_X1 U7142 ( .A(n5652), .ZN(n5655) );
  INV_X1 U7143 ( .A(n5653), .ZN(n5654) );
  INV_X1 U7144 ( .A(n5712), .ZN(n5656) );
  NAND2_X1 U7145 ( .A1(n5659), .A2(n5658), .ZN(n5661) );
  INV_X1 U7146 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5663) );
  INV_X1 U7147 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5662) );
  MUX2_X1 U7148 ( .A(n5663), .B(n5662), .S(n7775), .Z(n7655) );
  XNOR2_X1 U7149 ( .A(n7655), .B(SI_28_), .ZN(n7652) );
  NAND2_X1 U7150 ( .A1(n8643), .A2(n8736), .ZN(n5665) );
  NAND2_X1 U7151 ( .A1(n8733), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7152 ( .A1(n9333), .A2(n5666), .ZN(n5674) );
  NAND2_X1 U7153 ( .A1(n8092), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7154 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n5667), .ZN(n5682) );
  OAI21_X1 U7155 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n5667), .A(n5682), .ZN(
        n5691) );
  INV_X1 U7156 ( .A(n5691), .ZN(n9154) );
  NAND2_X1 U7157 ( .A1(n5683), .A2(n9154), .ZN(n5670) );
  NAND2_X1 U7158 ( .A1(n6217), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7159 ( .A1(n8093), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5668) );
  OR2_X1 U7160 ( .A1(n9173), .A2(n5672), .ZN(n5673) );
  NAND2_X1 U7161 ( .A1(n5674), .A2(n5673), .ZN(n5676) );
  XNOR2_X1 U7162 ( .A(n5676), .B(n5675), .ZN(n5679) );
  NAND2_X1 U7163 ( .A1(n9333), .A2(n5549), .ZN(n5677) );
  OAI21_X1 U7164 ( .B1(n9173), .B2(n5051), .A(n5677), .ZN(n5678) );
  XNOR2_X1 U7165 ( .A(n5679), .B(n5678), .ZN(n5681) );
  INV_X1 U7166 ( .A(n5681), .ZN(n5693) );
  NAND2_X1 U7167 ( .A1(n5680), .A2(n4377), .ZN(n5700) );
  AND2_X1 U7168 ( .A1(n5681), .A2(n8683), .ZN(n5698) );
  INV_X1 U7169 ( .A(n8726), .ZN(n7128) );
  NAND2_X1 U7170 ( .A1(n8092), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5687) );
  INV_X1 U7171 ( .A(n5682), .ZN(n8083) );
  NAND2_X1 U7172 ( .A1(n5683), .A2(n8083), .ZN(n5686) );
  NAND2_X1 U7173 ( .A1(n6217), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7174 ( .A1(n8093), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5684) );
  INV_X1 U7175 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5688) );
  OAI22_X1 U7176 ( .A1(n8706), .A2(n8860), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5688), .ZN(n5689) );
  AOI21_X1 U7177 ( .B1(n8664), .B2(n9190), .A(n5689), .ZN(n5690) );
  OAI21_X1 U7178 ( .B1(n7128), .B2(n5691), .A(n5690), .ZN(n5695) );
  NOR3_X1 U7179 ( .A1(n5693), .A2(n8716), .A3(n5692), .ZN(n5694) );
  AOI211_X1 U7180 ( .C1(n9333), .C2(n8709), .A(n5695), .B(n5694), .ZN(n5696)
         );
  INV_X1 U7181 ( .A(n5696), .ZN(n5697) );
  NAND2_X1 U7182 ( .A1(n5700), .A2(n5699), .ZN(P1_U3218) );
  AND2_X1 U7183 ( .A1(n5714), .A2(n8683), .ZN(n5704) );
  NAND2_X1 U7184 ( .A1(n5705), .A2(n5704), .ZN(n5711) );
  AOI22_X1 U7185 ( .A1(n8664), .A2(n9189), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n5706) );
  OAI21_X1 U7186 ( .B1(n8079), .B2(n8706), .A(n5706), .ZN(n5707) );
  AOI21_X1 U7187 ( .B1(n9183), .B2(n8726), .A(n5707), .ZN(n5708) );
  INV_X1 U7188 ( .A(n5709), .ZN(n5710) );
  NAND2_X1 U7189 ( .A1(n5711), .A2(n5710), .ZN(P1_U3238) );
  NOR2_X1 U7190 ( .A1(n8706), .A2(n9173), .ZN(n5719) );
  OAI22_X1 U7191 ( .A1(n8723), .A2(n10115), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5717), .ZN(n5718) );
  AOI211_X1 U7192 ( .C1(n9170), .C2(n8726), .A(n5719), .B(n5718), .ZN(n5720)
         );
  NAND3_X1 U7193 ( .A1(n5721), .A2(n5720), .A3(n4378), .ZN(P1_U3212) );
  INV_X1 U7194 ( .A(n7229), .ZN(n5722) );
  NAND2_X1 U7195 ( .A1(n5723), .A2(n5580), .ZN(n5724) );
  NAND2_X1 U7196 ( .A1(n5724), .A2(n7229), .ZN(n6162) );
  NAND2_X1 U7197 ( .A1(n5725), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U7198 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5729) );
  AND2_X2 U7199 ( .A1(n5806), .A2(n4630), .ZN(n5822) );
  NAND2_X1 U7200 ( .A1(n5735), .A2(n4856), .ZN(n5788) );
  NAND2_X1 U7201 ( .A1(n5787), .A2(n5786), .ZN(n5736) );
  NAND2_X1 U7202 ( .A1(n5755), .A2(n5754), .ZN(n5737) );
  NOR2_X1 U7203 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5743) );
  NOR2_X1 U7204 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5742) );
  NOR2_X1 U7205 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5741) );
  NAND2_X1 U7206 ( .A1(n5752), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5746) );
  MUX2_X1 U7207 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5746), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5747) );
  NAND2_X1 U7208 ( .A1(n5749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5751) );
  MUX2_X1 U7209 ( .A(n5751), .B(P2_IR_REG_31__SCAN_IN), .S(n5750), .Z(n5753)
         );
  NAND2_X1 U7210 ( .A1(n5753), .A2(n5752), .ZN(n7484) );
  INV_X1 U7211 ( .A(n6261), .ZN(n5756) );
  XNOR2_X1 U7212 ( .A(n5755), .B(n5754), .ZN(n6124) );
  NAND2_X1 U7213 ( .A1(n5912), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7214 ( .A1(n7764), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7215 ( .A1(n5816), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7216 ( .A1(n5800), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7217 ( .A1(n4914), .A2(SI_0_), .ZN(n5773) );
  INV_X1 U7218 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7219 ( .A1(n5773), .A2(n5772), .ZN(n5775) );
  AND2_X1 U7220 ( .A1(n5775), .A2(n5774), .ZN(n8648) );
  NAND2_X1 U7221 ( .A1(n5779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  MUX2_X1 U7222 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5777), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5778) );
  NAND2_X1 U7223 ( .A1(n5782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5783) );
  MUX2_X1 U7224 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8648), .S(n6263), .Z(n9804) );
  NAND2_X1 U7225 ( .A1(n6418), .A2(n9804), .ZN(n6846) );
  NAND2_X1 U7226 ( .A1(n5795), .A2(n5794), .ZN(n5792) );
  NAND2_X1 U7227 ( .A1(n5792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5793) );
  XNOR2_X2 U7228 ( .A(n5795), .B(n5794), .ZN(n8499) );
  OR2_X4 U7229 ( .A1(n9881), .A2(n9753), .ZN(n7985) );
  INV_X1 U7230 ( .A(n9804), .ZN(n8063) );
  NAND2_X1 U7231 ( .A1(n6052), .A2(n5796), .ZN(n5797) );
  NAND2_X4 U7232 ( .A1(n5797), .A2(n6742), .ZN(n7995) );
  NAND2_X1 U7233 ( .A1(n8063), .A2(n7593), .ZN(n5798) );
  INV_X1 U7234 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7235 ( .A1(n5816), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U7236 ( .A1(n7764), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7237 ( .A1(n5800), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7238 ( .A1(n6829), .A2(n7985), .ZN(n5813) );
  NAND2_X1 U7239 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5805) );
  MUX2_X1 U7240 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5805), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5808) );
  INV_X1 U7241 ( .A(n5821), .ZN(n5807) );
  NAND2_X1 U7242 ( .A1(n5808), .A2(n5807), .ZN(n6391) );
  INV_X1 U7243 ( .A(n6391), .ZN(n6270) );
  XNOR2_X1 U7244 ( .A(n7965), .B(n7995), .ZN(n5811) );
  XNOR2_X1 U7245 ( .A(n5813), .B(n5811), .ZN(n7967) );
  NAND2_X1 U7246 ( .A1(n7968), .A2(n7967), .ZN(n7966) );
  INV_X1 U7247 ( .A(n5811), .ZN(n5812) );
  NAND2_X1 U7248 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  NAND2_X1 U7249 ( .A1(n7966), .A2(n5814), .ZN(n8172) );
  INV_X1 U7250 ( .A(n8172), .ZN(n5828) );
  INV_X1 U7251 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6373) );
  OR2_X1 U7252 ( .A1(n7082), .A2(n6373), .ZN(n5820) );
  NAND2_X1 U7253 ( .A1(n7764), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5819) );
  INV_X1 U7254 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5815) );
  OR2_X1 U7255 ( .A1(n5850), .A2(n5815), .ZN(n5818) );
  NAND2_X1 U7256 ( .A1(n5816), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5817) );
  NOR2_X1 U7257 ( .A1(n6696), .A2(n5895), .ZN(n5823) );
  INV_X1 U7258 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  XNOR2_X1 U7259 ( .A(n8170), .B(n7995), .ZN(n5824) );
  NAND2_X1 U7260 ( .A1(n5823), .A2(n5824), .ZN(n5829) );
  INV_X1 U7261 ( .A(n5823), .ZN(n5825) );
  INV_X1 U7262 ( .A(n5824), .ZN(n6697) );
  NAND2_X1 U7263 ( .A1(n5825), .A2(n6697), .ZN(n5826) );
  NAND2_X1 U7264 ( .A1(n5829), .A2(n5826), .ZN(n8171) );
  NAND2_X1 U7265 ( .A1(n8173), .A2(n5829), .ZN(n5848) );
  INV_X1 U7266 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7267 ( .A1(n5816), .A2(n5830), .ZN(n5836) );
  NAND2_X1 U7268 ( .A1(n7764), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5835) );
  INV_X1 U7269 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5831) );
  OR2_X1 U7270 ( .A1(n5850), .A2(n5831), .ZN(n5834) );
  INV_X1 U7271 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5832) );
  OR2_X1 U7272 ( .A1(n7742), .A2(n5832), .ZN(n5833) );
  NOR2_X1 U7273 ( .A1(n6790), .A2(n7994), .ZN(n5844) );
  NAND2_X1 U7274 ( .A1(n7747), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5843) );
  NOR2_X1 U7275 ( .A1(n5822), .A2(n5838), .ZN(n5837) );
  MUX2_X1 U7276 ( .A(n5838), .B(n5837), .S(P2_IR_REG_3__SCAN_IN), .Z(n5841) );
  NAND2_X1 U7277 ( .A1(n5822), .A2(n5839), .ZN(n5859) );
  INV_X1 U7278 ( .A(n5859), .ZN(n5840) );
  NOR2_X1 U7279 ( .A1(n5841), .A2(n5840), .ZN(n6271) );
  NAND2_X1 U7280 ( .A1(n7515), .A2(n6271), .ZN(n5842) );
  OAI211_X1 U7281 ( .C1(n5856), .C2(n6091), .A(n5843), .B(n5842), .ZN(n6692)
         );
  XNOR2_X1 U7282 ( .A(n6692), .B(n7995), .ZN(n6708) );
  NAND2_X1 U7283 ( .A1(n5844), .A2(n6708), .ZN(n5863) );
  INV_X1 U7284 ( .A(n5844), .ZN(n5846) );
  INV_X1 U7285 ( .A(n6708), .ZN(n5845) );
  NAND2_X1 U7286 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  AND2_X1 U7287 ( .A1(n5863), .A2(n5847), .ZN(n6698) );
  NAND2_X1 U7288 ( .A1(n5848), .A2(n6698), .ZN(n6700) );
  NAND2_X1 U7289 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5888) );
  OAI21_X1 U7290 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5888), .ZN(n6793) );
  INV_X1 U7291 ( .A(n6793), .ZN(n5849) );
  NAND2_X1 U7292 ( .A1(n5816), .A2(n5849), .ZN(n5855) );
  NAND2_X1 U7293 ( .A1(n7764), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5854) );
  INV_X1 U7294 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6258) );
  OR2_X1 U7295 ( .A1(n7082), .A2(n6258), .ZN(n5853) );
  INV_X1 U7296 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5851) );
  OR2_X1 U7297 ( .A1(n5850), .A2(n5851), .ZN(n5852) );
  INV_X1 U7298 ( .A(n6849), .ZN(n8220) );
  NAND2_X1 U7299 ( .A1(n8220), .A2(n7985), .ZN(n5867) );
  INV_X1 U7300 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6090) );
  INV_X2 U7301 ( .A(n5856), .ZN(n5928) );
  NAND2_X1 U7302 ( .A1(n5928), .A2(n5857), .ZN(n5862) );
  NAND2_X1 U7303 ( .A1(n5859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  MUX2_X1 U7304 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5858), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5860) );
  AND2_X1 U7305 ( .A1(n5860), .A2(n5897), .ZN(n6341) );
  NAND2_X1 U7306 ( .A1(n7515), .A2(n6341), .ZN(n5861) );
  OAI211_X1 U7307 ( .C1(n5869), .C2(n6090), .A(n5862), .B(n5861), .ZN(n6783)
         );
  XNOR2_X1 U7308 ( .A(n6783), .B(n7995), .ZN(n5865) );
  XNOR2_X1 U7309 ( .A(n5867), .B(n5865), .ZN(n6707) );
  AND2_X1 U7310 ( .A1(n6707), .A2(n5863), .ZN(n5864) );
  NAND2_X1 U7311 ( .A1(n6700), .A2(n5864), .ZN(n6705) );
  INV_X1 U7312 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U7313 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  INV_X1 U7314 ( .A(n8106), .ZN(n5920) );
  NAND2_X1 U7315 ( .A1(n6103), .A2(n5928), .ZN(n5873) );
  INV_X2 U7316 ( .A(n5869), .ZN(n7747) );
  NAND2_X1 U7317 ( .A1(n5908), .A2(n5870), .ZN(n5929) );
  NAND2_X1 U7318 ( .A1(n5929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5871) );
  XNOR2_X1 U7319 ( .A(n5871), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6472) );
  AOI22_X1 U7320 ( .A1(n7747), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7515), .B2(
        n6472), .ZN(n5872) );
  XNOR2_X1 U7321 ( .A(n6854), .B(n7995), .ZN(n6553) );
  INV_X1 U7322 ( .A(n5888), .ZN(n5874) );
  NAND2_X1 U7323 ( .A1(n5874), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5913) );
  INV_X1 U7324 ( .A(n5913), .ZN(n5876) );
  AND2_X1 U7325 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5875) );
  NAND2_X1 U7326 ( .A1(n5876), .A2(n5875), .ZN(n5937) );
  INV_X1 U7327 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5877) );
  OAI21_X1 U7328 ( .B1(n5913), .B2(n5877), .A(n8115), .ZN(n5878) );
  AND2_X1 U7329 ( .A1(n5937), .A2(n5878), .ZN(n8113) );
  NAND2_X1 U7330 ( .A1(n5816), .A2(n8113), .ZN(n5884) );
  NAND2_X1 U7331 ( .A1(n7764), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5883) );
  INV_X1 U7332 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5879) );
  OR2_X1 U7333 ( .A1(n7742), .A2(n5879), .ZN(n5882) );
  INV_X1 U7334 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5880) );
  OR2_X1 U7335 ( .A1(n5850), .A2(n5880), .ZN(n5881) );
  NOR2_X1 U7336 ( .A1(n8179), .A2(n7994), .ZN(n5885) );
  NAND2_X1 U7337 ( .A1(n6553), .A2(n5885), .ZN(n5926) );
  INV_X1 U7338 ( .A(n8111), .ZN(n5925) );
  INV_X1 U7339 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7340 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  AND2_X1 U7341 ( .A1(n5913), .A2(n5889), .ZN(n9750) );
  NAND2_X1 U7342 ( .A1(n5816), .A2(n9750), .ZN(n5894) );
  NAND2_X1 U7343 ( .A1(n7764), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5893) );
  INV_X1 U7344 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5890) );
  INV_X1 U7345 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5891) );
  OR2_X1 U7346 ( .A1(n5850), .A2(n5891), .ZN(n5892) );
  NOR2_X1 U7347 ( .A1(n6860), .A2(n5895), .ZN(n5904) );
  NAND2_X1 U7348 ( .A1(n5896), .A2(n5928), .ZN(n5903) );
  NAND2_X1 U7349 ( .A1(n5897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5899) );
  MUX2_X1 U7350 ( .A(n5899), .B(P2_IR_REG_31__SCAN_IN), .S(n5898), .Z(n5901)
         );
  INV_X1 U7351 ( .A(n5908), .ZN(n5900) );
  AOI22_X1 U7352 ( .A1(n7747), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7515), .B2(
        n6355), .ZN(n5902) );
  XNOR2_X1 U7353 ( .A(n9831), .B(n7593), .ZN(n5905) );
  NAND2_X1 U7354 ( .A1(n5904), .A2(n5905), .ZN(n5923) );
  INV_X1 U7355 ( .A(n5904), .ZN(n5906) );
  INV_X1 U7356 ( .A(n5905), .ZN(n8188) );
  NAND2_X1 U7357 ( .A1(n5906), .A2(n8188), .ZN(n5907) );
  NAND2_X1 U7358 ( .A1(n5923), .A2(n5907), .ZN(n8148) );
  NAND2_X1 U7359 ( .A1(n6098), .A2(n5928), .ZN(n5911) );
  OR2_X1 U7360 ( .A1(n5908), .A2(n5838), .ZN(n5909) );
  XNOR2_X1 U7361 ( .A(n5909), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6398) );
  AOI22_X1 U7362 ( .A1(n7747), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7515), .B2(
        n6398), .ZN(n5910) );
  INV_X1 U7363 ( .A(n5922), .ZN(n5918) );
  INV_X1 U7364 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8512) );
  OR2_X1 U7365 ( .A1(n7082), .A2(n8512), .ZN(n5917) );
  NAND2_X1 U7366 ( .A1(n5912), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5916) );
  XNOR2_X1 U7367 ( .A(n5913), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U7368 ( .A1(n5816), .A2(n8513), .ZN(n5915) );
  NAND2_X1 U7369 ( .A1(n7764), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5914) );
  NAND4_X1 U7370 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n8219)
         );
  NAND2_X1 U7371 ( .A1(n8219), .A2(n7985), .ZN(n5921) );
  AND2_X1 U7372 ( .A1(n5918), .A2(n5921), .ZN(n5924) );
  OR2_X1 U7373 ( .A1(n8148), .A2(n5924), .ZN(n8107) );
  XNOR2_X1 U7374 ( .A(n5922), .B(n5921), .ZN(n8187) );
  AND2_X1 U7375 ( .A1(n8187), .A2(n5923), .ZN(n8182) );
  OR2_X1 U7376 ( .A1(n5925), .A2(n8108), .ZN(n6549) );
  AND2_X1 U7377 ( .A1(n6549), .A2(n5926), .ZN(n5927) );
  NAND2_X1 U7378 ( .A1(n6550), .A2(n5927), .ZN(n5948) );
  NAND2_X1 U7379 ( .A1(n6107), .A2(n5928), .ZN(n5935) );
  NAND2_X1 U7380 ( .A1(n5931), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5930) );
  MUX2_X1 U7381 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5930), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5933) );
  INV_X1 U7382 ( .A(n5967), .ZN(n5932) );
  AOI22_X1 U7383 ( .A1(n7747), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7515), .B2(
        n6601), .ZN(n5934) );
  NAND2_X1 U7384 ( .A1(n5935), .A2(n5934), .ZN(n6960) );
  XNOR2_X1 U7385 ( .A(n6960), .B(n7995), .ZN(n5944) );
  INV_X1 U7386 ( .A(n5937), .ZN(n5936) );
  NAND2_X1 U7387 ( .A1(n5936), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5953) );
  INV_X1 U7388 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U7389 ( .A1(n5937), .A2(n6546), .ZN(n5938) );
  AND2_X1 U7390 ( .A1(n5953), .A2(n5938), .ZN(n6545) );
  NAND2_X1 U7391 ( .A1(n5816), .A2(n6545), .ZN(n5943) );
  NAND2_X1 U7392 ( .A1(n7764), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5942) );
  INV_X1 U7393 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6870) );
  OR2_X1 U7394 ( .A1(n7742), .A2(n6870), .ZN(n5941) );
  INV_X1 U7395 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5939) );
  OR2_X1 U7396 ( .A1(n5850), .A2(n5939), .ZN(n5940) );
  NOR2_X1 U7397 ( .A1(n7042), .A2(n7994), .ZN(n5945) );
  NAND2_X1 U7398 ( .A1(n5944), .A2(n5945), .ZN(n5960) );
  INV_X1 U7399 ( .A(n5944), .ZN(n6638) );
  INV_X1 U7400 ( .A(n5945), .ZN(n5946) );
  NAND2_X1 U7401 ( .A1(n6638), .A2(n5946), .ZN(n5947) );
  AND2_X1 U7402 ( .A1(n5960), .A2(n5947), .ZN(n6551) );
  NAND2_X1 U7403 ( .A1(n5948), .A2(n6551), .ZN(n6637) );
  NAND2_X1 U7404 ( .A1(n6128), .A2(n5928), .ZN(n5951) );
  OR2_X1 U7405 ( .A1(n5967), .A2(n5838), .ZN(n5949) );
  XNOR2_X1 U7406 ( .A(n5949), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6771) );
  AOI22_X1 U7407 ( .A1(n7747), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7515), .B2(
        n6771), .ZN(n5950) );
  NAND2_X1 U7408 ( .A1(n5951), .A2(n5950), .ZN(n7055) );
  XNOR2_X1 U7409 ( .A(n7055), .B(n7995), .ZN(n5962) );
  NAND2_X1 U7410 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  AND2_X1 U7411 ( .A1(n5975), .A2(n5954), .ZN(n7047) );
  NAND2_X1 U7412 ( .A1(n5816), .A2(n7047), .ZN(n5959) );
  NAND2_X1 U7413 ( .A1(n7764), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5958) );
  INV_X1 U7414 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7049) );
  OR2_X1 U7415 ( .A1(n7742), .A2(n7049), .ZN(n5957) );
  INV_X1 U7416 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7417 ( .A1(n5850), .A2(n5955), .ZN(n5956) );
  INV_X1 U7418 ( .A(n7005), .ZN(n8217) );
  NAND2_X1 U7419 ( .A1(n8217), .A2(n7985), .ZN(n5963) );
  XNOR2_X1 U7420 ( .A(n5962), .B(n5963), .ZN(n6649) );
  AND2_X1 U7421 ( .A1(n6649), .A2(n5960), .ZN(n5961) );
  INV_X1 U7422 ( .A(n5962), .ZN(n5964) );
  NAND2_X1 U7423 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  NAND2_X1 U7424 ( .A1(n6184), .A2(n5928), .ZN(n5972) );
  INV_X1 U7425 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7426 ( .A1(n5967), .A2(n5966), .ZN(n6005) );
  NAND2_X1 U7427 ( .A1(n6005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5969) );
  INV_X1 U7428 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7429 ( .A1(n5969), .A2(n5968), .ZN(n5987) );
  OR2_X1 U7430 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  AOI22_X1 U7431 ( .A1(n7515), .A2(n7027), .B1(n7747), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5971) );
  NAND2_X2 U7432 ( .A1(n5972), .A2(n5971), .ZN(n9863) );
  XNOR2_X1 U7433 ( .A(n9863), .B(n7995), .ZN(n5981) );
  INV_X1 U7434 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7011) );
  OR2_X1 U7435 ( .A1(n7082), .A2(n7011), .ZN(n5980) );
  NAND2_X1 U7436 ( .A1(n5912), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5979) );
  INV_X1 U7437 ( .A(n5975), .ZN(n5973) );
  NAND2_X1 U7438 ( .A1(n5973), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5992) );
  INV_X1 U7439 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7440 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  AND2_X1 U7441 ( .A1(n5992), .A2(n5976), .ZN(n6755) );
  NAND2_X1 U7442 ( .A1(n5816), .A2(n6755), .ZN(n5978) );
  NAND2_X1 U7443 ( .A1(n7764), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5977) );
  NAND4_X1 U7444 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n8216)
         );
  AND2_X1 U7445 ( .A1(n8216), .A2(n7985), .ZN(n5982) );
  NAND2_X1 U7446 ( .A1(n5981), .A2(n5982), .ZN(n5986) );
  INV_X1 U7447 ( .A(n5981), .ZN(n6719) );
  INV_X1 U7448 ( .A(n5982), .ZN(n5983) );
  NAND2_X1 U7449 ( .A1(n6719), .A2(n5983), .ZN(n5984) );
  NAND2_X1 U7450 ( .A1(n5986), .A2(n5984), .ZN(n6760) );
  INV_X1 U7451 ( .A(n6760), .ZN(n5985) );
  NAND2_X1 U7452 ( .A1(n6757), .A2(n5986), .ZN(n6004) );
  NAND2_X1 U7453 ( .A1(n6182), .A2(n5928), .ZN(n5990) );
  NAND2_X1 U7454 ( .A1(n5987), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7455 ( .A(n5988), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7166) );
  AOI22_X1 U7456 ( .A1(n7166), .A2(n7515), .B1(n7747), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7457 ( .A1(n5990), .A2(n5989), .ZN(n6980) );
  XNOR2_X1 U7458 ( .A(n6980), .B(n7995), .ZN(n6000) );
  NAND2_X1 U7459 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  AND2_X1 U7460 ( .A1(n6010), .A2(n5993), .ZN(n6975) );
  NAND2_X1 U7461 ( .A1(n5816), .A2(n6975), .ZN(n5999) );
  NAND2_X1 U7462 ( .A1(n7764), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5998) );
  INV_X1 U7463 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5994) );
  OR2_X1 U7464 ( .A1(n7742), .A2(n5994), .ZN(n5997) );
  INV_X1 U7465 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5995) );
  OR2_X1 U7466 ( .A1(n5850), .A2(n5995), .ZN(n5996) );
  NOR2_X1 U7467 ( .A1(n7006), .A2(n7994), .ZN(n6001) );
  NAND2_X1 U7468 ( .A1(n6000), .A2(n6001), .ZN(n6018) );
  INV_X1 U7469 ( .A(n6000), .ZN(n6808) );
  INV_X1 U7470 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7471 ( .A1(n6808), .A2(n6002), .ZN(n6003) );
  AND2_X1 U7472 ( .A1(n6018), .A2(n6003), .ZN(n6717) );
  NAND2_X1 U7473 ( .A1(n6004), .A2(n6717), .ZN(n6720) );
  NAND2_X1 U7474 ( .A1(n6230), .A2(n5928), .ZN(n6008) );
  NAND2_X1 U7475 ( .A1(n6023), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U7476 ( .A(n6006), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7252) );
  AOI22_X1 U7477 ( .A1(n7252), .A2(n7515), .B1(n7747), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7478 ( .A1(n6008), .A2(n6007), .ZN(n7148) );
  XNOR2_X1 U7479 ( .A(n7148), .B(n7995), .ZN(n6020) );
  INV_X1 U7480 ( .A(n6010), .ZN(n6009) );
  NAND2_X1 U7481 ( .A1(n6009), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6026) );
  INV_X1 U7482 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7170) );
  NAND2_X1 U7483 ( .A1(n6010), .A2(n7170), .ZN(n6011) );
  AND2_X1 U7484 ( .A1(n6026), .A2(n6011), .ZN(n6993) );
  NAND2_X1 U7485 ( .A1(n5816), .A2(n6993), .ZN(n6017) );
  NAND2_X1 U7486 ( .A1(n7764), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6016) );
  INV_X1 U7487 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6012) );
  OR2_X1 U7488 ( .A1(n7082), .A2(n6012), .ZN(n6015) );
  INV_X1 U7489 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7490 ( .A1(n5850), .A2(n6013), .ZN(n6014) );
  NAND2_X1 U7491 ( .A1(n8214), .A2(n7985), .ZN(n6021) );
  XNOR2_X1 U7492 ( .A(n6020), .B(n6021), .ZN(n6817) );
  AND2_X1 U7493 ( .A1(n6817), .A2(n6018), .ZN(n6019) );
  INV_X1 U7494 ( .A(n6020), .ZN(n6022) );
  NAND2_X1 U7495 ( .A1(n6022), .A2(n6021), .ZN(n6055) );
  NAND2_X1 U7496 ( .A1(n6811), .A2(n6055), .ZN(n6059) );
  NAND2_X1 U7497 ( .A1(n6306), .A2(n5928), .ZN(n6025) );
  OAI21_X1 U7498 ( .B1(n6023), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6320) );
  XNOR2_X1 U7499 ( .A(n6320), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7376) );
  AOI22_X1 U7500 ( .A1(n7376), .A2(n7515), .B1(n7747), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6024) );
  XNOR2_X1 U7501 ( .A(n7881), .B(n7995), .ZN(n6032) );
  NAND2_X1 U7502 ( .A1(n5912), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6031) );
  INV_X1 U7503 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7154) );
  OR2_X1 U7504 ( .A1(n7742), .A2(n7154), .ZN(n6030) );
  NAND2_X1 U7505 ( .A1(n6026), .A2(n7247), .ZN(n6027) );
  AND2_X1 U7506 ( .A1(n6066), .A2(n6027), .ZN(n6064) );
  NAND2_X1 U7507 ( .A1(n5816), .A2(n6064), .ZN(n6029) );
  NAND2_X1 U7508 ( .A1(n7764), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6028) );
  NAND4_X1 U7509 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n8213)
         );
  AND2_X1 U7510 ( .A1(n8213), .A2(n7985), .ZN(n6033) );
  NAND2_X1 U7511 ( .A1(n6032), .A2(n6033), .ZN(n6919) );
  INV_X1 U7512 ( .A(n6032), .ZN(n6913) );
  INV_X1 U7513 ( .A(n6033), .ZN(n6034) );
  NAND2_X1 U7514 ( .A1(n6913), .A2(n6034), .ZN(n6035) );
  NAND2_X1 U7515 ( .A1(n6919), .A2(n6035), .ZN(n6058) );
  INV_X1 U7516 ( .A(P2_B_REG_SCAN_IN), .ZN(n8055) );
  XOR2_X1 U7517 ( .A(n7321), .B(n8055), .Z(n6036) );
  INV_X1 U7518 ( .A(n9766), .ZN(n6038) );
  NAND2_X1 U7519 ( .A1(n7484), .A2(n7533), .ZN(n9800) );
  INV_X1 U7520 ( .A(n6410), .ZN(n6741) );
  NOR4_X1 U7521 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6047) );
  INV_X1 U7522 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9781) );
  INV_X1 U7523 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10057) );
  INV_X1 U7524 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9796) );
  INV_X1 U7525 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9795) );
  NAND4_X1 U7526 ( .A1(n9781), .A2(n10057), .A3(n9796), .A4(n9795), .ZN(n6044)
         );
  NOR4_X1 U7527 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6042) );
  NOR4_X1 U7528 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6041) );
  NOR4_X1 U7529 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6040) );
  NOR4_X1 U7530 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6039) );
  NAND4_X1 U7531 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n6043)
         );
  NOR4_X1 U7532 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6044), .A4(n6043), .ZN(n6046) );
  NOR4_X1 U7533 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6045) );
  NAND3_X1 U7534 ( .A1(n6047), .A2(n6046), .A3(n6045), .ZN(n6048) );
  NAND2_X1 U7535 ( .A1(n7321), .A2(n7533), .ZN(n9798) );
  INV_X1 U7536 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7537 ( .A1(n9766), .A2(n6049), .ZN(n6050) );
  NOR2_X1 U7538 ( .A1(n6739), .A2(n6432), .ZN(n6051) );
  NAND2_X1 U7539 ( .A1(n6741), .A2(n6051), .ZN(n6078) );
  INV_X1 U7540 ( .A(n6052), .ZN(n9805) );
  INV_X1 U7541 ( .A(n6264), .ZN(n6076) );
  NOR2_X1 U7542 ( .A1(n9836), .A2(n6076), .ZN(n6053) );
  INV_X1 U7543 ( .A(n6058), .ZN(n6056) );
  AND2_X1 U7544 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  NAND2_X1 U7545 ( .A1(n6811), .A2(n6057), .ZN(n6921) );
  INV_X1 U7546 ( .A(n6921), .ZN(n6915) );
  AOI211_X1 U7547 ( .C1(n6059), .C2(n6058), .A(n8196), .B(n6915), .ZN(n6082)
         );
  INV_X1 U7548 ( .A(n7881), .ZN(n9472) );
  NOR2_X1 U7549 ( .A1(n6052), .A2(n7790), .ZN(n9749) );
  INV_X1 U7550 ( .A(n9749), .ZN(n6060) );
  NOR2_X1 U7551 ( .A1(n9472), .A2(n8207), .ZN(n6081) );
  NAND2_X1 U7552 ( .A1(n6078), .A2(n6407), .ZN(n6063) );
  OR2_X1 U7553 ( .A1(n6264), .A2(n6061), .ZN(n6735) );
  AND3_X1 U7554 ( .A1(n6261), .A2(n6124), .A3(n6735), .ZN(n6062) );
  NAND2_X1 U7555 ( .A1(n6063), .A2(n6062), .ZN(n8067) );
  INV_X1 U7556 ( .A(n6064), .ZN(n7153) );
  OAI22_X1 U7557 ( .A1(n8162), .A2(n7153), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7247), .ZN(n6080) );
  NAND2_X1 U7558 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  AND2_X1 U7559 ( .A1(n7071), .A2(n6067), .ZN(n7472) );
  NAND2_X1 U7560 ( .A1(n5816), .A2(n7472), .ZN(n6073) );
  NAND2_X1 U7561 ( .A1(n7764), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6072) );
  INV_X1 U7562 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7563 ( .A1(n7082), .A2(n6068), .ZN(n6071) );
  INV_X1 U7564 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6069) );
  OR2_X1 U7565 ( .A1(n5850), .A2(n6069), .ZN(n6070) );
  INV_X1 U7566 ( .A(n9765), .ZN(n6077) );
  NAND3_X1 U7567 ( .A1(n6077), .A2(n8506), .A3(n6735), .ZN(n7959) );
  OR2_X1 U7568 ( .A1(n6078), .A2(n7959), .ZN(n8200) );
  INV_X1 U7569 ( .A(n8200), .ZN(n8190) );
  OAI22_X1 U7570 ( .A1(n7451), .A2(n8202), .B1(n8200), .B2(n6985), .ZN(n6079)
         );
  OR4_X1 U7571 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(P2_U3236)
         );
  NOR2_X2 U7572 ( .A1(n7775), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9429) );
  INV_X1 U7573 ( .A(n9429), .ZN(n7481) );
  NAND2_X1 U7574 ( .A1(n7775), .A2(P1_U3084), .ZN(n7552) );
  CLKBUF_X1 U7575 ( .A(n7552), .Z(n9431) );
  INV_X1 U7576 ( .A(n9529), .ZN(n6135) );
  OAI222_X1 U7577 ( .A1(n7481), .A2(n6083), .B1(n9431), .B2(n6093), .C1(
        P1_U3084), .C2(n6135), .ZN(P1_U3351) );
  INV_X1 U7578 ( .A(n9072), .ZN(n9067) );
  OAI222_X1 U7579 ( .A1(n7481), .A2(n4918), .B1(n9431), .B2(n6095), .C1(
        P1_U3084), .C2(n9067), .ZN(P1_U3352) );
  INV_X1 U7580 ( .A(n9083), .ZN(n9081) );
  OAI222_X1 U7581 ( .A1(n7481), .A2(n6084), .B1(n9431), .B2(n6091), .C1(
        P1_U3084), .C2(n9081), .ZN(P1_U3350) );
  AOI22_X1 U7582 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n9429), .B1(n9541), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6085) );
  OAI21_X1 U7583 ( .B1(n6089), .B2(n9431), .A(n6085), .ZN(P1_U3349) );
  NAND2_X1 U7584 ( .A1(n4914), .A2(P2_U3152), .ZN(n8647) );
  AOI22_X1 U7585 ( .A1(n6355), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8644), .ZN(n6086) );
  OAI21_X1 U7586 ( .B1(n6088), .B2(n8647), .A(n6086), .ZN(P2_U3353) );
  AOI22_X1 U7587 ( .A1(n6178), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9429), .ZN(n6087) );
  OAI21_X1 U7588 ( .B1(n6088), .B2(n9431), .A(n6087), .ZN(P1_U3348) );
  INV_X1 U7589 ( .A(n8644), .ZN(n8641) );
  INV_X1 U7590 ( .A(n6341), .ZN(n6349) );
  OAI222_X1 U7591 ( .A1(n8641), .A2(n6090), .B1(n8016), .B2(n6089), .C1(
        P2_U3152), .C2(n6349), .ZN(P2_U3354) );
  INV_X1 U7592 ( .A(n6271), .ZN(n6335) );
  OAI222_X1 U7593 ( .A1(n8641), .A2(n6092), .B1(n8016), .B2(n6091), .C1(
        P2_U3152), .C2(n6335), .ZN(P2_U3355) );
  OAI222_X1 U7594 ( .A1(n8641), .A2(n6094), .B1(n8016), .B2(n6093), .C1(
        P2_U3152), .C2(n4478), .ZN(P2_U3356) );
  INV_X1 U7595 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6096) );
  OAI222_X1 U7596 ( .A1(n8641), .A2(n6096), .B1(n8016), .B2(n6095), .C1(
        P2_U3152), .C2(n6391), .ZN(P2_U3357) );
  NAND2_X1 U7597 ( .A1(n6212), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7598 ( .B1(n7112), .B2(n6212), .A(n6097), .ZN(P1_U3440) );
  INV_X1 U7599 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6099) );
  INV_X1 U7600 ( .A(n6098), .ZN(n6101) );
  INV_X1 U7601 ( .A(n6398), .ZN(n6365) );
  OAI222_X1 U7602 ( .A1(n8641), .A2(n6099), .B1(n8016), .B2(n6101), .C1(
        P2_U3152), .C2(n6365), .ZN(P2_U3352) );
  INV_X1 U7603 ( .A(n9558), .ZN(n6100) );
  OAI222_X1 U7604 ( .A1(n7481), .A2(n6102), .B1(n9431), .B2(n6101), .C1(
        P1_U3084), .C2(n6100), .ZN(P1_U3347) );
  INV_X1 U7605 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6104) );
  INV_X1 U7606 ( .A(n6103), .ZN(n6105) );
  INV_X1 U7607 ( .A(n6194), .ZN(n6159) );
  OAI222_X1 U7608 ( .A1(n7481), .A2(n6104), .B1(n9431), .B2(n6105), .C1(
        P1_U3084), .C2(n6159), .ZN(P1_U3346) );
  INV_X1 U7609 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6106) );
  INV_X1 U7610 ( .A(n6472), .ZN(n6406) );
  OAI222_X1 U7611 ( .A1(n8641), .A2(n6106), .B1(n8016), .B2(n6105), .C1(
        P2_U3152), .C2(n6406), .ZN(P2_U3351) );
  INV_X1 U7612 ( .A(n6107), .ZN(n6109) );
  INV_X1 U7613 ( .A(n6601), .ZN(n6609) );
  OAI222_X1 U7614 ( .A1(n8641), .A2(n6108), .B1(n8016), .B2(n6109), .C1(
        P2_U3152), .C2(n6609), .ZN(P2_U3350) );
  INV_X1 U7615 ( .A(n6292), .ZN(n6197) );
  OAI222_X1 U7616 ( .A1(n7481), .A2(n6110), .B1(n9431), .B2(n6109), .C1(
        P1_U3084), .C2(n6197), .ZN(P1_U3345) );
  INV_X1 U7617 ( .A(n6212), .ZN(n9038) );
  INV_X1 U7618 ( .A(n9650), .ZN(n9649) );
  OAI21_X1 U7619 ( .B1(n9649), .B2(P1_D_REG_1__SCAN_IN), .A(n6240), .ZN(n6111)
         );
  OAI21_X1 U7620 ( .B1(n6112), .B2(n9038), .A(n6111), .ZN(P1_U3441) );
  INV_X1 U7621 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8279) );
  AND2_X1 U7622 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n6113) );
  NAND2_X1 U7623 ( .A1(n6114), .A2(n6113), .ZN(n7080) );
  INV_X1 U7624 ( .A(n7080), .ZN(n6115) );
  INV_X1 U7625 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7447) );
  INV_X1 U7626 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7627 ( .B1(n7311), .B2(n7447), .A(n6116), .ZN(n6118) );
  NAND2_X1 U7628 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6117) );
  AND2_X1 U7629 ( .A1(n6118), .A2(n7522), .ZN(n8457) );
  NAND2_X1 U7630 ( .A1(n8457), .A2(n5816), .ZN(n6120) );
  AOI22_X1 U7631 ( .A1(n5800), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n5912), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n6119) );
  OAI211_X1 U7632 ( .C1(n7728), .C2(n8279), .A(n6120), .B(n6119), .ZN(n8476)
         );
  NAND2_X1 U7633 ( .A1(n8476), .A2(P2_U3966), .ZN(n6121) );
  OAI21_X1 U7634 ( .B1(n5394), .B2(P2_U3966), .A(n6121), .ZN(P2_U3571) );
  INV_X1 U7635 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7636 ( .A1(n6418), .A2(P2_U3966), .ZN(n6122) );
  OAI21_X1 U7637 ( .B1(n6123), .B2(P2_U3966), .A(n6122), .ZN(P2_U3552) );
  OR2_X1 U7638 ( .A1(n6124), .A2(P2_U3152), .ZN(n7963) );
  NAND2_X1 U7639 ( .A1(n9765), .A2(n7963), .ZN(n6125) );
  NAND2_X1 U7640 ( .A1(n6125), .A2(n7515), .ZN(n6127) );
  OR2_X1 U7641 ( .A1(n9765), .A2(n6264), .ZN(n6126) );
  AND2_X1 U7642 ( .A1(n6127), .A2(n6126), .ZN(n8291) );
  NOR2_X1 U7643 ( .A1(n9738), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7644 ( .A(n6128), .ZN(n6130) );
  OAI222_X1 U7645 ( .A1(n7481), .A2(n6129), .B1(n9431), .B2(n6130), .C1(n6289), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U7646 ( .A(n6771), .ZN(n6614) );
  OAI222_X1 U7647 ( .A1(n8641), .A2(n6131), .B1(n8016), .B2(n6130), .C1(n6614), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7648 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6168) );
  NOR2_X1 U7649 ( .A1(n9558), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6143) );
  INV_X1 U7650 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6133) );
  MUX2_X1 U7651 ( .A(n6133), .B(P1_REG1_REG_6__SCAN_IN), .S(n9558), .Z(n9560)
         );
  XNOR2_X1 U7652 ( .A(n9529), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9528) );
  NOR2_X1 U7653 ( .A1(n9515), .A2(n9510), .ZN(n9076) );
  NAND2_X1 U7654 ( .A1(n9072), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6134) );
  OAI211_X1 U7655 ( .C1(n9072), .C2(P1_REG1_REG_1__SCAN_IN), .A(n9076), .B(
        n6134), .ZN(n9074) );
  NAND2_X1 U7656 ( .A1(n9074), .A2(n6134), .ZN(n9527) );
  INV_X1 U7657 ( .A(n9527), .ZN(n6136) );
  INV_X1 U7658 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9716) );
  OAI22_X1 U7659 ( .A1(n9528), .A2(n6136), .B1(n9716), .B2(n6135), .ZN(n9090)
         );
  INV_X1 U7660 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6137) );
  MUX2_X1 U7661 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6137), .S(n9083), .Z(n9091)
         );
  NAND2_X1 U7662 ( .A1(n9090), .A2(n9091), .ZN(n9089) );
  NAND2_X1 U7663 ( .A1(n9083), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7664 ( .A1(n9089), .A2(n6138), .ZN(n9546) );
  INV_X1 U7665 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6139) );
  MUX2_X1 U7666 ( .A(n6139), .B(P1_REG1_REG_4__SCAN_IN), .S(n9541), .Z(n9547)
         );
  OR2_X1 U7667 ( .A1(n9546), .A2(n9547), .ZN(n9544) );
  OR2_X1 U7668 ( .A1(n9541), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7669 ( .A1(n9544), .A2(n6140), .ZN(n6171) );
  INV_X1 U7670 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9720) );
  MUX2_X1 U7671 ( .A(n9720), .B(P1_REG1_REG_5__SCAN_IN), .S(n6178), .Z(n6170)
         );
  INV_X1 U7672 ( .A(n6169), .ZN(n6142) );
  NAND2_X1 U7673 ( .A1(n6178), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7674 ( .A1(n6142), .A2(n6141), .ZN(n9561) );
  NOR2_X1 U7675 ( .A1(n9560), .A2(n9561), .ZN(n9559) );
  INV_X1 U7676 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6144) );
  MUX2_X1 U7677 ( .A(n6144), .B(P1_REG1_REG_7__SCAN_IN), .S(n6194), .Z(n6145)
         );
  NOR2_X1 U7678 ( .A1(n6146), .A2(n6145), .ZN(n6190) );
  AOI21_X1 U7679 ( .B1(n6146), .B2(n6145), .A(n6190), .ZN(n6164) );
  NAND2_X1 U7680 ( .A1(n6162), .A2(n4395), .ZN(n9521) );
  INV_X1 U7681 ( .A(n6147), .ZN(n9036) );
  NAND2_X1 U7682 ( .A1(n9558), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6157) );
  INV_X1 U7683 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6151) );
  NAND3_X1 U7684 ( .A1(n9071), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG2_REG_0__SCAN_IN), .ZN(n9070) );
  INV_X1 U7685 ( .A(n9070), .ZN(n6148) );
  AOI21_X1 U7686 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9072), .A(n6148), .ZN(
        n9536) );
  INV_X1 U7687 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6149) );
  MUX2_X1 U7688 ( .A(n6149), .B(P1_REG2_REG_2__SCAN_IN), .S(n9529), .Z(n9535)
         );
  AND2_X1 U7689 ( .A1(n9529), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9084) );
  MUX2_X1 U7690 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6151), .S(n9083), .Z(n6150)
         );
  INV_X1 U7691 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6629) );
  MUX2_X1 U7692 ( .A(n6629), .B(P1_REG2_REG_4__SCAN_IN), .S(n9541), .Z(n9551)
         );
  NOR2_X1 U7693 ( .A1(n9541), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6172) );
  INV_X1 U7694 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6152) );
  MUX2_X1 U7695 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6152), .S(n6178), .Z(n6173)
         );
  OAI21_X1 U7696 ( .B1(n9549), .B2(n6172), .A(n6173), .ZN(n6175) );
  INV_X1 U7697 ( .A(n6175), .ZN(n6154) );
  NOR2_X1 U7698 ( .A1(n6178), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6153) );
  NOR2_X1 U7699 ( .A1(n6154), .A2(n6153), .ZN(n9565) );
  INV_X1 U7700 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6155) );
  MUX2_X1 U7701 ( .A(n6155), .B(P1_REG2_REG_6__SCAN_IN), .S(n9558), .Z(n6156)
         );
  INV_X1 U7702 ( .A(n6156), .ZN(n9564) );
  NAND2_X1 U7703 ( .A1(n9565), .A2(n9564), .ZN(n9563) );
  INV_X1 U7704 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6158) );
  AOI22_X1 U7705 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6159), .B1(n6194), .B2(
        n6158), .ZN(n6160) );
  AOI21_X1 U7706 ( .B1(n6161), .B2(n6160), .A(n6195), .ZN(n6163) );
  NOR2_X1 U7707 ( .A1(n6147), .A2(P1_U3084), .ZN(n7550) );
  OAI22_X1 U7708 ( .A1(n6164), .A2(n9573), .B1(n6163), .B2(n9553), .ZN(n6165)
         );
  INV_X1 U7709 ( .A(n6165), .ZN(n6167) );
  AND2_X1 U7710 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6518) );
  AOI21_X1 U7711 ( .B1(n9578), .B2(n6194), .A(n6518), .ZN(n6166) );
  OAI211_X1 U7712 ( .C1(n9584), .C2(n6168), .A(n6167), .B(n6166), .ZN(P1_U3248) );
  INV_X1 U7713 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6181) );
  AOI211_X1 U7714 ( .C1(n6171), .C2(n6170), .A(n6169), .B(n9573), .ZN(n6177)
         );
  OR3_X1 U7715 ( .A1(n9549), .A2(n6173), .A3(n6172), .ZN(n6174) );
  AOI21_X1 U7716 ( .B1(n6175), .B2(n6174), .A(n9553), .ZN(n6176) );
  NOR2_X1 U7717 ( .A1(n6177), .A2(n6176), .ZN(n6180) );
  AND2_X1 U7718 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6459) );
  AOI21_X1 U7719 ( .B1(n9578), .B2(n6178), .A(n6459), .ZN(n6179) );
  OAI211_X1 U7720 ( .C1(n9584), .C2(n6181), .A(n6180), .B(n6179), .ZN(P1_U3246) );
  INV_X1 U7721 ( .A(n6182), .ZN(n6189) );
  AOI22_X1 U7722 ( .A1(n7166), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8644), .ZN(n6183) );
  OAI21_X1 U7723 ( .B1(n6189), .B2(n8647), .A(n6183), .ZN(P2_U3347) );
  INV_X1 U7724 ( .A(n6184), .ZN(n6186) );
  INV_X1 U7725 ( .A(n6578), .ZN(n6575) );
  OAI222_X1 U7726 ( .A1(n7481), .A2(n6185), .B1(n9431), .B2(n6186), .C1(n6575), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7727 ( .A(n7027), .ZN(n6779) );
  OAI222_X1 U7728 ( .A1(n8641), .A2(n6187), .B1(n8016), .B2(n6186), .C1(n6779), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7729 ( .A(n9591), .ZN(n9597) );
  OAI222_X1 U7730 ( .A1(P1_U3084), .A2(n9597), .B1(n9431), .B2(n6189), .C1(
        n6188), .C2(n7481), .ZN(P1_U3342) );
  NOR2_X1 U7731 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6194), .ZN(n6191) );
  NOR2_X1 U7732 ( .A1(n6191), .A2(n6190), .ZN(n6193) );
  INV_X1 U7733 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9724) );
  AOI22_X1 U7734 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6197), .B1(n6292), .B2(
        n9724), .ZN(n6192) );
  NOR2_X1 U7735 ( .A1(n6193), .A2(n6192), .ZN(n6285) );
  AOI21_X1 U7736 ( .B1(n6193), .B2(n6192), .A(n6285), .ZN(n6206) );
  INV_X1 U7737 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9454) );
  INV_X1 U7738 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6196) );
  AOI22_X1 U7739 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6197), .B1(n6292), .B2(
        n6196), .ZN(n6198) );
  AOI21_X1 U7740 ( .B1(n6199), .B2(n6198), .A(n6293), .ZN(n6200) );
  OR2_X1 U7741 ( .A1(n6200), .A2(n9553), .ZN(n6203) );
  INV_X1 U7742 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6201) );
  NOR2_X1 U7743 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6201), .ZN(n6594) );
  AOI21_X1 U7744 ( .B1(n9578), .B2(n6292), .A(n6594), .ZN(n6202) );
  OAI211_X1 U7745 ( .C1(n9454), .C2(n9584), .A(n6203), .B(n6202), .ZN(n6204)
         );
  INV_X1 U7746 ( .A(n6204), .ZN(n6205) );
  OAI21_X1 U7747 ( .B1(n6206), .B2(n9573), .A(n6205), .ZN(P1_U3249) );
  INV_X1 U7748 ( .A(n6509), .ZN(n9637) );
  OAI21_X1 U7749 ( .B1(n6207), .B2(n6209), .A(n6208), .ZN(n9523) );
  NAND2_X1 U7750 ( .A1(n9523), .A2(n8683), .ZN(n6216) );
  INV_X1 U7751 ( .A(n8706), .ZN(n8721) );
  INV_X1 U7752 ( .A(n6210), .ZN(n6214) );
  NOR2_X1 U7753 ( .A1(n5580), .A2(n9033), .ZN(n6211) );
  NAND3_X1 U7754 ( .A1(n6214), .A2(n6480), .A3(n6213), .ZN(n6236) );
  AOI22_X1 U7755 ( .A1(n8721), .A2(n6489), .B1(n6236), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7756 ( .C1(n8730), .C2(n9637), .A(n6216), .B(n6215), .ZN(P1_U3230) );
  INV_X1 U7757 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7758 ( .A1(n5024), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7759 ( .A1(n8093), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7760 ( .A1(n6217), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6218) );
  AND3_X1 U7761 ( .A1(n6220), .A2(n6219), .A3(n6218), .ZN(n8856) );
  INV_X1 U7762 ( .A(n8856), .ZN(n9139) );
  NAND2_X1 U7763 ( .A1(n9139), .A2(P1_U4006), .ZN(n6221) );
  OAI21_X1 U7764 ( .B1(P1_U4006), .B2(n6222), .A(n6221), .ZN(P1_U3586) );
  XNOR2_X1 U7765 ( .A(n6224), .B(n6223), .ZN(n6225) );
  XNOR2_X1 U7766 ( .A(n6226), .B(n6225), .ZN(n6229) );
  AOI22_X1 U7767 ( .A1(n8664), .A2(n6488), .B1(n8721), .B2(n9632), .ZN(n6228)
         );
  AOI22_X1 U7768 ( .A1(n8709), .A2(n4643), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6236), .ZN(n6227) );
  OAI211_X1 U7769 ( .C1(n6229), .C2(n8716), .A(n6228), .B(n6227), .ZN(P1_U3220) );
  INV_X1 U7770 ( .A(n6230), .ZN(n6232) );
  INV_X1 U7771 ( .A(n7252), .ZN(n7177) );
  OAI222_X1 U7772 ( .A1(n8641), .A2(n6231), .B1(n8016), .B2(n6232), .C1(
        P2_U3152), .C2(n7177), .ZN(P2_U3346) );
  OAI222_X1 U7773 ( .A1(n7481), .A2(n6233), .B1(n9431), .B2(n6232), .C1(
        P1_U3084), .C2(n4399), .ZN(P1_U3341) );
  XOR2_X1 U7774 ( .A(n6234), .B(n6235), .Z(n6239) );
  INV_X1 U7775 ( .A(n6620), .ZN(n9065) );
  AOI22_X1 U7776 ( .A1(n8664), .A2(n6489), .B1(n8721), .B2(n9065), .ZN(n6238)
         );
  AOI22_X1 U7777 ( .A1(n8709), .A2(n4970), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6236), .ZN(n6237) );
  OAI211_X1 U7778 ( .C1(n6239), .C2(n8716), .A(n6238), .B(n6237), .ZN(P1_U3235) );
  AND2_X1 U7779 ( .A1(n6480), .A2(n7112), .ZN(n6247) );
  OAI21_X1 U7780 ( .B1(n6241), .B2(P1_D_REG_1__SCAN_IN), .A(n6240), .ZN(n6245)
         );
  INV_X1 U7781 ( .A(n6241), .ZN(n6243) );
  NAND2_X1 U7782 ( .A1(n6243), .A2(n6242), .ZN(n6244) );
  OAI211_X1 U7783 ( .C1(n9706), .C2(n5579), .A(n6245), .B(n6244), .ZN(n6246)
         );
  INV_X1 U7784 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6253) );
  AND2_X1 U7785 ( .A1(n6488), .A2(n9637), .ZN(n8998) );
  NOR2_X1 U7786 ( .A1(n9629), .A2(n8998), .ZN(n8875) );
  INV_X1 U7787 ( .A(n6248), .ZN(n9037) );
  NOR3_X1 U7788 ( .A1(n8875), .A2(n6249), .A3(n9037), .ZN(n6250) );
  AOI21_X1 U7789 ( .B1(n9631), .B2(n6489), .A(n6250), .ZN(n6486) );
  OAI21_X1 U7790 ( .B1(n9637), .B2(n6251), .A(n6486), .ZN(n9405) );
  NAND2_X1 U7791 ( .A1(n9405), .A2(n9714), .ZN(n6252) );
  OAI21_X1 U7792 ( .B1(n9714), .B2(n6253), .A(n6252), .ZN(P1_U3454) );
  MUX2_X1 U7793 ( .A(n5890), .B(P2_REG2_REG_5__SCAN_IN), .S(n6355), .Z(n6356)
         );
  MUX2_X1 U7794 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6385), .S(n6391), .Z(n6255)
         );
  INV_X1 U7795 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6254) );
  INV_X1 U7796 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9740) );
  OR3_X1 U7797 ( .A1(n6255), .A2(n6254), .A3(n9740), .ZN(n6386) );
  INV_X1 U7798 ( .A(n6386), .ZN(n6256) );
  AOI21_X1 U7799 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n6270), .A(n6256), .ZN(
        n6374) );
  MUX2_X1 U7800 ( .A(n6373), .B(P2_REG2_REG_2__SCAN_IN), .S(n6372), .Z(n6257)
         );
  OR2_X1 U7801 ( .A1(n6374), .A2(n6257), .ZN(n6375) );
  NAND2_X1 U7802 ( .A1(n6372), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6331) );
  MUX2_X1 U7803 ( .A(n5832), .B(P2_REG2_REG_3__SCAN_IN), .S(n6271), .Z(n6330)
         );
  AOI21_X1 U7804 ( .B1(n6375), .B2(n6331), .A(n6330), .ZN(n6329) );
  NAND2_X1 U7805 ( .A1(n6271), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6343) );
  INV_X1 U7806 ( .A(n6343), .ZN(n6260) );
  MUX2_X1 U7807 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6258), .S(n6341), .Z(n6259)
         );
  OAI21_X1 U7808 ( .B1(n6329), .B2(n6260), .A(n6259), .ZN(n6346) );
  OAI21_X1 U7809 ( .B1(n6258), .B2(n6349), .A(n6346), .ZN(n6358) );
  XOR2_X1 U7810 ( .A(n6356), .B(n6358), .Z(n6284) );
  NAND2_X1 U7811 ( .A1(n6269), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8646) );
  OAI22_X1 U7812 ( .A1(n6261), .A2(n8646), .B1(n7515), .B2(n7963), .ZN(n6262)
         );
  INV_X1 U7813 ( .A(n6262), .ZN(n6267) );
  NAND2_X1 U7814 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  OR2_X1 U7815 ( .A1(n9765), .A2(n6265), .ZN(n6266) );
  NAND2_X1 U7816 ( .A1(n6274), .A2(n8222), .ZN(n6281) );
  INV_X1 U7817 ( .A(n8056), .ZN(n6268) );
  AND2_X1 U7818 ( .A1(n6281), .A2(n6268), .ZN(n9733) );
  AND2_X1 U7819 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6279) );
  XNOR2_X1 U7820 ( .A(n6270), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U7821 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6382) );
  NOR2_X1 U7822 ( .A1(n6381), .A2(n6382), .ZN(n6380) );
  AOI21_X1 U7823 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6270), .A(n6380), .ZN(
        n6369) );
  NOR2_X1 U7824 ( .A1(n6369), .A2(n6368), .ZN(n6367) );
  AOI21_X1 U7825 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n6372), .A(n6367), .ZN(
        n6326) );
  XNOR2_X1 U7826 ( .A(n6271), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6325) );
  INV_X1 U7827 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6272) );
  MUX2_X1 U7828 ( .A(n6272), .B(P2_REG1_REG_4__SCAN_IN), .S(n6341), .Z(n6337)
         );
  NAND2_X1 U7829 ( .A1(n6355), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6273) );
  OAI21_X1 U7830 ( .B1(n6355), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6273), .ZN(
        n6276) );
  INV_X1 U7831 ( .A(n6274), .ZN(n6275) );
  NOR2_X1 U7832 ( .A1(n6277), .A2(n6276), .ZN(n6350) );
  AOI211_X1 U7833 ( .C1(n6277), .C2(n6276), .A(n9731), .B(n6350), .ZN(n6278)
         );
  AOI211_X1 U7834 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9738), .A(n6279), .B(
        n6278), .ZN(n6283) );
  NAND2_X1 U7835 ( .A1(n8285), .A2(n6355), .ZN(n6282) );
  OAI211_X1 U7836 ( .C1(n6284), .C2(n8282), .A(n6283), .B(n6282), .ZN(P2_U3250) );
  INV_X1 U7837 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9727) );
  NOR2_X1 U7838 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6292), .ZN(n6286) );
  AOI22_X1 U7839 ( .A1(n9577), .A2(n9727), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6289), .ZN(n9571) );
  NOR2_X1 U7840 ( .A1(n9572), .A2(n9571), .ZN(n9570) );
  AOI21_X1 U7841 ( .B1(n6289), .B2(n9727), .A(n9570), .ZN(n6288) );
  INV_X1 U7842 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7117) );
  AOI22_X1 U7843 ( .A1(n6578), .A2(n7117), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6575), .ZN(n6287) );
  NOR2_X1 U7844 ( .A1(n6288), .A2(n6287), .ZN(n6574) );
  AOI21_X1 U7845 ( .B1(n6288), .B2(n6287), .A(n6574), .ZN(n6304) );
  INV_X1 U7846 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7847 ( .A1(n9577), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6295) );
  INV_X1 U7848 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6290) );
  MUX2_X1 U7849 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6290), .S(n6289), .Z(n6291)
         );
  INV_X1 U7850 ( .A(n6291), .ZN(n9580) );
  NOR2_X1 U7851 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6292), .ZN(n6294) );
  NOR2_X1 U7852 ( .A1(n6294), .A2(n6293), .ZN(n9581) );
  NAND2_X1 U7853 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  NAND2_X1 U7854 ( .A1(n6295), .A2(n9579), .ZN(n6297) );
  INV_X1 U7855 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7195) );
  MUX2_X1 U7856 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7195), .S(n6578), .Z(n6296)
         );
  NAND2_X1 U7857 ( .A1(n6296), .A2(n6297), .ZN(n6579) );
  OAI211_X1 U7858 ( .C1(n6297), .C2(n6296), .A(n9598), .B(n6579), .ZN(n6300)
         );
  NOR2_X1 U7859 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6298), .ZN(n6822) );
  AOI21_X1 U7860 ( .B1(n9578), .B2(n6578), .A(n6822), .ZN(n6299) );
  OAI211_X1 U7861 ( .C1(n9584), .C2(n6301), .A(n6300), .B(n6299), .ZN(n6302)
         );
  INV_X1 U7862 ( .A(n6302), .ZN(n6303) );
  OAI21_X1 U7863 ( .B1(n6304), .B2(n9573), .A(n6303), .ZN(P1_U3251) );
  INV_X1 U7864 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U7865 ( .A1(n9280), .A2(P1_U4006), .ZN(n6305) );
  OAI21_X1 U7866 ( .B1(n6959), .B2(P1_U4006), .A(n6305), .ZN(P1_U3576) );
  INV_X1 U7867 ( .A(n6306), .ZN(n6308) );
  AOI22_X1 U7868 ( .A1(n6904), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9429), .ZN(n6307) );
  OAI21_X1 U7869 ( .B1(n6308), .B2(n9431), .A(n6307), .ZN(P1_U3340) );
  INV_X1 U7870 ( .A(n7376), .ZN(n7250) );
  OAI222_X1 U7871 ( .A1(n8641), .A2(n6309), .B1(n8016), .B2(n6308), .C1(n7250), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  XNOR2_X1 U7872 ( .A(n6311), .B(n6310), .ZN(n6312) );
  NAND2_X1 U7873 ( .A1(n6312), .A2(n8683), .ZN(n6317) );
  NAND2_X1 U7874 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9080) );
  INV_X1 U7875 ( .A(n9080), .ZN(n6315) );
  OAI22_X1 U7876 ( .A1(n8730), .A2(n6313), .B1(n6676), .B2(n8706), .ZN(n6314)
         );
  AOI211_X1 U7877 ( .C1(n8664), .C2(n9632), .A(n6315), .B(n6314), .ZN(n6316)
         );
  OAI211_X1 U7878 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n7128), .A(n6317), .B(
        n6316), .ZN(P1_U3216) );
  INV_X1 U7879 ( .A(n6916), .ZN(n6322) );
  AOI22_X1 U7880 ( .A1(n7210), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9429), .ZN(n6318) );
  OAI21_X1 U7881 ( .B1(n6322), .B2(n9431), .A(n6318), .ZN(P1_U3339) );
  INV_X1 U7882 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7883 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  NAND2_X1 U7884 ( .A1(n6321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6448) );
  XNOR2_X1 U7885 ( .A(n6448), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7577) );
  INV_X1 U7886 ( .A(n7577), .ZN(n7572) );
  OAI222_X1 U7887 ( .A1(n8641), .A2(n6323), .B1(n8016), .B2(n6322), .C1(n7572), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NOR2_X1 U7888 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5830), .ZN(n6328) );
  AOI211_X1 U7889 ( .C1(n6326), .C2(n6325), .A(n6324), .B(n9731), .ZN(n6327)
         );
  AOI211_X1 U7890 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9738), .A(n6328), .B(
        n6327), .ZN(n6334) );
  INV_X1 U7891 ( .A(n6329), .ZN(n6344) );
  NAND3_X1 U7892 ( .A1(n6375), .A2(n6331), .A3(n6330), .ZN(n6332) );
  NAND3_X1 U7893 ( .A1(n9735), .A2(n6344), .A3(n6332), .ZN(n6333) );
  OAI211_X1 U7894 ( .C1(n9730), .C2(n6335), .A(n6334), .B(n6333), .ZN(P2_U3248) );
  NAND2_X1 U7895 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6711) );
  INV_X1 U7896 ( .A(n6711), .ZN(n6340) );
  AOI211_X1 U7897 ( .C1(n6338), .C2(n6337), .A(n6336), .B(n9731), .ZN(n6339)
         );
  AOI211_X1 U7898 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9738), .A(n6340), .B(
        n6339), .ZN(n6348) );
  MUX2_X1 U7899 ( .A(n6258), .B(P2_REG2_REG_4__SCAN_IN), .S(n6341), .Z(n6342)
         );
  NAND3_X1 U7900 ( .A1(n6344), .A2(n6343), .A3(n6342), .ZN(n6345) );
  NAND3_X1 U7901 ( .A1(n9735), .A2(n6346), .A3(n6345), .ZN(n6347) );
  OAI211_X1 U7902 ( .C1(n9730), .C2(n6349), .A(n6348), .B(n6347), .ZN(P2_U3249) );
  AND2_X1 U7903 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8181) );
  AOI21_X1 U7904 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n6355), .A(n6350), .ZN(
        n6353) );
  NAND2_X1 U7905 ( .A1(n6398), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7906 ( .B1(n6398), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6351), .ZN(
        n6352) );
  NOR2_X1 U7907 ( .A1(n6353), .A2(n6352), .ZN(n6392) );
  AOI211_X1 U7908 ( .C1(n6353), .C2(n6352), .A(n6392), .B(n9731), .ZN(n6354)
         );
  AOI211_X1 U7909 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9738), .A(n8181), .B(
        n6354), .ZN(n6364) );
  NAND2_X1 U7910 ( .A1(n6355), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6360) );
  INV_X1 U7911 ( .A(n6356), .ZN(n6357) );
  NAND2_X1 U7912 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X1 U7913 ( .A1(n6360), .A2(n6359), .ZN(n6362) );
  MUX2_X1 U7914 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n8512), .S(n6398), .Z(n6361)
         );
  NAND2_X1 U7915 ( .A1(n6361), .A2(n6362), .ZN(n6399) );
  OAI211_X1 U7916 ( .C1(n6362), .C2(n6361), .A(n9735), .B(n6399), .ZN(n6363)
         );
  OAI211_X1 U7917 ( .C1(n9730), .C2(n6365), .A(n6364), .B(n6363), .ZN(P2_U3251) );
  INV_X1 U7918 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6366) );
  NOR2_X1 U7919 ( .A1(n6366), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6371) );
  AOI211_X1 U7920 ( .C1(n6369), .C2(n6368), .A(n6367), .B(n9731), .ZN(n6370)
         );
  AOI211_X1 U7921 ( .C1(P2_ADDR_REG_2__SCAN_IN), .C2(n9738), .A(n6371), .B(
        n6370), .ZN(n6379) );
  MUX2_X1 U7922 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6373), .S(n6372), .Z(n6377)
         );
  INV_X1 U7923 ( .A(n6374), .ZN(n6376) );
  OAI211_X1 U7924 ( .C1(n6377), .C2(n6376), .A(n9735), .B(n6375), .ZN(n6378)
         );
  OAI211_X1 U7925 ( .C1(n9730), .C2(n4478), .A(n6379), .B(n6378), .ZN(P2_U3247) );
  INV_X1 U7926 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U7927 ( .A1(n6841), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6384) );
  AOI211_X1 U7928 ( .C1(n6382), .C2(n6381), .A(n6380), .B(n9731), .ZN(n6383)
         );
  AOI211_X1 U7929 ( .C1(P2_ADDR_REG_1__SCAN_IN), .C2(n9738), .A(n6384), .B(
        n6383), .ZN(n6390) );
  NOR2_X1 U7930 ( .A1(n9740), .A2(n6254), .ZN(n6388) );
  INV_X1 U7931 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6385) );
  MUX2_X1 U7932 ( .A(n6385), .B(P2_REG2_REG_1__SCAN_IN), .S(n6391), .Z(n6387)
         );
  OAI211_X1 U7933 ( .C1(n6388), .C2(n6387), .A(n9735), .B(n6386), .ZN(n6389)
         );
  OAI211_X1 U7934 ( .C1(n9730), .C2(n6391), .A(n6390), .B(n6389), .ZN(P2_U3246) );
  INV_X1 U7935 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8115) );
  NOR2_X1 U7936 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8115), .ZN(n6397) );
  AOI21_X1 U7937 ( .B1(n6398), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6392), .ZN(
        n6395) );
  NAND2_X1 U7938 ( .A1(n6472), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6393) );
  OAI21_X1 U7939 ( .B1(n6472), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6393), .ZN(
        n6394) );
  NOR2_X1 U7940 ( .A1(n6395), .A2(n6394), .ZN(n6466) );
  AOI211_X1 U7941 ( .C1(n6395), .C2(n6394), .A(n6466), .B(n9731), .ZN(n6396)
         );
  AOI211_X1 U7942 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9738), .A(n6397), .B(
        n6396), .ZN(n6405) );
  NAND2_X1 U7943 ( .A1(n6398), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U7944 ( .A1(n6400), .A2(n6399), .ZN(n6403) );
  MUX2_X1 U7945 ( .A(n5879), .B(P2_REG2_REG_7__SCAN_IN), .S(n6472), .Z(n6401)
         );
  INV_X1 U7946 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U7947 ( .A1(n6402), .A2(n6403), .ZN(n6473) );
  OAI211_X1 U7948 ( .C1(n6403), .C2(n6402), .A(n9735), .B(n6473), .ZN(n6404)
         );
  OAI211_X1 U7949 ( .C1(n9730), .C2(n6406), .A(n6405), .B(n6404), .ZN(P2_U3252) );
  NAND2_X1 U7950 ( .A1(n6407), .A2(n6735), .ZN(n6408) );
  OR2_X1 U7951 ( .A1(n6408), .A2(n9765), .ZN(n6409) );
  NOR2_X1 U7952 ( .A1(n6739), .A2(n6409), .ZN(n6411) );
  INV_X1 U7953 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U7954 ( .A1(n6412), .A2(n7965), .ZN(n7836) );
  NAND2_X1 U7955 ( .A1(n6419), .A2(n7836), .ZN(n6835) );
  NAND2_X1 U7956 ( .A1(n6835), .A2(n6846), .ZN(n6845) );
  INV_X1 U7957 ( .A(n7965), .ZN(n9813) );
  NAND2_X1 U7958 ( .A1(n6412), .A2(n9813), .ZN(n6413) );
  NAND2_X1 U7959 ( .A1(n6845), .A2(n6413), .ZN(n6744) );
  NAND2_X1 U7960 ( .A1(n6696), .A2(n8170), .ZN(n7838) );
  NAND2_X1 U7961 ( .A1(n7838), .A2(n7839), .ZN(n7789) );
  NAND2_X1 U7962 ( .A1(n6744), .A2(n7789), .ZN(n6743) );
  NAND2_X1 U7963 ( .A1(n6696), .A2(n9820), .ZN(n6414) );
  NAND2_X1 U7964 ( .A1(n6743), .A2(n6414), .ZN(n6415) );
  NAND2_X1 U7965 ( .A1(n6790), .A2(n6692), .ZN(n6858) );
  INV_X1 U7966 ( .A(n6790), .ZN(n8221) );
  INV_X1 U7967 ( .A(n6692), .ZN(n6802) );
  NAND2_X1 U7968 ( .A1(n8221), .A2(n6802), .ZN(n7842) );
  NAND2_X1 U7969 ( .A1(n6858), .A2(n7842), .ZN(n6422) );
  NAND2_X1 U7970 ( .A1(n6415), .A2(n6422), .ZN(n6781) );
  OR2_X1 U7971 ( .A1(n6415), .A2(n6422), .ZN(n6416) );
  NAND2_X1 U7972 ( .A1(n6781), .A2(n6416), .ZN(n6426) );
  INV_X1 U7973 ( .A(n6426), .ZN(n6803) );
  OR3_X1 U7974 ( .A1(n7960), .A2(n7956), .A3(n8499), .ZN(n9849) );
  XNOR2_X1 U7975 ( .A(n7960), .B(n6742), .ZN(n6417) );
  NAND2_X1 U7976 ( .A1(n6417), .A2(n8499), .ZN(n8532) );
  INV_X1 U7977 ( .A(n8532), .ZN(n6427) );
  OAI22_X1 U7978 ( .A1(n6696), .A2(n8498), .B1(n6849), .B2(n8496), .ZN(n6425)
         );
  NAND2_X1 U7979 ( .A1(n7831), .A2(n6419), .ZN(n6750) );
  INV_X1 U7980 ( .A(n6750), .ZN(n6421) );
  INV_X1 U7981 ( .A(n7789), .ZN(n6420) );
  INV_X1 U7982 ( .A(n6422), .ZN(n7834) );
  NAND3_X1 U7983 ( .A1(n6748), .A2(n6422), .A3(n7838), .ZN(n6423) );
  NAND2_X1 U7984 ( .A1(n7960), .A2(n9753), .ZN(n7957) );
  NAND2_X1 U7985 ( .A1(n7956), .A2(n7829), .ZN(n7786) );
  INV_X1 U7986 ( .A(n8511), .ZN(n9759) );
  AOI21_X1 U7987 ( .B1(n6859), .B2(n6423), .A(n9759), .ZN(n6424) );
  AOI211_X1 U7988 ( .C1(n6427), .C2(n6426), .A(n6425), .B(n6424), .ZN(n6807)
         );
  NAND2_X1 U7989 ( .A1(n9817), .A2(n6692), .ZN(n6428) );
  AND2_X1 U7990 ( .A1(n6784), .A2(n6428), .ZN(n6798) );
  AOI22_X1 U7991 ( .A1(n6798), .A2(n9837), .B1(n9836), .B2(n6692), .ZN(n6429)
         );
  OAI211_X1 U7992 ( .C1(n6803), .C2(n9849), .A(n6807), .B(n6429), .ZN(n6434)
         );
  NAND2_X1 U7993 ( .A1(n6434), .A2(n9906), .ZN(n6430) );
  OAI21_X1 U7994 ( .B1(n9906), .B2(n6431), .A(n6430), .ZN(P2_U3523) );
  NAND2_X1 U7995 ( .A1(n6434), .A2(n9888), .ZN(n6435) );
  OAI21_X1 U7996 ( .B1(n9888), .B2(n5831), .A(n6435), .ZN(P2_U3460) );
  XOR2_X1 U7997 ( .A(n6438), .B(n6437), .Z(n6439) );
  XNOR2_X1 U7998 ( .A(n6436), .B(n6439), .ZN(n6446) );
  NAND2_X1 U7999 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9568) );
  INV_X1 U8000 ( .A(n9568), .ZN(n6440) );
  AOI21_X1 U8001 ( .B1(n8664), .B2(n9064), .A(n6440), .ZN(n6443) );
  NAND2_X1 U8002 ( .A1(n8726), .A2(n6441), .ZN(n6442) );
  OAI211_X1 U8003 ( .C1(n9617), .C2(n8706), .A(n6443), .B(n6442), .ZN(n6444)
         );
  AOI21_X1 U8004 ( .B1(n6672), .B2(n8709), .A(n6444), .ZN(n6445) );
  OAI21_X1 U8005 ( .B1(n6446), .B2(n8716), .A(n6445), .ZN(P1_U3237) );
  INV_X1 U8006 ( .A(n7063), .ZN(n6452) );
  INV_X1 U8007 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8008 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND2_X1 U8009 ( .A1(n6449), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6450) );
  XNOR2_X1 U8010 ( .A(n6450), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8230) );
  INV_X1 U8011 ( .A(n8230), .ZN(n8224) );
  OAI222_X1 U8012 ( .A1(n8641), .A2(n6451), .B1(n8016), .B2(n6452), .C1(
        P2_U3152), .C2(n8224), .ZN(P2_U3343) );
  OAI222_X1 U8013 ( .A1(n7481), .A2(n6453), .B1(n9431), .B2(n6452), .C1(
        P1_U3084), .C2(n7359), .ZN(P1_U3338) );
  NAND2_X1 U8014 ( .A1(n6564), .A2(n6454), .ZN(n6458) );
  XNOR2_X1 U8015 ( .A(n6456), .B(n6455), .ZN(n6457) );
  XNOR2_X1 U8016 ( .A(n6458), .B(n6457), .ZN(n6465) );
  OR2_X1 U8017 ( .A1(n6676), .A2(n8723), .ZN(n6461) );
  INV_X1 U8018 ( .A(n6459), .ZN(n6460) );
  OAI211_X1 U8019 ( .C1(n8706), .C2(n6681), .A(n6461), .B(n6460), .ZN(n6462)
         );
  AOI21_X1 U8020 ( .B1(n9676), .B2(n8709), .A(n6462), .ZN(n6464) );
  NAND2_X1 U8021 ( .A1(n8726), .A2(n9315), .ZN(n6463) );
  OAI211_X1 U8022 ( .C1(n6465), .C2(n8716), .A(n6464), .B(n6463), .ZN(P1_U3225) );
  NOR2_X1 U8023 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6546), .ZN(n6471) );
  INV_X1 U8024 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6467) );
  MUX2_X1 U8025 ( .A(n6467), .B(P2_REG1_REG_8__SCAN_IN), .S(n6601), .Z(n6468)
         );
  AOI211_X1 U8026 ( .C1(n6469), .C2(n6468), .A(n6600), .B(n9731), .ZN(n6470)
         );
  AOI211_X1 U8027 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9738), .A(n6471), .B(
        n6470), .ZN(n6478) );
  NAND2_X1 U8028 ( .A1(n6472), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U8029 ( .A1(n6474), .A2(n6473), .ZN(n6476) );
  MUX2_X1 U8030 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6870), .S(n6601), .Z(n6475)
         );
  NAND2_X1 U8031 ( .A1(n6476), .A2(n6475), .ZN(n6608) );
  OAI211_X1 U8032 ( .C1(n6476), .C2(n6475), .A(n9735), .B(n6608), .ZN(n6477)
         );
  OAI211_X1 U8033 ( .C1(n9730), .C2(n6609), .A(n6478), .B(n6477), .ZN(P2_U3253) );
  INV_X1 U8034 ( .A(n6479), .ZN(n6481) );
  NAND3_X1 U8035 ( .A1(n6481), .A2(n6480), .A3(n7112), .ZN(n6685) );
  AOI22_X1 U8036 ( .A1(n9648), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9314), .ZN(n6485) );
  NOR2_X1 U8037 ( .A1(n9706), .A2(n5398), .ZN(n6483) );
  OAI21_X1 U8038 ( .B1(n9316), .B2(n9612), .A(n6509), .ZN(n6484) );
  OAI211_X1 U8039 ( .C1(n6486), .C2(n9648), .A(n6485), .B(n6484), .ZN(P1_U3291) );
  NAND2_X1 U8040 ( .A1(n6488), .A2(n6509), .ZN(n9628) );
  NAND2_X1 U8041 ( .A1(n6496), .A2(n9628), .ZN(n6491) );
  INV_X1 U8042 ( .A(n6489), .ZN(n6497) );
  NAND2_X1 U8043 ( .A1(n6497), .A2(n6487), .ZN(n6490) );
  NAND2_X1 U8044 ( .A1(n6491), .A2(n6490), .ZN(n6525) );
  NAND2_X1 U8045 ( .A1(n6525), .A2(n6526), .ZN(n6494) );
  INV_X1 U8046 ( .A(n9632), .ZN(n6505) );
  NAND2_X1 U8047 ( .A1(n6505), .A2(n6492), .ZN(n6493) );
  NAND2_X1 U8048 ( .A1(n6494), .A2(n6493), .ZN(n6616) );
  NAND2_X1 U8049 ( .A1(n6620), .A2(n6513), .ZN(n9003) );
  NAND2_X1 U8050 ( .A1(n9065), .A2(n6313), .ZN(n8953) );
  NAND2_X1 U8051 ( .A1(n9003), .A2(n8953), .ZN(n6615) );
  XNOR2_X1 U8052 ( .A(n6616), .B(n8876), .ZN(n9660) );
  NAND2_X1 U8053 ( .A1(n6495), .A2(n5398), .ZN(n6683) );
  INV_X1 U8054 ( .A(n6683), .ZN(n9645) );
  NAND2_X1 U8055 ( .A1(n9646), .A2(n9645), .ZN(n7299) );
  NAND2_X1 U8056 ( .A1(n8874), .A2(n9629), .ZN(n6499) );
  NAND2_X1 U8057 ( .A1(n6497), .A2(n4643), .ZN(n6498) );
  NAND2_X1 U8058 ( .A1(n6499), .A2(n6498), .ZN(n6530) );
  INV_X1 U8059 ( .A(n6526), .ZN(n8877) );
  NAND2_X1 U8060 ( .A1(n6530), .A2(n8877), .ZN(n6501) );
  NAND2_X1 U8061 ( .A1(n6505), .A2(n4970), .ZN(n6500) );
  NAND2_X1 U8062 ( .A1(n6501), .A2(n6500), .ZN(n6621) );
  XNOR2_X1 U8063 ( .A(n6621), .B(n8876), .ZN(n6507) );
  NAND2_X1 U8064 ( .A1(n6502), .A2(n5398), .ZN(n6503) );
  OR2_X1 U8065 ( .A1(n4926), .A2(n8912), .ZN(n8868) );
  INV_X1 U8066 ( .A(n9633), .ZN(n9618) );
  OAI22_X1 U8067 ( .A1(n6505), .A2(n9618), .B1(n6676), .B2(n9616), .ZN(n6506)
         );
  AOI21_X1 U8068 ( .B1(n6507), .B2(n9313), .A(n6506), .ZN(n6508) );
  OAI21_X1 U8069 ( .B1(n9660), .B2(n7290), .A(n6508), .ZN(n9662) );
  NAND2_X1 U8070 ( .A1(n9662), .A2(n9646), .ZN(n6515) );
  OAI22_X1 U8071 ( .A1(n9646), .A2(n6151), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9641), .ZN(n6512) );
  OR2_X1 U8072 ( .A1(n6528), .A2(n6313), .ZN(n6510) );
  NAND2_X1 U8073 ( .A1(n6631), .A2(n6510), .ZN(n9661) );
  INV_X1 U8074 ( .A(n9612), .ZN(n9148) );
  NOR2_X1 U8075 ( .A1(n9661), .A2(n9148), .ZN(n6511) );
  AOI211_X1 U8076 ( .C1(n9316), .C2(n6513), .A(n6512), .B(n6511), .ZN(n6514)
         );
  OAI211_X1 U8077 ( .C1(n9660), .C2(n7299), .A(n6515), .B(n6514), .ZN(P1_U3288) );
  XNOR2_X1 U8078 ( .A(n6516), .B(n6517), .ZN(n6523) );
  AOI21_X1 U8079 ( .B1(n8664), .B2(n9311), .A(n6518), .ZN(n6520) );
  NAND2_X1 U8080 ( .A1(n8726), .A2(n6686), .ZN(n6519) );
  OAI211_X1 U8081 ( .C1(n7225), .C2(n8706), .A(n6520), .B(n6519), .ZN(n6521)
         );
  AOI21_X1 U8082 ( .B1(n6889), .B2(n8709), .A(n6521), .ZN(n6522) );
  OAI21_X1 U8083 ( .B1(n6523), .B2(n8716), .A(n6522), .ZN(P1_U3211) );
  INV_X1 U8084 ( .A(n7304), .ZN(n6572) );
  AOI22_X1 U8085 ( .A1(n9113), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9429), .ZN(n6524) );
  OAI21_X1 U8086 ( .B1(n6572), .B2(n9431), .A(n6524), .ZN(P1_U3336) );
  XNOR2_X1 U8087 ( .A(n6525), .B(n6526), .ZN(n9658) );
  INV_X1 U8088 ( .A(n7299), .ZN(n9613) );
  NOR2_X1 U8089 ( .A1(n9639), .A2(n6492), .ZN(n6527) );
  OR2_X1 U8090 ( .A1(n6528), .A2(n6527), .ZN(n9655) );
  AOI22_X1 U8091 ( .A1(n9316), .A2(n4970), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9314), .ZN(n6529) );
  OAI21_X1 U8092 ( .B1(n9148), .B2(n9655), .A(n6529), .ZN(n6537) );
  XNOR2_X1 U8093 ( .A(n6530), .B(n8877), .ZN(n6533) );
  NAND2_X1 U8094 ( .A1(n6489), .A2(n9633), .ZN(n6531) );
  OAI21_X1 U8095 ( .B1(n6620), .B2(n9616), .A(n6531), .ZN(n6532) );
  AOI21_X1 U8096 ( .B1(n6533), .B2(n9313), .A(n6532), .ZN(n6535) );
  INV_X1 U8097 ( .A(n7290), .ZN(n9630) );
  NAND2_X1 U8098 ( .A1(n9658), .A2(n9630), .ZN(n6534) );
  NAND2_X1 U8099 ( .A1(n6535), .A2(n6534), .ZN(n9656) );
  MUX2_X1 U8100 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9656), .S(n9646), .Z(n6536)
         );
  AOI211_X1 U8101 ( .C1(n9658), .C2(n9613), .A(n6537), .B(n6536), .ZN(n6538)
         );
  INV_X1 U8102 ( .A(n6538), .ZN(P1_U3289) );
  INV_X1 U8103 ( .A(n9100), .ZN(n7366) );
  INV_X1 U8104 ( .A(n7067), .ZN(n6544) );
  OAI222_X1 U8105 ( .A1(P1_U3084), .A2(n7366), .B1(n7552), .B2(n6544), .C1(
        n10072), .C2(n7481), .ZN(P1_U3337) );
  NAND2_X1 U8106 ( .A1(n6539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6540) );
  MUX2_X1 U8107 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6540), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6543) );
  AND2_X1 U8108 ( .A1(n6543), .A2(n6542), .ZN(n8250) );
  INV_X1 U8109 ( .A(n8250), .ZN(n8240) );
  OAI222_X1 U8110 ( .A1(n8641), .A2(n10103), .B1(n8016), .B2(n6544), .C1(n8240), .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8111 ( .A(n6545), .ZN(n6869) );
  OAI22_X1 U8112 ( .A1(n8162), .A2(n6869), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6546), .ZN(n6548) );
  OAI22_X1 U8113 ( .A1(n8179), .A2(n8200), .B1(n8202), .B2(n7005), .ZN(n6547)
         );
  AOI211_X1 U8114 ( .C1(n6960), .C2(n4315), .A(n6548), .B(n6547), .ZN(n6558)
         );
  AND2_X1 U8115 ( .A1(n6550), .A2(n6549), .ZN(n8110) );
  INV_X1 U8116 ( .A(n6551), .ZN(n6552) );
  AOI21_X1 U8117 ( .B1(n8110), .B2(n6552), .A(n8196), .ZN(n6556) );
  INV_X1 U8118 ( .A(n6553), .ZN(n6554) );
  NOR3_X1 U8119 ( .A1(n8189), .A2(n6554), .A3(n8179), .ZN(n6555) );
  OAI21_X1 U8120 ( .B1(n6556), .B2(n6555), .A(n6637), .ZN(n6557) );
  NAND2_X1 U8121 ( .A1(n6558), .A2(n6557), .ZN(P2_U3223) );
  AOI22_X1 U8122 ( .A1(n8709), .A2(n9666), .B1(n8721), .B2(n9064), .ZN(n6560)
         );
  NAND2_X1 U8123 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n9556) );
  OAI211_X1 U8124 ( .C1(n6620), .C2(n8723), .A(n6560), .B(n9556), .ZN(n6568)
         );
  NAND2_X1 U8125 ( .A1(n6562), .A2(n6563), .ZN(n6566) );
  INV_X1 U8126 ( .A(n6564), .ZN(n6565) );
  AOI211_X1 U8127 ( .C1(n6561), .C2(n6566), .A(n8716), .B(n6565), .ZN(n6567)
         );
  AOI211_X1 U8128 ( .C1(n6632), .C2(n8726), .A(n6568), .B(n6567), .ZN(n6569)
         );
  INV_X1 U8129 ( .A(n6569), .ZN(P1_U3228) );
  NAND2_X1 U8130 ( .A1(n6542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U8131 ( .A(n6570), .B(P2_IR_REG_31__SCAN_IN), .S(n10083), .Z(n6571)
         );
  NAND2_X1 U8132 ( .A1(n6571), .A2(n6652), .ZN(n8258) );
  OAI222_X1 U8133 ( .A1(n8641), .A2(n6573), .B1(n8016), .B2(n6572), .C1(n8258), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  AOI21_X1 U8134 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9591), .A(n9596), .ZN(
        n6576) );
  NOR2_X1 U8135 ( .A1(n9591), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9592) );
  MUX2_X1 U8136 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n4398), .S(n6661), .Z(n6577)
         );
  NAND2_X1 U8137 ( .A1(n6577), .A2(n9594), .ZN(n6657) );
  OAI21_X1 U8138 ( .B1(n9594), .B2(n6577), .A(n6657), .ZN(n6588) );
  NAND2_X1 U8139 ( .A1(n6578), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8140 ( .A1(n6580), .A2(n6579), .ZN(n9601) );
  INV_X1 U8141 ( .A(n9601), .ZN(n6581) );
  INV_X1 U8142 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10068) );
  NOR2_X1 U8143 ( .A1(n6581), .A2(n10068), .ZN(n6582) );
  NAND2_X1 U8144 ( .A1(n6661), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6583) );
  OAI21_X1 U8145 ( .B1(n6661), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6583), .ZN(
        n6584) );
  AOI211_X1 U8146 ( .C1(n9599), .C2(n6584), .A(n6660), .B(n9553), .ZN(n6587)
         );
  INV_X1 U8147 ( .A(n9584), .ZN(n9589) );
  NAND2_X1 U8148 ( .A1(n9589), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U8149 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7139) );
  OAI211_X1 U8150 ( .C1(n9587), .C2(n4399), .A(n6585), .B(n7139), .ZN(n6586)
         );
  AOI211_X1 U8151 ( .C1(n6588), .C2(n9593), .A(n6587), .B(n6586), .ZN(n6589)
         );
  INV_X1 U8152 ( .A(n6589), .ZN(P1_U3253) );
  XOR2_X1 U8153 ( .A(n6592), .B(n6591), .Z(n6593) );
  XNOR2_X1 U8154 ( .A(n6590), .B(n6593), .ZN(n6599) );
  INV_X1 U8155 ( .A(n9061), .ZN(n7104) );
  INV_X1 U8156 ( .A(n9617), .ZN(n9063) );
  AOI21_X1 U8157 ( .B1(n8664), .B2(n9063), .A(n6594), .ZN(n6596) );
  NAND2_X1 U8158 ( .A1(n8726), .A2(n6886), .ZN(n6595) );
  OAI211_X1 U8159 ( .C1(n7104), .C2(n8706), .A(n6596), .B(n6595), .ZN(n6597)
         );
  AOI21_X1 U8160 ( .B1(n7096), .B2(n8709), .A(n6597), .ZN(n6598) );
  OAI21_X1 U8161 ( .B1(n6599), .B2(n8716), .A(n6598), .ZN(P1_U3219) );
  NAND2_X1 U8162 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6642) );
  INV_X1 U8163 ( .A(n6642), .ZN(n6606) );
  INV_X1 U8164 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6602) );
  MUX2_X1 U8165 ( .A(n6602), .B(P2_REG1_REG_9__SCAN_IN), .S(n6771), .Z(n6603)
         );
  AOI211_X1 U8166 ( .C1(n6604), .C2(n6603), .A(n6765), .B(n9731), .ZN(n6605)
         );
  AOI211_X1 U8167 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9738), .A(n6606), .B(
        n6605), .ZN(n6613) );
  MUX2_X1 U8168 ( .A(n7049), .B(P2_REG2_REG_9__SCAN_IN), .S(n6771), .Z(n6607)
         );
  INV_X1 U8169 ( .A(n6607), .ZN(n6611) );
  OAI21_X1 U8170 ( .B1(n6870), .B2(n6609), .A(n6608), .ZN(n6610) );
  NAND2_X1 U8171 ( .A1(n6611), .A2(n6610), .ZN(n6772) );
  OAI211_X1 U8172 ( .C1(n6611), .C2(n6610), .A(n9735), .B(n6772), .ZN(n6612)
         );
  OAI211_X1 U8173 ( .C1(n9730), .C2(n6614), .A(n6613), .B(n6612), .ZN(P2_U3254) );
  NAND2_X1 U8174 ( .A1(n6616), .A2(n6615), .ZN(n6618) );
  NAND2_X1 U8175 ( .A1(n6620), .A2(n6313), .ZN(n6617) );
  NAND2_X1 U8176 ( .A1(n6618), .A2(n6617), .ZN(n6674) );
  NAND2_X1 U8177 ( .A1(n6676), .A2(n9666), .ZN(n8944) );
  INV_X1 U8178 ( .A(n6676), .ZN(n9310) );
  NAND2_X1 U8179 ( .A1(n8944), .A2(n9307), .ZN(n8873) );
  XNOR2_X1 U8180 ( .A(n6674), .B(n8873), .ZN(n6628) );
  INV_X1 U8181 ( .A(n6628), .ZN(n9672) );
  OAI22_X1 U8182 ( .A1(n6620), .A2(n9618), .B1(n6619), .B2(n9616), .ZN(n6627)
         );
  NAND2_X1 U8183 ( .A1(n6621), .A2(n8876), .ZN(n6622) );
  INV_X1 U8184 ( .A(n8873), .ZN(n6624) );
  INV_X1 U8185 ( .A(n9308), .ZN(n6625) );
  AOI211_X1 U8186 ( .C1(n8873), .C2(n6623), .A(n8091), .B(n6625), .ZN(n6626)
         );
  AOI211_X1 U8187 ( .C1(n9630), .C2(n6628), .A(n6627), .B(n6626), .ZN(n9670)
         );
  MUX2_X1 U8188 ( .A(n6629), .B(n9670), .S(n9646), .Z(n6636) );
  OR2_X1 U8189 ( .A1(n6631), .A2(n9666), .ZN(n9321) );
  INV_X1 U8190 ( .A(n9321), .ZN(n6630) );
  AOI21_X1 U8191 ( .B1(n9666), .B2(n6631), .A(n6630), .ZN(n9668) );
  INV_X1 U8192 ( .A(n6632), .ZN(n6633) );
  OAI22_X1 U8193 ( .A1(n9623), .A2(n6675), .B1(n9641), .B2(n6633), .ZN(n6634)
         );
  AOI21_X1 U8194 ( .B1(n9668), .B2(n9612), .A(n6634), .ZN(n6635) );
  OAI211_X1 U8195 ( .C1(n9672), .C2(n7299), .A(n6636), .B(n6635), .ZN(P1_U3287) );
  INV_X1 U8196 ( .A(n6637), .ZN(n6640) );
  NOR3_X1 U8197 ( .A1(n8189), .A2(n6638), .A3(n7042), .ZN(n6639) );
  AOI21_X1 U8198 ( .B1(n6640), .B2(n8185), .A(n6639), .ZN(n6650) );
  INV_X1 U8199 ( .A(n7042), .ZN(n8218) );
  NAND2_X1 U8200 ( .A1(n8190), .A2(n8218), .ZN(n6644) );
  NAND2_X1 U8201 ( .A1(n8168), .A2(n8216), .ZN(n6643) );
  NAND2_X1 U8202 ( .A1(n8205), .A2(n7047), .ZN(n6641) );
  NAND4_X1 U8203 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6647)
         );
  NOR2_X1 U8204 ( .A1(n6645), .A2(n8196), .ZN(n6646) );
  AOI211_X1 U8205 ( .C1(n7055), .C2(n4315), .A(n6647), .B(n6646), .ZN(n6648)
         );
  OAI21_X1 U8206 ( .B1(n6650), .B2(n6649), .A(n6648), .ZN(P2_U3233) );
  INV_X1 U8207 ( .A(n7436), .ZN(n6655) );
  AOI22_X1 U8208 ( .A1(n9126), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9429), .ZN(n6651) );
  OAI21_X1 U8209 ( .B1(n6655), .B2(n9431), .A(n6651), .ZN(P1_U3335) );
  NAND2_X1 U8210 ( .A1(n6652), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6653) );
  XNOR2_X1 U8211 ( .A(n6653), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8276) );
  AOI22_X1 U8212 ( .A1(n8276), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8644), .ZN(n6654) );
  OAI21_X1 U8213 ( .B1(n6655), .B2(n8647), .A(n6654), .ZN(P2_U3340) );
  INV_X1 U8214 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6669) );
  INV_X1 U8215 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6656) );
  MUX2_X1 U8216 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6656), .S(n6904), .Z(n6659)
         );
  OAI21_X1 U8217 ( .B1(n6659), .B2(n6658), .A(n6900), .ZN(n6666) );
  NAND2_X1 U8218 ( .A1(n6904), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U8219 ( .B1(n6904), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6662), .ZN(
        n6663) );
  AOI211_X1 U8220 ( .C1(n6664), .C2(n6663), .A(n6903), .B(n9553), .ZN(n6665)
         );
  AOI21_X1 U8221 ( .B1(n9593), .B2(n6666), .A(n6665), .ZN(n6668) );
  AND2_X1 U8222 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7125) );
  AOI21_X1 U8223 ( .B1(n9578), .B2(n6904), .A(n7125), .ZN(n6667) );
  OAI211_X1 U8224 ( .C1(n9584), .C2(n6669), .A(n6668), .B(n6667), .ZN(P1_U3254) );
  NAND2_X1 U8225 ( .A1(n9064), .A2(n6670), .ZN(n8948) );
  NAND2_X1 U8226 ( .A1(n6681), .A2(n6672), .ZN(n8949) );
  NAND2_X1 U8227 ( .A1(n9311), .A2(n9683), .ZN(n8762) );
  NAND2_X1 U8228 ( .A1(n9617), .A2(n6889), .ZN(n6878) );
  NAND2_X1 U8229 ( .A1(n9063), .A2(n9692), .ZN(n8763) );
  NAND2_X1 U8230 ( .A1(n6878), .A2(n8763), .ZN(n8880) );
  XNOR2_X1 U8231 ( .A(n6876), .B(n8880), .ZN(n6673) );
  AOI222_X1 U8232 ( .A1(n9313), .A2(n6673), .B1(n9062), .B2(n9631), .C1(n9311), 
        .C2(n9633), .ZN(n9691) );
  NAND2_X1 U8233 ( .A1(n6674), .A2(n8873), .ZN(n6678) );
  NAND2_X1 U8234 ( .A1(n6676), .A2(n6675), .ZN(n6677) );
  NAND2_X1 U8235 ( .A1(n6678), .A2(n6677), .ZN(n9319) );
  NAND2_X1 U8236 ( .A1(n9064), .A2(n9676), .ZN(n6679) );
  NAND2_X1 U8237 ( .A1(n6681), .A2(n9683), .ZN(n6682) );
  NAND2_X1 U8238 ( .A1(n9606), .A2(n6682), .ZN(n6891) );
  XNOR2_X1 U8239 ( .A(n6891), .B(n8880), .ZN(n9694) );
  NAND2_X1 U8240 ( .A1(n7290), .A2(n6683), .ZN(n6684) );
  INV_X1 U8241 ( .A(n9306), .ZN(n9320) );
  AND2_X1 U8242 ( .A1(n9608), .A2(n9683), .ZN(n9610) );
  NAND2_X1 U8243 ( .A1(n9610), .A2(n9692), .ZN(n6884) );
  OAI211_X1 U8244 ( .C1(n9610), .C2(n9692), .A(n9667), .B(n6884), .ZN(n9690)
         );
  OR2_X1 U8245 ( .A1(n6685), .A2(n5398), .ZN(n7392) );
  AOI22_X1 U8246 ( .A1(n9648), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6686), .B2(
        n9314), .ZN(n6688) );
  NAND2_X1 U8247 ( .A1(n9316), .A2(n6889), .ZN(n6687) );
  OAI211_X1 U8248 ( .C1(n9690), .C2(n7392), .A(n6688), .B(n6687), .ZN(n6689)
         );
  AOI21_X1 U8249 ( .B1(n9694), .B2(n9320), .A(n6689), .ZN(n6690) );
  OAI21_X1 U8250 ( .B1(n9691), .B2(n9648), .A(n6690), .ZN(P1_U3284) );
  NAND2_X1 U8251 ( .A1(n4315), .A2(n6692), .ZN(n6693) );
  OAI21_X1 U8252 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5830), .A(n6693), .ZN(n6695) );
  OAI22_X1 U8253 ( .A1(n8202), .A2(n6849), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8162), .ZN(n6694) );
  AOI211_X1 U8254 ( .C1(n8190), .C2(n6691), .A(n6695), .B(n6694), .ZN(n6704)
         );
  NOR3_X1 U8255 ( .A1(n8189), .A2(n6697), .A3(n6696), .ZN(n6702) );
  INV_X1 U8256 ( .A(n6698), .ZN(n6699) );
  AOI21_X1 U8257 ( .B1(n8173), .B2(n6699), .A(n8196), .ZN(n6701) );
  OAI21_X1 U8258 ( .B1(n6702), .B2(n6701), .A(n6700), .ZN(n6703) );
  NAND2_X1 U8259 ( .A1(n6704), .A2(n6703), .ZN(P2_U3220) );
  OAI21_X1 U8260 ( .B1(n6707), .B2(n6700), .A(n6705), .ZN(n6715) );
  INV_X1 U8261 ( .A(n8189), .ZN(n8156) );
  INV_X1 U8262 ( .A(n6707), .ZN(n6709) );
  NAND3_X1 U8263 ( .A1(n8156), .A2(n6709), .A3(n6708), .ZN(n6710) );
  AOI21_X1 U8264 ( .B1(n6710), .B2(n8200), .A(n6790), .ZN(n6714) );
  AOI22_X1 U8265 ( .A1(n8168), .A2(n8507), .B1(n6783), .B2(n4315), .ZN(n6712)
         );
  OAI211_X1 U8266 ( .C1(n6793), .C2(n8162), .A(n6712), .B(n6711), .ZN(n6713)
         );
  AOI211_X1 U8267 ( .C1(n8185), .C2(n6715), .A(n6714), .B(n6713), .ZN(n6716)
         );
  INV_X1 U8268 ( .A(n6716), .ZN(P2_U3232) );
  INV_X1 U8269 ( .A(n6980), .ZN(n9873) );
  INV_X1 U8270 ( .A(n6717), .ZN(n6718) );
  AOI21_X1 U8271 ( .B1(n6757), .B2(n6718), .A(n8196), .ZN(n6722) );
  INV_X1 U8272 ( .A(n8216), .ZN(n7043) );
  NOR3_X1 U8273 ( .A1(n8189), .A2(n6719), .A3(n7043), .ZN(n6721) );
  OAI21_X1 U8274 ( .B1(n6722), .B2(n6721), .A(n6720), .ZN(n6725) );
  AND2_X1 U8275 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7031) );
  OAI22_X1 U8276 ( .A1(n7043), .A2(n8200), .B1(n8202), .B2(n6985), .ZN(n6723)
         );
  AOI211_X1 U8277 ( .C1(n8205), .C2(n6975), .A(n7031), .B(n6723), .ZN(n6724)
         );
  OAI211_X1 U8278 ( .C1(n9873), .C2(n8207), .A(n6725), .B(n6724), .ZN(P2_U3238) );
  INV_X1 U8279 ( .A(n6726), .ZN(n6727) );
  AOI21_X1 U8280 ( .B1(n6729), .B2(n6728), .A(n6727), .ZN(n6734) );
  AND2_X1 U8281 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9576) );
  AOI21_X1 U8282 ( .B1(n8664), .B2(n9062), .A(n9576), .ZN(n6731) );
  NAND2_X1 U8283 ( .A1(n8726), .A2(n7221), .ZN(n6730) );
  OAI211_X1 U8284 ( .C1(n7261), .C2(n8706), .A(n6731), .B(n6730), .ZN(n6732)
         );
  AOI21_X1 U8285 ( .B1(n9704), .B2(n8709), .A(n6732), .ZN(n6733) );
  OAI21_X1 U8286 ( .B1(n6734), .B2(n8716), .A(n6733), .ZN(P1_U3229) );
  INV_X1 U8287 ( .A(n6735), .ZN(n6736) );
  OR3_X1 U8288 ( .A1(n9765), .A2(n6737), .A3(n6736), .ZN(n6738) );
  NOR2_X1 U8289 ( .A1(n6739), .A2(n6738), .ZN(n6740) );
  NAND2_X1 U8290 ( .A1(n6741), .A2(n6740), .ZN(n6745) );
  OR2_X1 U8291 ( .A1(n6742), .A2(n8499), .ZN(n6800) );
  NAND2_X1 U8292 ( .A1(n8532), .A2(n6800), .ZN(n9762) );
  OAI21_X1 U8293 ( .B1(n6744), .B2(n7789), .A(n6743), .ZN(n9823) );
  OR2_X1 U8294 ( .A1(n6840), .A2(n9820), .ZN(n9818) );
  NAND3_X1 U8295 ( .A1(n8521), .A2(n9817), .A3(n9818), .ZN(n6747) );
  NAND2_X1 U8296 ( .A1(n9751), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6746) );
  OAI211_X1 U8297 ( .C1(n8469), .C2(n9820), .A(n6747), .B(n6746), .ZN(n6753)
         );
  INV_X1 U8298 ( .A(n6748), .ZN(n6749) );
  AOI21_X1 U8299 ( .B1(n7789), .B2(n6750), .A(n6749), .ZN(n6751) );
  OAI222_X1 U8300 ( .A1(n8498), .A2(n6412), .B1(n8496), .B2(n6790), .C1(n9759), 
        .C2(n6751), .ZN(n9821) );
  MUX2_X1 U8301 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9821), .S(n9763), .Z(n6752)
         );
  AOI211_X1 U8302 ( .C1(n8518), .C2(n9823), .A(n6753), .B(n6752), .ZN(n6754)
         );
  INV_X1 U8303 ( .A(n6754), .ZN(P2_U3294) );
  INV_X1 U8304 ( .A(n7514), .ZN(n6828) );
  OAI222_X1 U8305 ( .A1(n8641), .A2(n9961), .B1(n8016), .B2(n6828), .C1(n8499), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U8306 ( .A(n6755), .ZN(n7010) );
  INV_X1 U8307 ( .A(n7006), .ZN(n8215) );
  AOI22_X1 U8308 ( .A1(n8168), .A2(n8215), .B1(n8190), .B2(n8217), .ZN(n6756)
         );
  NAND2_X1 U8309 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n6764) );
  OAI211_X1 U8310 ( .C1(n7010), .C2(n8162), .A(n6756), .B(n6764), .ZN(n6762)
         );
  INV_X1 U8311 ( .A(n6757), .ZN(n6758) );
  AOI211_X1 U8312 ( .C1(n6760), .C2(n6759), .A(n8196), .B(n6758), .ZN(n6761)
         );
  AOI211_X1 U8313 ( .C1(n9863), .C2(n4315), .A(n6762), .B(n6761), .ZN(n6763)
         );
  INV_X1 U8314 ( .A(n6763), .ZN(P2_U3219) );
  INV_X1 U8315 ( .A(n6764), .ZN(n6770) );
  AOI21_X1 U8316 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n6771), .A(n6765), .ZN(
        n6768) );
  INV_X1 U8317 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6766) );
  MUX2_X1 U8318 ( .A(n6766), .B(P2_REG1_REG_10__SCAN_IN), .S(n7027), .Z(n6767)
         );
  NOR2_X1 U8319 ( .A1(n6768), .A2(n6767), .ZN(n7026) );
  AOI211_X1 U8320 ( .C1(n6768), .C2(n6767), .A(n7026), .B(n9731), .ZN(n6769)
         );
  AOI211_X1 U8321 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9738), .A(n6770), .B(
        n6769), .ZN(n6778) );
  NAND2_X1 U8322 ( .A1(n6771), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U8323 ( .A1(n6773), .A2(n6772), .ZN(n6776) );
  MUX2_X1 U8324 ( .A(n7011), .B(P2_REG2_REG_10__SCAN_IN), .S(n7027), .Z(n6774)
         );
  INV_X1 U8325 ( .A(n6774), .ZN(n6775) );
  NAND2_X1 U8326 ( .A1(n6775), .A2(n6776), .ZN(n7020) );
  OAI211_X1 U8327 ( .C1(n6776), .C2(n6775), .A(n9735), .B(n7020), .ZN(n6777)
         );
  OAI211_X1 U8328 ( .C1(n9730), .C2(n6779), .A(n6778), .B(n6777), .ZN(P2_U3255) );
  NAND2_X1 U8329 ( .A1(n6790), .A2(n6802), .ZN(n6780) );
  NAND2_X1 U8330 ( .A1(n6781), .A2(n6780), .ZN(n6782) );
  NAND2_X1 U8331 ( .A1(n6849), .A2(n6783), .ZN(n7791) );
  INV_X1 U8332 ( .A(n6783), .ZN(n9824) );
  NAND2_X1 U8333 ( .A1(n8220), .A2(n9824), .ZN(n9754) );
  NAND2_X1 U8334 ( .A1(n7791), .A2(n9754), .ZN(n6787) );
  OAI21_X1 U8335 ( .B1(n6782), .B2(n6787), .A(n6851), .ZN(n9829) );
  INV_X1 U8336 ( .A(n6784), .ZN(n6786) );
  INV_X1 U8337 ( .A(n9746), .ZN(n6785) );
  OAI21_X1 U8338 ( .B1(n9824), .B2(n6786), .A(n6785), .ZN(n9825) );
  OAI22_X1 U8339 ( .A1(n8469), .A2(n9824), .B1(n9825), .B2(n8400), .ZN(n6796)
         );
  NAND2_X1 U8340 ( .A1(n6859), .A2(n6858), .ZN(n6789) );
  INV_X1 U8341 ( .A(n6787), .ZN(n6788) );
  XNOR2_X1 U8342 ( .A(n6789), .B(n6788), .ZN(n6792) );
  OAI22_X1 U8343 ( .A1(n6790), .A2(n8498), .B1(n6860), .B2(n8496), .ZN(n6791)
         );
  AOI21_X1 U8344 ( .B1(n6792), .B2(n8511), .A(n6791), .ZN(n9826) );
  OAI21_X1 U8345 ( .B1(n6793), .B2(n8485), .A(n9826), .ZN(n6794) );
  MUX2_X1 U8346 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6794), .S(n9763), .Z(n6795)
         );
  AOI211_X1 U8347 ( .C1(n8518), .C2(n9829), .A(n6796), .B(n6795), .ZN(n6797)
         );
  INV_X1 U8348 ( .A(n6797), .ZN(P2_U3292) );
  INV_X1 U8349 ( .A(n6798), .ZN(n6799) );
  OAI22_X1 U8350 ( .A1(n8400), .A2(n6799), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8485), .ZN(n6805) );
  INV_X1 U8351 ( .A(n6800), .ZN(n6801) );
  NAND2_X1 U8352 ( .A1(n9763), .A2(n6801), .ZN(n7546) );
  OAI22_X1 U8353 ( .A1(n6803), .A2(n7546), .B1(n8469), .B2(n6802), .ZN(n6804)
         );
  AOI211_X1 U8354 ( .C1(n8467), .C2(P2_REG2_REG_3__SCAN_IN), .A(n6805), .B(
        n6804), .ZN(n6806) );
  OAI21_X1 U8355 ( .B1(n8467), .B2(n6807), .A(n6806), .ZN(P2_U3293) );
  INV_X1 U8356 ( .A(n6720), .ZN(n6810) );
  NOR3_X1 U8357 ( .A1(n6808), .A2(n8189), .A3(n7006), .ZN(n6809) );
  AOI21_X1 U8358 ( .B1(n6810), .B2(n8185), .A(n6809), .ZN(n6818) );
  OR2_X1 U8359 ( .A1(n6811), .A2(n8196), .ZN(n6815) );
  AOI22_X1 U8360 ( .A1(n8205), .A2(n6993), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n6814) );
  AOI22_X1 U8361 ( .A1(n8168), .A2(n8213), .B1(n8190), .B2(n8215), .ZN(n6813)
         );
  NAND2_X1 U8362 ( .A1(n4315), .A2(n7148), .ZN(n6812) );
  AND4_X1 U8363 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6816)
         );
  OAI21_X1 U8364 ( .B1(n6818), .B2(n6817), .A(n6816), .ZN(P2_U3226) );
  OAI21_X1 U8365 ( .B1(n6820), .B2(n6819), .A(n6938), .ZN(n6821) );
  NAND2_X1 U8366 ( .A1(n6821), .A2(n8683), .ZN(n6827) );
  INV_X1 U8367 ( .A(n9059), .ZN(n7285) );
  AOI21_X1 U8368 ( .B1(n8664), .B2(n9061), .A(n6822), .ZN(n6824) );
  NAND2_X1 U8369 ( .A1(n8726), .A2(n7192), .ZN(n6823) );
  OAI211_X1 U8370 ( .C1(n7285), .C2(n8706), .A(n6824), .B(n6823), .ZN(n6825)
         );
  AOI21_X1 U8371 ( .B1(n7262), .B2(n8709), .A(n6825), .ZN(n6826) );
  NAND2_X1 U8372 ( .A1(n6827), .A2(n6826), .ZN(P1_U3215) );
  OAI222_X1 U8373 ( .A1(P1_U3084), .A2(n5579), .B1(n7552), .B2(n6828), .C1(
        n7481), .C2(n5394), .ZN(P1_U3334) );
  NAND2_X1 U8374 ( .A1(n6418), .A2(n8063), .ZN(n7835) );
  NAND2_X1 U8375 ( .A1(n6836), .A2(n7835), .ZN(n9806) );
  INV_X1 U8376 ( .A(n9806), .ZN(n6834) );
  AOI22_X1 U8377 ( .A1(n9806), .A2(n8511), .B1(n8508), .B2(n6829), .ZN(n9808)
         );
  INV_X1 U8378 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6830) );
  OAI22_X1 U8379 ( .A1(n8467), .A2(n9808), .B1(n6830), .B2(n8485), .ZN(n6831)
         );
  AOI21_X1 U8380 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8467), .A(n6831), .ZN(
        n6833) );
  OAI21_X1 U8381 ( .B1(n8514), .B2(n8521), .A(n9804), .ZN(n6832) );
  OAI211_X1 U8382 ( .C1(n6834), .C2(n8504), .A(n6833), .B(n6832), .ZN(P2_U3296) );
  XNOR2_X1 U8383 ( .A(n6835), .B(n6836), .ZN(n6837) );
  NAND2_X1 U8384 ( .A1(n6837), .A2(n8511), .ZN(n6839) );
  AOI22_X1 U8385 ( .A1(n6691), .A2(n8508), .B1(n8506), .B2(n6418), .ZN(n6838)
         );
  NAND2_X1 U8386 ( .A1(n6839), .A2(n6838), .ZN(n9814) );
  NOR2_X1 U8387 ( .A1(n9763), .A2(n6385), .ZN(n6844) );
  INV_X1 U8388 ( .A(n6840), .ZN(n9811) );
  NAND2_X1 U8389 ( .A1(n9804), .A2(n7965), .ZN(n9810) );
  NAND2_X1 U8390 ( .A1(n9811), .A2(n9810), .ZN(n6842) );
  OAI22_X1 U8391 ( .A1(n8400), .A2(n6842), .B1(n6841), .B2(n8485), .ZN(n6843)
         );
  AOI211_X1 U8392 ( .C1(n9763), .C2(n9814), .A(n6844), .B(n6843), .ZN(n6848)
         );
  OAI21_X1 U8393 ( .B1(n6835), .B2(n6846), .A(n6845), .ZN(n9816) );
  AOI22_X1 U8394 ( .A1(n8518), .A2(n9816), .B1(n8514), .B2(n7965), .ZN(n6847)
         );
  NAND2_X1 U8395 ( .A1(n6848), .A2(n6847), .ZN(P2_U3295) );
  NAND2_X1 U8396 ( .A1(n6849), .A2(n9824), .ZN(n6850) );
  NAND2_X1 U8397 ( .A1(n8178), .A2(n8219), .ZN(n7846) );
  INV_X1 U8398 ( .A(n8219), .ZN(n6955) );
  NAND2_X1 U8399 ( .A1(n6955), .A2(n9835), .ZN(n7848) );
  NAND2_X1 U8400 ( .A1(n6852), .A2(n7795), .ZN(n8515) );
  NAND2_X1 U8401 ( .A1(n9835), .A2(n8219), .ZN(n6853) );
  NAND2_X1 U8402 ( .A1(n8515), .A2(n6853), .ZN(n6947) );
  OR2_X1 U8403 ( .A1(n6854), .A2(n8179), .ZN(n7851) );
  NAND2_X1 U8404 ( .A1(n6854), .A2(n8179), .ZN(n7850) );
  INV_X1 U8405 ( .A(n8179), .ZN(n8509) );
  OR2_X1 U8406 ( .A1(n6854), .A2(n8509), .ZN(n6855) );
  NAND2_X1 U8407 ( .A1(n4336), .A2(n6855), .ZN(n6856) );
  OR2_X1 U8408 ( .A1(n6960), .A2(n7042), .ZN(n7854) );
  NAND2_X1 U8409 ( .A1(n6960), .A2(n7042), .ZN(n7858) );
  NAND2_X1 U8410 ( .A1(n6856), .A2(n7853), .ZN(n6857) );
  NAND2_X1 U8411 ( .A1(n6962), .A2(n6857), .ZN(n9850) );
  AND2_X1 U8412 ( .A1(n7791), .A2(n6858), .ZN(n7826) );
  NAND2_X1 U8413 ( .A1(n9755), .A2(n7843), .ZN(n6861) );
  INV_X1 U8414 ( .A(n9831), .ZN(n9748) );
  NAND2_X1 U8415 ( .A1(n6860), .A2(n9748), .ZN(n9744) );
  NAND2_X1 U8416 ( .A1(n6861), .A2(n9744), .ZN(n8505) );
  NAND2_X1 U8417 ( .A1(n8505), .A2(n8516), .ZN(n6862) );
  INV_X1 U8418 ( .A(n7850), .ZN(n6863) );
  INV_X1 U8419 ( .A(n7853), .ZN(n6864) );
  OAI21_X1 U8420 ( .B1(n6865), .B2(n7853), .A(n6969), .ZN(n6867) );
  OAI22_X1 U8421 ( .A1(n8179), .A2(n8498), .B1(n7005), .B2(n8496), .ZN(n6866)
         );
  AOI21_X1 U8422 ( .B1(n6867), .B2(n8511), .A(n6866), .ZN(n6868) );
  OAI21_X1 U8423 ( .B1(n9850), .B2(n8532), .A(n6868), .ZN(n9853) );
  NAND2_X1 U8424 ( .A1(n9853), .A2(n9763), .ZN(n6875) );
  OAI22_X1 U8425 ( .A1(n9763), .A2(n6870), .B1(n6869), .B2(n8485), .ZN(n6873)
         );
  NAND2_X1 U8426 ( .A1(n9746), .A2(n9831), .ZN(n8520) );
  OR2_X1 U8427 ( .A1(n8520), .A2(n9835), .ZN(n6949) );
  INV_X1 U8428 ( .A(n6960), .ZN(n9851) );
  AND2_X1 U8429 ( .A1(n6950), .A2(n9851), .ZN(n7050) );
  NOR2_X1 U8430 ( .A1(n6950), .A2(n9851), .ZN(n6871) );
  OR2_X1 U8431 ( .A1(n7050), .A2(n6871), .ZN(n9852) );
  NOR2_X1 U8432 ( .A1(n9852), .A2(n8400), .ZN(n6872) );
  AOI211_X1 U8433 ( .C1(n8514), .C2(n6960), .A(n6873), .B(n6872), .ZN(n6874)
         );
  OAI211_X1 U8434 ( .C1(n9850), .C2(n7546), .A(n6875), .B(n6874), .ZN(P2_U3288) );
  NAND2_X1 U8435 ( .A1(n7225), .A2(n7096), .ZN(n8752) );
  AND2_X1 U8436 ( .A1(n8752), .A2(n6878), .ZN(n8955) );
  INV_X1 U8437 ( .A(n7103), .ZN(n6881) );
  INV_X1 U8438 ( .A(n7096), .ZN(n9698) );
  NAND2_X1 U8439 ( .A1(n9698), .A2(n9062), .ZN(n8751) );
  NAND2_X1 U8440 ( .A1(n8752), .A2(n8751), .ZN(n6892) );
  INV_X1 U8441 ( .A(n6892), .ZN(n8881) );
  AOI21_X1 U8442 ( .B1(n6879), .B2(n6878), .A(n8881), .ZN(n6880) );
  AOI211_X1 U8443 ( .C1(n6881), .C2(n8751), .A(n8091), .B(n6880), .ZN(n6883)
         );
  OAI22_X1 U8444 ( .A1(n7104), .A2(n9616), .B1(n9617), .B2(n9618), .ZN(n6882)
         );
  OR2_X1 U8445 ( .A1(n6883), .A2(n6882), .ZN(n9700) );
  NAND2_X1 U8446 ( .A1(n6884), .A2(n7096), .ZN(n6885) );
  NAND2_X1 U8447 ( .A1(n7218), .A2(n6885), .ZN(n9699) );
  AOI22_X1 U8448 ( .A1(n9648), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6886), .B2(
        n9314), .ZN(n6888) );
  NAND2_X1 U8449 ( .A1(n9316), .A2(n7096), .ZN(n6887) );
  OAI211_X1 U8450 ( .C1(n9699), .C2(n9148), .A(n6888), .B(n6887), .ZN(n6896)
         );
  NOR2_X1 U8451 ( .A1(n9063), .A2(n6889), .ZN(n6890) );
  AOI21_X1 U8452 ( .B1(n6891), .B2(n8880), .A(n6890), .ZN(n6893) );
  NOR2_X1 U8453 ( .A1(n6893), .A2(n6892), .ZN(n9697) );
  NAND2_X1 U8454 ( .A1(n6893), .A2(n6892), .ZN(n9702) );
  INV_X1 U8455 ( .A(n9702), .ZN(n6894) );
  NOR3_X1 U8456 ( .A1(n9697), .A2(n6894), .A3(n9306), .ZN(n6895) );
  AOI211_X1 U8457 ( .C1(n9646), .C2(n9700), .A(n6896), .B(n6895), .ZN(n6897)
         );
  INV_X1 U8458 ( .A(n6897), .ZN(P1_U3283) );
  INV_X1 U8459 ( .A(n7555), .ZN(n6936) );
  OAI222_X1 U8460 ( .A1(n8647), .A2(n6936), .B1(P2_U3152), .B2(n7790), .C1(
        n6898), .C2(n8641), .ZN(P2_U3338) );
  INV_X1 U8461 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6912) );
  INV_X1 U8462 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6899) );
  MUX2_X1 U8463 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6899), .S(n7210), .Z(n6902)
         );
  OAI21_X1 U8464 ( .B1(n6904), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6900), .ZN(
        n6901) );
  NAND2_X1 U8465 ( .A1(n6902), .A2(n6901), .ZN(n7209) );
  OAI21_X1 U8466 ( .B1(n6902), .B2(n6901), .A(n7209), .ZN(n6908) );
  INV_X1 U8467 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6906) );
  AOI21_X1 U8468 ( .B1(n6904), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6903), .ZN(
        n7204) );
  XNOR2_X1 U8469 ( .A(n7204), .B(n7210), .ZN(n6905) );
  NAND2_X1 U8470 ( .A1(n6905), .A2(n6906), .ZN(n7205) );
  OAI21_X1 U8471 ( .B1(n6906), .B2(n6905), .A(n7205), .ZN(n6907) );
  AOI22_X1 U8472 ( .A1(n9593), .A2(n6908), .B1(n9598), .B2(n6907), .ZN(n6911)
         );
  NAND2_X1 U8473 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7237) );
  INV_X1 U8474 ( .A(n7237), .ZN(n6909) );
  AOI21_X1 U8475 ( .B1(n9578), .B2(n7210), .A(n6909), .ZN(n6910) );
  OAI211_X1 U8476 ( .C1(n9584), .C2(n6912), .A(n6911), .B(n6910), .ZN(P1_U3255) );
  INV_X1 U8477 ( .A(n8213), .ZN(n7882) );
  NOR3_X1 U8478 ( .A1(n6913), .A2(n7882), .A3(n8189), .ZN(n6914) );
  AOI21_X1 U8479 ( .B1(n6915), .B2(n8185), .A(n6914), .ZN(n6934) );
  NAND2_X1 U8480 ( .A1(n6916), .A2(n5928), .ZN(n6918) );
  AOI22_X1 U8481 ( .A1(n7577), .A2(n7515), .B1(n7747), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6917) );
  XNOR2_X1 U8482 ( .A(n8612), .B(n7995), .ZN(n7058) );
  INV_X1 U8483 ( .A(n7451), .ZN(n8212) );
  NAND2_X1 U8484 ( .A1(n8212), .A2(n7985), .ZN(n7059) );
  XNOR2_X1 U8485 ( .A(n7058), .B(n7059), .ZN(n6933) );
  AND2_X1 U8486 ( .A1(n6933), .A2(n6919), .ZN(n6920) );
  INV_X1 U8487 ( .A(n7062), .ZN(n6931) );
  NAND2_X1 U8488 ( .A1(n7764), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6926) );
  XNOR2_X1 U8489 ( .A(n7071), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U8490 ( .A1(n5816), .A2(n7462), .ZN(n6925) );
  INV_X1 U8491 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6922) );
  OR2_X1 U8492 ( .A1(n5850), .A2(n6922), .ZN(n6924) );
  INV_X1 U8493 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7454) );
  OR2_X1 U8494 ( .A1(n7082), .A2(n7454), .ZN(n6923) );
  INV_X1 U8495 ( .A(n7535), .ZN(n8211) );
  AOI22_X1 U8496 ( .A1(n8168), .A2(n8211), .B1(n8190), .B2(n8213), .ZN(n6929)
         );
  NAND2_X1 U8497 ( .A1(n8612), .A2(n4315), .ZN(n6928) );
  NAND2_X1 U8498 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7379) );
  NAND2_X1 U8499 ( .A1(n8205), .A2(n7472), .ZN(n6927) );
  NAND4_X1 U8500 ( .A1(n6929), .A2(n6928), .A3(n7379), .A4(n6927), .ZN(n6930)
         );
  AOI21_X1 U8501 ( .B1(n6931), .B2(n8185), .A(n6930), .ZN(n6932) );
  OAI21_X1 U8502 ( .B1(n6934), .B2(n6933), .A(n6932), .ZN(P2_U3217) );
  OAI222_X1 U8503 ( .A1(P1_U3084), .A2(n8912), .B1(n7552), .B2(n6936), .C1(
        n6935), .C2(n7481), .ZN(P1_U3333) );
  INV_X1 U8504 ( .A(n7426), .ZN(n7272) );
  AND2_X1 U8505 ( .A1(n6938), .A2(n6937), .ZN(n6941) );
  OAI211_X1 U8506 ( .C1(n6941), .C2(n6940), .A(n8683), .B(n6939), .ZN(n6946)
         );
  INV_X1 U8507 ( .A(n7261), .ZN(n9060) );
  NAND2_X1 U8508 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9604) );
  INV_X1 U8509 ( .A(n9604), .ZN(n6942) );
  AOI21_X1 U8510 ( .B1(n8664), .B2(n9060), .A(n6942), .ZN(n6943) );
  OAI21_X1 U8511 ( .B1(n7322), .B2(n8706), .A(n6943), .ZN(n6944) );
  AOI21_X1 U8512 ( .B1(n7270), .B2(n8726), .A(n6944), .ZN(n6945) );
  OAI211_X1 U8513 ( .C1(n7272), .C2(n8730), .A(n6946), .B(n6945), .ZN(P1_U3234) );
  INV_X1 U8514 ( .A(n6947), .ZN(n6948) );
  INV_X1 U8515 ( .A(n7847), .ZN(n7797) );
  OAI21_X1 U8516 ( .B1(n6948), .B2(n7797), .A(n4336), .ZN(n9848) );
  INV_X1 U8517 ( .A(n6854), .ZN(n9844) );
  INV_X1 U8518 ( .A(n6949), .ZN(n8519) );
  INV_X1 U8519 ( .A(n6950), .ZN(n6951) );
  OAI21_X1 U8520 ( .B1(n9844), .B2(n8519), .A(n6951), .ZN(n9845) );
  AOI22_X1 U8521 ( .A1(n8514), .A2(n6854), .B1(n9751), .B2(n8113), .ZN(n6952)
         );
  OAI21_X1 U8522 ( .B1(n8400), .B2(n9845), .A(n6952), .ZN(n6957) );
  XNOR2_X1 U8523 ( .A(n6953), .B(n7797), .ZN(n6954) );
  OAI222_X1 U8524 ( .A1(n8498), .A2(n6955), .B1(n8496), .B2(n7042), .C1(n6954), 
        .C2(n9759), .ZN(n9846) );
  MUX2_X1 U8525 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9846), .S(n9763), .Z(n6956)
         );
  AOI211_X1 U8526 ( .C1(n8518), .C2(n9848), .A(n6957), .B(n6956), .ZN(n6958)
         );
  INV_X1 U8527 ( .A(n6958), .ZN(P2_U3289) );
  INV_X1 U8528 ( .A(n7590), .ZN(n7019) );
  OAI222_X1 U8529 ( .A1(n8647), .A2(n7019), .B1(n8641), .B2(n6959), .C1(n7953), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8530 ( .A1(n6960), .A2(n8218), .ZN(n6961) );
  OR2_X1 U8531 ( .A1(n7055), .A2(n7005), .ZN(n7862) );
  NAND2_X1 U8532 ( .A1(n7055), .A2(n7005), .ZN(n7859) );
  AND2_X1 U8533 ( .A1(n9863), .A2(n8216), .ZN(n6964) );
  OR2_X1 U8534 ( .A1(n7799), .A2(n6964), .ZN(n6981) );
  OR2_X1 U8535 ( .A1(n7040), .A2(n6981), .ZN(n6966) );
  XNOR2_X1 U8536 ( .A(n9863), .B(n8216), .ZN(n7861) );
  INV_X1 U8537 ( .A(n7861), .ZN(n6963) );
  OR2_X1 U8538 ( .A1(n7055), .A2(n8217), .ZN(n7000) );
  AND2_X1 U8539 ( .A1(n6963), .A2(n7000), .ZN(n6999) );
  AND2_X1 U8540 ( .A1(n6966), .A2(n6965), .ZN(n6968) );
  OR2_X1 U8541 ( .A1(n6980), .A2(n7006), .ZN(n7875) );
  NAND2_X1 U8542 ( .A1(n6980), .A2(n7006), .ZN(n7872) );
  NAND2_X1 U8543 ( .A1(n7875), .A2(n7872), .ZN(n6970) );
  NAND2_X1 U8544 ( .A1(n6966), .A2(n6982), .ZN(n6967) );
  OAI21_X1 U8545 ( .B1(n6968), .B2(n6970), .A(n6967), .ZN(n9872) );
  OR2_X1 U8546 ( .A1(n9863), .A2(n7043), .ZN(n7867) );
  NAND2_X1 U8547 ( .A1(n9863), .A2(n7043), .ZN(n7866) );
  INV_X1 U8548 ( .A(n6970), .ZN(n7800) );
  XNOR2_X1 U8549 ( .A(n6987), .B(n7800), .ZN(n6971) );
  NAND2_X1 U8550 ( .A1(n6971), .A2(n8511), .ZN(n6973) );
  AOI22_X1 U8551 ( .A1(n8214), .A2(n8508), .B1(n8506), .B2(n8216), .ZN(n6972)
         );
  NAND2_X1 U8552 ( .A1(n6973), .A2(n6972), .ZN(n9876) );
  INV_X1 U8553 ( .A(n7055), .ZN(n9857) );
  NAND2_X1 U8554 ( .A1(n7050), .A2(n9857), .ZN(n7052) );
  OR2_X1 U8555 ( .A1(n7052), .A2(n9863), .ZN(n7013) );
  AND2_X1 U8556 ( .A1(n7013), .A2(n6980), .ZN(n6974) );
  OR2_X1 U8557 ( .A1(n6974), .A2(n6992), .ZN(n9874) );
  AOI22_X1 U8558 ( .A1(n8467), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n6975), .B2(
        n9751), .ZN(n6977) );
  NAND2_X1 U8559 ( .A1(n8514), .A2(n6980), .ZN(n6976) );
  OAI211_X1 U8560 ( .C1(n9874), .C2(n8400), .A(n6977), .B(n6976), .ZN(n6978)
         );
  AOI21_X1 U8561 ( .B1(n9876), .B2(n9763), .A(n6978), .ZN(n6979) );
  OAI21_X1 U8562 ( .B1(n9872), .B2(n8504), .A(n6979), .ZN(P2_U3285) );
  AND2_X1 U8563 ( .A1(n6980), .A2(n8215), .ZN(n6983) );
  OR2_X1 U8564 ( .A1(n6981), .A2(n6983), .ZN(n6984) );
  OR2_X1 U8565 ( .A1(n7148), .A2(n6985), .ZN(n7876) );
  NAND2_X1 U8566 ( .A1(n7148), .A2(n6985), .ZN(n7878) );
  NAND2_X1 U8567 ( .A1(n7876), .A2(n7878), .ZN(n7802) );
  NAND2_X1 U8568 ( .A1(n6986), .A2(n7802), .ZN(n7150) );
  OAI21_X1 U8569 ( .B1(n6986), .B2(n7802), .A(n7150), .ZN(n9886) );
  INV_X1 U8570 ( .A(n9886), .ZN(n6998) );
  OAI211_X1 U8571 ( .C1(n4863), .C2(n6988), .A(n7145), .B(n8511), .ZN(n6990)
         );
  AOI22_X1 U8572 ( .A1(n8215), .A2(n8506), .B1(n8508), .B2(n8213), .ZN(n6989)
         );
  NAND2_X1 U8573 ( .A1(n6990), .A2(n6989), .ZN(n9884) );
  INV_X1 U8574 ( .A(n7148), .ZN(n9880) );
  INV_X1 U8575 ( .A(n7155), .ZN(n6991) );
  OAI21_X1 U8576 ( .B1(n9880), .B2(n6992), .A(n6991), .ZN(n9882) );
  AOI22_X1 U8577 ( .A1(n8467), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n6993), .B2(
        n9751), .ZN(n6995) );
  NAND2_X1 U8578 ( .A1(n8514), .A2(n7148), .ZN(n6994) );
  OAI211_X1 U8579 ( .C1(n9882), .C2(n8400), .A(n6995), .B(n6994), .ZN(n6996)
         );
  AOI21_X1 U8580 ( .B1(n9884), .B2(n9763), .A(n6996), .ZN(n6997) );
  OAI21_X1 U8581 ( .B1(n6998), .B2(n8504), .A(n6997), .ZN(P2_U3284) );
  NAND2_X1 U8582 ( .A1(n7038), .A2(n6999), .ZN(n7003) );
  NAND2_X1 U8583 ( .A1(n7038), .A2(n7000), .ZN(n7001) );
  NAND2_X1 U8584 ( .A1(n7001), .A2(n7861), .ZN(n7002) );
  NAND2_X1 U8585 ( .A1(n7003), .A2(n7002), .ZN(n9862) );
  XNOR2_X1 U8586 ( .A(n7004), .B(n7861), .ZN(n7008) );
  OAI22_X1 U8587 ( .A1(n7006), .A2(n8496), .B1(n7005), .B2(n8498), .ZN(n7007)
         );
  AOI21_X1 U8588 ( .B1(n7008), .B2(n8511), .A(n7007), .ZN(n7009) );
  OAI21_X1 U8589 ( .B1(n9862), .B2(n8532), .A(n7009), .ZN(n9866) );
  NAND2_X1 U8590 ( .A1(n9866), .A2(n9763), .ZN(n7017) );
  OAI22_X1 U8591 ( .A1(n9763), .A2(n7011), .B1(n7010), .B2(n8485), .ZN(n7015)
         );
  NAND2_X1 U8592 ( .A1(n7052), .A2(n9863), .ZN(n7012) );
  NAND2_X1 U8593 ( .A1(n7013), .A2(n7012), .ZN(n9865) );
  NOR2_X1 U8594 ( .A1(n9865), .A2(n8400), .ZN(n7014) );
  AOI211_X1 U8595 ( .C1(n8514), .C2(n9863), .A(n7015), .B(n7014), .ZN(n7016)
         );
  OAI211_X1 U8596 ( .C1(n9862), .C2(n7546), .A(n7017), .B(n7016), .ZN(P2_U3286) );
  INV_X1 U8597 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7018) );
  OAI222_X1 U8598 ( .A1(P1_U3084), .A2(n4926), .B1(n7552), .B2(n7019), .C1(
        n7018), .C2(n7481), .ZN(P1_U3332) );
  NAND2_X1 U8599 ( .A1(n7027), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8600 ( .A1(n7021), .A2(n7020), .ZN(n7024) );
  MUX2_X1 U8601 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n5994), .S(n7166), .Z(n7022)
         );
  INV_X1 U8602 ( .A(n7022), .ZN(n7023) );
  NOR2_X1 U8603 ( .A1(n7024), .A2(n7023), .ZN(n7160) );
  AOI21_X1 U8604 ( .B1(n7024), .B2(n7023), .A(n7160), .ZN(n7037) );
  INV_X1 U8605 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7034) );
  INV_X1 U8606 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7025) );
  MUX2_X1 U8607 ( .A(n7025), .B(P2_REG1_REG_11__SCAN_IN), .S(n7166), .Z(n7029)
         );
  AOI21_X1 U8608 ( .B1(n7029), .B2(n7028), .A(n7165), .ZN(n7030) );
  NAND2_X1 U8609 ( .A1(n9734), .A2(n7030), .ZN(n7033) );
  INV_X1 U8610 ( .A(n7031), .ZN(n7032) );
  OAI211_X1 U8611 ( .C1(n8291), .C2(n7034), .A(n7033), .B(n7032), .ZN(n7035)
         );
  AOI21_X1 U8612 ( .B1(n7166), .B2(n8285), .A(n7035), .ZN(n7036) );
  OAI21_X1 U8613 ( .B1(n7037), .B2(n8282), .A(n7036), .ZN(P2_U3256) );
  INV_X1 U8614 ( .A(n7038), .ZN(n7039) );
  AOI21_X1 U8615 ( .B1(n7799), .B2(n7040), .A(n7039), .ZN(n9856) );
  XNOR2_X1 U8616 ( .A(n7041), .B(n7799), .ZN(n7045) );
  OAI22_X1 U8617 ( .A1(n7043), .A2(n8496), .B1(n7042), .B2(n8498), .ZN(n7044)
         );
  AOI21_X1 U8618 ( .B1(n7045), .B2(n8511), .A(n7044), .ZN(n7046) );
  OAI21_X1 U8619 ( .B1(n9856), .B2(n8532), .A(n7046), .ZN(n9859) );
  NAND2_X1 U8620 ( .A1(n9859), .A2(n9763), .ZN(n7057) );
  INV_X1 U8621 ( .A(n7047), .ZN(n7048) );
  OAI22_X1 U8622 ( .A1(n9763), .A2(n7049), .B1(n7048), .B2(n8485), .ZN(n7054)
         );
  OR2_X1 U8623 ( .A1(n7050), .A2(n9857), .ZN(n7051) );
  NAND2_X1 U8624 ( .A1(n7052), .A2(n7051), .ZN(n9858) );
  NOR2_X1 U8625 ( .A1(n9858), .A2(n8400), .ZN(n7053) );
  AOI211_X1 U8626 ( .C1(n8514), .C2(n7055), .A(n7054), .B(n7053), .ZN(n7056)
         );
  OAI211_X1 U8627 ( .C1(n9856), .C2(n7546), .A(n7057), .B(n7056), .ZN(P2_U3287) );
  INV_X1 U8628 ( .A(n7058), .ZN(n7060) );
  NAND2_X1 U8629 ( .A1(n7060), .A2(n7059), .ZN(n7061) );
  NAND2_X1 U8630 ( .A1(n7063), .A2(n5928), .ZN(n7065) );
  AOI22_X1 U8631 ( .A1(n8230), .A2(n7515), .B1(n7747), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7064) );
  NAND2_X1 U8632 ( .A1(n8211), .A2(n7985), .ZN(n7181) );
  NAND2_X1 U8633 ( .A1(n7179), .A2(n7181), .ZN(n7079) );
  NAND2_X1 U8634 ( .A1(n7066), .A2(n4355), .ZN(n7178) );
  NAND2_X1 U8635 ( .A1(n7067), .A2(n5928), .ZN(n7069) );
  AOI22_X1 U8636 ( .A1(n7747), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7515), .B2(
        n8250), .ZN(n7068) );
  XNOR2_X1 U8637 ( .A(n8602), .B(n7593), .ZN(n7301) );
  INV_X1 U8638 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7184) );
  INV_X1 U8639 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7070) );
  OAI21_X1 U8640 ( .B1(n7071), .B2(n7184), .A(n7070), .ZN(n7072) );
  AND2_X1 U8641 ( .A1(n7080), .A2(n7072), .ZN(n7543) );
  NAND2_X1 U8642 ( .A1(n5816), .A2(n7543), .ZN(n7078) );
  NAND2_X1 U8643 ( .A1(n7764), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7077) );
  INV_X1 U8644 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7073) );
  OR2_X1 U8645 ( .A1(n7742), .A2(n7073), .ZN(n7076) );
  INV_X1 U8646 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7074) );
  OR2_X1 U8647 ( .A1(n5850), .A2(n7074), .ZN(n7075) );
  INV_X1 U8648 ( .A(n8497), .ZN(n8210) );
  NAND2_X1 U8649 ( .A1(n8210), .A2(n7985), .ZN(n7300) );
  XNOR2_X1 U8650 ( .A(n7301), .B(n7300), .ZN(n7091) );
  AOI21_X1 U8651 ( .B1(n7079), .B2(n7178), .A(n7091), .ZN(n7303) );
  INV_X1 U8652 ( .A(n7303), .ZN(n7095) );
  INV_X1 U8653 ( .A(n7543), .ZN(n7089) );
  INV_X1 U8654 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U8655 ( .A1(n7080), .A2(n8248), .ZN(n7081) );
  NAND2_X1 U8656 ( .A1(n7311), .A2(n7081), .ZN(n8486) );
  OR2_X1 U8657 ( .A1(n7763), .A2(n8486), .ZN(n7087) );
  NAND2_X1 U8658 ( .A1(n7764), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7086) );
  INV_X1 U8659 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8487) );
  OR2_X1 U8660 ( .A1(n7082), .A2(n8487), .ZN(n7085) );
  INV_X1 U8661 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7083) );
  OR2_X1 U8662 ( .A1(n5850), .A2(n7083), .ZN(n7084) );
  INV_X1 U8663 ( .A(n7673), .ZN(n8477) );
  AOI22_X1 U8664 ( .A1(n8190), .A2(n8211), .B1(n8168), .B2(n8477), .ZN(n7088)
         );
  NAND2_X1 U8665 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8236) );
  OAI211_X1 U8666 ( .C1(n7089), .C2(n8162), .A(n7088), .B(n8236), .ZN(n7090)
         );
  AOI21_X1 U8667 ( .B1(n8602), .B2(n4315), .A(n7090), .ZN(n7094) );
  NOR2_X1 U8668 ( .A1(n7179), .A2(n8196), .ZN(n7092) );
  NOR2_X1 U8669 ( .A1(n8189), .A2(n7535), .ZN(n7180) );
  OAI211_X1 U8670 ( .C1(n7092), .C2(n7180), .A(n7091), .B(n7178), .ZN(n7093)
         );
  OAI211_X1 U8671 ( .C1(n7095), .C2(n8196), .A(n7094), .B(n7093), .ZN(P2_U3228) );
  INV_X1 U8672 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7110) );
  OR2_X1 U8673 ( .A1(n7262), .A2(n7261), .ZN(n8926) );
  NAND2_X1 U8674 ( .A1(n7262), .A2(n7261), .ZN(n8768) );
  NAND2_X1 U8675 ( .A1(n7096), .A2(n9062), .ZN(n7097) );
  NAND2_X1 U8676 ( .A1(n9702), .A2(n7097), .ZN(n7217) );
  OR2_X1 U8677 ( .A1(n9704), .A2(n9061), .ZN(n7098) );
  NAND2_X1 U8678 ( .A1(n7217), .A2(n7098), .ZN(n7100) );
  NAND2_X1 U8679 ( .A1(n9704), .A2(n9061), .ZN(n7099) );
  NAND2_X1 U8680 ( .A1(n7100), .A2(n7099), .ZN(n7102) );
  INV_X1 U8681 ( .A(n7264), .ZN(n7101) );
  AOI21_X1 U8682 ( .B1(n8887), .B2(n7102), .A(n7101), .ZN(n7196) );
  NAND2_X1 U8683 ( .A1(n7118), .A2(n5398), .ZN(n8859) );
  OR2_X1 U8684 ( .A1(n8859), .A2(n9032), .ZN(n9671) );
  OR2_X1 U8685 ( .A1(n9704), .A2(n7104), .ZN(n8757) );
  AND2_X1 U8686 ( .A1(n8757), .A2(n8751), .ZN(n8927) );
  NAND2_X1 U8687 ( .A1(n9704), .A2(n7104), .ZN(n8767) );
  XNOR2_X1 U8688 ( .A(n7259), .B(n8887), .ZN(n7105) );
  AOI222_X1 U8689 ( .A1(n9313), .A2(n7105), .B1(n9061), .B2(n9633), .C1(n9059), 
        .C2(n9631), .ZN(n7202) );
  NAND2_X1 U8690 ( .A1(n7220), .A2(n7262), .ZN(n7106) );
  NAND2_X1 U8691 ( .A1(n7106), .A2(n9667), .ZN(n7107) );
  NOR2_X1 U8692 ( .A1(n7268), .A2(n7107), .ZN(n7200) );
  AOI21_X1 U8693 ( .B1(n9677), .B2(n7262), .A(n7200), .ZN(n7108) );
  OAI211_X1 U8694 ( .C1(n7196), .C2(n9696), .A(n7202), .B(n7108), .ZN(n7115)
         );
  NAND2_X1 U8695 ( .A1(n7115), .A2(n9714), .ZN(n7109) );
  OAI21_X1 U8696 ( .B1(n9714), .B2(n7110), .A(n7109), .ZN(P1_U3484) );
  NOR2_X1 U8697 ( .A1(n7112), .A2(n7111), .ZN(n7113) );
  NAND2_X1 U8698 ( .A1(n7115), .A2(n9729), .ZN(n7116) );
  OAI21_X1 U8699 ( .B1(n9729), .B2(n7117), .A(n7116), .ZN(P1_U3533) );
  INV_X1 U8700 ( .A(n7678), .ZN(n8015) );
  OAI222_X1 U8701 ( .A1(n7481), .A2(n7119), .B1(n9431), .B2(n8015), .C1(
        P1_U3084), .C2(n7118), .ZN(P1_U3331) );
  XOR2_X1 U8702 ( .A(n7121), .B(n7120), .Z(n7122) );
  XNOR2_X1 U8703 ( .A(n7123), .B(n7122), .ZN(n7131) );
  NOR2_X1 U8704 ( .A1(n8723), .A2(n7322), .ZN(n7124) );
  AOI211_X1 U8705 ( .C1(n8721), .C2(n9056), .A(n7125), .B(n7124), .ZN(n7126)
         );
  OAI21_X1 U8706 ( .B1(n7128), .B2(n7127), .A(n7126), .ZN(n7129) );
  AOI21_X1 U8707 ( .B1(n9400), .B2(n8709), .A(n7129), .ZN(n7130) );
  OAI21_X1 U8708 ( .B1(n7131), .B2(n8716), .A(n7130), .ZN(P1_U3232) );
  INV_X1 U8709 ( .A(n7323), .ZN(n9499) );
  INV_X1 U8710 ( .A(n7134), .ZN(n7138) );
  AOI21_X1 U8711 ( .B1(n7134), .B2(n7133), .A(n7132), .ZN(n7135) );
  NOR2_X1 U8712 ( .A1(n7135), .A2(n8716), .ZN(n7136) );
  OAI21_X1 U8713 ( .B1(n7138), .B2(n7137), .A(n7136), .ZN(n7144) );
  NAND2_X1 U8714 ( .A1(n8721), .A2(n9057), .ZN(n7140) );
  OAI211_X1 U8715 ( .C1(n7285), .C2(n8723), .A(n7140), .B(n7139), .ZN(n7141)
         );
  AOI21_X1 U8716 ( .B1(n7142), .B2(n8726), .A(n7141), .ZN(n7143) );
  OAI211_X1 U8717 ( .C1(n9499), .C2(n8730), .A(n7144), .B(n7143), .ZN(P1_U3222) );
  XNOR2_X1 U8718 ( .A(n7881), .B(n8213), .ZN(n7879) );
  OAI21_X1 U8719 ( .B1(n7146), .B2(n7879), .A(n7455), .ZN(n7147) );
  AOI222_X1 U8720 ( .A1(n8511), .A2(n7147), .B1(n8214), .B2(n8506), .C1(n8212), 
        .C2(n8508), .ZN(n9474) );
  OR2_X1 U8721 ( .A1(n7148), .A2(n8214), .ZN(n7149) );
  AND2_X1 U8722 ( .A1(n7151), .A2(n7879), .ZN(n9471) );
  INV_X1 U8723 ( .A(n9471), .ZN(n7152) );
  NAND3_X1 U8724 ( .A1(n7152), .A2(n8518), .A3(n4747), .ZN(n7159) );
  OAI22_X1 U8725 ( .A1(n9763), .A2(n7154), .B1(n7153), .B2(n8485), .ZN(n7157)
         );
  OAI21_X1 U8726 ( .B1(n7155), .B2(n9472), .A(n7471), .ZN(n9473) );
  NOR2_X1 U8727 ( .A1(n9473), .A2(n8400), .ZN(n7156) );
  AOI211_X1 U8728 ( .C1(n8514), .C2(n7881), .A(n7157), .B(n7156), .ZN(n7158)
         );
  OAI211_X1 U8729 ( .C1(n8467), .C2(n9474), .A(n7159), .B(n7158), .ZN(P2_U3283) );
  NOR2_X1 U8730 ( .A1(n7166), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7161) );
  NOR2_X1 U8731 ( .A1(n7161), .A2(n7160), .ZN(n7164) );
  MUX2_X1 U8732 ( .A(n6012), .B(P2_REG2_REG_12__SCAN_IN), .S(n7252), .Z(n7162)
         );
  INV_X1 U8733 ( .A(n7162), .ZN(n7163) );
  NAND2_X1 U8734 ( .A1(n7163), .A2(n7164), .ZN(n7243) );
  OAI211_X1 U8735 ( .C1(n7164), .C2(n7163), .A(n9735), .B(n7243), .ZN(n7176)
         );
  INV_X1 U8736 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7167) );
  MUX2_X1 U8737 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7167), .S(n7252), .Z(n7168)
         );
  OAI21_X1 U8738 ( .B1(n7169), .B2(n7168), .A(n7251), .ZN(n7174) );
  NOR2_X1 U8739 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7170), .ZN(n7173) );
  INV_X1 U8740 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7171) );
  NOR2_X1 U8741 ( .A1(n8291), .A2(n7171), .ZN(n7172) );
  AOI211_X1 U8742 ( .C1(n9734), .C2(n7174), .A(n7173), .B(n7172), .ZN(n7175)
         );
  OAI211_X1 U8743 ( .C1(n9730), .C2(n7177), .A(n7176), .B(n7175), .ZN(P2_U3257) );
  AND2_X1 U8744 ( .A1(n7179), .A2(n7178), .ZN(n7191) );
  INV_X1 U8745 ( .A(n7180), .ZN(n7190) );
  NAND3_X1 U8746 ( .A1(n7191), .A2(n8185), .A3(n7181), .ZN(n7189) );
  INV_X1 U8747 ( .A(n8152), .ZN(n7185) );
  NAND2_X1 U8748 ( .A1(n8210), .A2(n8508), .ZN(n7183) );
  NAND2_X1 U8749 ( .A1(n8212), .A2(n8506), .ZN(n7182) );
  AND2_X1 U8750 ( .A1(n7183), .A2(n7182), .ZN(n7460) );
  OAI22_X1 U8751 ( .A1(n7185), .A2(n7460), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7184), .ZN(n7187) );
  NOR2_X1 U8752 ( .A1(n4675), .A2(n8207), .ZN(n7186) );
  AOI211_X1 U8753 ( .C1(n8205), .C2(n7462), .A(n7187), .B(n7186), .ZN(n7188)
         );
  OAI211_X1 U8754 ( .C1(n7191), .C2(n7190), .A(n7189), .B(n7188), .ZN(P2_U3243) );
  INV_X1 U8755 ( .A(n7392), .ZN(n9322) );
  NAND2_X1 U8756 ( .A1(n7262), .A2(n9316), .ZN(n7194) );
  NAND2_X1 U8757 ( .A1(n9314), .A2(n7192), .ZN(n7193) );
  OAI211_X1 U8758 ( .C1(n9646), .C2(n7195), .A(n7194), .B(n7193), .ZN(n7199)
         );
  NAND2_X1 U8759 ( .A1(n9646), .A2(n9630), .ZN(n7197) );
  AOI21_X1 U8760 ( .B1(n7299), .B2(n7197), .A(n7196), .ZN(n7198) );
  AOI211_X1 U8761 ( .C1(n7200), .C2(n9322), .A(n7199), .B(n7198), .ZN(n7201)
         );
  OAI21_X1 U8762 ( .B1(n9648), .B2(n7202), .A(n7201), .ZN(P1_U3281) );
  INV_X1 U8763 ( .A(n7210), .ZN(n7203) );
  NAND2_X1 U8764 ( .A1(n7204), .A2(n7203), .ZN(n7206) );
  NAND2_X1 U8765 ( .A1(n7206), .A2(n7205), .ZN(n7353) );
  INV_X1 U8766 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7207) );
  AOI211_X1 U8767 ( .C1(n7208), .C2(n7207), .A(n7354), .B(n9553), .ZN(n7216)
         );
  INV_X1 U8768 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7212) );
  OAI21_X1 U8769 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n7210), .A(n7209), .ZN(
        n7358) );
  NOR2_X1 U8770 ( .A1(n7212), .A2(n7211), .ZN(n7360) );
  AOI211_X1 U8771 ( .C1(n7212), .C2(n7211), .A(n7360), .B(n9573), .ZN(n7215)
         );
  NAND2_X1 U8772 ( .A1(n9589), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7213) );
  NAND2_X1 U8773 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7346) );
  OAI211_X1 U8774 ( .C1(n9587), .C2(n7359), .A(n7213), .B(n7346), .ZN(n7214)
         );
  OR3_X1 U8775 ( .A1(n7216), .A2(n7215), .A3(n7214), .ZN(P1_U3256) );
  NAND2_X1 U8776 ( .A1(n8757), .A2(n8767), .ZN(n8883) );
  XOR2_X1 U8777 ( .A(n7217), .B(n8883), .Z(n9711) );
  NAND2_X1 U8778 ( .A1(n7218), .A2(n9704), .ZN(n7219) );
  NAND2_X1 U8779 ( .A1(n7220), .A2(n7219), .ZN(n9707) );
  AOI22_X1 U8780 ( .A1(n9316), .A2(n9704), .B1(n7221), .B2(n9314), .ZN(n7222)
         );
  OAI21_X1 U8781 ( .B1(n9707), .B2(n9148), .A(n7222), .ZN(n7227) );
  NAND2_X1 U8782 ( .A1(n7103), .A2(n8751), .ZN(n7223) );
  XOR2_X1 U8783 ( .A(n8883), .B(n7223), .Z(n7224) );
  OAI222_X1 U8784 ( .A1(n9616), .A2(n7261), .B1(n9618), .B2(n7225), .C1(n8091), 
        .C2(n7224), .ZN(n9708) );
  MUX2_X1 U8785 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9708), .S(n9646), .Z(n7226)
         );
  AOI211_X1 U8786 ( .C1(n9320), .C2(n9711), .A(n7227), .B(n7226), .ZN(n7228)
         );
  INV_X1 U8787 ( .A(n7228), .ZN(P1_U3282) );
  INV_X1 U8788 ( .A(n7683), .ZN(n7232) );
  OR2_X1 U8789 ( .A1(n7229), .A2(P1_U3084), .ZN(n9040) );
  INV_X1 U8790 ( .A(n9040), .ZN(n9034) );
  AOI21_X1 U8791 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9429), .A(n9034), .ZN(
        n7230) );
  OAI21_X1 U8792 ( .B1(n7232), .B2(n9431), .A(n7230), .ZN(P1_U3330) );
  NAND2_X1 U8793 ( .A1(n8644), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7231) );
  OAI211_X1 U8794 ( .C1(n7232), .C2(n8647), .A(n7963), .B(n7231), .ZN(P2_U3335) );
  XOR2_X1 U8795 ( .A(n7235), .B(n7234), .Z(n7236) );
  XNOR2_X1 U8796 ( .A(n7233), .B(n7236), .ZN(n7242) );
  INV_X1 U8797 ( .A(n9055), .ZN(n7409) );
  NAND2_X1 U8798 ( .A1(n8664), .A2(n9057), .ZN(n7238) );
  OAI211_X1 U8799 ( .C1(n7409), .C2(n8706), .A(n7238), .B(n7237), .ZN(n7240)
         );
  NOR2_X1 U8800 ( .A1(n9493), .A2(n8730), .ZN(n7239) );
  AOI211_X1 U8801 ( .C1(n7336), .C2(n8726), .A(n7240), .B(n7239), .ZN(n7241)
         );
  OAI21_X1 U8802 ( .B1(n7242), .B2(n8716), .A(n7241), .ZN(P1_U3213) );
  NAND2_X1 U8803 ( .A1(n7252), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7244) );
  NAND2_X1 U8804 ( .A1(n7244), .A2(n7243), .ZN(n7246) );
  AOI22_X1 U8805 ( .A1(n7376), .A2(n7154), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7250), .ZN(n7245) );
  NOR2_X1 U8806 ( .A1(n7246), .A2(n7245), .ZN(n7370) );
  AOI21_X1 U8807 ( .B1(n7246), .B2(n7245), .A(n7370), .ZN(n7258) );
  INV_X1 U8808 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7248) );
  OAI22_X1 U8809 ( .A1(n8291), .A2(n7248), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7247), .ZN(n7249) );
  AOI21_X1 U8810 ( .B1(n8285), .B2(n7376), .A(n7249), .ZN(n7257) );
  INV_X1 U8811 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9478) );
  AOI22_X1 U8812 ( .A1(n7376), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9478), .B2(
        n7250), .ZN(n7254) );
  OAI21_X1 U8813 ( .B1(n7252), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7251), .ZN(
        n7253) );
  OAI21_X1 U8814 ( .B1(n7254), .B2(n7253), .A(n7375), .ZN(n7255) );
  NAND2_X1 U8815 ( .A1(n7255), .A2(n9734), .ZN(n7256) );
  OAI211_X1 U8816 ( .C1(n7258), .C2(n8282), .A(n7257), .B(n7256), .ZN(P2_U3258) );
  NAND2_X1 U8817 ( .A1(n7259), .A2(n8887), .ZN(n7260) );
  XNOR2_X1 U8818 ( .A(n7426), .B(n7285), .ZN(n8773) );
  INV_X1 U8819 ( .A(n8773), .ZN(n8885) );
  XNOR2_X1 U8820 ( .A(n7283), .B(n8885), .ZN(n7267) );
  OAI22_X1 U8821 ( .A1(n7261), .A2(n9618), .B1(n7322), .B2(n9616), .ZN(n7266)
         );
  OR2_X1 U8822 ( .A1(n7262), .A2(n9060), .ZN(n7263) );
  XNOR2_X1 U8823 ( .A(n7276), .B(n8885), .ZN(n7430) );
  NOR2_X1 U8824 ( .A1(n7430), .A2(n7290), .ZN(n7265) );
  AOI211_X1 U8825 ( .C1(n9313), .C2(n7267), .A(n7266), .B(n7265), .ZN(n7429)
         );
  INV_X1 U8826 ( .A(n7268), .ZN(n7269) );
  INV_X1 U8827 ( .A(n7293), .ZN(n7294) );
  AOI21_X1 U8828 ( .B1(n7426), .B2(n7269), .A(n7294), .ZN(n7427) );
  AOI22_X1 U8829 ( .A1(n9648), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7270), .B2(
        n9314), .ZN(n7271) );
  OAI21_X1 U8830 ( .B1(n7272), .B2(n9623), .A(n7271), .ZN(n7274) );
  NOR2_X1 U8831 ( .A1(n7430), .A2(n7299), .ZN(n7273) );
  AOI211_X1 U8832 ( .C1(n7427), .C2(n9612), .A(n7274), .B(n7273), .ZN(n7275)
         );
  OAI21_X1 U8833 ( .B1(n7429), .B2(n9648), .A(n7275), .ZN(P1_U3280) );
  OR2_X1 U8834 ( .A1(n7426), .A2(n9059), .ZN(n7277) );
  INV_X1 U8835 ( .A(n7281), .ZN(n7280) );
  OR2_X1 U8836 ( .A1(n7323), .A2(n7322), .ZN(n8776) );
  NAND2_X1 U8837 ( .A1(n7323), .A2(n7322), .ZN(n8791) );
  NAND2_X1 U8838 ( .A1(n7281), .A2(n8888), .ZN(n7282) );
  NAND2_X1 U8839 ( .A1(n7402), .A2(n7282), .ZN(n9497) );
  AOI22_X1 U8840 ( .A1(n9631), .A2(n9057), .B1(n9059), .B2(n9633), .ZN(n7289)
         );
  AND2_X1 U8841 ( .A1(n7426), .A2(n7285), .ZN(n8775) );
  OR2_X1 U8842 ( .A1(n7426), .A2(n7285), .ZN(n7326) );
  NAND2_X1 U8843 ( .A1(n7419), .A2(n7326), .ZN(n7286) );
  XOR2_X1 U8844 ( .A(n8888), .B(n7286), .Z(n7287) );
  NAND2_X1 U8845 ( .A1(n7287), .A2(n9313), .ZN(n7288) );
  OAI211_X1 U8846 ( .C1(n9497), .C2(n7290), .A(n7289), .B(n7288), .ZN(n9500)
         );
  NAND2_X1 U8847 ( .A1(n9500), .A2(n9646), .ZN(n7298) );
  INV_X1 U8848 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7292) );
  OAI22_X1 U8849 ( .A1(n9646), .A2(n7292), .B1(n7291), .B2(n9641), .ZN(n7296)
         );
  OAI211_X1 U8850 ( .C1(n7294), .C2(n9499), .A(n9667), .B(n7415), .ZN(n9498)
         );
  NOR2_X1 U8851 ( .A1(n9498), .A2(n7392), .ZN(n7295) );
  AOI211_X1 U8852 ( .C1(n9316), .C2(n7323), .A(n7296), .B(n7295), .ZN(n7297)
         );
  OAI211_X1 U8853 ( .C1(n9497), .C2(n7299), .A(n7298), .B(n7297), .ZN(P1_U3279) );
  NOR2_X1 U8854 ( .A1(n7303), .A2(n7302), .ZN(n7308) );
  INV_X1 U8855 ( .A(n8258), .ZN(n8264) );
  AOI22_X1 U8856 ( .A1(n7747), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7515), .B2(
        n8264), .ZN(n7305) );
  NAND2_X1 U8857 ( .A1(n8477), .A2(n7985), .ZN(n7306) );
  AOI21_X1 U8858 ( .B1(n7439), .B2(n7306), .A(n7440), .ZN(n7307) );
  OAI211_X1 U8859 ( .C1(n7308), .C2(n7307), .A(n7443), .B(n8185), .ZN(n7317)
         );
  OAI22_X1 U8860 ( .A1(n8162), .A2(n8486), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8248), .ZN(n7315) );
  INV_X1 U8861 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U8862 ( .A1(n5800), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7310) );
  NAND2_X1 U8863 ( .A1(n5912), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7309) );
  AND2_X1 U8864 ( .A1(n7310), .A2(n7309), .ZN(n7313) );
  XNOR2_X1 U8865 ( .A(n7311), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U8866 ( .A1(n8466), .A2(n5816), .ZN(n7312) );
  OAI211_X1 U8867 ( .C1(n7728), .C2(n8262), .A(n7313), .B(n7312), .ZN(n8453)
         );
  INV_X1 U8868 ( .A(n8453), .ZN(n8495) );
  OAI22_X1 U8869 ( .A1(n8495), .A2(n8202), .B1(n8200), .B2(n8497), .ZN(n7314)
         );
  AOI211_X1 U8870 ( .C1(n8599), .C2(n4315), .A(n7315), .B(n7314), .ZN(n7316)
         );
  NAND2_X1 U8871 ( .A1(n7317), .A2(n7316), .ZN(P2_U3230) );
  INV_X1 U8872 ( .A(n7697), .ZN(n7320) );
  OAI222_X1 U8873 ( .A1(P1_U3084), .A2(n7318), .B1(n7552), .B2(n7320), .C1(
        n10071), .C2(n7481), .ZN(P1_U3329) );
  OAI222_X1 U8874 ( .A1(n7321), .A2(P2_U3152), .B1(n8016), .B2(n7320), .C1(
        n7319), .C2(n8641), .ZN(P2_U3334) );
  INV_X1 U8875 ( .A(n7322), .ZN(n9058) );
  NAND2_X1 U8876 ( .A1(n7323), .A2(n9058), .ZN(n7400) );
  NAND2_X1 U8877 ( .A1(n7402), .A2(n7400), .ZN(n7413) );
  OR2_X1 U8878 ( .A1(n9400), .A2(n9057), .ZN(n7405) );
  NAND2_X1 U8879 ( .A1(n7413), .A2(n7405), .ZN(n7324) );
  NAND2_X1 U8880 ( .A1(n9400), .A2(n9057), .ZN(n7396) );
  NAND2_X1 U8881 ( .A1(n7324), .A2(n7396), .ZN(n7325) );
  INV_X1 U8882 ( .A(n9056), .ZN(n8783) );
  OR2_X1 U8883 ( .A1(n7395), .A2(n8783), .ZN(n8934) );
  NAND2_X1 U8884 ( .A1(n7395), .A2(n8783), .ZN(n8923) );
  NAND2_X1 U8885 ( .A1(n8934), .A2(n8923), .ZN(n7331) );
  XNOR2_X1 U8886 ( .A(n7325), .B(n7328), .ZN(n9496) );
  INV_X1 U8887 ( .A(n9496), .ZN(n7341) );
  AND2_X1 U8888 ( .A1(n8776), .A2(n7326), .ZN(n8792) );
  INV_X1 U8889 ( .A(n9057), .ZN(n8779) );
  OR2_X1 U8890 ( .A1(n9400), .A2(n8779), .ZN(n8933) );
  NAND2_X1 U8891 ( .A1(n9400), .A2(n8779), .ZN(n8959) );
  AND2_X1 U8892 ( .A1(n8792), .A2(n8890), .ZN(n7327) );
  INV_X1 U8893 ( .A(n7331), .ZN(n7328) );
  AND2_X1 U8894 ( .A1(n8959), .A2(n7328), .ZN(n7329) );
  NAND2_X1 U8895 ( .A1(n7330), .A2(n7329), .ZN(n7386) );
  NAND2_X1 U8896 ( .A1(n7330), .A2(n8959), .ZN(n7332) );
  NAND2_X1 U8897 ( .A1(n7332), .A2(n7331), .ZN(n7333) );
  NAND3_X1 U8898 ( .A1(n7386), .A2(n9313), .A3(n7333), .ZN(n7335) );
  AOI22_X1 U8899 ( .A1(n9633), .A2(n9057), .B1(n9055), .B2(n9631), .ZN(n7334)
         );
  NAND2_X1 U8900 ( .A1(n7335), .A2(n7334), .ZN(n9495) );
  AND2_X2 U8901 ( .A1(n7414), .A2(n9493), .ZN(n7391) );
  INV_X1 U8902 ( .A(n7391), .ZN(n7487) );
  OAI211_X1 U8903 ( .C1(n9493), .C2(n7414), .A(n7487), .B(n9667), .ZN(n9492)
         );
  AOI22_X1 U8904 ( .A1(n9648), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7336), .B2(
        n9314), .ZN(n7338) );
  NAND2_X1 U8905 ( .A1(n7395), .A2(n9316), .ZN(n7337) );
  OAI211_X1 U8906 ( .C1(n9492), .C2(n7392), .A(n7338), .B(n7337), .ZN(n7339)
         );
  AOI21_X1 U8907 ( .B1(n9495), .B2(n9646), .A(n7339), .ZN(n7340) );
  OAI21_X1 U8908 ( .B1(n7341), .B2(n9306), .A(n7340), .ZN(P1_U3277) );
  XNOR2_X1 U8909 ( .A(n7344), .B(n7343), .ZN(n7345) );
  XNOR2_X1 U8910 ( .A(n7342), .B(n7345), .ZN(n7352) );
  INV_X1 U8911 ( .A(n7346), .ZN(n7347) );
  AOI21_X1 U8912 ( .B1(n8664), .B2(n9056), .A(n7347), .ZN(n7349) );
  NAND2_X1 U8913 ( .A1(n8726), .A2(n7488), .ZN(n7348) );
  OAI211_X1 U8914 ( .C1(n7492), .C2(n8706), .A(n7349), .B(n7348), .ZN(n7350)
         );
  AOI21_X1 U8915 ( .B1(n9395), .B2(n8709), .A(n7350), .ZN(n7351) );
  OAI21_X1 U8916 ( .B1(n7352), .B2(n8716), .A(n7351), .ZN(P1_U3239) );
  NOR2_X1 U8917 ( .A1(n7359), .A2(n7353), .ZN(n7355) );
  NAND2_X1 U8918 ( .A1(n9100), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7356) );
  OAI21_X1 U8919 ( .B1(n9100), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7356), .ZN(
        n7357) );
  AOI211_X1 U8920 ( .C1(n4379), .C2(n7357), .A(n9095), .B(n9553), .ZN(n7369)
         );
  NOR2_X1 U8921 ( .A1(n7359), .A2(n7358), .ZN(n7361) );
  NOR2_X1 U8922 ( .A1(n7361), .A2(n7360), .ZN(n7364) );
  INV_X1 U8923 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7362) );
  MUX2_X1 U8924 ( .A(n7362), .B(P1_REG1_REG_16__SCAN_IN), .S(n9100), .Z(n7363)
         );
  NOR2_X1 U8925 ( .A1(n7364), .A2(n7363), .ZN(n9099) );
  AOI211_X1 U8926 ( .C1(n7364), .C2(n7363), .A(n9099), .B(n9573), .ZN(n7368)
         );
  NAND2_X1 U8927 ( .A1(n9589), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7365) );
  NAND2_X1 U8928 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7501) );
  OAI211_X1 U8929 ( .C1(n9587), .C2(n7366), .A(n7365), .B(n7501), .ZN(n7367)
         );
  OR3_X1 U8930 ( .A1(n7369), .A2(n7368), .A3(n7367), .ZN(P1_U3257) );
  NOR2_X1 U8931 ( .A1(n7376), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7371) );
  NOR2_X1 U8932 ( .A1(n7371), .A2(n7370), .ZN(n7373) );
  AOI22_X1 U8933 ( .A1(n7577), .A2(n6068), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7572), .ZN(n7372) );
  NOR2_X1 U8934 ( .A1(n7373), .A2(n7372), .ZN(n7571) );
  AOI21_X1 U8935 ( .B1(n7373), .B2(n7372), .A(n7571), .ZN(n7385) );
  INV_X1 U8936 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7374) );
  AOI22_X1 U8937 ( .A1(n7577), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7374), .B2(
        n7572), .ZN(n7378) );
  OAI21_X1 U8938 ( .B1(n7378), .B2(n7377), .A(n7576), .ZN(n7383) );
  INV_X1 U8939 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7381) );
  NAND2_X1 U8940 ( .A1(n8285), .A2(n7577), .ZN(n7380) );
  OAI211_X1 U8941 ( .C1(n8291), .C2(n7381), .A(n7380), .B(n7379), .ZN(n7382)
         );
  AOI21_X1 U8942 ( .B1(n7383), .B2(n9734), .A(n7382), .ZN(n7384) );
  OAI21_X1 U8943 ( .B1(n7385), .B2(n8282), .A(n7384), .ZN(P2_U3259) );
  OR2_X1 U8944 ( .A1(n7623), .A2(n7492), .ZN(n8940) );
  NAND2_X1 U8945 ( .A1(n7623), .A2(n7492), .ZN(n8920) );
  NAND2_X1 U8946 ( .A1(n8940), .A2(n8920), .ZN(n8893) );
  NOR2_X1 U8947 ( .A1(n9395), .A2(n7409), .ZN(n8938) );
  NAND2_X1 U8948 ( .A1(n9395), .A2(n7409), .ZN(n8924) );
  OAI21_X1 U8949 ( .B1(n7410), .B2(n7387), .A(n7628), .ZN(n7388) );
  AOI222_X1 U8950 ( .A1(n9313), .A2(n7388), .B1(n9053), .B2(n9631), .C1(n9055), 
        .C2(n9633), .ZN(n9488) );
  INV_X1 U8951 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7390) );
  INV_X1 U8952 ( .A(n7503), .ZN(n7389) );
  OAI22_X1 U8953 ( .A1(n9646), .A2(n7390), .B1(n7389), .B2(n9641), .ZN(n7394)
         );
  INV_X1 U8954 ( .A(n9395), .ZN(n7490) );
  INV_X1 U8955 ( .A(n7623), .ZN(n9489) );
  OAI211_X1 U8956 ( .C1(n4375), .C2(n9489), .A(n9667), .B(n7626), .ZN(n9487)
         );
  NOR2_X1 U8957 ( .A1(n9487), .A2(n7392), .ZN(n7393) );
  AOI211_X1 U8958 ( .C1(n9316), .C2(n7623), .A(n7394), .B(n7393), .ZN(n7412)
         );
  OR2_X1 U8959 ( .A1(n7395), .A2(n9056), .ZN(n7404) );
  INV_X1 U8960 ( .A(n7404), .ZN(n7399) );
  NAND2_X1 U8961 ( .A1(n7395), .A2(n9056), .ZN(n7397) );
  AND2_X1 U8962 ( .A1(n7397), .A2(n7396), .ZN(n7398) );
  AND2_X1 U8963 ( .A1(n7400), .A2(n7403), .ZN(n7401) );
  INV_X1 U8964 ( .A(n7403), .ZN(n7407) );
  AND2_X1 U8965 ( .A1(n7405), .A2(n7404), .ZN(n7406) );
  XNOR2_X1 U8966 ( .A(n7622), .B(n7410), .ZN(n9491) );
  NAND2_X1 U8967 ( .A1(n9491), .A2(n9320), .ZN(n7411) );
  OAI211_X1 U8968 ( .C1(n9488), .C2(n9648), .A(n7412), .B(n7411), .ZN(P1_U3275) );
  XOR2_X1 U8969 ( .A(n8890), .B(n7413), .Z(n9404) );
  AOI21_X1 U8970 ( .B1(n9400), .B2(n7415), .A(n7414), .ZN(n9401) );
  INV_X1 U8971 ( .A(n9400), .ZN(n7418) );
  AOI22_X1 U8972 ( .A1(n9648), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7416), .B2(
        n9314), .ZN(n7417) );
  OAI21_X1 U8973 ( .B1(n7418), .B2(n9623), .A(n7417), .ZN(n7424) );
  NAND2_X1 U8974 ( .A1(n7419), .A2(n8792), .ZN(n7420) );
  NAND2_X1 U8975 ( .A1(n7420), .A2(n8791), .ZN(n7421) );
  XNOR2_X1 U8976 ( .A(n7421), .B(n8890), .ZN(n7422) );
  AOI222_X1 U8977 ( .A1(n9313), .A2(n7422), .B1(n9056), .B2(n9631), .C1(n9058), 
        .C2(n9633), .ZN(n9403) );
  NOR2_X1 U8978 ( .A1(n9403), .A2(n9648), .ZN(n7423) );
  AOI211_X1 U8979 ( .C1(n9401), .C2(n9612), .A(n7424), .B(n7423), .ZN(n7425)
         );
  OAI21_X1 U8980 ( .B1(n9306), .B2(n9404), .A(n7425), .ZN(P1_U3278) );
  INV_X1 U8981 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7432) );
  AOI22_X1 U8982 ( .A1(n7427), .A2(n9667), .B1(n9677), .B2(n7426), .ZN(n7428)
         );
  OAI211_X1 U8983 ( .C1(n9671), .C2(n7430), .A(n7429), .B(n7428), .ZN(n7433)
         );
  NAND2_X1 U8984 ( .A1(n7433), .A2(n9714), .ZN(n7431) );
  OAI21_X1 U8985 ( .B1(n9714), .B2(n7432), .A(n7431), .ZN(P1_U3487) );
  INV_X1 U8986 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U8987 ( .A1(n7433), .A2(n9729), .ZN(n7434) );
  OAI21_X1 U8988 ( .B1(n9729), .B2(n7435), .A(n7434), .ZN(P1_U3534) );
  NAND2_X1 U8989 ( .A1(n7436), .A2(n5928), .ZN(n7438) );
  AOI22_X1 U8990 ( .A1(n7747), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7515), .B2(
        n8276), .ZN(n7437) );
  INV_X1 U8991 ( .A(n8592), .ZN(n8470) );
  NOR3_X1 U8992 ( .A1(n7439), .A2(n7673), .A3(n8189), .ZN(n7446) );
  XNOR2_X1 U8993 ( .A(n8592), .B(n7593), .ZN(n7509) );
  NAND2_X1 U8994 ( .A1(n8453), .A2(n7985), .ZN(n7510) );
  XNOR2_X1 U8995 ( .A(n7509), .B(n7510), .ZN(n7441) );
  AOI21_X1 U8996 ( .B1(n7443), .B2(n7441), .A(n8196), .ZN(n7445) );
  INV_X1 U8997 ( .A(n7440), .ZN(n7442) );
  INV_X1 U8998 ( .A(n7513), .ZN(n7444) );
  OAI21_X1 U8999 ( .B1(n7446), .B2(n7445), .A(n7444), .ZN(n7450) );
  NOR2_X1 U9000 ( .A1(n7447), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8266) );
  INV_X1 U9001 ( .A(n8476), .ZN(n7675) );
  OAI22_X1 U9002 ( .A1(n7675), .A2(n8202), .B1(n8200), .B2(n7673), .ZN(n7448)
         );
  AOI211_X1 U9003 ( .C1(n8205), .C2(n8466), .A(n8266), .B(n7448), .ZN(n7449)
         );
  OAI211_X1 U9004 ( .C1(n8470), .C2(n8207), .A(n7450), .B(n7449), .ZN(P2_U3240) );
  NAND2_X1 U9005 ( .A1(n8612), .A2(n7451), .ZN(n7884) );
  NAND2_X1 U9006 ( .A1(n7883), .A2(n7884), .ZN(n7886) );
  OR2_X1 U9007 ( .A1(n8612), .A2(n8212), .ZN(n7452) );
  NAND2_X1 U9008 ( .A1(n7467), .A2(n7452), .ZN(n7538) );
  NAND2_X1 U9009 ( .A1(n8607), .A2(n7535), .ZN(n7890) );
  NAND2_X1 U9010 ( .A1(n7889), .A2(n7890), .ZN(n7537) );
  XNOR2_X1 U9011 ( .A(n7538), .B(n7887), .ZN(n8611) );
  INV_X1 U9012 ( .A(n8045), .ZN(n7453) );
  AOI21_X1 U9013 ( .B1(n8607), .B2(n7469), .A(n7453), .ZN(n8608) );
  OAI22_X1 U9014 ( .A1(n4675), .A2(n8469), .B1(n9763), .B2(n7454), .ZN(n7465)
         );
  NAND2_X1 U9015 ( .A1(n7881), .A2(n7882), .ZN(n7874) );
  INV_X1 U9016 ( .A(n7886), .ZN(n7456) );
  NAND2_X1 U9017 ( .A1(n7458), .A2(n7883), .ZN(n7457) );
  NAND3_X1 U9018 ( .A1(n7458), .A2(n7537), .A3(n7883), .ZN(n7459) );
  NAND3_X1 U9019 ( .A1(n7534), .A2(n8511), .A3(n7459), .ZN(n7461) );
  AND2_X1 U9020 ( .A1(n7461), .A2(n7460), .ZN(n8610) );
  NAND2_X1 U9021 ( .A1(n9751), .A2(n7462), .ZN(n7463) );
  AOI21_X1 U9022 ( .B1(n8610), .B2(n7463), .A(n8467), .ZN(n7464) );
  AOI211_X1 U9023 ( .C1(n8608), .C2(n8521), .A(n7465), .B(n7464), .ZN(n7466)
         );
  OAI21_X1 U9024 ( .B1(n8611), .B2(n8504), .A(n7466), .ZN(P2_U3281) );
  OAI21_X1 U9025 ( .B1(n4385), .B2(n7886), .A(n7467), .ZN(n7468) );
  INV_X1 U9026 ( .A(n7468), .ZN(n8616) );
  INV_X1 U9027 ( .A(n7469), .ZN(n7470) );
  AOI21_X1 U9028 ( .B1(n8612), .B2(n7471), .A(n7470), .ZN(n8613) );
  AOI22_X1 U9029 ( .A1(n8467), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7472), .B2(
        n9751), .ZN(n7473) );
  OAI21_X1 U9030 ( .B1(n4676), .B2(n8469), .A(n7473), .ZN(n7477) );
  XOR2_X1 U9031 ( .A(n7474), .B(n7886), .Z(n7475) );
  AOI222_X1 U9032 ( .A1(n8511), .A2(n7475), .B1(n8213), .B2(n8506), .C1(n8211), 
        .C2(n8508), .ZN(n8615) );
  NOR2_X1 U9033 ( .A1(n8615), .A2(n8467), .ZN(n7476) );
  AOI211_X1 U9034 ( .C1(n8613), .C2(n8521), .A(n7477), .B(n7476), .ZN(n7478)
         );
  OAI21_X1 U9035 ( .B1(n8616), .B2(n8504), .A(n7478), .ZN(P2_U3282) );
  INV_X1 U9036 ( .A(n7709), .ZN(n7483) );
  OAI222_X1 U9037 ( .A1(n7481), .A2(n7480), .B1(n9431), .B2(n7483), .C1(
        P1_U3084), .C2(n7479), .ZN(P1_U3328) );
  OAI222_X1 U9038 ( .A1(P2_U3152), .A2(n7484), .B1(n8647), .B2(n7483), .C1(
        n7482), .C2(n8641), .ZN(P2_U3333) );
  INV_X1 U9039 ( .A(n7721), .ZN(n7532) );
  AOI22_X1 U9040 ( .A1(n5554), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9429), .ZN(n7485) );
  OAI21_X1 U9041 ( .B1(n7532), .B2(n9431), .A(n7485), .ZN(P1_U3327) );
  XNOR2_X1 U9042 ( .A(n9395), .B(n9055), .ZN(n8798) );
  XNOR2_X1 U9043 ( .A(n7486), .B(n8798), .ZN(n9399) );
  AOI21_X1 U9044 ( .B1(n9395), .B2(n7487), .A(n4375), .ZN(n9396) );
  AOI22_X1 U9045 ( .A1(n9648), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7488), .B2(
        n9314), .ZN(n7489) );
  OAI21_X1 U9046 ( .B1(n7490), .B2(n9623), .A(n7489), .ZN(n7495) );
  INV_X1 U9047 ( .A(n8798), .ZN(n8892) );
  XNOR2_X1 U9048 ( .A(n7491), .B(n8892), .ZN(n7493) );
  INV_X1 U9049 ( .A(n7492), .ZN(n9054) );
  AOI222_X1 U9050 ( .A1(n9313), .A2(n7493), .B1(n9054), .B2(n9631), .C1(n9056), 
        .C2(n9633), .ZN(n9398) );
  NOR2_X1 U9051 ( .A1(n9398), .A2(n9648), .ZN(n7494) );
  AOI211_X1 U9052 ( .C1(n9396), .C2(n9612), .A(n7495), .B(n7494), .ZN(n7496)
         );
  OAI21_X1 U9053 ( .B1(n9306), .B2(n9399), .A(n7496), .ZN(P1_U3276) );
  INV_X1 U9054 ( .A(n7497), .ZN(n7498) );
  AOI21_X1 U9055 ( .B1(n7500), .B2(n7499), .A(n7498), .ZN(n7508) );
  INV_X1 U9056 ( .A(n9053), .ZN(n8724) );
  INV_X1 U9057 ( .A(n7501), .ZN(n7502) );
  AOI21_X1 U9058 ( .B1(n8664), .B2(n9055), .A(n7502), .ZN(n7505) );
  NAND2_X1 U9059 ( .A1(n8726), .A2(n7503), .ZN(n7504) );
  OAI211_X1 U9060 ( .C1(n8724), .C2(n8706), .A(n7505), .B(n7504), .ZN(n7506)
         );
  AOI21_X1 U9061 ( .B1(n7623), .B2(n8709), .A(n7506), .ZN(n7507) );
  OAI21_X1 U9062 ( .B1(n7508), .B2(n8716), .A(n7507), .ZN(P1_U3224) );
  INV_X1 U9063 ( .A(n7509), .ZN(n7512) );
  INV_X1 U9064 ( .A(n7510), .ZN(n7511) );
  NAND2_X1 U9065 ( .A1(n7514), .A2(n5928), .ZN(n7517) );
  AOI22_X1 U9066 ( .A1(n7747), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7515), .B2(
        n9753), .ZN(n7516) );
  XNOR2_X1 U9067 ( .A(n8588), .B(n7995), .ZN(n7519) );
  AND2_X1 U9068 ( .A1(n8476), .A2(n7985), .ZN(n7518) );
  NAND2_X1 U9069 ( .A1(n7519), .A2(n7518), .ZN(n7553) );
  NAND2_X1 U9070 ( .A1(n4390), .A2(n7553), .ZN(n7520) );
  XNOR2_X1 U9071 ( .A(n7554), .B(n7520), .ZN(n7531) );
  INV_X1 U9072 ( .A(n8457), .ZN(n7528) );
  INV_X1 U9073 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9074 ( .A1(n7522), .A2(n7558), .ZN(n7523) );
  NAND2_X1 U9075 ( .A1(n7598), .A2(n7523), .ZN(n8441) );
  OR2_X1 U9076 ( .A1(n8441), .A2(n7763), .ZN(n7526) );
  AOI22_X1 U9077 ( .A1(n5800), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n5912), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n7525) );
  NAND2_X1 U9078 ( .A1(n7764), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7524) );
  AOI22_X1 U9079 ( .A1(n8190), .A2(n8453), .B1(n8168), .B2(n8454), .ZN(n7527)
         );
  NAND2_X1 U9080 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8289) );
  OAI211_X1 U9081 ( .C1(n8162), .C2(n7528), .A(n7527), .B(n8289), .ZN(n7529)
         );
  AOI21_X1 U9082 ( .B1(n8588), .B2(n4315), .A(n7529), .ZN(n7530) );
  OAI21_X1 U9083 ( .B1(n7531), .B2(n8196), .A(n7530), .ZN(P2_U3221) );
  OAI222_X1 U9084 ( .A1(n7533), .A2(P2_U3152), .B1(n8641), .B2(n10116), .C1(
        n8016), .C2(n7532), .ZN(P2_U3332) );
  NAND2_X1 U9085 ( .A1(n8602), .A2(n8497), .ZN(n7894) );
  NAND2_X1 U9086 ( .A1(n7895), .A2(n7894), .ZN(n7788) );
  XNOR2_X1 U9087 ( .A(n7672), .B(n7788), .ZN(n7542) );
  OAI22_X1 U9088 ( .A1(n7673), .A2(n8496), .B1(n7535), .B2(n8498), .ZN(n7541)
         );
  NOR2_X1 U9089 ( .A1(n8607), .A2(n8211), .ZN(n7536) );
  AOI21_X1 U9090 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(n7539) );
  OAI21_X1 U9091 ( .B1(n7539), .B2(n7788), .A(n8026), .ZN(n8606) );
  NOR2_X1 U9092 ( .A1(n8606), .A2(n8532), .ZN(n7540) );
  AOI211_X1 U9093 ( .C1(n8511), .C2(n7542), .A(n7541), .B(n7540), .ZN(n8605)
         );
  XOR2_X1 U9094 ( .A(n8045), .B(n8602), .Z(n8603) );
  INV_X1 U9095 ( .A(n8602), .ZN(n7545) );
  AOI22_X1 U9096 ( .A1(n8467), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7543), .B2(
        n9751), .ZN(n7544) );
  OAI21_X1 U9097 ( .B1(n7545), .B2(n8469), .A(n7544), .ZN(n7548) );
  NOR2_X1 U9098 ( .A1(n8606), .A2(n7546), .ZN(n7547) );
  AOI211_X1 U9099 ( .C1(n8603), .C2(n8521), .A(n7548), .B(n7547), .ZN(n7549)
         );
  OAI21_X1 U9100 ( .B1(n8605), .B2(n8467), .A(n7549), .ZN(P2_U3280) );
  INV_X1 U9101 ( .A(n7733), .ZN(n7570) );
  AOI21_X1 U9102 ( .B1(n9429), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7550), .ZN(
        n7551) );
  OAI21_X1 U9103 ( .B1(n7570), .B2(n7552), .A(n7551), .ZN(P1_U3326) );
  NAND2_X1 U9104 ( .A1(n7555), .A2(n5928), .ZN(n7557) );
  NAND2_X1 U9105 ( .A1(n7747), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7556) );
  XNOR2_X1 U9106 ( .A(n8582), .B(n7995), .ZN(n7586) );
  NAND2_X1 U9107 ( .A1(n8454), .A2(n7985), .ZN(n7585) );
  XNOR2_X1 U9108 ( .A(n7586), .B(n7585), .ZN(n7588) );
  XNOR2_X1 U9109 ( .A(n7589), .B(n7588), .ZN(n7568) );
  OAI22_X1 U9110 ( .A1(n8162), .A2(n8441), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7558), .ZN(n7566) );
  XNOR2_X1 U9111 ( .A(n7598), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U9112 ( .A1(n8424), .A2(n5816), .ZN(n7564) );
  INV_X1 U9113 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n7561) );
  NAND2_X1 U9114 ( .A1(n5912), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9115 ( .A1(n5800), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7559) );
  OAI211_X1 U9116 ( .C1(n7561), .C2(n7728), .A(n7560), .B(n7559), .ZN(n7562)
         );
  INV_X1 U9117 ( .A(n7562), .ZN(n7563) );
  NAND2_X1 U9118 ( .A1(n7564), .A2(n7563), .ZN(n8434) );
  INV_X1 U9119 ( .A(n8434), .ZN(n8412) );
  OAI22_X1 U9120 ( .A1(n7675), .A2(n8200), .B1(n8202), .B2(n8412), .ZN(n7565)
         );
  AOI211_X1 U9121 ( .C1(n8582), .C2(n4315), .A(n7566), .B(n7565), .ZN(n7567)
         );
  OAI21_X1 U9122 ( .B1(n7568), .B2(n8196), .A(n7567), .ZN(P2_U3235) );
  OAI222_X1 U9123 ( .A1(n8647), .A2(n7570), .B1(P2_U3152), .B2(n8056), .C1(
        n7569), .C2(n8641), .ZN(P2_U3331) );
  AOI21_X1 U9124 ( .B1(n7572), .B2(n6068), .A(n7571), .ZN(n8229) );
  XNOR2_X1 U9125 ( .A(n8229), .B(n8230), .ZN(n7573) );
  NOR2_X1 U9126 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7573), .ZN(n8231) );
  AOI21_X1 U9127 ( .B1(n7573), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8231), .ZN(
        n7584) );
  AND2_X1 U9128 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7575) );
  NOR2_X1 U9129 ( .A1(n9730), .A2(n8224), .ZN(n7574) );
  AOI211_X1 U9130 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9738), .A(n7575), .B(
        n7574), .ZN(n7583) );
  XNOR2_X1 U9131 ( .A(n8223), .B(n8224), .ZN(n7578) );
  INV_X1 U9132 ( .A(n7578), .ZN(n7581) );
  INV_X1 U9133 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7579) );
  NOR2_X1 U9134 ( .A1(n7579), .A2(n7578), .ZN(n8225) );
  INV_X1 U9135 ( .A(n8225), .ZN(n7580) );
  OAI211_X1 U9136 ( .C1(n7581), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9734), .B(
        n7580), .ZN(n7582) );
  OAI211_X1 U9137 ( .C1(n7584), .C2(n8282), .A(n7583), .B(n7582), .ZN(P2_U3260) );
  INV_X1 U9138 ( .A(n7585), .ZN(n7587) );
  NAND2_X1 U9139 ( .A1(n7590), .A2(n5928), .ZN(n7592) );
  NAND2_X1 U9140 ( .A1(n7747), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7591) );
  XNOR2_X1 U9141 ( .A(n8576), .B(n7593), .ZN(n7973) );
  NAND2_X1 U9142 ( .A1(n8434), .A2(n7985), .ZN(n7972) );
  XNOR2_X1 U9143 ( .A(n7973), .B(n7972), .ZN(n7974) );
  XNOR2_X1 U9144 ( .A(n4384), .B(n7974), .ZN(n7609) );
  INV_X1 U9145 ( .A(n8424), .ZN(n7594) );
  INV_X1 U9146 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7596) );
  OAI22_X1 U9147 ( .A1(n8162), .A2(n7594), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7596), .ZN(n7607) );
  INV_X1 U9148 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7595) );
  OAI21_X1 U9149 ( .B1(n7598), .B2(n7596), .A(n7595), .ZN(n7599) );
  NAND2_X1 U9150 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n7597) );
  AND2_X1 U9151 ( .A1(n7599), .A2(n7688), .ZN(n8405) );
  NAND2_X1 U9152 ( .A1(n8405), .A2(n5816), .ZN(n7605) );
  INV_X1 U9153 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9154 ( .A1(n7764), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7601) );
  NAND2_X1 U9155 ( .A1(n5912), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7600) );
  OAI211_X1 U9156 ( .C1(n7742), .C2(n7602), .A(n7601), .B(n7600), .ZN(n7603)
         );
  INV_X1 U9157 ( .A(n7603), .ZN(n7604) );
  OAI22_X1 U9158 ( .A1(n7676), .A2(n8200), .B1(n8202), .B2(n8038), .ZN(n7606)
         );
  AOI211_X1 U9159 ( .C1(n8576), .C2(n4315), .A(n7607), .B(n7606), .ZN(n7608)
         );
  OAI21_X1 U9160 ( .B1(n7609), .B2(n8196), .A(n7608), .ZN(P2_U3225) );
  INV_X1 U9161 ( .A(n7614), .ZN(n7610) );
  NOR2_X1 U9162 ( .A1(n7611), .A2(n7610), .ZN(n7616) );
  AOI21_X1 U9163 ( .B1(n7614), .B2(n7613), .A(n7612), .ZN(n7615) );
  OAI21_X1 U9164 ( .B1(n7616), .B2(n7615), .A(n8683), .ZN(n7621) );
  NAND2_X1 U9165 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9103) );
  INV_X1 U9166 ( .A(n9103), .ZN(n7617) );
  AOI21_X1 U9167 ( .B1(n8664), .B2(n9054), .A(n7617), .ZN(n7618) );
  OAI21_X1 U9168 ( .B1(n7633), .B2(n8706), .A(n7618), .ZN(n7619) );
  AOI21_X1 U9169 ( .B1(n4859), .B2(n8726), .A(n7619), .ZN(n7620) );
  OAI211_X1 U9170 ( .C1(n4613), .C2(n8730), .A(n7621), .B(n7620), .ZN(P1_U3226) );
  NAND2_X1 U9171 ( .A1(n7622), .A2(n8893), .ZN(n7625) );
  NAND2_X1 U9172 ( .A1(n7623), .A2(n9054), .ZN(n7624) );
  NAND2_X1 U9173 ( .A1(n7625), .A2(n7624), .ZN(n7643) );
  AND2_X1 U9174 ( .A1(n9391), .A2(n8724), .ZN(n8921) );
  INV_X1 U9175 ( .A(n8921), .ZN(n8747) );
  OR2_X1 U9176 ( .A1(n9391), .A2(n8724), .ZN(n8085) );
  XOR2_X1 U9177 ( .A(n7643), .B(n8895), .Z(n9394) );
  AOI211_X1 U9178 ( .C1(n9391), .C2(n7626), .A(n9706), .B(n4374), .ZN(n9390)
         );
  AOI22_X1 U9179 ( .A1(n9648), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n4859), .B2(
        n9314), .ZN(n7627) );
  OAI21_X1 U9180 ( .B1(n4613), .B2(n9623), .A(n7627), .ZN(n7631) );
  XNOR2_X1 U9181 ( .A(n7634), .B(n8895), .ZN(n7629) );
  AOI222_X1 U9182 ( .A1(n9313), .A2(n7629), .B1(n9300), .B2(n9631), .C1(n9054), 
        .C2(n9633), .ZN(n9393) );
  NOR2_X1 U9183 ( .A1(n9393), .A2(n9648), .ZN(n7630) );
  AOI211_X1 U9184 ( .C1(n9390), .C2(n9322), .A(n7631), .B(n7630), .ZN(n7632)
         );
  OAI21_X1 U9185 ( .B1(n9306), .B2(n9394), .A(n7632), .ZN(P1_U3274) );
  OR2_X1 U9186 ( .A1(n9386), .A2(n7633), .ZN(n8809) );
  NAND2_X1 U9187 ( .A1(n9386), .A2(n7633), .ZN(n9297) );
  NAND2_X1 U9188 ( .A1(n9295), .A2(n8085), .ZN(n7635) );
  XOR2_X1 U9189 ( .A(n8896), .B(n7635), .Z(n7636) );
  AOI222_X1 U9190 ( .A1(n9313), .A2(n7636), .B1(n9053), .B2(n9633), .C1(n9279), 
        .C2(n9631), .ZN(n9388) );
  INV_X1 U9191 ( .A(n9386), .ZN(n8731) );
  OAI21_X1 U9192 ( .B1(n4374), .B2(n8731), .A(n9667), .ZN(n7637) );
  NOR2_X1 U9193 ( .A1(n7637), .A2(n9287), .ZN(n9385) );
  INV_X1 U9194 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U9195 ( .A1(n9386), .A2(n9316), .ZN(n7639) );
  NAND2_X1 U9196 ( .A1(n9314), .A2(n8727), .ZN(n7638) );
  OAI211_X1 U9197 ( .C1(n9646), .C2(n7640), .A(n7639), .B(n7638), .ZN(n7648)
         );
  AND2_X1 U9198 ( .A1(n9391), .A2(n9053), .ZN(n7642) );
  OR2_X1 U9199 ( .A1(n9391), .A2(n9053), .ZN(n7641) );
  OAI21_X1 U9200 ( .B1(n7643), .B2(n7642), .A(n7641), .ZN(n7644) );
  INV_X1 U9201 ( .A(n7644), .ZN(n7646) );
  INV_X1 U9202 ( .A(n8896), .ZN(n7645) );
  OAI21_X1 U9203 ( .B1(n7646), .B2(n7645), .A(n8073), .ZN(n9389) );
  NOR2_X1 U9204 ( .A1(n9389), .A2(n9306), .ZN(n7647) );
  AOI211_X1 U9205 ( .C1(n9385), .C2(n9322), .A(n7648), .B(n7647), .ZN(n7649)
         );
  OAI21_X1 U9206 ( .B1(n9648), .B2(n9388), .A(n7649), .ZN(P1_U3273) );
  INV_X1 U9207 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10069) );
  INV_X1 U9208 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10060) );
  OR2_X1 U9209 ( .A1(n5850), .A2(n10060), .ZN(n7651) );
  NAND2_X1 U9210 ( .A1(n7764), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7650) );
  OAI211_X1 U9211 ( .C1(n7742), .C2(n10069), .A(n7651), .B(n7650), .ZN(n8294)
         );
  INV_X1 U9212 ( .A(n8294), .ZN(n7780) );
  NAND2_X1 U9213 ( .A1(n7780), .A2(n7829), .ZN(n7771) );
  INV_X1 U9214 ( .A(SI_28_), .ZN(n7654) );
  NAND2_X1 U9215 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  INV_X1 U9216 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9947) );
  INV_X1 U9217 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7657) );
  MUX2_X1 U9218 ( .A(n9947), .B(n7657), .S(n7775), .Z(n7759) );
  INV_X1 U9219 ( .A(SI_29_), .ZN(n7658) );
  AND2_X1 U9220 ( .A1(n7759), .A2(n7658), .ZN(n7661) );
  INV_X1 U9221 ( .A(n7759), .ZN(n7659) );
  NAND2_X1 U9222 ( .A1(n7659), .A2(SI_29_), .ZN(n7660) );
  INV_X1 U9223 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7663) );
  INV_X1 U9224 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7662) );
  MUX2_X1 U9225 ( .A(n7663), .B(n7662), .S(n7775), .Z(n7665) );
  INV_X1 U9226 ( .A(SI_30_), .ZN(n7664) );
  NAND2_X1 U9227 ( .A1(n7665), .A2(n7664), .ZN(n7772) );
  INV_X1 U9228 ( .A(n7665), .ZN(n7666) );
  NAND2_X1 U9229 ( .A1(n7666), .A2(SI_30_), .ZN(n7667) );
  NAND2_X1 U9230 ( .A1(n7772), .A2(n7667), .ZN(n7773) );
  NAND2_X1 U9231 ( .A1(n8737), .A2(n5928), .ZN(n7669) );
  NAND2_X1 U9232 ( .A1(n7747), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7668) );
  INV_X1 U9233 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U9234 ( .A1(n5912), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9235 ( .A1(n7764), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7670) );
  OAI211_X1 U9236 ( .C1(n7742), .C2(n8300), .A(n7671), .B(n7670), .ZN(n8208)
         );
  AND2_X1 U9237 ( .A1(n8299), .A2(n8208), .ZN(n7787) );
  INV_X1 U9238 ( .A(n7787), .ZN(n7944) );
  NAND2_X1 U9239 ( .A1(n8599), .A2(n7673), .ZN(n7822) );
  NAND2_X1 U9240 ( .A1(n8493), .A2(n8492), .ZN(n7674) );
  NAND2_X1 U9241 ( .A1(n7674), .A2(n7824), .ZN(n8471) );
  OR2_X1 U9242 ( .A1(n8592), .A2(n8495), .ZN(n7900) );
  NAND2_X1 U9243 ( .A1(n8592), .A2(n8495), .ZN(n7902) );
  NAND2_X1 U9244 ( .A1(n7900), .A2(n7902), .ZN(n8472) );
  NAND2_X1 U9245 ( .A1(n8473), .A2(n7902), .ZN(n8451) );
  OR2_X1 U9246 ( .A1(n8588), .A2(n7675), .ZN(n7901) );
  NAND2_X1 U9247 ( .A1(n8588), .A2(n7675), .ZN(n8432) );
  NAND2_X1 U9248 ( .A1(n8582), .A2(n7676), .ZN(n7911) );
  INV_X1 U9249 ( .A(n8432), .ZN(n7907) );
  OR2_X1 U9250 ( .A1(n8576), .A2(n8412), .ZN(n7915) );
  NAND2_X1 U9251 ( .A1(n8576), .A2(n8412), .ZN(n8409) );
  NAND2_X1 U9252 ( .A1(n7915), .A2(n8409), .ZN(n8419) );
  NAND2_X1 U9253 ( .A1(n7678), .A2(n5928), .ZN(n7680) );
  NAND2_X1 U9254 ( .A1(n7747), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U9255 ( .A1(n8571), .A2(n8038), .ZN(n7917) );
  INV_X1 U9256 ( .A(n8409), .ZN(n7681) );
  NOR2_X1 U9257 ( .A1(n4746), .A2(n7681), .ZN(n7682) );
  NAND2_X1 U9258 ( .A1(n7683), .A2(n5928), .ZN(n7685) );
  NAND2_X1 U9259 ( .A1(n7747), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7684) );
  INV_X1 U9260 ( .A(n7688), .ZN(n7686) );
  NAND2_X1 U9261 ( .A1(n7686), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7700) );
  INV_X1 U9262 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9263 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  NAND2_X1 U9264 ( .A1(n7700), .A2(n7689), .ZN(n8395) );
  OR2_X1 U9265 ( .A1(n8395), .A2(n7763), .ZN(n7694) );
  INV_X1 U9266 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U9267 ( .A1(n5912), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9268 ( .A1(n5800), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7690) );
  OAI211_X1 U9269 ( .C1(n7728), .C2(n8569), .A(n7691), .B(n7690), .ZN(n7692)
         );
  INV_X1 U9270 ( .A(n7692), .ZN(n7693) );
  OR2_X1 U9271 ( .A1(n8397), .A2(n8413), .ZN(n7919) );
  NAND2_X1 U9272 ( .A1(n8397), .A2(n8413), .ZN(n7918) );
  INV_X1 U9273 ( .A(n8379), .ZN(n8385) );
  INV_X1 U9274 ( .A(n8384), .ZN(n7695) );
  NOR2_X1 U9275 ( .A1(n8385), .A2(n7695), .ZN(n7696) );
  INV_X1 U9276 ( .A(n8371), .ZN(n7708) );
  NAND2_X1 U9277 ( .A1(n7697), .A2(n5928), .ZN(n7699) );
  NAND2_X1 U9278 ( .A1(n7747), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7698) );
  INV_X1 U9279 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U9280 ( .A1(n7700), .A2(n8161), .ZN(n7701) );
  NAND2_X1 U9281 ( .A1(n7714), .A2(n7701), .ZN(n8367) );
  OR2_X1 U9282 ( .A1(n8367), .A2(n7763), .ZN(n7707) );
  INV_X1 U9283 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U9284 ( .A1(n7764), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U9285 ( .A1(n5912), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7702) );
  OAI211_X1 U9286 ( .C1(n7742), .C2(n7704), .A(n7703), .B(n7702), .ZN(n7705)
         );
  INV_X1 U9287 ( .A(n7705), .ZN(n7706) );
  NAND2_X1 U9288 ( .A1(n7707), .A2(n7706), .ZN(n8390) );
  XNOR2_X1 U9289 ( .A(n8558), .B(n8390), .ZN(n8039) );
  INV_X1 U9290 ( .A(n8390), .ZN(n8142) );
  OR2_X1 U9291 ( .A1(n8558), .A2(n8142), .ZN(n7922) );
  NAND2_X1 U9292 ( .A1(n7709), .A2(n5928), .ZN(n7711) );
  NAND2_X1 U9293 ( .A1(n7747), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7710) );
  INV_X1 U9294 ( .A(n7714), .ZN(n7712) );
  NAND2_X1 U9295 ( .A1(n7712), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7724) );
  INV_X1 U9296 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U9297 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  NAND2_X1 U9298 ( .A1(n7724), .A2(n7715), .ZN(n8353) );
  OR2_X1 U9299 ( .A1(n8353), .A2(n7763), .ZN(n7720) );
  INV_X1 U9300 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U9301 ( .A1(n5800), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9302 ( .A1(n5912), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7716) );
  OAI211_X1 U9303 ( .C1(n10061), .C2(n7728), .A(n7717), .B(n7716), .ZN(n7718)
         );
  INV_X1 U9304 ( .A(n7718), .ZN(n7719) );
  NAND2_X1 U9305 ( .A1(n8554), .A2(n8372), .ZN(n7928) );
  NAND2_X1 U9306 ( .A1(n7927), .A2(n7928), .ZN(n8355) );
  INV_X1 U9307 ( .A(n8355), .ZN(n7926) );
  NAND2_X1 U9308 ( .A1(n7721), .A2(n5928), .ZN(n7723) );
  NAND2_X1 U9309 ( .A1(n7747), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7722) );
  INV_X1 U9310 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U9311 ( .A1(n7724), .A2(n8199), .ZN(n7725) );
  NAND2_X1 U9312 ( .A1(n8345), .A2(n5816), .ZN(n7732) );
  INV_X1 U9313 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U9314 ( .A1(n5800), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7727) );
  NAND2_X1 U9315 ( .A1(n5912), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7726) );
  OAI211_X1 U9316 ( .C1(n7729), .C2(n7728), .A(n7727), .B(n7726), .ZN(n7730)
         );
  INV_X1 U9317 ( .A(n7730), .ZN(n7731) );
  NAND2_X1 U9318 ( .A1(n8549), .A2(n8143), .ZN(n7930) );
  NAND2_X1 U9319 ( .A1(n7931), .A2(n7930), .ZN(n8337) );
  INV_X1 U9320 ( .A(n8337), .ZN(n7810) );
  NAND2_X1 U9321 ( .A1(n7733), .A2(n5928), .ZN(n7735) );
  NAND2_X1 U9322 ( .A1(n7747), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7734) );
  INV_X1 U9323 ( .A(n7738), .ZN(n7736) );
  NAND2_X1 U9324 ( .A1(n7736), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7751) );
  INV_X1 U9325 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U9326 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  NAND2_X1 U9327 ( .A1(n7751), .A2(n7739), .ZN(n8327) );
  INV_X1 U9328 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U9329 ( .A1(n5912), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U9330 ( .A1(n7764), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7740) );
  OAI211_X1 U9331 ( .C1(n8328), .C2(n7742), .A(n7741), .B(n7740), .ZN(n7743)
         );
  INV_X1 U9332 ( .A(n7743), .ZN(n7744) );
  XNOR2_X1 U9333 ( .A(n8543), .B(n8201), .ZN(n8323) );
  INV_X1 U9334 ( .A(n8323), .ZN(n7808) );
  OR2_X1 U9335 ( .A1(n8543), .A2(n8201), .ZN(n7819) );
  NAND2_X1 U9336 ( .A1(n7746), .A2(n7819), .ZN(n8304) );
  NAND2_X1 U9337 ( .A1(n8643), .A2(n5928), .ZN(n7749) );
  NAND2_X1 U9338 ( .A1(n7747), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7748) );
  INV_X1 U9339 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U9340 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U9341 ( .A1(n8048), .A2(n7752), .ZN(n8313) );
  INV_X1 U9342 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U9343 ( .A1(n7764), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U9344 ( .A1(n5912), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7753) );
  OAI211_X1 U9345 ( .C1(n7742), .C2(n8312), .A(n7754), .B(n7753), .ZN(n7755)
         );
  INV_X1 U9346 ( .A(n7755), .ZN(n7756) );
  NAND2_X1 U9347 ( .A1(n8537), .A2(n8126), .ZN(n7935) );
  NAND2_X1 U9348 ( .A1(n7934), .A2(n7935), .ZN(n8308) );
  INV_X1 U9349 ( .A(n8308), .ZN(n7811) );
  XNOR2_X1 U9350 ( .A(n7759), .B(SI_29_), .ZN(n7760) );
  NAND2_X1 U9351 ( .A1(n8640), .A2(n5928), .ZN(n7762) );
  NAND2_X1 U9352 ( .A1(n7747), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7761) );
  OR2_X1 U9353 ( .A1(n8048), .A2(n7763), .ZN(n7770) );
  INV_X1 U9354 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U9355 ( .A1(n7764), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U9356 ( .A1(n5800), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7765) );
  OAI211_X1 U9357 ( .C1(n5850), .C2(n7767), .A(n7766), .B(n7765), .ZN(n7768)
         );
  INV_X1 U9358 ( .A(n7768), .ZN(n7769) );
  NAND2_X1 U9359 ( .A1(n8533), .A2(n8007), .ZN(n7941) );
  INV_X1 U9360 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7776) );
  MUX2_X1 U9361 ( .A(n6222), .B(n7776), .S(n7775), .Z(n7777) );
  XNOR2_X1 U9362 ( .A(n7777), .B(SI_31_), .ZN(n7778) );
  XNOR2_X1 U9363 ( .A(n7779), .B(n7778), .ZN(n8732) );
  INV_X1 U9364 ( .A(n8292), .ZN(n7781) );
  INV_X1 U9365 ( .A(n8208), .ZN(n7782) );
  NAND2_X1 U9366 ( .A1(n8528), .A2(n7782), .ZN(n7943) );
  XNOR2_X1 U9367 ( .A(n7784), .B(n9753), .ZN(n7785) );
  INV_X1 U9368 ( .A(n7818), .ZN(n7814) );
  NOR2_X1 U9369 ( .A1(n7949), .A2(n7787), .ZN(n7817) );
  INV_X1 U9370 ( .A(n7817), .ZN(n7813) );
  INV_X1 U9371 ( .A(n8452), .ZN(n8448) );
  INV_X1 U9372 ( .A(n8492), .ZN(n7805) );
  INV_X1 U9373 ( .A(n7788), .ZN(n7892) );
  NOR2_X1 U9374 ( .A1(n7789), .A2(n6835), .ZN(n7793) );
  NOR2_X1 U9375 ( .A1(n9806), .A2(n7790), .ZN(n7792) );
  AND2_X1 U9376 ( .A1(n9744), .A2(n7791), .ZN(n7825) );
  NAND4_X1 U9377 ( .A1(n7793), .A2(n7834), .A3(n7792), .A4(n7825), .ZN(n7796)
         );
  INV_X1 U9378 ( .A(n8516), .ZN(n7795) );
  INV_X1 U9379 ( .A(n7843), .ZN(n7794) );
  NOR4_X1 U9380 ( .A1(n7797), .A2(n7796), .A3(n7795), .A4(n7794), .ZN(n7798)
         );
  NAND4_X1 U9381 ( .A1(n7800), .A2(n7799), .A3(n7853), .A4(n7798), .ZN(n7801)
         );
  NOR4_X1 U9382 ( .A1(n7886), .A2(n6963), .A3(n7802), .A4(n7801), .ZN(n7803)
         );
  NAND4_X1 U9383 ( .A1(n7892), .A2(n7887), .A3(n7803), .A4(n7879), .ZN(n7804)
         );
  NOR4_X1 U9384 ( .A1(n8448), .A2(n7805), .A3(n8472), .A4(n7804), .ZN(n7806)
         );
  NAND4_X1 U9385 ( .A1(n8408), .A2(n8437), .A3(n7677), .A4(n7806), .ZN(n7807)
         );
  NOR4_X1 U9386 ( .A1(n8355), .A2(n8370), .A3(n8385), .A4(n7807), .ZN(n7809)
         );
  NAND4_X1 U9387 ( .A1(n7811), .A2(n7810), .A3(n7809), .A4(n7808), .ZN(n7812)
         );
  XNOR2_X1 U9388 ( .A(n7815), .B(n8499), .ZN(n7954) );
  NOR2_X1 U9389 ( .A1(n7953), .A2(n8499), .ZN(n7816) );
  MUX2_X1 U9390 ( .A(n7818), .B(n7817), .S(n7947), .Z(n7952) );
  INV_X1 U9391 ( .A(n7819), .ZN(n7821) );
  INV_X1 U9392 ( .A(n8543), .ZN(n8326) );
  OAI21_X1 U9393 ( .B1(n8326), .B2(n8340), .A(n7935), .ZN(n7820) );
  MUX2_X1 U9394 ( .A(n7821), .B(n7820), .S(n7947), .Z(n7938) );
  AND2_X1 U9395 ( .A1(n7902), .A2(n7822), .ZN(n7823) );
  INV_X1 U9396 ( .A(n7947), .ZN(n7939) );
  MUX2_X1 U9397 ( .A(n7824), .B(n7823), .S(n7939), .Z(n7899) );
  MUX2_X1 U9398 ( .A(n7825), .B(n7843), .S(n7947), .Z(n7845) );
  INV_X1 U9399 ( .A(n7826), .ZN(n7828) );
  NAND2_X1 U9400 ( .A1(n7848), .A2(n9744), .ZN(n7827) );
  AND2_X1 U9401 ( .A1(n7835), .A2(n7829), .ZN(n7830) );
  OAI211_X1 U9402 ( .C1(n7831), .C2(n7830), .A(n7839), .B(n6419), .ZN(n7832)
         );
  NAND3_X1 U9403 ( .A1(n7832), .A2(n7838), .A3(n7947), .ZN(n7833) );
  NAND2_X1 U9404 ( .A1(n6419), .A2(n7835), .ZN(n7837) );
  NAND3_X1 U9405 ( .A1(n7838), .A2(n7837), .A3(n7836), .ZN(n7840) );
  NAND3_X1 U9406 ( .A1(n7840), .A2(n7939), .A3(n7839), .ZN(n7841) );
  INV_X1 U9407 ( .A(n9743), .ZN(n7844) );
  OAI21_X1 U9408 ( .B1(n7848), .B2(n7947), .A(n7847), .ZN(n7849) );
  MUX2_X1 U9409 ( .A(n7851), .B(n7850), .S(n7947), .Z(n7852) );
  NAND2_X1 U9410 ( .A1(n7853), .A2(n7852), .ZN(n7855) );
  OAI22_X1 U9411 ( .A1(n7856), .A2(n7855), .B1(n7939), .B2(n7854), .ZN(n7857)
         );
  NAND2_X1 U9412 ( .A1(n7857), .A2(n7859), .ZN(n7865) );
  AND2_X1 U9413 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  MUX2_X1 U9414 ( .A(n7862), .B(n7860), .S(n7939), .Z(n7864) );
  OAI21_X1 U9415 ( .B1(n7862), .B2(n7947), .A(n7861), .ZN(n7863) );
  AOI21_X1 U9416 ( .B1(n7865), .B2(n7864), .A(n7863), .ZN(n7871) );
  NAND2_X1 U9417 ( .A1(n7872), .A2(n7866), .ZN(n7869) );
  NAND2_X1 U9418 ( .A1(n7875), .A2(n7867), .ZN(n7868) );
  MUX2_X1 U9419 ( .A(n7869), .B(n7868), .S(n7947), .Z(n7870) );
  OR2_X1 U9420 ( .A1(n7871), .A2(n7870), .ZN(n7877) );
  NAND3_X1 U9421 ( .A1(n7877), .A2(n7878), .A3(n7872), .ZN(n7873) );
  NAND3_X1 U9422 ( .A1(n7877), .A2(n7876), .A3(n7875), .ZN(n7880) );
  MUX2_X1 U9423 ( .A(n7884), .B(n7883), .S(n7947), .Z(n7885) );
  NAND2_X1 U9424 ( .A1(n7888), .A2(n7887), .ZN(n7893) );
  MUX2_X1 U9425 ( .A(n7890), .B(n7889), .S(n7947), .Z(n7891) );
  NAND3_X1 U9426 ( .A1(n7893), .A2(n7892), .A3(n7891), .ZN(n7897) );
  MUX2_X1 U9427 ( .A(n7895), .B(n7894), .S(n7947), .Z(n7896) );
  NAND3_X1 U9428 ( .A1(n7897), .A2(n8492), .A3(n7896), .ZN(n7898) );
  NAND2_X1 U9429 ( .A1(n7899), .A2(n7898), .ZN(n7909) );
  NAND2_X1 U9430 ( .A1(n7901), .A2(n7900), .ZN(n7906) );
  AOI21_X1 U9431 ( .B1(n7909), .B2(n7902), .A(n7906), .ZN(n7904) );
  NAND2_X1 U9432 ( .A1(n7911), .A2(n8432), .ZN(n7903) );
  OAI211_X1 U9433 ( .C1(n7904), .C2(n7903), .A(n7910), .B(n7915), .ZN(n7905)
         );
  INV_X1 U9434 ( .A(n7906), .ZN(n7908) );
  AOI21_X1 U9435 ( .B1(n7909), .B2(n7908), .A(n7907), .ZN(n7913) );
  INV_X1 U9436 ( .A(n7910), .ZN(n7912) );
  OAI211_X1 U9437 ( .C1(n7913), .C2(n7912), .A(n8409), .B(n7911), .ZN(n7914)
         );
  NAND3_X1 U9438 ( .A1(n8384), .A2(n7915), .A3(n7914), .ZN(n7916) );
  MUX2_X1 U9439 ( .A(n7919), .B(n7918), .S(n7947), .Z(n7920) );
  NAND3_X1 U9440 ( .A1(n7921), .A2(n8039), .A3(n7920), .ZN(n7925) );
  NAND2_X1 U9441 ( .A1(n8558), .A2(n8142), .ZN(n7923) );
  MUX2_X1 U9442 ( .A(n7923), .B(n7922), .S(n7947), .Z(n7924) );
  NAND2_X1 U9443 ( .A1(n7930), .A2(n7928), .ZN(n7929) );
  NOR2_X1 U9444 ( .A1(n7931), .A2(n7939), .ZN(n7932) );
  NAND2_X1 U9445 ( .A1(n7933), .A2(n7934), .ZN(n7937) );
  MUX2_X1 U9446 ( .A(n7935), .B(n7934), .S(n7947), .Z(n7936) );
  OAI211_X1 U9447 ( .C1(n7938), .C2(n7937), .A(n8053), .B(n7936), .ZN(n7945)
         );
  MUX2_X1 U9448 ( .A(n7941), .B(n7940), .S(n7939), .Z(n7942) );
  NAND4_X1 U9449 ( .A1(n7945), .A2(n7944), .A3(n7943), .A4(n7942), .ZN(n7951)
         );
  INV_X1 U9450 ( .A(n7946), .ZN(n7948) );
  MUX2_X1 U9451 ( .A(n7949), .B(n7948), .S(n7947), .Z(n7950) );
  AOI211_X1 U9452 ( .C1(n6052), .C2(n7957), .A(n7956), .B(n7955), .ZN(n7958)
         );
  NOR2_X1 U9453 ( .A1(n7959), .A2(n8056), .ZN(n7962) );
  OAI21_X1 U9454 ( .B1(n7963), .B2(n7960), .A(P2_B_REG_SCAN_IN), .ZN(n7961) );
  OAI22_X1 U9455 ( .A1(n7964), .A2(n7963), .B1(n7962), .B2(n7961), .ZN(
        P2_U3244) );
  AOI22_X1 U9456 ( .A1(n8168), .A2(n6691), .B1(n7965), .B2(n4315), .ZN(n7971)
         );
  OAI21_X1 U9457 ( .B1(n7968), .B2(n7967), .A(n7966), .ZN(n7969) );
  OR2_X1 U9458 ( .A1(n8067), .A2(P2_U3152), .ZN(n8169) );
  AOI22_X1 U9459 ( .A1(n8185), .A2(n7969), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8169), .ZN(n7970) );
  OAI211_X1 U9460 ( .C1(n8200), .C2(n8064), .A(n7971), .B(n7970), .ZN(P2_U3224) );
  XNOR2_X1 U9461 ( .A(n8571), .B(n7995), .ZN(n7978) );
  INV_X1 U9462 ( .A(n7978), .ZN(n7975) );
  NAND2_X1 U9463 ( .A1(n7976), .A2(n7985), .ZN(n7977) );
  NAND2_X1 U9464 ( .A1(n8018), .A2(n7977), .ZN(n8024) );
  OR2_X1 U9465 ( .A1(n7979), .A2(n7978), .ZN(n7980) );
  XNOR2_X1 U9466 ( .A(n8397), .B(n7995), .ZN(n7982) );
  NOR2_X1 U9467 ( .A1(n8413), .A2(n7994), .ZN(n8131) );
  INV_X1 U9468 ( .A(n7981), .ZN(n7983) );
  XNOR2_X1 U9469 ( .A(n8558), .B(n7995), .ZN(n7984) );
  NOR2_X1 U9470 ( .A1(n8142), .A2(n7994), .ZN(n8157) );
  XOR2_X1 U9471 ( .A(n7995), .B(n8554), .Z(n8140) );
  NAND2_X1 U9472 ( .A1(n8339), .A2(n7985), .ZN(n8139) );
  XNOR2_X1 U9473 ( .A(n8549), .B(n7995), .ZN(n8121) );
  NOR2_X1 U9474 ( .A1(n8143), .A2(n7994), .ZN(n7986) );
  NAND2_X1 U9475 ( .A1(n8121), .A2(n7986), .ZN(n7987) );
  OAI21_X1 U9476 ( .B1(n8121), .B2(n7986), .A(n7987), .ZN(n8198) );
  XNOR2_X1 U9477 ( .A(n8543), .B(n7995), .ZN(n7988) );
  NOR2_X1 U9478 ( .A1(n8201), .A2(n7994), .ZN(n7989) );
  NAND2_X1 U9479 ( .A1(n7988), .A2(n7989), .ZN(n7993) );
  INV_X1 U9480 ( .A(n7988), .ZN(n7991) );
  INV_X1 U9481 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U9482 ( .A1(n7991), .A2(n7990), .ZN(n7992) );
  AND2_X1 U9483 ( .A1(n7993), .A2(n7992), .ZN(n8120) );
  NAND2_X1 U9484 ( .A1(n8124), .A2(n7993), .ZN(n8006) );
  NOR2_X1 U9485 ( .A1(n8126), .A2(n7994), .ZN(n7996) );
  XNOR2_X1 U9486 ( .A(n7996), .B(n7995), .ZN(n7998) );
  INV_X1 U9487 ( .A(n7998), .ZN(n7999) );
  NOR3_X1 U9488 ( .A1(n8047), .A2(n4315), .A3(n7999), .ZN(n7997) );
  AOI21_X1 U9489 ( .B1(n8047), .B2(n7999), .A(n7997), .ZN(n8005) );
  OAI21_X1 U9490 ( .B1(n8047), .B2(n8207), .A(n8196), .ZN(n8004) );
  NOR3_X1 U9491 ( .A1(n8047), .A2(n7998), .A3(n4315), .ZN(n8001) );
  NOR2_X1 U9492 ( .A1(n8537), .A2(n7999), .ZN(n8000) );
  NAND2_X1 U9493 ( .A1(n8006), .A2(n8002), .ZN(n8003) );
  OAI211_X1 U9494 ( .C1(n8006), .C2(n8005), .A(n8004), .B(n8003), .ZN(n8012)
         );
  INV_X1 U9495 ( .A(n8007), .ZN(n8305) );
  AOI22_X1 U9496 ( .A1(n8168), .A2(n8305), .B1(n8190), .B2(n8340), .ZN(n8010)
         );
  INV_X1 U9497 ( .A(n8313), .ZN(n8008) );
  AOI22_X1 U9498 ( .A1(n8205), .A2(n8008), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8009) );
  AND2_X1 U9499 ( .A1(n8010), .A2(n8009), .ZN(n8011) );
  NAND2_X1 U9500 ( .A1(n8012), .A2(n8011), .ZN(P2_U3222) );
  OAI222_X1 U9501 ( .A1(n8641), .A2(n8017), .B1(n8016), .B2(n8015), .C1(n8014), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NOR3_X1 U9502 ( .A1(n8018), .A2(n8038), .A3(n8189), .ZN(n8022) );
  AOI22_X1 U9503 ( .A1(n8205), .A2(n8405), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8020) );
  INV_X1 U9504 ( .A(n8413), .ZN(n8209) );
  AOI22_X1 U9505 ( .A1(n8168), .A2(n8209), .B1(n8190), .B2(n8434), .ZN(n8019)
         );
  OAI211_X1 U9506 ( .C1(n4745), .C2(n8207), .A(n8020), .B(n8019), .ZN(n8021)
         );
  NOR2_X1 U9507 ( .A1(n8022), .A2(n8021), .ZN(n8023) );
  OAI21_X1 U9508 ( .B1(n8024), .B2(n8196), .A(n8023), .ZN(P2_U3237) );
  NAND2_X1 U9509 ( .A1(n8602), .A2(n8210), .ZN(n8025) );
  OR2_X1 U9510 ( .A1(n8592), .A2(n8453), .ZN(n8027) );
  OR2_X1 U9511 ( .A1(n8599), .A2(n8477), .ZN(n8462) );
  AND2_X1 U9512 ( .A1(n8027), .A2(n8462), .ZN(n8028) );
  NAND2_X1 U9513 ( .A1(n8592), .A2(n8453), .ZN(n8029) );
  NAND2_X1 U9514 ( .A1(n8030), .A2(n8029), .ZN(n8449) );
  AND2_X1 U9515 ( .A1(n8588), .A2(n8476), .ZN(n8032) );
  OAI21_X2 U9516 ( .B1(n8449), .B2(n8032), .A(n8031), .ZN(n8438) );
  NAND2_X1 U9517 ( .A1(n8582), .A2(n8454), .ZN(n8034) );
  OR2_X1 U9518 ( .A1(n8576), .A2(n8434), .ZN(n8035) );
  NAND2_X1 U9519 ( .A1(n8576), .A2(n8434), .ZN(n8036) );
  NAND2_X1 U9520 ( .A1(n8037), .A2(n8036), .ZN(n8404) );
  NAND2_X1 U9521 ( .A1(n8351), .A2(n8355), .ZN(n8350) );
  NAND2_X1 U9522 ( .A1(n8350), .A2(n8040), .ZN(n8334) );
  NAND2_X1 U9523 ( .A1(n8334), .A2(n8337), .ZN(n8333) );
  NAND2_X1 U9524 ( .A1(n8333), .A2(n8041), .ZN(n8324) );
  NAND2_X1 U9525 ( .A1(n8324), .A2(n8323), .ZN(n8322) );
  NAND2_X1 U9526 ( .A1(n8322), .A2(n8042), .ZN(n8309) );
  NAND2_X1 U9527 ( .A1(n8309), .A2(n8308), .ZN(n8307) );
  INV_X1 U9528 ( .A(n8549), .ZN(n8336) );
  INV_X1 U9529 ( .A(n8576), .ZN(n8426) );
  INV_X1 U9530 ( .A(n8582), .ZN(n8444) );
  INV_X1 U9531 ( .A(n8599), .ZN(n8046) );
  NAND2_X1 U9532 ( .A1(n8488), .A2(n8046), .ZN(n8489) );
  NOR2_X2 U9533 ( .A1(n8588), .A2(n8464), .ZN(n8456) );
  NOR2_X2 U9534 ( .A1(n8554), .A2(n8365), .ZN(n8359) );
  NAND2_X1 U9535 ( .A1(n8336), .A2(n8359), .ZN(n8342) );
  NOR2_X2 U9536 ( .A1(n8342), .A2(n8543), .ZN(n8310) );
  NOR2_X2 U9537 ( .A1(n8533), .A2(n8311), .ZN(n8298) );
  INV_X1 U9538 ( .A(n8048), .ZN(n8049) );
  AOI22_X1 U9539 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(n8467), .B1(n8049), .B2(
        n9751), .ZN(n8050) );
  OAI21_X1 U9540 ( .B1(n4673), .B2(n8469), .A(n8050), .ZN(n8061) );
  OAI21_X1 U9541 ( .B1(n8053), .B2(n8052), .A(n8051), .ZN(n8054) );
  NAND2_X1 U9542 ( .A1(n8054), .A2(n8511), .ZN(n8059) );
  NOR2_X1 U9543 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  NOR2_X1 U9544 ( .A1(n8496), .A2(n8057), .ZN(n8293) );
  NOR2_X1 U9545 ( .A1(n4322), .A2(n8467), .ZN(n8060) );
  OAI21_X1 U9546 ( .B1(n8535), .B2(n8504), .A(n8062), .ZN(P2_U3267) );
  OAI22_X1 U9547 ( .A1(n8189), .A2(n8064), .B1(n8063), .B2(n8196), .ZN(n8066)
         );
  NAND2_X1 U9548 ( .A1(n8066), .A2(n8065), .ZN(n8071) );
  NAND2_X1 U9549 ( .A1(n8067), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U9550 ( .A1(P2_U3152), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U9551 ( .A1(n8068), .A2(n9736), .ZN(n8069) );
  AOI21_X1 U9552 ( .B1(n4315), .B2(n9804), .A(n8069), .ZN(n8070) );
  OAI211_X1 U9553 ( .C1(n8202), .C2(n6412), .A(n8071), .B(n8070), .ZN(P2_U3234) );
  INV_X1 U9554 ( .A(n9173), .ZN(n9052) );
  NAND2_X1 U9555 ( .A1(n9386), .A2(n9300), .ZN(n8072) );
  OR2_X1 U9556 ( .A1(n9381), .A2(n9279), .ZN(n8075) );
  AND2_X1 U9557 ( .A1(n9381), .A2(n9279), .ZN(n8074) );
  NAND2_X1 U9558 ( .A1(n9375), .A2(n9301), .ZN(n8076) );
  NAND2_X1 U9559 ( .A1(n9264), .A2(n8703), .ZN(n8826) );
  NAND2_X1 U9560 ( .A1(n9240), .A2(n8826), .ZN(n9254) );
  INV_X1 U9561 ( .A(n9260), .ZN(n8676) );
  INV_X1 U9562 ( .A(n9364), .ZN(n9239) );
  NAND2_X1 U9563 ( .A1(n9222), .A2(n8077), .ZN(n8078) );
  INV_X1 U9564 ( .A(n9354), .ZN(n9213) );
  NAND2_X1 U9565 ( .A1(n9348), .A2(n9214), .ZN(n8835) );
  NOR2_X1 U9566 ( .A1(n9343), .A2(n9203), .ZN(n8839) );
  OAI22_X1 U9567 ( .A1(n9180), .A2(n8839), .B1(n10115), .B2(n9185), .ZN(n9166)
         );
  NAND2_X1 U9568 ( .A1(n9339), .A2(n8079), .ZN(n8917) );
  OAI22_X1 U9569 ( .A1(n9166), .A2(n8901), .B1(n9190), .B2(n9339), .ZN(n9150)
         );
  NAND2_X1 U9570 ( .A1(n9333), .A2(n9173), .ZN(n8918) );
  NOR2_X1 U9571 ( .A1(n9150), .A2(n9158), .ZN(n9149) );
  NAND2_X1 U9572 ( .A1(n8640), .A2(n8080), .ZN(n8082) );
  NAND2_X1 U9573 ( .A1(n5399), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8081) );
  NOR2_X1 U9574 ( .A1(n9327), .A2(n8860), .ZN(n8989) );
  INV_X1 U9575 ( .A(n9381), .ZN(n9293) );
  NAND2_X1 U9576 ( .A1(n9287), .A2(n9293), .ZN(n9288) );
  NOR2_X1 U9577 ( .A1(n9265), .A2(n9364), .ZN(n9248) );
  NAND2_X1 U9578 ( .A1(n9248), .A2(n9228), .ZN(n9223) );
  NOR2_X2 U9579 ( .A1(n9209), .A2(n9348), .ZN(n9196) );
  AND2_X2 U9580 ( .A1(n9185), .A2(n9196), .ZN(n9181) );
  AOI21_X1 U9581 ( .B1(n9327), .B2(n9152), .A(n9143), .ZN(n9328) );
  INV_X1 U9582 ( .A(n9327), .ZN(n8861) );
  AOI22_X1 U9583 ( .A1(n9648), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8083), .B2(
        n9314), .ZN(n8084) );
  OAI21_X1 U9584 ( .B1(n8861), .B2(n9623), .A(n8084), .ZN(n8104) );
  AND2_X1 U9585 ( .A1(n8809), .A2(n8085), .ZN(n9294) );
  INV_X1 U9586 ( .A(n9279), .ZN(n8692) );
  OR2_X1 U9587 ( .A1(n9381), .A2(n8692), .ZN(n8815) );
  OR2_X1 U9588 ( .A1(n9296), .A2(n9297), .ZN(n8086) );
  INV_X1 U9589 ( .A(n9301), .ZN(n8674) );
  AND2_X1 U9590 ( .A1(n9375), .A2(n8674), .ZN(n8871) );
  OR2_X1 U9591 ( .A1(n9375), .A2(n8674), .ZN(n8872) );
  INV_X1 U9592 ( .A(n9254), .ZN(n9259) );
  NAND2_X1 U9593 ( .A1(n9364), .A2(n8676), .ZN(n8828) );
  NAND3_X1 U9594 ( .A1(n9257), .A2(n9244), .A3(n9240), .ZN(n9243) );
  NAND2_X1 U9595 ( .A1(n9243), .A2(n8828), .ZN(n9232) );
  NAND2_X1 U9596 ( .A1(n9358), .A2(n8705), .ZN(n8976) );
  NAND2_X1 U9597 ( .A1(n8829), .A2(n8976), .ZN(n9231) );
  INV_X1 U9598 ( .A(n8829), .ZN(n8087) );
  OR2_X1 U9599 ( .A1(n9354), .A2(n9229), .ZN(n8743) );
  NAND2_X1 U9600 ( .A1(n9354), .A2(n9229), .ZN(n8978) );
  NAND2_X1 U9601 ( .A1(n8743), .A2(n8978), .ZN(n9215) );
  NAND2_X1 U9602 ( .A1(n8743), .A2(n8829), .ZN(n8919) );
  INV_X1 U9603 ( .A(n8835), .ZN(n8979) );
  OR2_X1 U9604 ( .A1(n9343), .A2(n10115), .ZN(n8088) );
  NAND2_X1 U9605 ( .A1(n8088), .A2(n9186), .ZN(n8982) );
  NAND2_X1 U9606 ( .A1(n9343), .A2(n10115), .ZN(n8914) );
  INV_X1 U9607 ( .A(n8984), .ZN(n8089) );
  NAND2_X1 U9608 ( .A1(n9157), .A2(n8918), .ZN(n8090) );
  XNOR2_X1 U9609 ( .A(n8090), .B(n8870), .ZN(n8102) );
  INV_X1 U9610 ( .A(n9313), .ZN(n8091) );
  OR2_X1 U9611 ( .A1(n9173), .A2(n9618), .ZN(n8101) );
  INV_X1 U9612 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U9613 ( .A1(n8092), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U9614 ( .A1(n8093), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8094) );
  OAI211_X1 U9615 ( .C1(n8097), .C2(n8096), .A(n8095), .B(n8094), .ZN(n9051)
         );
  INV_X1 U9616 ( .A(n9051), .ZN(n8100) );
  AND2_X1 U9617 ( .A1(n9036), .A2(P1_B_REG_SCAN_IN), .ZN(n8098) );
  NOR2_X1 U9618 ( .A1(n9616), .A2(n8098), .ZN(n9138) );
  INV_X1 U9619 ( .A(n9138), .ZN(n8099) );
  NOR2_X1 U9620 ( .A1(n9330), .A2(n9648), .ZN(n8103) );
  OAI21_X1 U9621 ( .B1(n9332), .B2(n9306), .A(n8105), .ZN(P1_U3355) );
  OR2_X1 U9622 ( .A1(n8149), .A2(n8107), .ZN(n8109) );
  NAND2_X1 U9623 ( .A1(n8109), .A2(n8108), .ZN(n8112) );
  OAI211_X1 U9624 ( .C1(n8112), .C2(n8111), .A(n8110), .B(n8185), .ZN(n8119)
         );
  AOI22_X1 U9625 ( .A1(n8168), .A2(n8218), .B1(n8113), .B2(n8205), .ZN(n8118)
         );
  NAND2_X1 U9626 ( .A1(n4315), .A2(n6854), .ZN(n8114) );
  OAI21_X1 U9627 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8115), .A(n8114), .ZN(n8116) );
  AOI21_X1 U9628 ( .B1(n8190), .B2(n8219), .A(n8116), .ZN(n8117) );
  NAND3_X1 U9629 ( .A1(n8119), .A2(n8118), .A3(n8117), .ZN(P2_U3215) );
  NOR2_X1 U9630 ( .A1(n8195), .A2(n8120), .ZN(n8123) );
  NAND3_X1 U9631 ( .A1(n8121), .A2(n8156), .A3(n8320), .ZN(n8122) );
  OAI21_X1 U9632 ( .B1(n8123), .B2(n8196), .A(n8122), .ZN(n8125) );
  NAND2_X1 U9633 ( .A1(n8125), .A2(n8124), .ZN(n8130) );
  NOR2_X1 U9634 ( .A1(n8162), .A2(n8327), .ZN(n8128) );
  OAI22_X1 U9635 ( .A1(n8126), .A2(n8202), .B1(n8200), .B2(n8143), .ZN(n8127)
         );
  AOI211_X1 U9636 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n8128), 
        .B(n8127), .ZN(n8129) );
  OAI211_X1 U9637 ( .C1(n8326), .C2(n8207), .A(n8130), .B(n8129), .ZN(P2_U3216) );
  NAND2_X1 U9638 ( .A1(n8156), .A2(n8209), .ZN(n8134) );
  OR2_X1 U9639 ( .A1(n8196), .A2(n8131), .ZN(n8133) );
  MUX2_X1 U9640 ( .A(n8134), .B(n8133), .S(n8132), .Z(n8138) );
  AOI22_X1 U9641 ( .A1(n8190), .A2(n7976), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8135) );
  OAI21_X1 U9642 ( .B1(n8162), .B2(n8395), .A(n8135), .ZN(n8136) );
  AOI21_X1 U9643 ( .B1(n8168), .B2(n8390), .A(n8136), .ZN(n8137) );
  OAI211_X1 U9644 ( .C1(n8563), .C2(n8207), .A(n8138), .B(n8137), .ZN(P2_U3218) );
  XNOR2_X1 U9645 ( .A(n8140), .B(n8139), .ZN(n8141) );
  XNOR2_X1 U9646 ( .A(n4342), .B(n8141), .ZN(n8147) );
  OAI22_X1 U9647 ( .A1(n8143), .A2(n8496), .B1(n8142), .B2(n8498), .ZN(n8357)
         );
  AOI22_X1 U9648 ( .A1(n8357), .A2(n8152), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8144) );
  OAI21_X1 U9649 ( .B1(n8353), .B2(n8162), .A(n8144), .ZN(n8145) );
  AOI21_X1 U9650 ( .B1(n8554), .B2(n4315), .A(n8145), .ZN(n8146) );
  OAI21_X1 U9651 ( .B1(n8147), .B2(n8196), .A(n8146), .ZN(P2_U3227) );
  AOI21_X1 U9652 ( .B1(n8149), .B2(n8148), .A(n8196), .ZN(n8150) );
  OR2_X1 U9653 ( .A1(n8149), .A2(n8148), .ZN(n8184) );
  NAND2_X1 U9654 ( .A1(n8150), .A2(n8184), .ZN(n8155) );
  AOI22_X1 U9655 ( .A1(n8220), .A2(n8506), .B1(n8508), .B2(n8219), .ZN(n9758)
         );
  INV_X1 U9656 ( .A(n9758), .ZN(n8151) );
  AOI22_X1 U9657 ( .A1(n8152), .A2(n8151), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8154) );
  AOI22_X1 U9658 ( .A1(n4315), .A2(n9748), .B1(n8205), .B2(n9750), .ZN(n8153)
         );
  NAND3_X1 U9659 ( .A1(n8155), .A2(n8154), .A3(n8153), .ZN(P2_U3229) );
  NAND2_X1 U9660 ( .A1(n8156), .A2(n8390), .ZN(n8160) );
  OR2_X1 U9661 ( .A1(n8196), .A2(n8157), .ZN(n8159) );
  MUX2_X1 U9662 ( .A(n8160), .B(n8159), .S(n8158), .Z(n8167) );
  OAI22_X1 U9663 ( .A1(n8162), .A2(n8367), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8161), .ZN(n8164) );
  OAI22_X1 U9664 ( .A1(n8413), .A2(n8200), .B1(n8202), .B2(n8372), .ZN(n8163)
         );
  AOI211_X1 U9665 ( .C1(n8558), .C2(n4315), .A(n8164), .B(n8163), .ZN(n8166)
         );
  NAND2_X1 U9666 ( .A1(n8167), .A2(n8166), .ZN(P2_U3231) );
  AOI22_X1 U9667 ( .A1(n8168), .A2(n8221), .B1(n8190), .B2(n6829), .ZN(n8177)
         );
  AOI22_X1 U9668 ( .A1(n4315), .A2(n8170), .B1(n8169), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8176) );
  AOI21_X1 U9669 ( .B1(n8172), .B2(n8171), .A(n8196), .ZN(n8174) );
  NAND2_X1 U9670 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  NAND3_X1 U9671 ( .A1(n8177), .A2(n8176), .A3(n8175), .ZN(P2_U3239) );
  OAI22_X1 U9672 ( .A1(n8202), .A2(n8179), .B1(n8178), .B2(n8207), .ZN(n8180)
         );
  AOI211_X1 U9673 ( .C1(n8513), .C2(n8205), .A(n8181), .B(n8180), .ZN(n8194)
         );
  NAND2_X1 U9674 ( .A1(n8184), .A2(n8182), .ZN(n8183) );
  OAI21_X1 U9675 ( .B1(n8187), .B2(n8184), .A(n8183), .ZN(n8186) );
  NAND2_X1 U9676 ( .A1(n8186), .A2(n8185), .ZN(n8193) );
  NOR3_X1 U9677 ( .A1(n8189), .A2(n8188), .A3(n8187), .ZN(n8191) );
  OAI21_X1 U9678 ( .B1(n8191), .B2(n8190), .A(n8507), .ZN(n8192) );
  NAND3_X1 U9679 ( .A1(n8194), .A2(n8193), .A3(n8192), .ZN(P2_U3241) );
  OAI22_X1 U9680 ( .A1(n8200), .A2(n8372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8199), .ZN(n8204) );
  NOR2_X1 U9681 ( .A1(n8202), .A2(n8201), .ZN(n8203) );
  AOI211_X1 U9682 ( .C1(n8205), .C2(n8345), .A(n8204), .B(n8203), .ZN(n8206)
         );
  MUX2_X1 U9683 ( .A(n8294), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8222), .Z(
        P2_U3583) );
  MUX2_X1 U9684 ( .A(n8208), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8222), .Z(
        P2_U3582) );
  MUX2_X1 U9685 ( .A(n8305), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8222), .Z(
        P2_U3581) );
  MUX2_X1 U9686 ( .A(n8319), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8222), .Z(
        P2_U3580) );
  MUX2_X1 U9687 ( .A(n8340), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8222), .Z(
        P2_U3579) );
  MUX2_X1 U9688 ( .A(n8320), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8222), .Z(
        P2_U3578) );
  MUX2_X1 U9689 ( .A(n8339), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8222), .Z(
        P2_U3577) );
  MUX2_X1 U9690 ( .A(n8390), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8222), .Z(
        P2_U3576) );
  MUX2_X1 U9691 ( .A(n8209), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8222), .Z(
        P2_U3575) );
  MUX2_X1 U9692 ( .A(n7976), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8222), .Z(
        P2_U3574) );
  MUX2_X1 U9693 ( .A(n8434), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8222), .Z(
        P2_U3573) );
  MUX2_X1 U9694 ( .A(n8454), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8222), .Z(
        P2_U3572) );
  MUX2_X1 U9695 ( .A(n8453), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8222), .Z(
        P2_U3570) );
  MUX2_X1 U9696 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8477), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9697 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8210), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9698 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8211), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9699 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8212), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9700 ( .A(n8213), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8222), .Z(
        P2_U3565) );
  MUX2_X1 U9701 ( .A(n8214), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8222), .Z(
        P2_U3564) );
  MUX2_X1 U9702 ( .A(n8215), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8222), .Z(
        P2_U3563) );
  MUX2_X1 U9703 ( .A(n8216), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8222), .Z(
        P2_U3562) );
  MUX2_X1 U9704 ( .A(n8217), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8222), .Z(
        P2_U3561) );
  MUX2_X1 U9705 ( .A(n8218), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8222), .Z(
        P2_U3560) );
  MUX2_X1 U9706 ( .A(n8509), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8222), .Z(
        P2_U3559) );
  MUX2_X1 U9707 ( .A(n8219), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8222), .Z(
        P2_U3558) );
  MUX2_X1 U9708 ( .A(n8507), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8222), .Z(
        P2_U3557) );
  MUX2_X1 U9709 ( .A(n8220), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8222), .Z(
        P2_U3556) );
  MUX2_X1 U9710 ( .A(n8221), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8222), .Z(
        P2_U3555) );
  MUX2_X1 U9711 ( .A(n6691), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8222), .Z(
        P2_U3554) );
  MUX2_X1 U9712 ( .A(n6829), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8222), .Z(
        P2_U3553) );
  NOR2_X1 U9713 ( .A1(n8224), .A2(n8223), .ZN(n8226) );
  NOR2_X1 U9714 ( .A1(n8226), .A2(n8225), .ZN(n8228) );
  XOR2_X1 U9715 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8250), .Z(n8227) );
  NAND2_X1 U9716 ( .A1(n8227), .A2(n8228), .ZN(n8249) );
  OAI21_X1 U9717 ( .B1(n8228), .B2(n8227), .A(n8249), .ZN(n8242) );
  NOR2_X1 U9718 ( .A1(n8230), .A2(n8229), .ZN(n8232) );
  NOR2_X1 U9719 ( .A1(n8232), .A2(n8231), .ZN(n8235) );
  NAND2_X1 U9720 ( .A1(n8250), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8245) );
  INV_X1 U9721 ( .A(n8245), .ZN(n8233) );
  AOI21_X1 U9722 ( .B1(n7073), .B2(n8240), .A(n8233), .ZN(n8234) );
  NAND2_X1 U9723 ( .A1(n8234), .A2(n8235), .ZN(n8244) );
  OAI211_X1 U9724 ( .C1(n8235), .C2(n8234), .A(n9735), .B(n8244), .ZN(n8239)
         );
  INV_X1 U9725 ( .A(n8236), .ZN(n8237) );
  AOI21_X1 U9726 ( .B1(n9738), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8237), .ZN(
        n8238) );
  OAI211_X1 U9727 ( .C1(n9730), .C2(n8240), .A(n8239), .B(n8238), .ZN(n8241)
         );
  AOI21_X1 U9728 ( .B1(n9734), .B2(n8242), .A(n8241), .ZN(n8243) );
  INV_X1 U9729 ( .A(n8243), .ZN(P2_U3261) );
  NAND2_X1 U9730 ( .A1(n8245), .A2(n8244), .ZN(n8247) );
  XNOR2_X1 U9731 ( .A(n8258), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U9732 ( .A1(n8246), .A2(n8247), .ZN(n8257) );
  OAI211_X1 U9733 ( .C1(n8247), .C2(n8246), .A(n9735), .B(n8257), .ZN(n8256)
         );
  NOR2_X1 U9734 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8248), .ZN(n8254) );
  XNOR2_X1 U9735 ( .A(n8264), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8251) );
  AOI211_X1 U9736 ( .C1(n8252), .C2(n8251), .A(n8263), .B(n9731), .ZN(n8253)
         );
  AOI211_X1 U9737 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9738), .A(n8254), .B(
        n8253), .ZN(n8255) );
  OAI211_X1 U9738 ( .C1(n9730), .C2(n8258), .A(n8256), .B(n8255), .ZN(P2_U3262) );
  OAI21_X1 U9739 ( .B1(n8258), .B2(n8487), .A(n8257), .ZN(n8259) );
  NOR2_X1 U9740 ( .A1(n8259), .A2(n8276), .ZN(n8271) );
  AOI21_X1 U9741 ( .B1(n8276), .B2(n8259), .A(n8271), .ZN(n8260) );
  INV_X1 U9742 ( .A(n8260), .ZN(n8261) );
  NOR2_X1 U9743 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8261), .ZN(n8272) );
  AOI21_X1 U9744 ( .B1(n8261), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8272), .ZN(
        n8270) );
  XNOR2_X1 U9745 ( .A(n8276), .B(n8262), .ZN(n8275) );
  XNOR2_X1 U9746 ( .A(n8275), .B(n8274), .ZN(n8267) );
  INV_X1 U9747 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U9748 ( .A1(n8291), .A2(n10125), .ZN(n8265) );
  AOI211_X1 U9749 ( .C1(n9734), .C2(n8267), .A(n8266), .B(n8265), .ZN(n8269)
         );
  NAND2_X1 U9750 ( .A1(n8285), .A2(n8276), .ZN(n8268) );
  OAI211_X1 U9751 ( .C1(n8270), .C2(n8282), .A(n8269), .B(n8268), .ZN(P2_U3263) );
  NOR2_X1 U9752 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  XOR2_X1 U9753 ( .A(n8273), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8283) );
  OR2_X1 U9754 ( .A1(n8276), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U9755 ( .A1(n8278), .A2(n8277), .ZN(n8280) );
  XNOR2_X1 U9756 ( .A(n8280), .B(n8279), .ZN(n8286) );
  INV_X1 U9757 ( .A(n8286), .ZN(n8281) );
  AOI22_X1 U9758 ( .A1(n8283), .A2(n9735), .B1(n8281), .B2(n9734), .ZN(n8288)
         );
  NOR2_X1 U9759 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  AOI211_X1 U9760 ( .C1(n9734), .C2(n8286), .A(n8285), .B(n8284), .ZN(n8287)
         );
  MUX2_X1 U9761 ( .A(n8288), .B(n8287), .S(n9753), .Z(n8290) );
  OAI211_X1 U9762 ( .C1(n4912), .C2(n8291), .A(n8290), .B(n8289), .ZN(P2_U3264) );
  NAND2_X1 U9763 ( .A1(n8299), .A2(n8298), .ZN(n8297) );
  XNOR2_X1 U9764 ( .A(n8292), .B(n8297), .ZN(n8526) );
  NAND2_X1 U9765 ( .A1(n8526), .A2(n8521), .ZN(n8296) );
  NAND2_X1 U9766 ( .A1(n8294), .A2(n8293), .ZN(n8530) );
  NOR2_X1 U9767 ( .A1(n8467), .A2(n8530), .ZN(n8301) );
  AOI21_X1 U9768 ( .B1(n8467), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8301), .ZN(
        n8295) );
  OAI211_X1 U9769 ( .C1(n8292), .C2(n8469), .A(n8296), .B(n8295), .ZN(P2_U3265) );
  OAI21_X1 U9770 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8531) );
  NOR2_X1 U9771 ( .A1(n9763), .A2(n8300), .ZN(n8302) );
  AOI211_X1 U9772 ( .C1(n8528), .C2(n8514), .A(n8302), .B(n8301), .ZN(n8303)
         );
  OAI21_X1 U9773 ( .B1(n8400), .B2(n8531), .A(n8303), .ZN(P2_U3266) );
  XNOR2_X1 U9774 ( .A(n8304), .B(n8308), .ZN(n8306) );
  AOI222_X1 U9775 ( .A1(n8511), .A2(n8306), .B1(n8340), .B2(n8506), .C1(n8305), 
        .C2(n8508), .ZN(n8540) );
  OAI21_X1 U9776 ( .B1(n8309), .B2(n8308), .A(n8307), .ZN(n8536) );
  NAND2_X1 U9777 ( .A1(n8536), .A2(n8518), .ZN(n8317) );
  AOI21_X1 U9778 ( .B1(n8537), .B2(n8325), .A(n4674), .ZN(n8538) );
  NOR2_X1 U9779 ( .A1(n8047), .A2(n8469), .ZN(n8315) );
  OAI22_X1 U9780 ( .A1(n8313), .A2(n8485), .B1(n9763), .B2(n8312), .ZN(n8314)
         );
  AOI211_X1 U9781 ( .C1(n8538), .C2(n8521), .A(n8315), .B(n8314), .ZN(n8316)
         );
  OAI211_X1 U9782 ( .C1(n8467), .C2(n8540), .A(n8317), .B(n8316), .ZN(P2_U3268) );
  XNOR2_X1 U9783 ( .A(n8318), .B(n8323), .ZN(n8321) );
  AOI222_X1 U9784 ( .A1(n8511), .A2(n8321), .B1(n8320), .B2(n8506), .C1(n8319), 
        .C2(n8508), .ZN(n8546) );
  OAI21_X1 U9785 ( .B1(n8324), .B2(n8323), .A(n8322), .ZN(n8542) );
  NAND2_X1 U9786 ( .A1(n8542), .A2(n8518), .ZN(n8332) );
  AOI21_X1 U9787 ( .B1(n8543), .B2(n8342), .A(n8310), .ZN(n8544) );
  NOR2_X1 U9788 ( .A1(n8326), .A2(n8469), .ZN(n8330) );
  OAI22_X1 U9789 ( .A1(n8328), .A2(n9763), .B1(n8327), .B2(n8485), .ZN(n8329)
         );
  AOI211_X1 U9790 ( .C1(n8544), .C2(n8521), .A(n8330), .B(n8329), .ZN(n8331)
         );
  OAI211_X1 U9791 ( .C1(n8467), .C2(n8546), .A(n8332), .B(n8331), .ZN(P2_U3269) );
  OAI21_X1 U9792 ( .B1(n8334), .B2(n8337), .A(n8333), .ZN(n8335) );
  INV_X1 U9793 ( .A(n8335), .ZN(n8552) );
  NOR2_X1 U9794 ( .A1(n8336), .A2(n8469), .ZN(n8348) );
  XNOR2_X1 U9795 ( .A(n8338), .B(n8337), .ZN(n8341) );
  AOI222_X1 U9796 ( .A1(n8511), .A2(n8341), .B1(n8340), .B2(n8508), .C1(n8339), 
        .C2(n8506), .ZN(n8551) );
  INV_X1 U9797 ( .A(n8359), .ZN(n8344) );
  INV_X1 U9798 ( .A(n8342), .ZN(n8343) );
  AOI211_X1 U9799 ( .C1(n8549), .C2(n8344), .A(n9881), .B(n8343), .ZN(n8548)
         );
  AOI22_X1 U9800 ( .A1(n8548), .A2(n8499), .B1(n9751), .B2(n8345), .ZN(n8346)
         );
  AOI21_X1 U9801 ( .B1(n8551), .B2(n8346), .A(n8467), .ZN(n8347) );
  AOI211_X1 U9802 ( .C1(n8467), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8348), .B(
        n8347), .ZN(n8349) );
  OAI21_X1 U9803 ( .B1(n8552), .B2(n8504), .A(n8349), .ZN(P2_U3270) );
  OAI21_X1 U9804 ( .B1(n8351), .B2(n8355), .A(n8350), .ZN(n8352) );
  INV_X1 U9805 ( .A(n8352), .ZN(n8557) );
  INV_X1 U9806 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8354) );
  OAI22_X1 U9807 ( .A1(n9763), .A2(n8354), .B1(n8353), .B2(n8485), .ZN(n8362)
         );
  XNOR2_X1 U9808 ( .A(n8356), .B(n8355), .ZN(n8358) );
  AOI21_X1 U9809 ( .B1(n8358), .B2(n8511), .A(n8357), .ZN(n8556) );
  AOI211_X1 U9810 ( .C1(n8554), .C2(n8365), .A(n9881), .B(n8359), .ZN(n8553)
         );
  NAND2_X1 U9811 ( .A1(n8553), .A2(n8499), .ZN(n8360) );
  AOI21_X1 U9812 ( .B1(n8556), .B2(n8360), .A(n8467), .ZN(n8361) );
  AOI211_X1 U9813 ( .C1(n8514), .C2(n8554), .A(n8362), .B(n8361), .ZN(n8363)
         );
  OAI21_X1 U9814 ( .B1(n8557), .B2(n8504), .A(n8363), .ZN(P2_U3271) );
  XNOR2_X1 U9815 ( .A(n8364), .B(n8370), .ZN(n8562) );
  INV_X1 U9816 ( .A(n8365), .ZN(n8366) );
  AOI21_X1 U9817 ( .B1(n8558), .B2(n8393), .A(n8366), .ZN(n8559) );
  INV_X1 U9818 ( .A(n8367), .ZN(n8368) );
  AOI22_X1 U9819 ( .A1(n8467), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8368), .B2(
        n9751), .ZN(n8369) );
  OAI21_X1 U9820 ( .B1(n4678), .B2(n8469), .A(n8369), .ZN(n8377) );
  AOI21_X1 U9821 ( .B1(n8371), .B2(n8370), .A(n9759), .ZN(n8375) );
  OAI22_X1 U9822 ( .A1(n8372), .A2(n8496), .B1(n8413), .B2(n8498), .ZN(n8373)
         );
  AOI21_X1 U9823 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8561) );
  NOR2_X1 U9824 ( .A1(n8561), .A2(n8467), .ZN(n8376) );
  AOI211_X1 U9825 ( .C1(n8559), .C2(n8521), .A(n8377), .B(n8376), .ZN(n8378)
         );
  OAI21_X1 U9826 ( .B1(n8562), .B2(n8504), .A(n8378), .ZN(P2_U3272) );
  NAND2_X1 U9827 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  INV_X1 U9828 ( .A(n8568), .ZN(n8403) );
  NAND2_X1 U9829 ( .A1(n8383), .A2(n8384), .ZN(n8386) );
  NAND2_X1 U9830 ( .A1(n8386), .A2(n8385), .ZN(n8388) );
  NAND2_X1 U9831 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  NAND2_X1 U9832 ( .A1(n8389), .A2(n8511), .ZN(n8392) );
  AOI22_X1 U9833 ( .A1(n8390), .A2(n8508), .B1(n7976), .B2(n8506), .ZN(n8391)
         );
  NAND2_X1 U9834 ( .A1(n8392), .A2(n8391), .ZN(n8566) );
  OR2_X1 U9835 ( .A1(n8563), .A2(n4338), .ZN(n8394) );
  NAND2_X1 U9836 ( .A1(n8394), .A2(n8393), .ZN(n8564) );
  INV_X1 U9837 ( .A(n8395), .ZN(n8396) );
  AOI22_X1 U9838 ( .A1(n8467), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8396), .B2(
        n9751), .ZN(n8399) );
  NAND2_X1 U9839 ( .A1(n8397), .A2(n8514), .ZN(n8398) );
  OAI211_X1 U9840 ( .C1(n8564), .C2(n8400), .A(n8399), .B(n8398), .ZN(n8401)
         );
  AOI21_X1 U9841 ( .B1(n8566), .B2(n9763), .A(n8401), .ZN(n8402) );
  OAI21_X1 U9842 ( .B1(n8403), .B2(n8504), .A(n8402), .ZN(P2_U3273) );
  XNOR2_X1 U9843 ( .A(n8404), .B(n4746), .ZN(n8575) );
  AOI21_X1 U9844 ( .B1(n8571), .B2(n8421), .A(n4338), .ZN(n8572) );
  AOI22_X1 U9845 ( .A1(n8467), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8405), .B2(
        n9751), .ZN(n8406) );
  OAI21_X1 U9846 ( .B1(n4745), .B2(n8469), .A(n8406), .ZN(n8417) );
  INV_X1 U9847 ( .A(n8383), .ZN(n8411) );
  AOI21_X1 U9848 ( .B1(n8407), .B2(n8409), .A(n8408), .ZN(n8410) );
  NOR3_X1 U9849 ( .A1(n8411), .A2(n8410), .A3(n9759), .ZN(n8415) );
  OAI22_X1 U9850 ( .A1(n8413), .A2(n8496), .B1(n8412), .B2(n8498), .ZN(n8414)
         );
  NOR2_X1 U9851 ( .A1(n8415), .A2(n8414), .ZN(n8574) );
  NOR2_X1 U9852 ( .A1(n8574), .A2(n8467), .ZN(n8416) );
  AOI211_X1 U9853 ( .C1(n8572), .C2(n8521), .A(n8417), .B(n8416), .ZN(n8418)
         );
  OAI21_X1 U9854 ( .B1(n8575), .B2(n8504), .A(n8418), .ZN(P2_U3274) );
  XNOR2_X1 U9855 ( .A(n8420), .B(n8419), .ZN(n8580) );
  INV_X1 U9856 ( .A(n8439), .ZN(n8423) );
  INV_X1 U9857 ( .A(n8421), .ZN(n8422) );
  AOI21_X1 U9858 ( .B1(n8576), .B2(n8423), .A(n8422), .ZN(n8577) );
  AOI22_X1 U9859 ( .A1(n8467), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8424), .B2(
        n9751), .ZN(n8425) );
  OAI21_X1 U9860 ( .B1(n8426), .B2(n8469), .A(n8425), .ZN(n8430) );
  OAI21_X1 U9861 ( .B1(n8427), .B2(n7677), .A(n8407), .ZN(n8428) );
  AOI222_X1 U9862 ( .A1(n8511), .A2(n8428), .B1(n7976), .B2(n8508), .C1(n8454), 
        .C2(n8506), .ZN(n8579) );
  NOR2_X1 U9863 ( .A1(n8579), .A2(n8467), .ZN(n8429) );
  AOI211_X1 U9864 ( .C1(n8577), .C2(n8521), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI21_X1 U9865 ( .B1(n8504), .B2(n8580), .A(n8431), .ZN(P2_U3275) );
  NAND2_X1 U9866 ( .A1(n8450), .A2(n8432), .ZN(n8433) );
  XNOR2_X1 U9867 ( .A(n8433), .B(n8437), .ZN(n8435) );
  AOI222_X1 U9868 ( .A1(n8511), .A2(n8435), .B1(n8434), .B2(n8508), .C1(n8476), 
        .C2(n8506), .ZN(n8585) );
  NAND2_X1 U9869 ( .A1(n8438), .A2(n8437), .ZN(n8581) );
  NAND3_X1 U9870 ( .A1(n8436), .A2(n8581), .A3(n8518), .ZN(n8447) );
  INV_X1 U9871 ( .A(n8456), .ZN(n8440) );
  AOI21_X1 U9872 ( .B1(n8582), .B2(n8440), .A(n8439), .ZN(n8583) );
  INV_X1 U9873 ( .A(n8441), .ZN(n8442) );
  AOI22_X1 U9874 ( .A1(n8467), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8442), .B2(
        n9751), .ZN(n8443) );
  OAI21_X1 U9875 ( .B1(n8444), .B2(n8469), .A(n8443), .ZN(n8445) );
  AOI21_X1 U9876 ( .B1(n8583), .B2(n8521), .A(n8445), .ZN(n8446) );
  OAI211_X1 U9877 ( .C1(n8467), .C2(n8585), .A(n8447), .B(n8446), .ZN(P2_U3276) );
  XNOR2_X1 U9878 ( .A(n8449), .B(n8448), .ZN(n8591) );
  AOI22_X1 U9879 ( .A1(n8588), .A2(n8514), .B1(n8467), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8461) );
  OAI21_X1 U9880 ( .B1(n8452), .B2(n8451), .A(n8450), .ZN(n8455) );
  AOI222_X1 U9881 ( .A1(n8511), .A2(n8455), .B1(n8454), .B2(n8508), .C1(n8453), 
        .C2(n8506), .ZN(n8590) );
  AOI211_X1 U9882 ( .C1(n8588), .C2(n8464), .A(n9881), .B(n8456), .ZN(n8587)
         );
  AOI22_X1 U9883 ( .A1(n8587), .A2(n8499), .B1(n9751), .B2(n8457), .ZN(n8458)
         );
  AOI21_X1 U9884 ( .B1(n8590), .B2(n8458), .A(n8467), .ZN(n8459) );
  INV_X1 U9885 ( .A(n8459), .ZN(n8460) );
  OAI211_X1 U9886 ( .C1(n8591), .C2(n8504), .A(n8461), .B(n8460), .ZN(P2_U3277) );
  NAND2_X1 U9887 ( .A1(n8482), .A2(n8462), .ZN(n8463) );
  XOR2_X1 U9888 ( .A(n8472), .B(n8463), .Z(n8596) );
  INV_X1 U9889 ( .A(n8464), .ZN(n8465) );
  AOI21_X1 U9890 ( .B1(n8592), .B2(n8489), .A(n8465), .ZN(n8593) );
  AOI22_X1 U9891 ( .A1(n8467), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8466), .B2(
        n9751), .ZN(n8468) );
  OAI21_X1 U9892 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8480) );
  INV_X1 U9893 ( .A(n8471), .ZN(n8475) );
  INV_X1 U9894 ( .A(n8472), .ZN(n8474) );
  OAI21_X1 U9895 ( .B1(n8475), .B2(n8474), .A(n8473), .ZN(n8478) );
  AOI222_X1 U9896 ( .A1(n8511), .A2(n8478), .B1(n8477), .B2(n8506), .C1(n8476), 
        .C2(n8508), .ZN(n8595) );
  NOR2_X1 U9897 ( .A1(n8595), .A2(n8467), .ZN(n8479) );
  AOI211_X1 U9898 ( .C1(n8593), .C2(n8521), .A(n8480), .B(n8479), .ZN(n8481)
         );
  OAI21_X1 U9899 ( .B1(n8596), .B2(n8504), .A(n8481), .ZN(P2_U3278) );
  INV_X1 U9900 ( .A(n8482), .ZN(n8483) );
  AOI21_X1 U9901 ( .B1(n8492), .B2(n8484), .A(n8483), .ZN(n8601) );
  OAI22_X1 U9902 ( .A1(n9763), .A2(n8487), .B1(n8486), .B2(n8485), .ZN(n8502)
         );
  INV_X1 U9903 ( .A(n8488), .ZN(n8491) );
  INV_X1 U9904 ( .A(n8489), .ZN(n8490) );
  AOI211_X1 U9905 ( .C1(n8599), .C2(n8491), .A(n9881), .B(n8490), .ZN(n8598)
         );
  XNOR2_X1 U9906 ( .A(n8493), .B(n8492), .ZN(n8494) );
  OAI222_X1 U9907 ( .A1(n8498), .A2(n8497), .B1(n8496), .B2(n8495), .C1(n9759), 
        .C2(n8494), .ZN(n8597) );
  AOI21_X1 U9908 ( .B1(n8598), .B2(n8499), .A(n8597), .ZN(n8500) );
  NOR2_X1 U9909 ( .A1(n8500), .A2(n8467), .ZN(n8501) );
  AOI211_X1 U9910 ( .C1(n8514), .C2(n8599), .A(n8502), .B(n8501), .ZN(n8503)
         );
  OAI21_X1 U9911 ( .B1(n8601), .B2(n8504), .A(n8503), .ZN(P2_U3279) );
  XNOR2_X1 U9912 ( .A(n8505), .B(n8516), .ZN(n8510) );
  AOI222_X1 U9913 ( .A1(n8511), .A2(n8510), .B1(n8509), .B2(n8508), .C1(n8507), 
        .C2(n8506), .ZN(n9842) );
  MUX2_X1 U9914 ( .A(n8512), .B(n9842), .S(n9763), .Z(n8525) );
  AOI22_X1 U9915 ( .A1(n8514), .A2(n9835), .B1(n9751), .B2(n8513), .ZN(n8524)
         );
  NAND2_X1 U9916 ( .A1(n8517), .A2(n8516), .ZN(n9839) );
  NAND3_X1 U9917 ( .A1(n8515), .A2(n9839), .A3(n8518), .ZN(n8523) );
  AOI21_X1 U9918 ( .B1(n9835), .B2(n8520), .A(n8519), .ZN(n9838) );
  NAND2_X1 U9919 ( .A1(n9838), .A2(n8521), .ZN(n8522) );
  NAND4_X1 U9920 ( .A1(n8525), .A2(n8524), .A3(n8523), .A4(n8522), .ZN(
        P2_U3290) );
  NAND2_X1 U9921 ( .A1(n8526), .A2(n9837), .ZN(n8527) );
  OAI211_X1 U9922 ( .C1(n8292), .C2(n9879), .A(n8527), .B(n8530), .ZN(n8617)
         );
  MUX2_X1 U9923 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8617), .S(n9906), .Z(
        P2_U3551) );
  NAND2_X1 U9924 ( .A1(n8528), .A2(n9836), .ZN(n8529) );
  OAI211_X1 U9925 ( .C1(n8531), .C2(n9881), .A(n8530), .B(n8529), .ZN(n8618)
         );
  MUX2_X1 U9926 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8618), .S(n9906), .Z(
        P2_U3550) );
  MUX2_X1 U9927 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8619), .S(n9906), .Z(
        P2_U3549) );
  INV_X1 U9928 ( .A(n8536), .ZN(n8541) );
  AOI22_X1 U9929 ( .A1(n8538), .A2(n9837), .B1(n9836), .B2(n8537), .ZN(n8539)
         );
  OAI211_X1 U9930 ( .C1(n8541), .C2(n9871), .A(n8540), .B(n8539), .ZN(n8620)
         );
  MUX2_X1 U9931 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8620), .S(n9906), .Z(
        P2_U3548) );
  INV_X1 U9932 ( .A(n8542), .ZN(n8547) );
  AOI22_X1 U9933 ( .A1(n8544), .A2(n9837), .B1(n9836), .B2(n8543), .ZN(n8545)
         );
  OAI211_X1 U9934 ( .C1(n8547), .C2(n9871), .A(n8546), .B(n8545), .ZN(n8621)
         );
  MUX2_X1 U9935 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8621), .S(n9906), .Z(
        P2_U3547) );
  AOI21_X1 U9936 ( .B1(n9836), .B2(n8549), .A(n8548), .ZN(n8550) );
  OAI211_X1 U9937 ( .C1(n8552), .C2(n9871), .A(n8551), .B(n8550), .ZN(n8622)
         );
  MUX2_X1 U9938 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8622), .S(n9906), .Z(
        P2_U3546) );
  AOI21_X1 U9939 ( .B1(n9836), .B2(n8554), .A(n8553), .ZN(n8555) );
  OAI211_X1 U9940 ( .C1(n8557), .C2(n9871), .A(n8556), .B(n8555), .ZN(n8623)
         );
  MUX2_X1 U9941 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8623), .S(n9906), .Z(
        P2_U3545) );
  AOI22_X1 U9942 ( .A1(n8559), .A2(n9837), .B1(n9836), .B2(n8558), .ZN(n8560)
         );
  OAI211_X1 U9943 ( .C1(n8562), .C2(n9871), .A(n8561), .B(n8560), .ZN(n8624)
         );
  MUX2_X1 U9944 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8624), .S(n9906), .Z(
        P2_U3544) );
  OAI22_X1 U9945 ( .A1(n8564), .A2(n9881), .B1(n8563), .B2(n9879), .ZN(n8565)
         );
  OR2_X1 U9946 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  AOI21_X1 U9947 ( .B1(n8568), .B2(n9885), .A(n8567), .ZN(n8625) );
  MUX2_X1 U9948 ( .A(n8569), .B(n8625), .S(n9906), .Z(n8570) );
  INV_X1 U9949 ( .A(n8570), .ZN(P2_U3543) );
  AOI22_X1 U9950 ( .A1(n8572), .A2(n9837), .B1(n9836), .B2(n8571), .ZN(n8573)
         );
  OAI211_X1 U9951 ( .C1(n8575), .C2(n9871), .A(n8574), .B(n8573), .ZN(n8628)
         );
  MUX2_X1 U9952 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8628), .S(n9906), .Z(
        P2_U3542) );
  AOI22_X1 U9953 ( .A1(n8577), .A2(n9837), .B1(n9836), .B2(n8576), .ZN(n8578)
         );
  OAI211_X1 U9954 ( .C1(n8580), .C2(n9871), .A(n8579), .B(n8578), .ZN(n8629)
         );
  MUX2_X1 U9955 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8629), .S(n9906), .Z(
        P2_U3541) );
  NAND3_X1 U9956 ( .A1(n8436), .A2(n9885), .A3(n8581), .ZN(n8586) );
  AOI22_X1 U9957 ( .A1(n8583), .A2(n9837), .B1(n9836), .B2(n8582), .ZN(n8584)
         );
  NAND3_X1 U9958 ( .A1(n8586), .A2(n8585), .A3(n8584), .ZN(n8630) );
  MUX2_X1 U9959 ( .A(n8630), .B(P2_REG1_REG_20__SCAN_IN), .S(n9904), .Z(
        P2_U3540) );
  AOI21_X1 U9960 ( .B1(n9836), .B2(n8588), .A(n8587), .ZN(n8589) );
  OAI211_X1 U9961 ( .C1(n8591), .C2(n9871), .A(n8590), .B(n8589), .ZN(n8631)
         );
  MUX2_X1 U9962 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8631), .S(n9906), .Z(
        P2_U3539) );
  AOI22_X1 U9963 ( .A1(n8593), .A2(n9837), .B1(n9836), .B2(n8592), .ZN(n8594)
         );
  OAI211_X1 U9964 ( .C1(n8596), .C2(n9871), .A(n8595), .B(n8594), .ZN(n8632)
         );
  MUX2_X1 U9965 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8632), .S(n9906), .Z(
        P2_U3538) );
  AOI211_X1 U9966 ( .C1(n9836), .C2(n8599), .A(n8598), .B(n8597), .ZN(n8600)
         );
  OAI21_X1 U9967 ( .B1(n8601), .B2(n9871), .A(n8600), .ZN(n8633) );
  MUX2_X1 U9968 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8633), .S(n9906), .Z(
        P2_U3537) );
  AOI22_X1 U9969 ( .A1(n8603), .A2(n9837), .B1(n9836), .B2(n8602), .ZN(n8604)
         );
  OAI211_X1 U9970 ( .C1(n9849), .C2(n8606), .A(n8605), .B(n8604), .ZN(n8634)
         );
  MUX2_X1 U9971 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8634), .S(n9906), .Z(
        P2_U3536) );
  AOI22_X1 U9972 ( .A1(n8608), .A2(n9837), .B1(n9836), .B2(n8607), .ZN(n8609)
         );
  OAI211_X1 U9973 ( .C1(n8611), .C2(n9871), .A(n8610), .B(n8609), .ZN(n8635)
         );
  MUX2_X1 U9974 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8635), .S(n9906), .Z(
        P2_U3535) );
  AOI22_X1 U9975 ( .A1(n8613), .A2(n9837), .B1(n9836), .B2(n8612), .ZN(n8614)
         );
  OAI211_X1 U9976 ( .C1(n8616), .C2(n9871), .A(n8615), .B(n8614), .ZN(n8636)
         );
  MUX2_X1 U9977 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8636), .S(n9906), .Z(
        P2_U3534) );
  MUX2_X1 U9978 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8617), .S(n9888), .Z(
        P2_U3519) );
  MUX2_X1 U9979 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8618), .S(n9888), .Z(
        P2_U3518) );
  MUX2_X1 U9980 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8620), .S(n9888), .Z(
        P2_U3516) );
  MUX2_X1 U9981 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8621), .S(n9888), .Z(
        P2_U3515) );
  MUX2_X1 U9982 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8622), .S(n9888), .Z(
        P2_U3514) );
  MUX2_X1 U9983 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8623), .S(n9888), .Z(
        P2_U3513) );
  MUX2_X1 U9984 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8624), .S(n9888), .Z(
        P2_U3512) );
  INV_X1 U9985 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8626) );
  MUX2_X1 U9986 ( .A(n8626), .B(n8625), .S(n9888), .Z(n8627) );
  INV_X1 U9987 ( .A(n8627), .ZN(P2_U3511) );
  MUX2_X1 U9988 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8628), .S(n9888), .Z(
        P2_U3510) );
  MUX2_X1 U9989 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8629), .S(n9888), .Z(
        P2_U3509) );
  MUX2_X1 U9990 ( .A(n8630), .B(P2_REG0_REG_20__SCAN_IN), .S(n9887), .Z(
        P2_U3508) );
  MUX2_X1 U9991 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8631), .S(n9888), .Z(
        P2_U3507) );
  MUX2_X1 U9992 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8632), .S(n9888), .Z(
        P2_U3505) );
  MUX2_X1 U9993 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8633), .S(n9888), .Z(
        P2_U3502) );
  MUX2_X1 U9994 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8634), .S(n9888), .Z(
        P2_U3499) );
  MUX2_X1 U9995 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8635), .S(n9888), .Z(
        P2_U3496) );
  MUX2_X1 U9996 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8636), .S(n9888), .Z(
        P2_U3493) );
  INV_X1 U9997 ( .A(n8732), .ZN(n9422) );
  NOR4_X1 U9998 ( .A1(n4786), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5838), .A4(
        P2_U3152), .ZN(n8637) );
  AOI21_X1 U9999 ( .B1(n8644), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8637), .ZN(
        n8638) );
  OAI21_X1 U10000 ( .B1(n9422), .B2(n8647), .A(n8638), .ZN(P2_U3327) );
  INV_X1 U10001 ( .A(n8737), .ZN(n9425) );
  AOI22_X1 U10002 ( .A1(n5767), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8644), .ZN(n8639) );
  OAI21_X1 U10003 ( .B1(n9425), .B2(n8647), .A(n8639), .ZN(P2_U3328) );
  INV_X1 U10004 ( .A(n8640), .ZN(n9428) );
  OAI222_X1 U10005 ( .A1(n8647), .A2(n9428), .B1(P2_U3152), .B2(n8642), .C1(
        n9947), .C2(n8641), .ZN(P2_U3329) );
  INV_X1 U10006 ( .A(n8643), .ZN(n9432) );
  NAND2_X1 U10007 ( .A1(n8644), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8645) );
  OAI211_X1 U10008 ( .C1(n9432), .C2(n8647), .A(n8646), .B(n8645), .ZN(
        P2_U3330) );
  MUX2_X1 U10009 ( .A(n8648), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10010 ( .A(n8682), .ZN(n8650) );
  NOR2_X1 U10011 ( .A1(n8649), .A2(n8650), .ZN(n8654) );
  AOI21_X1 U10012 ( .B1(n8652), .B2(n8682), .A(n8651), .ZN(n8653) );
  OAI21_X1 U10013 ( .B1(n8654), .B2(n8653), .A(n8683), .ZN(n8658) );
  AOI22_X1 U10014 ( .A1(n8721), .A2(n9202), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8655) );
  OAI21_X1 U10015 ( .B1(n8676), .B2(n8723), .A(n8655), .ZN(n8656) );
  AOI21_X1 U10016 ( .B1(n9226), .B2(n8726), .A(n8656), .ZN(n8657) );
  OAI211_X1 U10017 ( .C1(n9228), .C2(n8730), .A(n8658), .B(n8657), .ZN(
        P1_U3214) );
  XOR2_X1 U10018 ( .A(n8661), .B(n8660), .Z(n8662) );
  XNOR2_X1 U10019 ( .A(n8663), .B(n8662), .ZN(n8669) );
  NAND2_X1 U10020 ( .A1(n8664), .A2(n9300), .ZN(n8665) );
  NAND2_X1 U10021 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9134) );
  OAI211_X1 U10022 ( .C1(n8674), .C2(n8706), .A(n8665), .B(n9134), .ZN(n8667)
         );
  NOR2_X1 U10023 ( .A1(n9293), .A2(n8730), .ZN(n8666) );
  AOI211_X1 U10024 ( .C1(n9291), .C2(n8726), .A(n8667), .B(n8666), .ZN(n8668)
         );
  OAI21_X1 U10025 ( .B1(n8669), .B2(n8716), .A(n8668), .ZN(P1_U3217) );
  INV_X1 U10026 ( .A(n9264), .ZN(n9370) );
  OAI21_X1 U10027 ( .B1(n8672), .B2(n8671), .A(n8670), .ZN(n8673) );
  NAND2_X1 U10028 ( .A1(n8673), .A2(n8683), .ZN(n8680) );
  NOR2_X1 U10029 ( .A1(n8723), .A2(n8674), .ZN(n8678) );
  OAI22_X1 U10030 ( .A1(n8706), .A2(n8676), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8675), .ZN(n8677) );
  AOI211_X1 U10031 ( .C1(n9267), .C2(n8726), .A(n8678), .B(n8677), .ZN(n8679)
         );
  OAI211_X1 U10032 ( .C1(n9370), .C2(n8730), .A(n8680), .B(n8679), .ZN(
        P1_U3221) );
  AND3_X1 U10033 ( .A1(n8649), .A2(n8682), .A3(n8681), .ZN(n8684) );
  OAI21_X1 U10034 ( .B1(n8685), .B2(n8684), .A(n8683), .ZN(n8689) );
  AOI22_X1 U10035 ( .A1(n8721), .A2(n9189), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8686) );
  OAI21_X1 U10036 ( .B1(n8705), .B2(n8723), .A(n8686), .ZN(n8687) );
  AOI21_X1 U10037 ( .B1(n9211), .B2(n8726), .A(n8687), .ZN(n8688) );
  OAI211_X1 U10038 ( .C1(n9213), .C2(n8730), .A(n8689), .B(n8688), .ZN(
        P1_U3227) );
  AOI21_X1 U10039 ( .B1(n8691), .B2(n8690), .A(n4347), .ZN(n8698) );
  NOR2_X1 U10040 ( .A1(n8723), .A2(n8692), .ZN(n8695) );
  OAI22_X1 U10041 ( .A1(n8706), .A2(n8703), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8693), .ZN(n8694) );
  AOI211_X1 U10042 ( .C1(n9274), .C2(n8726), .A(n8695), .B(n8694), .ZN(n8697)
         );
  NAND2_X1 U10043 ( .A1(n9375), .A2(n8709), .ZN(n8696) );
  OAI211_X1 U10044 ( .C1(n8698), .C2(n8716), .A(n8697), .B(n8696), .ZN(
        P1_U3231) );
  NAND2_X1 U10045 ( .A1(n8700), .A2(n8699), .ZN(n8702) );
  XNOR2_X1 U10046 ( .A(n8702), .B(n8701), .ZN(n8712) );
  NOR2_X1 U10047 ( .A1(n8723), .A2(n8703), .ZN(n8708) );
  INV_X1 U10048 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8704) );
  OAI22_X1 U10049 ( .A1(n8706), .A2(n8705), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8704), .ZN(n8707) );
  AOI211_X1 U10050 ( .C1(n9249), .C2(n8726), .A(n8708), .B(n8707), .ZN(n8711)
         );
  NAND2_X1 U10051 ( .A1(n9364), .A2(n8709), .ZN(n8710) );
  OAI211_X1 U10052 ( .C1(n8712), .C2(n8716), .A(n8711), .B(n8710), .ZN(
        P1_U3233) );
  INV_X1 U10053 ( .A(n8715), .ZN(n8720) );
  AOI21_X1 U10054 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8717) );
  NOR2_X1 U10055 ( .A1(n8717), .A2(n8716), .ZN(n8718) );
  OAI21_X1 U10056 ( .B1(n8720), .B2(n8719), .A(n8718), .ZN(n8729) );
  NAND2_X1 U10057 ( .A1(n8721), .A2(n9279), .ZN(n8722) );
  NAND2_X1 U10058 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9119) );
  OAI211_X1 U10059 ( .C1(n8724), .C2(n8723), .A(n8722), .B(n9119), .ZN(n8725)
         );
  AOI21_X1 U10060 ( .B1(n8727), .B2(n8726), .A(n8725), .ZN(n8728) );
  OAI211_X1 U10061 ( .C1(n8731), .C2(n8730), .A(n8729), .B(n8728), .ZN(
        P1_U3236) );
  NAND2_X1 U10062 ( .A1(n8732), .A2(n8736), .ZN(n8735) );
  NAND2_X1 U10063 ( .A1(n8733), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U10064 ( .A1(n8735), .A2(n8734), .ZN(n8857) );
  NAND2_X1 U10065 ( .A1(n8857), .A2(n8856), .ZN(n8852) );
  NAND2_X1 U10066 ( .A1(n8737), .A2(n8736), .ZN(n8739) );
  NAND2_X1 U10067 ( .A1(n5399), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8738) );
  OR2_X1 U10068 ( .A1(n9485), .A2(n8100), .ZN(n8740) );
  NOR2_X1 U10069 ( .A1(n9029), .A2(n9465), .ZN(n8995) );
  OAI21_X1 U10070 ( .B1(n9343), .B2(n9186), .A(n10115), .ZN(n8741) );
  INV_X1 U10071 ( .A(n8859), .ZN(n8845) );
  MUX2_X1 U10072 ( .A(n9343), .B(n8741), .S(n8845), .Z(n8840) );
  NAND2_X1 U10073 ( .A1(n4351), .A2(n9186), .ZN(n8746) );
  INV_X1 U10074 ( .A(n8976), .ZN(n8742) );
  NAND2_X1 U10075 ( .A1(n8743), .A2(n8742), .ZN(n8744) );
  AND2_X1 U10076 ( .A1(n8744), .A2(n8978), .ZN(n8745) );
  NAND2_X1 U10077 ( .A1(n8745), .A2(n8835), .ZN(n9018) );
  MUX2_X1 U10078 ( .A(n8746), .B(n9018), .S(n8845), .Z(n8837) );
  AND2_X1 U10079 ( .A1(n9297), .A2(n8747), .ZN(n8748) );
  MUX2_X1 U10080 ( .A(n8748), .B(n9294), .S(n8859), .Z(n8808) );
  MUX2_X1 U10081 ( .A(n8940), .B(n8920), .S(n8859), .Z(n8806) );
  INV_X1 U10082 ( .A(n8926), .ZN(n8761) );
  NAND3_X1 U10083 ( .A1(n6623), .A2(n9318), .A3(n9307), .ZN(n8750) );
  NAND2_X1 U10084 ( .A1(n8945), .A2(n8944), .ZN(n9007) );
  NAND2_X1 U10085 ( .A1(n9007), .A2(n8948), .ZN(n8749) );
  AOI21_X1 U10086 ( .B1(n8750), .B2(n8749), .A(n6680), .ZN(n8756) );
  NAND2_X1 U10087 ( .A1(n8955), .A2(n8949), .ZN(n8755) );
  NAND2_X1 U10088 ( .A1(n8751), .A2(n8763), .ZN(n8753) );
  NAND2_X1 U10089 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  OAI21_X1 U10090 ( .B1(n8756), .B2(n8755), .A(n8754), .ZN(n8759) );
  NAND2_X1 U10091 ( .A1(n8926), .A2(n8757), .ZN(n8758) );
  AOI21_X1 U10092 ( .B1(n8759), .B2(n8767), .A(n8758), .ZN(n8760) );
  MUX2_X1 U10093 ( .A(n8761), .B(n8760), .S(n8859), .Z(n8774) );
  INV_X1 U10094 ( .A(n8768), .ZN(n8771) );
  NAND3_X1 U10095 ( .A1(n9318), .A2(n8949), .A3(n8944), .ZN(n8765) );
  AND2_X1 U10096 ( .A1(n8763), .A2(n8762), .ZN(n8951) );
  NAND2_X1 U10097 ( .A1(n8948), .A2(n9307), .ZN(n8943) );
  NAND3_X1 U10098 ( .A1(n8943), .A2(n8949), .A3(n8945), .ZN(n8764) );
  OAI211_X1 U10099 ( .C1(n6623), .C2(n8765), .A(n8951), .B(n8764), .ZN(n8766)
         );
  NAND2_X1 U10100 ( .A1(n8766), .A2(n8955), .ZN(n8769) );
  NAND2_X1 U10101 ( .A1(n8768), .A2(n8767), .ZN(n8947) );
  AOI21_X1 U10102 ( .B1(n8769), .B2(n8927), .A(n8947), .ZN(n8770) );
  MUX2_X1 U10103 ( .A(n8771), .B(n8770), .S(n8845), .Z(n8772) );
  OR3_X1 U10104 ( .A1(n8774), .A2(n8773), .A3(n8772), .ZN(n8796) );
  AND2_X1 U10105 ( .A1(n8791), .A2(n7284), .ZN(n8957) );
  NAND2_X1 U10106 ( .A1(n8796), .A2(n8957), .ZN(n8777) );
  NAND2_X1 U10107 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  NAND4_X1 U10108 ( .A1(n8778), .A2(n8845), .A3(n8923), .A4(n8959), .ZN(n8800)
         );
  NAND2_X1 U10109 ( .A1(n8779), .A2(n8859), .ZN(n8784) );
  INV_X1 U10110 ( .A(n8784), .ZN(n8780) );
  AOI22_X1 U10111 ( .A1(n9400), .A2(n8780), .B1(n8783), .B2(n8859), .ZN(n8789)
         );
  NAND2_X1 U10112 ( .A1(n9057), .A2(n8845), .ZN(n8782) );
  OAI22_X1 U10113 ( .A1(n9400), .A2(n8782), .B1(n8783), .B2(n8859), .ZN(n8781)
         );
  NAND2_X1 U10114 ( .A1(n9493), .A2(n8781), .ZN(n8788) );
  NOR2_X1 U10115 ( .A1(n8783), .A2(n8782), .ZN(n8786) );
  OAI21_X1 U10116 ( .B1(n9056), .B2(n8784), .A(n9400), .ZN(n8785) );
  OAI21_X1 U10117 ( .B1(n8786), .B2(n9400), .A(n8785), .ZN(n8787) );
  OAI211_X1 U10118 ( .C1(n9493), .C2(n8789), .A(n8788), .B(n8787), .ZN(n8790)
         );
  INV_X1 U10119 ( .A(n8790), .ZN(n8799) );
  INV_X1 U10120 ( .A(n8791), .ZN(n8795) );
  OR2_X1 U10121 ( .A1(n8792), .A2(n8795), .ZN(n8793) );
  AND2_X1 U10122 ( .A1(n8934), .A2(n8793), .ZN(n8925) );
  AND2_X1 U10123 ( .A1(n8933), .A2(n8859), .ZN(n8794) );
  OAI211_X1 U10124 ( .C1(n8796), .C2(n8795), .A(n8925), .B(n8794), .ZN(n8797)
         );
  NAND4_X1 U10125 ( .A1(n8800), .A2(n8799), .A3(n8798), .A4(n8797), .ZN(n8804)
         );
  INV_X1 U10126 ( .A(n8924), .ZN(n8801) );
  MUX2_X1 U10127 ( .A(n8938), .B(n8801), .S(n8845), .Z(n8802) );
  NOR2_X1 U10128 ( .A1(n8893), .A2(n8802), .ZN(n8803) );
  NAND2_X1 U10129 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  NAND3_X1 U10130 ( .A1(n8895), .A2(n8806), .A3(n8805), .ZN(n8807) );
  NAND2_X1 U10131 ( .A1(n8808), .A2(n8807), .ZN(n8814) );
  AND2_X1 U10132 ( .A1(n8815), .A2(n8809), .ZN(n8810) );
  NAND2_X1 U10133 ( .A1(n8814), .A2(n8810), .ZN(n8813) );
  INV_X1 U10134 ( .A(n8966), .ZN(n8811) );
  NOR2_X1 U10135 ( .A1(n8871), .A2(n8811), .ZN(n8812) );
  NAND2_X1 U10136 ( .A1(n8813), .A2(n8812), .ZN(n8818) );
  AND2_X1 U10137 ( .A1(n8966), .A2(n9297), .ZN(n8969) );
  NAND2_X1 U10138 ( .A1(n8814), .A2(n8969), .ZN(n8816) );
  AND2_X1 U10139 ( .A1(n8872), .A2(n8815), .ZN(n8970) );
  NAND2_X1 U10140 ( .A1(n8816), .A2(n8970), .ZN(n8817) );
  MUX2_X1 U10141 ( .A(n8818), .B(n8817), .S(n8859), .Z(n8824) );
  INV_X1 U10142 ( .A(n8824), .ZN(n8821) );
  NAND2_X1 U10143 ( .A1(n9240), .A2(n8871), .ZN(n8819) );
  AND2_X1 U10144 ( .A1(n8819), .A2(n8826), .ZN(n8820) );
  NAND2_X1 U10145 ( .A1(n8828), .A2(n8820), .ZN(n8975) );
  AOI21_X1 U10146 ( .B1(n8821), .B2(n9240), .A(n8975), .ZN(n8823) );
  INV_X1 U10147 ( .A(n8973), .ZN(n8822) );
  OAI21_X1 U10148 ( .B1(n8823), .B2(n8822), .A(n8976), .ZN(n8833) );
  NAND2_X1 U10149 ( .A1(n8824), .A2(n8872), .ZN(n8827) );
  NAND2_X1 U10150 ( .A1(n8973), .A2(n9240), .ZN(n8825) );
  AOI21_X1 U10151 ( .B1(n8827), .B2(n8826), .A(n8825), .ZN(n8831) );
  INV_X1 U10152 ( .A(n8828), .ZN(n8830) );
  OAI21_X1 U10153 ( .B1(n8831), .B2(n8830), .A(n8829), .ZN(n8832) );
  MUX2_X1 U10154 ( .A(n8833), .B(n8832), .S(n8845), .Z(n8834) );
  NOR2_X1 U10155 ( .A1(n8834), .A2(n9215), .ZN(n8836) );
  OAI22_X1 U10156 ( .A1(n8837), .A2(n8836), .B1(n8845), .B2(n8835), .ZN(n8838)
         );
  OAI21_X1 U10157 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8843) );
  AOI21_X1 U10158 ( .B1(n9343), .B2(n9186), .A(n8859), .ZN(n8841) );
  OAI21_X1 U10159 ( .B1(n10115), .B2(n8841), .A(n8840), .ZN(n8842) );
  NAND2_X1 U10160 ( .A1(n8843), .A2(n8842), .ZN(n8844) );
  NAND2_X1 U10161 ( .A1(n8844), .A2(n8901), .ZN(n8847) );
  MUX2_X1 U10162 ( .A(n8917), .B(n8984), .S(n8845), .Z(n8846) );
  NAND3_X1 U10163 ( .A1(n8847), .A2(n9158), .A3(n8846), .ZN(n8849) );
  MUX2_X1 U10164 ( .A(n8918), .B(n8987), .S(n8859), .Z(n8848) );
  NAND2_X1 U10165 ( .A1(n8849), .A2(n8848), .ZN(n8862) );
  NAND2_X1 U10166 ( .A1(n9485), .A2(n8100), .ZN(n9024) );
  NAND2_X1 U10167 ( .A1(n9485), .A2(n8856), .ZN(n8850) );
  NAND2_X1 U10168 ( .A1(n9024), .A2(n8850), .ZN(n8992) );
  NOR3_X1 U10169 ( .A1(n8862), .A2(n8992), .A3(n8860), .ZN(n8851) );
  NOR2_X1 U10170 ( .A1(n8995), .A2(n8851), .ZN(n8855) );
  NOR3_X1 U10171 ( .A1(n8995), .A2(n8861), .A3(n8862), .ZN(n8853) );
  OAI21_X1 U10172 ( .B1(n8853), .B2(n8992), .A(n8852), .ZN(n8854) );
  MUX2_X1 U10173 ( .A(n8855), .B(n8854), .S(n8859), .Z(n8867) );
  OR2_X1 U10174 ( .A1(n8857), .A2(n8856), .ZN(n9030) );
  INV_X1 U10175 ( .A(n8860), .ZN(n9160) );
  NOR2_X1 U10176 ( .A1(n8861), .A2(n8859), .ZN(n8858) );
  AOI211_X1 U10177 ( .C1(n9160), .C2(n8859), .A(n8858), .B(n8992), .ZN(n8865)
         );
  INV_X1 U10178 ( .A(n8995), .ZN(n8864) );
  NAND3_X1 U10179 ( .A1(n8862), .A2(n8861), .A3(n8860), .ZN(n8863) );
  NAND3_X1 U10180 ( .A1(n8865), .A2(n8864), .A3(n8863), .ZN(n8866) );
  NAND3_X1 U10181 ( .A1(n8867), .A2(n9030), .A3(n8866), .ZN(n8909) );
  INV_X1 U10182 ( .A(n8909), .ZN(n9050) );
  INV_X1 U10183 ( .A(n9030), .ZN(n8869) );
  OR4_X1 U10184 ( .A1(n8869), .A2(n6502), .A3(n8868), .A4(n9040), .ZN(n9049)
         );
  INV_X1 U10185 ( .A(n8870), .ZN(n8905) );
  XNOR2_X1 U10186 ( .A(n9343), .B(n9203), .ZN(n9188) );
  INV_X1 U10187 ( .A(n9188), .ZN(n8904) );
  INV_X1 U10188 ( .A(n9158), .ZN(n8903) );
  NAND2_X1 U10189 ( .A1(n4443), .A2(n8872), .ZN(n9278) );
  NAND4_X1 U10190 ( .A1(n8876), .A2(n8875), .A3(n6624), .A4(n8874), .ZN(n8879)
         );
  NAND2_X1 U10191 ( .A1(n9318), .A2(n8877), .ZN(n8878) );
  NOR2_X1 U10192 ( .A1(n8879), .A2(n8878), .ZN(n8882) );
  NAND4_X1 U10193 ( .A1(n8882), .A2(n8881), .A3(n6877), .A4(n9614), .ZN(n8884)
         );
  NOR2_X1 U10194 ( .A1(n8884), .A2(n8883), .ZN(n8886) );
  AND4_X1 U10195 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n8889)
         );
  NAND3_X1 U10196 ( .A1(n7328), .A2(n8890), .A3(n8889), .ZN(n8891) );
  NOR3_X1 U10197 ( .A1(n8893), .A2(n8892), .A3(n8891), .ZN(n8894) );
  NAND4_X1 U10198 ( .A1(n9285), .A2(n8896), .A3(n8895), .A4(n8894), .ZN(n8897)
         );
  NOR2_X1 U10199 ( .A1(n9278), .A2(n8897), .ZN(n8898) );
  NAND3_X1 U10200 ( .A1(n9244), .A2(n9259), .A3(n8898), .ZN(n8899) );
  NOR2_X1 U10201 ( .A1(n9231), .A2(n8899), .ZN(n8900) );
  NAND4_X1 U10202 ( .A1(n8901), .A2(n9200), .A3(n4813), .A4(n8900), .ZN(n8902)
         );
  NOR4_X1 U10203 ( .A1(n8905), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(n8906)
         );
  NAND3_X1 U10204 ( .A1(n8906), .A2(n9030), .A3(n9024), .ZN(n8908) );
  INV_X1 U10205 ( .A(n9029), .ZN(n8907) );
  OAI21_X1 U10206 ( .B1(n8908), .B2(n8907), .A(n4926), .ZN(n8911) );
  OAI21_X1 U10207 ( .B1(n8909), .B2(n5580), .A(n8911), .ZN(n8910) );
  NAND4_X1 U10208 ( .A1(n8910), .A2(n9032), .A3(n5398), .A4(n9034), .ZN(n9048)
         );
  INV_X1 U10209 ( .A(n8911), .ZN(n8913) );
  NOR4_X1 U10210 ( .A1(n8913), .A2(n5398), .A3(n8912), .A4(n9040), .ZN(n9046)
         );
  INV_X1 U10211 ( .A(n8914), .ZN(n8915) );
  NAND2_X1 U10212 ( .A1(n8984), .A2(n8915), .ZN(n8916) );
  NAND3_X1 U10213 ( .A1(n8918), .A2(n8917), .A3(n8916), .ZN(n8986) );
  INV_X1 U10214 ( .A(n8986), .ZN(n9022) );
  INV_X1 U10215 ( .A(n8919), .ZN(n9020) );
  NOR2_X1 U10216 ( .A1(n8921), .A2(n4432), .ZN(n8922) );
  NAND2_X1 U10217 ( .A1(n8922), .A2(n9297), .ZN(n8962) );
  NAND2_X1 U10218 ( .A1(n8924), .A2(n8923), .ZN(n8961) );
  INV_X1 U10219 ( .A(n8961), .ZN(n8937) );
  INV_X1 U10220 ( .A(n8925), .ZN(n8932) );
  INV_X1 U10221 ( .A(n8957), .ZN(n8930) );
  OAI21_X1 U10222 ( .B1(n8947), .B2(n8927), .A(n8926), .ZN(n8928) );
  INV_X1 U10223 ( .A(n8928), .ZN(n8929) );
  NOR2_X1 U10224 ( .A1(n8930), .A2(n8929), .ZN(n8931) );
  OAI21_X1 U10225 ( .B1(n8932), .B2(n8931), .A(n8959), .ZN(n8935) );
  NAND3_X1 U10226 ( .A1(n8935), .A2(n8934), .A3(n8933), .ZN(n8936) );
  NAND2_X1 U10227 ( .A1(n8937), .A2(n8936), .ZN(n8941) );
  INV_X1 U10228 ( .A(n8938), .ZN(n8939) );
  AND3_X1 U10229 ( .A1(n8941), .A2(n8940), .A3(n8939), .ZN(n8942) );
  OR2_X1 U10230 ( .A1(n8962), .A2(n8942), .ZN(n9012) );
  AOI21_X1 U10231 ( .B1(n8944), .B2(n9003), .A(n8943), .ZN(n8946) );
  INV_X1 U10232 ( .A(n8949), .ZN(n9008) );
  NOR3_X1 U10233 ( .A1(n8946), .A2(n9008), .A3(n6671), .ZN(n8965) );
  INV_X1 U10234 ( .A(n8951), .ZN(n8964) );
  INV_X1 U10235 ( .A(n8947), .ZN(n8958) );
  INV_X1 U10236 ( .A(n8948), .ZN(n8950) );
  NAND2_X1 U10237 ( .A1(n8950), .A2(n8949), .ZN(n8952) );
  NAND2_X1 U10238 ( .A1(n8952), .A2(n8951), .ZN(n9005) );
  NAND2_X1 U10239 ( .A1(n9307), .A2(n8953), .ZN(n8954) );
  NOR2_X1 U10240 ( .A1(n9005), .A2(n8954), .ZN(n8997) );
  AOI21_X1 U10241 ( .B1(n6621), .B2(n8997), .A(n4428), .ZN(n8956) );
  NAND4_X1 U10242 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8960)
         );
  OR3_X1 U10243 ( .A1(n8962), .A2(n8961), .A3(n8960), .ZN(n9014) );
  INV_X1 U10244 ( .A(n9014), .ZN(n8963) );
  OAI21_X1 U10245 ( .B1(n8965), .B2(n8964), .A(n8963), .ZN(n8968) );
  INV_X1 U10246 ( .A(n8975), .ZN(n8967) );
  NAND2_X1 U10247 ( .A1(n8967), .A2(n8966), .ZN(n8996) );
  AOI21_X1 U10248 ( .B1(n9012), .B2(n8968), .A(n8996), .ZN(n8977) );
  INV_X1 U10249 ( .A(n8969), .ZN(n8971) );
  OAI211_X1 U10250 ( .C1(n9294), .C2(n8971), .A(n9240), .B(n8970), .ZN(n8972)
         );
  INV_X1 U10251 ( .A(n8972), .ZN(n8974) );
  OAI21_X1 U10252 ( .B1(n8975), .B2(n8974), .A(n8973), .ZN(n9015) );
  OAI21_X1 U10253 ( .B1(n8977), .B2(n9015), .A(n8976), .ZN(n8981) );
  INV_X1 U10254 ( .A(n8978), .ZN(n8980) );
  AOI211_X1 U10255 ( .C1(n9020), .C2(n8981), .A(n8980), .B(n8979), .ZN(n8991)
         );
  INV_X1 U10256 ( .A(n8982), .ZN(n8983) );
  AND2_X1 U10257 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  NOR2_X1 U10258 ( .A1(n8986), .A2(n8985), .ZN(n8990) );
  INV_X1 U10259 ( .A(n8987), .ZN(n8988) );
  OR3_X1 U10260 ( .A1(n8990), .A2(n8989), .A3(n8988), .ZN(n9027) );
  AOI21_X1 U10261 ( .B1(n9022), .B2(n8991), .A(n9027), .ZN(n8993) );
  NOR3_X1 U10262 ( .A1(n8993), .A2(n9023), .A3(n8992), .ZN(n8994) );
  OAI211_X1 U10263 ( .C1(n8995), .C2(n8994), .A(n8999), .B(n9030), .ZN(n9045)
         );
  INV_X1 U10264 ( .A(n8996), .ZN(n9017) );
  INV_X1 U10265 ( .A(n8997), .ZN(n9011) );
  INV_X1 U10266 ( .A(n8998), .ZN(n9002) );
  NAND2_X1 U10267 ( .A1(n6489), .A2(n6487), .ZN(n9001) );
  NAND2_X1 U10268 ( .A1(n9632), .A2(n6492), .ZN(n9000) );
  NAND4_X1 U10269 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n9004)
         );
  AND2_X1 U10270 ( .A1(n9004), .A2(n9003), .ZN(n9010) );
  INV_X1 U10271 ( .A(n9005), .ZN(n9006) );
  OAI21_X1 U10272 ( .B1(n9008), .B2(n9007), .A(n9006), .ZN(n9009) );
  OAI21_X1 U10273 ( .B1(n9011), .B2(n9010), .A(n9009), .ZN(n9013) );
  OAI21_X1 U10274 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9016) );
  AOI21_X1 U10275 ( .B1(n9017), .B2(n9016), .A(n9015), .ZN(n9019) );
  AOI21_X1 U10276 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n9021) );
  AND2_X1 U10277 ( .A1(n9022), .A2(n9021), .ZN(n9026) );
  INV_X1 U10278 ( .A(n9023), .ZN(n9025) );
  OAI211_X1 U10279 ( .C1(n9027), .C2(n9026), .A(n9025), .B(n9024), .ZN(n9028)
         );
  NAND2_X1 U10280 ( .A1(n9029), .A2(n9028), .ZN(n9031) );
  NAND2_X1 U10281 ( .A1(n9031), .A2(n9030), .ZN(n9035) );
  OR4_X1 U10282 ( .A1(n9035), .A2(n9032), .A3(n5579), .A4(n9040), .ZN(n9043)
         );
  NAND3_X1 U10283 ( .A1(n9035), .A2(n9034), .A3(n9033), .ZN(n9042) );
  NAND4_X1 U10284 ( .A1(n9038), .A2(n9037), .A3(n9512), .A4(n9036), .ZN(n9039)
         );
  OAI211_X1 U10285 ( .C1(n6502), .C2(n9040), .A(n9039), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9041) );
  NAND3_X1 U10286 ( .A1(n9043), .A2(n9042), .A3(n9041), .ZN(n9044) );
  AOI21_X1 U10287 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9047) );
  OAI211_X1 U10288 ( .C1(n9050), .C2(n9049), .A(n9048), .B(n9047), .ZN(
        P1_U3240) );
  MUX2_X1 U10289 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9051), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10290 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9160), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10291 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9052), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10292 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9190), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10293 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9189), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10294 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9202), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10295 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9246), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10296 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9260), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10297 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9301), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10298 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9279), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10299 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9300), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10300 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9053), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10301 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9054), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10302 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9055), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10303 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9056), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10304 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9057), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10305 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9058), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10306 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9059), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10307 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9060), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10308 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9061), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10309 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9062), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10310 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9063), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10311 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9311), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10312 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9064), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10313 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9310), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10314 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9065), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10315 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9632), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10316 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6489), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10317 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6488), .S(P1_U4006), .Z(
        P1_U3555) );
  NAND2_X1 U10318 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n9066) );
  OAI21_X1 U10319 ( .B1(n9587), .B2(n9067), .A(n9066), .ZN(n9068) );
  AOI21_X1 U10320 ( .B1(n9589), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n9068), .ZN(
        n9079) );
  INV_X1 U10321 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9069) );
  NOR2_X1 U10322 ( .A1(n9515), .A2(n9069), .ZN(n9522) );
  OAI211_X1 U10323 ( .C1(n9071), .C2(n9522), .A(n9598), .B(n9070), .ZN(n9078)
         );
  INV_X1 U10324 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9073) );
  MUX2_X1 U10325 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9073), .S(n9072), .Z(n9075)
         );
  OAI211_X1 U10326 ( .C1(n9076), .C2(n9075), .A(n9593), .B(n9074), .ZN(n9077)
         );
  NAND3_X1 U10327 ( .A1(n9079), .A2(n9078), .A3(n9077), .ZN(P1_U3242) );
  OAI21_X1 U10328 ( .B1(n9587), .B2(n9081), .A(n9080), .ZN(n9082) );
  AOI21_X1 U10329 ( .B1(n9589), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9082), .ZN(
        n9094) );
  MUX2_X1 U10330 ( .A(n6151), .B(P1_REG2_REG_3__SCAN_IN), .S(n9083), .Z(n9086)
         );
  INV_X1 U10331 ( .A(n9084), .ZN(n9085) );
  NAND2_X1 U10332 ( .A1(n9086), .A2(n9085), .ZN(n9088) );
  OAI211_X1 U10333 ( .C1(n9534), .C2(n9088), .A(n9598), .B(n9087), .ZN(n9093)
         );
  OAI211_X1 U10334 ( .C1(n9091), .C2(n9090), .A(n9593), .B(n9089), .ZN(n9092)
         );
  NAND3_X1 U10335 ( .A1(n9094), .A2(n9093), .A3(n9092), .ZN(P1_U3244) );
  AOI21_X1 U10336 ( .B1(n9100), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9095), .ZN(
        n9098) );
  NAND2_X1 U10337 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9113), .ZN(n9096) );
  OAI21_X1 U10338 ( .B1(n9113), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9096), .ZN(
        n9097) );
  NOR2_X1 U10339 ( .A1(n9098), .A2(n9097), .ZN(n9112) );
  AOI211_X1 U10340 ( .C1(n9098), .C2(n9097), .A(n9112), .B(n9553), .ZN(n9108)
         );
  XNOR2_X1 U10341 ( .A(n9113), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9101) );
  NOR2_X1 U10342 ( .A1(n9102), .A2(n9101), .ZN(n9109) );
  AOI211_X1 U10343 ( .C1(n9102), .C2(n9101), .A(n9109), .B(n9573), .ZN(n9107)
         );
  INV_X1 U10344 ( .A(n9113), .ZN(n9105) );
  NAND2_X1 U10345 ( .A1(n9589), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9104) );
  OAI211_X1 U10346 ( .C1(n9587), .C2(n9105), .A(n9104), .B(n9103), .ZN(n9106)
         );
  OR3_X1 U10347 ( .A1(n9108), .A2(n9107), .A3(n9106), .ZN(P1_U3258) );
  INV_X1 U10348 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9123) );
  XOR2_X1 U10349 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9126), .Z(n9111) );
  AOI21_X1 U10350 ( .B1(n9113), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9109), .ZN(
        n9110) );
  NAND2_X1 U10351 ( .A1(n9111), .A2(n9110), .ZN(n9125) );
  OAI21_X1 U10352 ( .B1(n9111), .B2(n9110), .A(n9125), .ZN(n9118) );
  NAND2_X1 U10353 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9126), .ZN(n9114) );
  OAI21_X1 U10354 ( .B1(n9126), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9114), .ZN(
        n9115) );
  AOI211_X1 U10355 ( .C1(n9116), .C2(n9115), .A(n9124), .B(n9553), .ZN(n9117)
         );
  AOI21_X1 U10356 ( .B1(n9593), .B2(n9118), .A(n9117), .ZN(n9122) );
  INV_X1 U10357 ( .A(n9119), .ZN(n9120) );
  AOI21_X1 U10358 ( .B1(n9578), .B2(n9126), .A(n9120), .ZN(n9121) );
  OAI211_X1 U10359 ( .C1(n9584), .C2(n9123), .A(n9122), .B(n9121), .ZN(
        P1_U3259) );
  NAND2_X1 U10360 ( .A1(n9131), .A2(n9598), .ZN(n9129) );
  OAI21_X1 U10361 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9126), .A(n9125), .ZN(
        n9127) );
  XOR2_X1 U10362 ( .A(n9127), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9130) );
  AOI21_X1 U10363 ( .B1(n9130), .B2(n9593), .A(n9578), .ZN(n9128) );
  NAND2_X1 U10364 ( .A1(n9129), .A2(n9128), .ZN(n9133) );
  OAI22_X1 U10365 ( .A1(n9131), .A2(n9553), .B1(n9130), .B2(n9573), .ZN(n9132)
         );
  MUX2_X1 U10366 ( .A(n9133), .B(n9132), .S(n5579), .Z(n9137) );
  OAI21_X1 U10367 ( .B1(n9584), .B2(n9135), .A(n9134), .ZN(n9136) );
  XNOR2_X1 U10368 ( .A(n9465), .B(n9142), .ZN(n9467) );
  NAND2_X1 U10369 ( .A1(n9467), .A2(n9612), .ZN(n9141) );
  NAND2_X1 U10370 ( .A1(n9139), .A2(n9138), .ZN(n9481) );
  NOR2_X1 U10371 ( .A1(n9481), .A2(n9648), .ZN(n9146) );
  AOI21_X1 U10372 ( .B1(n9648), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9146), .ZN(
        n9140) );
  OAI211_X1 U10373 ( .C1(n9465), .C2(n9623), .A(n9141), .B(n9140), .ZN(
        P1_U3261) );
  OAI21_X1 U10374 ( .B1(n9144), .B2(n9143), .A(n9142), .ZN(n9482) );
  NOR2_X1 U10375 ( .A1(n9144), .A2(n9623), .ZN(n9145) );
  AOI211_X1 U10376 ( .C1(n9648), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9146), .B(
        n9145), .ZN(n9147) );
  OAI21_X1 U10377 ( .B1(n9148), .B2(n9482), .A(n9147), .ZN(P1_U3262) );
  AOI21_X1 U10378 ( .B1(n9158), .B2(n9150), .A(n9149), .ZN(n9151) );
  INV_X1 U10379 ( .A(n9151), .ZN(n9337) );
  INV_X1 U10380 ( .A(n9152), .ZN(n9153) );
  AOI21_X1 U10381 ( .B1(n9333), .B2(n9167), .A(n9153), .ZN(n9334) );
  INV_X1 U10382 ( .A(n9333), .ZN(n9156) );
  AOI22_X1 U10383 ( .A1(n9648), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9154), .B2(
        n9314), .ZN(n9155) );
  OAI21_X1 U10384 ( .B1(n9156), .B2(n9623), .A(n9155), .ZN(n9164) );
  OAI21_X1 U10385 ( .B1(n9158), .B2(n4352), .A(n9157), .ZN(n9159) );
  AOI211_X1 U10386 ( .C1(n9334), .C2(n9612), .A(n9164), .B(n9163), .ZN(n9165)
         );
  OAI21_X1 U10387 ( .B1(n9337), .B2(n9306), .A(n9165), .ZN(P1_U3263) );
  XNOR2_X1 U10388 ( .A(n9166), .B(n9176), .ZN(n9342) );
  INV_X1 U10389 ( .A(n9181), .ZN(n9169) );
  INV_X1 U10390 ( .A(n9167), .ZN(n9168) );
  AOI211_X1 U10391 ( .C1(n9339), .C2(n9169), .A(n9706), .B(n9168), .ZN(n9338)
         );
  AOI22_X1 U10392 ( .A1(n9648), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9170), .B2(
        n9314), .ZN(n9171) );
  OAI21_X1 U10393 ( .B1(n9172), .B2(n9623), .A(n9171), .ZN(n9178) );
  NOR2_X1 U10394 ( .A1(n9173), .A2(n9616), .ZN(n9177) );
  OAI21_X1 U10395 ( .B1(n9342), .B2(n9306), .A(n9179), .ZN(P1_U3264) );
  XNOR2_X1 U10396 ( .A(n9180), .B(n9188), .ZN(n9347) );
  INV_X1 U10397 ( .A(n9196), .ZN(n9182) );
  AOI21_X1 U10398 ( .B1(n9343), .B2(n9182), .A(n9181), .ZN(n9344) );
  AOI22_X1 U10399 ( .A1(n9648), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9183), .B2(
        n9314), .ZN(n9184) );
  OAI21_X1 U10400 ( .B1(n9185), .B2(n9623), .A(n9184), .ZN(n9193) );
  AOI222_X1 U10401 ( .A1(n9313), .A2(n9191), .B1(n9190), .B2(n9631), .C1(n9189), .C2(n9633), .ZN(n9346) );
  NOR2_X1 U10402 ( .A1(n9346), .A2(n9648), .ZN(n9192) );
  AOI211_X1 U10403 ( .C1(n9344), .C2(n9612), .A(n9193), .B(n9192), .ZN(n9194)
         );
  OAI21_X1 U10404 ( .B1(n9306), .B2(n9347), .A(n9194), .ZN(P1_U3265) );
  XOR2_X1 U10405 ( .A(n9200), .B(n9195), .Z(n9352) );
  AOI21_X1 U10406 ( .B1(n9348), .B2(n9209), .A(n9196), .ZN(n9349) );
  INV_X1 U10407 ( .A(n9348), .ZN(n9199) );
  AOI22_X1 U10408 ( .A1(n9648), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9197), .B2(
        n9314), .ZN(n9198) );
  OAI21_X1 U10409 ( .B1(n9199), .B2(n9623), .A(n9198), .ZN(n9206) );
  XNOR2_X1 U10410 ( .A(n9201), .B(n9200), .ZN(n9204) );
  AOI222_X1 U10411 ( .A1(n9313), .A2(n9204), .B1(n9203), .B2(n9631), .C1(n9202), .C2(n9633), .ZN(n9351) );
  NOR2_X1 U10412 ( .A1(n9351), .A2(n9648), .ZN(n9205) );
  AOI211_X1 U10413 ( .C1(n9349), .C2(n9612), .A(n9206), .B(n9205), .ZN(n9207)
         );
  OAI21_X1 U10414 ( .B1(n9352), .B2(n9306), .A(n9207), .ZN(P1_U3266) );
  XNOR2_X1 U10415 ( .A(n9208), .B(n9215), .ZN(n9357) );
  INV_X1 U10416 ( .A(n9209), .ZN(n9210) );
  AOI211_X1 U10417 ( .C1(n9354), .C2(n9223), .A(n9706), .B(n9210), .ZN(n9353)
         );
  AOI22_X1 U10418 ( .A1(n9648), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9211), .B2(
        n9314), .ZN(n9212) );
  OAI21_X1 U10419 ( .B1(n9213), .B2(n9623), .A(n9212), .ZN(n9220) );
  NOR2_X1 U10420 ( .A1(n9214), .A2(n9616), .ZN(n9218) );
  AOI211_X1 U10421 ( .C1(n9216), .C2(n9215), .A(n8091), .B(n4349), .ZN(n9217)
         );
  AOI211_X1 U10422 ( .C1(n9633), .C2(n9246), .A(n9218), .B(n9217), .ZN(n9356)
         );
  NOR2_X1 U10423 ( .A1(n9356), .A2(n9648), .ZN(n9219) );
  AOI211_X1 U10424 ( .C1(n9353), .C2(n9322), .A(n9220), .B(n9219), .ZN(n9221)
         );
  OAI21_X1 U10425 ( .B1(n9306), .B2(n9357), .A(n9221), .ZN(P1_U3267) );
  XNOR2_X1 U10426 ( .A(n9222), .B(n9231), .ZN(n9362) );
  INV_X1 U10427 ( .A(n9248), .ZN(n9225) );
  INV_X1 U10428 ( .A(n9223), .ZN(n9224) );
  AOI21_X1 U10429 ( .B1(n9358), .B2(n9225), .A(n9224), .ZN(n9359) );
  AOI22_X1 U10430 ( .A1(n9648), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9226), .B2(
        n9314), .ZN(n9227) );
  OAI21_X1 U10431 ( .B1(n9228), .B2(n9623), .A(n9227), .ZN(n9236) );
  NOR2_X1 U10432 ( .A1(n9229), .A2(n9616), .ZN(n9234) );
  AOI211_X1 U10433 ( .C1(n9232), .C2(n9231), .A(n8091), .B(n9230), .ZN(n9233)
         );
  AOI211_X1 U10434 ( .C1(n9633), .C2(n9260), .A(n9234), .B(n9233), .ZN(n9361)
         );
  NOR2_X1 U10435 ( .A1(n9361), .A2(n9648), .ZN(n9235) );
  AOI211_X1 U10436 ( .C1(n9359), .C2(n9612), .A(n9236), .B(n9235), .ZN(n9237)
         );
  OAI21_X1 U10437 ( .B1(n9306), .B2(n9362), .A(n9237), .ZN(P1_U3268) );
  XNOR2_X1 U10438 ( .A(n9238), .B(n9244), .ZN(n9367) );
  NOR2_X1 U10439 ( .A1(n9239), .A2(n9623), .ZN(n9252) );
  INV_X1 U10440 ( .A(n9257), .ZN(n9242) );
  INV_X1 U10441 ( .A(n9240), .ZN(n9241) );
  NOR2_X1 U10442 ( .A1(n9242), .A2(n9241), .ZN(n9245) );
  OAI21_X1 U10443 ( .B1(n9245), .B2(n9244), .A(n9243), .ZN(n9247) );
  AOI222_X1 U10444 ( .A1(n9313), .A2(n9247), .B1(n9280), .B2(n9633), .C1(n9246), .C2(n9631), .ZN(n9366) );
  AOI211_X1 U10445 ( .C1(n9364), .C2(n9265), .A(n9706), .B(n9248), .ZN(n9363)
         );
  AOI22_X1 U10446 ( .A1(n9363), .A2(n5579), .B1(n9314), .B2(n9249), .ZN(n9250)
         );
  AOI21_X1 U10447 ( .B1(n9366), .B2(n9250), .A(n9648), .ZN(n9251) );
  AOI211_X1 U10448 ( .C1(n9648), .C2(P1_REG2_REG_22__SCAN_IN), .A(n9252), .B(
        n9251), .ZN(n9253) );
  OAI21_X1 U10449 ( .B1(n9306), .B2(n9367), .A(n9253), .ZN(P1_U3269) );
  NOR2_X1 U10450 ( .A1(n4386), .A2(n9254), .ZN(n9255) );
  AOI22_X1 U10451 ( .A1(n9264), .A2(n9316), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9648), .ZN(n9271) );
  OAI211_X1 U10452 ( .C1(n9259), .C2(n9258), .A(n9257), .B(n9313), .ZN(n9262)
         );
  AOI22_X1 U10453 ( .A1(n9631), .A2(n9260), .B1(n9301), .B2(n9633), .ZN(n9261)
         );
  NAND2_X1 U10454 ( .A1(n9262), .A2(n9261), .ZN(n9372) );
  INV_X1 U10455 ( .A(n9263), .ZN(n9273) );
  AOI21_X1 U10456 ( .B1(n9273), .B2(n9264), .A(n9706), .ZN(n9266) );
  NAND2_X1 U10457 ( .A1(n9266), .A2(n9265), .ZN(n9369) );
  INV_X1 U10458 ( .A(n9267), .ZN(n9268) );
  OAI22_X1 U10459 ( .A1(n9369), .A2(n5398), .B1(n9268), .B2(n9641), .ZN(n9269)
         );
  OAI21_X1 U10460 ( .B1(n9372), .B2(n9269), .A(n9646), .ZN(n9270) );
  OAI211_X1 U10461 ( .C1(n9368), .C2(n9306), .A(n9271), .B(n9270), .ZN(
        P1_U3270) );
  XOR2_X1 U10462 ( .A(n9272), .B(n9278), .Z(n9379) );
  AOI21_X1 U10463 ( .B1(n9375), .B2(n9288), .A(n9263), .ZN(n9376) );
  INV_X1 U10464 ( .A(n9375), .ZN(n9276) );
  AOI22_X1 U10465 ( .A1(n9648), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9274), .B2(
        n9314), .ZN(n9275) );
  OAI21_X1 U10466 ( .B1(n9276), .B2(n9623), .A(n9275), .ZN(n9283) );
  XOR2_X1 U10467 ( .A(n9278), .B(n9277), .Z(n9281) );
  AOI222_X1 U10468 ( .A1(n9313), .A2(n9281), .B1(n9280), .B2(n9631), .C1(n9279), .C2(n9633), .ZN(n9378) );
  NOR2_X1 U10469 ( .A1(n9378), .A2(n9648), .ZN(n9282) );
  AOI211_X1 U10470 ( .C1(n9376), .C2(n9612), .A(n9283), .B(n9282), .ZN(n9284)
         );
  OAI21_X1 U10471 ( .B1(n9306), .B2(n9379), .A(n9284), .ZN(P1_U3271) );
  XOR2_X1 U10472 ( .A(n9286), .B(n9285), .Z(n9384) );
  INV_X1 U10473 ( .A(n9287), .ZN(n9290) );
  INV_X1 U10474 ( .A(n9288), .ZN(n9289) );
  AOI211_X1 U10475 ( .C1(n9381), .C2(n9290), .A(n9706), .B(n9289), .ZN(n9380)
         );
  AOI22_X1 U10476 ( .A1(n9648), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9291), .B2(
        n9314), .ZN(n9292) );
  OAI21_X1 U10477 ( .B1(n9293), .B2(n9623), .A(n9292), .ZN(n9304) );
  NAND2_X1 U10478 ( .A1(n9295), .A2(n9294), .ZN(n9298) );
  NAND3_X1 U10479 ( .A1(n9298), .A2(n9297), .A3(n9296), .ZN(n9299) );
  NAND2_X1 U10480 ( .A1(n4387), .A2(n9299), .ZN(n9302) );
  AOI222_X1 U10481 ( .A1(n9313), .A2(n9302), .B1(n9301), .B2(n9631), .C1(n9300), .C2(n9633), .ZN(n9383) );
  NOR2_X1 U10482 ( .A1(n9383), .A2(n9648), .ZN(n9303) );
  AOI211_X1 U10483 ( .C1(n9380), .C2(n9322), .A(n9304), .B(n9303), .ZN(n9305)
         );
  OAI21_X1 U10484 ( .B1(n9306), .B2(n9384), .A(n9305), .ZN(P1_U3272) );
  NAND2_X1 U10485 ( .A1(n9308), .A2(n9307), .ZN(n9309) );
  XOR2_X1 U10486 ( .A(n9318), .B(n9309), .Z(n9312) );
  AOI222_X1 U10487 ( .A1(n9313), .A2(n9312), .B1(n9311), .B2(n9631), .C1(n9310), .C2(n9633), .ZN(n9681) );
  MUX2_X1 U10488 ( .A(n6152), .B(n9681), .S(n9646), .Z(n9326) );
  AOI22_X1 U10489 ( .A1(n9316), .A2(n9676), .B1(n9315), .B2(n9314), .ZN(n9325)
         );
  NAND2_X1 U10490 ( .A1(n9319), .A2(n9318), .ZN(n9678) );
  NAND3_X1 U10491 ( .A1(n9317), .A2(n9678), .A3(n9320), .ZN(n9324) );
  AOI211_X1 U10492 ( .C1(n9676), .C2(n9321), .A(n9706), .B(n9608), .ZN(n9675)
         );
  NAND2_X1 U10493 ( .A1(n9675), .A2(n9322), .ZN(n9323) );
  NAND4_X1 U10494 ( .A1(n9326), .A2(n9325), .A3(n9324), .A4(n9323), .ZN(
        P1_U3286) );
  AOI22_X1 U10495 ( .A1(n9328), .A2(n9667), .B1(n9677), .B2(n9327), .ZN(n9329)
         );
  AOI22_X1 U10496 ( .A1(n9334), .A2(n9667), .B1(n9677), .B2(n9333), .ZN(n9335)
         );
  OAI211_X1 U10497 ( .C1(n9337), .C2(n9696), .A(n9336), .B(n9335), .ZN(n9406)
         );
  MUX2_X1 U10498 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9406), .S(n9729), .Z(
        P1_U3551) );
  AOI21_X1 U10499 ( .B1(n9677), .B2(n9339), .A(n9338), .ZN(n9340) );
  OAI211_X1 U10500 ( .C1(n9342), .C2(n9696), .A(n9341), .B(n9340), .ZN(n9407)
         );
  MUX2_X1 U10501 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9407), .S(n9729), .Z(
        P1_U3550) );
  AOI22_X1 U10502 ( .A1(n9344), .A2(n9667), .B1(n9677), .B2(n9343), .ZN(n9345)
         );
  OAI211_X1 U10503 ( .C1(n9347), .C2(n9696), .A(n9346), .B(n9345), .ZN(n9408)
         );
  MUX2_X1 U10504 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9408), .S(n9729), .Z(
        P1_U3549) );
  AOI22_X1 U10505 ( .A1(n9349), .A2(n9667), .B1(n9677), .B2(n9348), .ZN(n9350)
         );
  OAI211_X1 U10506 ( .C1(n9352), .C2(n9696), .A(n9351), .B(n9350), .ZN(n9409)
         );
  MUX2_X1 U10507 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9409), .S(n9729), .Z(
        P1_U3548) );
  AOI21_X1 U10508 ( .B1(n9677), .B2(n9354), .A(n9353), .ZN(n9355) );
  OAI211_X1 U10509 ( .C1(n9696), .C2(n9357), .A(n9356), .B(n9355), .ZN(n9410)
         );
  MUX2_X1 U10510 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9410), .S(n9729), .Z(
        P1_U3547) );
  AOI22_X1 U10511 ( .A1(n9359), .A2(n9667), .B1(n9677), .B2(n9358), .ZN(n9360)
         );
  OAI211_X1 U10512 ( .C1(n9362), .C2(n9696), .A(n9361), .B(n9360), .ZN(n9411)
         );
  MUX2_X1 U10513 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9411), .S(n9729), .Z(
        P1_U3546) );
  AOI21_X1 U10514 ( .B1(n9677), .B2(n9364), .A(n9363), .ZN(n9365) );
  OAI211_X1 U10515 ( .C1(n9367), .C2(n9696), .A(n9366), .B(n9365), .ZN(n9412)
         );
  MUX2_X1 U10516 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9412), .S(n9729), .Z(
        P1_U3545) );
  OAI21_X1 U10517 ( .B1(n9370), .B2(n9705), .A(n9369), .ZN(n9371) );
  NOR2_X1 U10518 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  NAND2_X1 U10519 ( .A1(n9374), .A2(n9373), .ZN(n9413) );
  MUX2_X1 U10520 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9413), .S(n9729), .Z(
        P1_U3544) );
  AOI22_X1 U10521 ( .A1(n9376), .A2(n9667), .B1(n9677), .B2(n9375), .ZN(n9377)
         );
  OAI211_X1 U10522 ( .C1(n9379), .C2(n9696), .A(n9378), .B(n9377), .ZN(n9414)
         );
  MUX2_X1 U10523 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9414), .S(n9729), .Z(
        P1_U3543) );
  AOI21_X1 U10524 ( .B1(n9677), .B2(n9381), .A(n9380), .ZN(n9382) );
  OAI211_X1 U10525 ( .C1(n9384), .C2(n9696), .A(n9383), .B(n9382), .ZN(n9415)
         );
  MUX2_X1 U10526 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9415), .S(n9729), .Z(
        P1_U3542) );
  AOI21_X1 U10527 ( .B1(n9677), .B2(n9386), .A(n9385), .ZN(n9387) );
  OAI211_X1 U10528 ( .C1(n9696), .C2(n9389), .A(n9388), .B(n9387), .ZN(n9416)
         );
  MUX2_X1 U10529 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9416), .S(n9729), .Z(
        P1_U3541) );
  AOI21_X1 U10530 ( .B1(n9677), .B2(n9391), .A(n9390), .ZN(n9392) );
  OAI211_X1 U10531 ( .C1(n9394), .C2(n9696), .A(n9393), .B(n9392), .ZN(n9417)
         );
  MUX2_X1 U10532 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9417), .S(n9729), .Z(
        P1_U3540) );
  AOI22_X1 U10533 ( .A1(n9396), .A2(n9667), .B1(n9677), .B2(n9395), .ZN(n9397)
         );
  OAI211_X1 U10534 ( .C1(n9399), .C2(n9696), .A(n9398), .B(n9397), .ZN(n9418)
         );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9418), .S(n9729), .Z(
        P1_U3538) );
  AOI22_X1 U10536 ( .A1(n9401), .A2(n9667), .B1(n9677), .B2(n9400), .ZN(n9402)
         );
  OAI211_X1 U10537 ( .C1(n9404), .C2(n9696), .A(n9403), .B(n9402), .ZN(n9419)
         );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9419), .S(n9729), .Z(
        P1_U3536) );
  MUX2_X1 U10539 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9405), .S(n9729), .Z(
        P1_U3523) );
  MUX2_X1 U10540 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9406), .S(n9714), .Z(
        P1_U3519) );
  MUX2_X1 U10541 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9407), .S(n9714), .Z(
        P1_U3518) );
  MUX2_X1 U10542 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9408), .S(n9714), .Z(
        P1_U3517) );
  MUX2_X1 U10543 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9409), .S(n9714), .Z(
        P1_U3516) );
  MUX2_X1 U10544 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9410), .S(n9714), .Z(
        P1_U3515) );
  MUX2_X1 U10545 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9411), .S(n9714), .Z(
        P1_U3514) );
  MUX2_X1 U10546 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9412), .S(n9714), .Z(
        P1_U3513) );
  MUX2_X1 U10547 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9413), .S(n9714), .Z(
        P1_U3512) );
  MUX2_X1 U10548 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9414), .S(n9714), .Z(
        P1_U3511) );
  MUX2_X1 U10549 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9415), .S(n9714), .Z(
        P1_U3510) );
  MUX2_X1 U10550 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9416), .S(n9714), .Z(
        P1_U3508) );
  MUX2_X1 U10551 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9417), .S(n9714), .Z(
        P1_U3505) );
  MUX2_X1 U10552 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9418), .S(n9714), .Z(
        P1_U3499) );
  MUX2_X1 U10553 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9419), .S(n9714), .Z(
        P1_U3493) );
  NOR4_X1 U10554 ( .A1(n4879), .A2(P1_IR_REG_30__SCAN_IN), .A3(n4880), .A4(
        P1_U3084), .ZN(n9420) );
  AOI21_X1 U10555 ( .B1(n9429), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9420), .ZN(
        n9421) );
  OAI21_X1 U10556 ( .B1(n9422), .B2(n9431), .A(n9421), .ZN(P1_U3322) );
  AOI22_X1 U10557 ( .A1(n9423), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9429), .ZN(n9424) );
  OAI21_X1 U10558 ( .B1(n9425), .B2(n9431), .A(n9424), .ZN(P1_U3323) );
  AOI22_X1 U10559 ( .A1(n9426), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9429), .ZN(n9427) );
  OAI21_X1 U10560 ( .B1(n9428), .B2(n9431), .A(n9427), .ZN(P1_U3324) );
  AOI22_X1 U10561 ( .A1(n9512), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9429), .ZN(n9430) );
  OAI21_X1 U10562 ( .B1(n9432), .B2(n9431), .A(n9430), .ZN(P1_U3325) );
  MUX2_X1 U10563 ( .A(n9433), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  MUX2_X1 U10564 ( .A(n4912), .B(P2_ADDR_REG_19__SCAN_IN), .S(
        P1_ADDR_REG_19__SCAN_IN), .Z(n9464) );
  NOR2_X1 U10565 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9434) );
  AOI21_X1 U10566 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9434), .ZN(n9913) );
  NOR2_X1 U10567 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9435) );
  AOI21_X1 U10568 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9435), .ZN(n9916) );
  NOR2_X1 U10569 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9436) );
  AOI21_X1 U10570 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9436), .ZN(n9919) );
  NOR2_X1 U10571 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9437) );
  AOI21_X1 U10572 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9437), .ZN(n9922) );
  NOR2_X1 U10573 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9438) );
  AOI21_X1 U10574 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9438), .ZN(n9925) );
  NOR2_X1 U10575 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9444) );
  XNOR2_X1 U10576 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10137) );
  NAND2_X1 U10577 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9442) );
  XOR2_X1 U10578 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10135) );
  NAND2_X1 U10579 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9440) );
  XOR2_X1 U10580 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10133) );
  AOI21_X1 U10581 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9907) );
  INV_X1 U10582 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10081) );
  NAND3_X1 U10583 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9909) );
  OAI21_X1 U10584 ( .B1(n9907), .B2(n10081), .A(n9909), .ZN(n10132) );
  NAND2_X1 U10585 ( .A1(n10133), .A2(n10132), .ZN(n9439) );
  NAND2_X1 U10586 ( .A1(n9440), .A2(n9439), .ZN(n10134) );
  NAND2_X1 U10587 ( .A1(n10135), .A2(n10134), .ZN(n9441) );
  NAND2_X1 U10588 ( .A1(n9442), .A2(n9441), .ZN(n10136) );
  NOR2_X1 U10589 ( .A1(n10137), .A2(n10136), .ZN(n9443) );
  NOR2_X1 U10590 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  NOR2_X1 U10591 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9445), .ZN(n10121) );
  AND2_X1 U10592 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9445), .ZN(n10120) );
  NOR2_X1 U10593 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10120), .ZN(n9446) );
  NOR2_X1 U10594 ( .A1(n10121), .A2(n9446), .ZN(n9447) );
  NAND2_X1 U10595 ( .A1(n9447), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9449) );
  XOR2_X1 U10596 ( .A(n9447), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10119) );
  NAND2_X1 U10597 ( .A1(n10119), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U10598 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  NAND2_X1 U10599 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9450), .ZN(n9452) );
  XOR2_X1 U10600 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9450), .Z(n10131) );
  NAND2_X1 U10601 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10131), .ZN(n9451) );
  NAND2_X1 U10602 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  NAND2_X1 U10603 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9453), .ZN(n9456) );
  XNOR2_X1 U10604 ( .A(n9454), .B(n9453), .ZN(n10130) );
  NAND2_X1 U10605 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10130), .ZN(n9455) );
  NAND2_X1 U10606 ( .A1(n9456), .A2(n9455), .ZN(n9457) );
  AND2_X1 U10607 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9457), .ZN(n9458) );
  INV_X1 U10608 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10129) );
  XNOR2_X1 U10609 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9457), .ZN(n10128) );
  NOR2_X1 U10610 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  NAND2_X1 U10611 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9459) );
  OAI21_X1 U10612 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9459), .ZN(n9933) );
  NAND2_X1 U10613 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9460) );
  OAI21_X1 U10614 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9460), .ZN(n9930) );
  NOR2_X1 U10615 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9461) );
  AOI21_X1 U10616 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9461), .ZN(n9927) );
  NAND2_X1 U10617 ( .A1(n9928), .A2(n9927), .ZN(n9926) );
  NAND2_X1 U10618 ( .A1(n9925), .A2(n9924), .ZN(n9923) );
  OAI21_X1 U10619 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9923), .ZN(n9921) );
  NAND2_X1 U10620 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  OAI21_X1 U10621 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9920), .ZN(n9918) );
  NAND2_X1 U10622 ( .A1(n9919), .A2(n9918), .ZN(n9917) );
  OAI21_X1 U10623 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9917), .ZN(n9915) );
  NAND2_X1 U10624 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  OAI21_X1 U10625 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9914), .ZN(n9912) );
  NAND2_X1 U10626 ( .A1(n9913), .A2(n9912), .ZN(n9911) );
  OAI21_X1 U10627 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9911), .ZN(n10124) );
  NOR2_X1 U10628 ( .A1(n10125), .A2(n10124), .ZN(n9462) );
  NAND2_X1 U10629 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  OAI21_X1 U10630 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9462), .A(n10123), .ZN(
        n9463) );
  XOR2_X1 U10631 ( .A(n9464), .B(n9463), .Z(ADD_1071_U4) );
  OAI21_X1 U10632 ( .B1(n9465), .B2(n9705), .A(n9481), .ZN(n9466) );
  AOI21_X1 U10633 ( .B1(n9467), .B2(n9667), .A(n9466), .ZN(n9470) );
  INV_X1 U10634 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9468) );
  AOI22_X1 U10635 ( .A1(n9729), .A2(n9470), .B1(n9468), .B2(n9726), .ZN(
        P1_U3554) );
  INV_X1 U10636 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U10637 ( .A1(n9714), .A2(n9470), .B1(n9469), .B2(n9712), .ZN(
        P1_U3522) );
  NOR2_X1 U10638 ( .A1(n9471), .A2(n9871), .ZN(n9477) );
  OAI22_X1 U10639 ( .A1(n9473), .A2(n9881), .B1(n9472), .B2(n9879), .ZN(n9476)
         );
  INV_X1 U10640 ( .A(n9474), .ZN(n9475) );
  AOI211_X1 U10641 ( .C1(n9477), .C2(n4747), .A(n9476), .B(n9475), .ZN(n9480)
         );
  AOI22_X1 U10642 ( .A1(n9906), .A2(n9480), .B1(n9478), .B2(n9904), .ZN(
        P2_U3533) );
  INV_X1 U10643 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9479) );
  AOI22_X1 U10644 ( .A1(n9888), .A2(n9480), .B1(n9479), .B2(n9887), .ZN(
        P2_U3490) );
  INV_X1 U10645 ( .A(n9481), .ZN(n9484) );
  NOR2_X1 U10646 ( .A1(n9482), .A2(n9706), .ZN(n9483) );
  INV_X1 U10647 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9486) );
  AOI22_X1 U10648 ( .A1(n9729), .A2(n9503), .B1(n9486), .B2(n9726), .ZN(
        P1_U3553) );
  OAI211_X1 U10649 ( .C1(n9489), .C2(n9705), .A(n9488), .B(n9487), .ZN(n9490)
         );
  AOI21_X1 U10650 ( .B1(n9491), .B2(n9710), .A(n9490), .ZN(n9505) );
  AOI22_X1 U10651 ( .A1(n9729), .A2(n9505), .B1(n7362), .B2(n9726), .ZN(
        P1_U3539) );
  OAI21_X1 U10652 ( .B1(n9493), .B2(n9705), .A(n9492), .ZN(n9494) );
  AOI211_X1 U10653 ( .C1(n9496), .C2(n9710), .A(n9495), .B(n9494), .ZN(n9507)
         );
  AOI22_X1 U10654 ( .A1(n9729), .A2(n9507), .B1(n6899), .B2(n9726), .ZN(
        P1_U3537) );
  INV_X1 U10655 ( .A(n9671), .ZN(n9688) );
  INV_X1 U10656 ( .A(n9497), .ZN(n9502) );
  OAI21_X1 U10657 ( .B1(n9499), .B2(n9705), .A(n9498), .ZN(n9501) );
  AOI211_X1 U10658 ( .C1(n9688), .C2(n9502), .A(n9501), .B(n9500), .ZN(n9509)
         );
  AOI22_X1 U10659 ( .A1(n9729), .A2(n9509), .B1(n4398), .B2(n9726), .ZN(
        P1_U3535) );
  AOI22_X1 U10660 ( .A1(n9714), .A2(n9503), .B1(n8096), .B2(n9712), .ZN(
        P1_U3521) );
  INV_X1 U10661 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9504) );
  AOI22_X1 U10662 ( .A1(n9714), .A2(n9505), .B1(n9504), .B2(n9712), .ZN(
        P1_U3502) );
  INV_X1 U10663 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9506) );
  AOI22_X1 U10664 ( .A1(n9714), .A2(n9507), .B1(n9506), .B2(n9712), .ZN(
        P1_U3496) );
  INV_X1 U10665 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9508) );
  AOI22_X1 U10666 ( .A1(n9714), .A2(n9509), .B1(n9508), .B2(n9712), .ZN(
        P1_U3490) );
  XNOR2_X1 U10667 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10668 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U10669 ( .A1(n6147), .A2(n9510), .ZN(n9514) );
  OR2_X1 U10670 ( .A1(n6147), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U10671 ( .A1(n9512), .A2(n9511), .ZN(n9516) );
  NOR2_X1 U10672 ( .A1(n9516), .A2(n9514), .ZN(n9513) );
  MUX2_X1 U10673 ( .A(n9514), .B(n9513), .S(P1_IR_REG_0__SCAN_IN), .Z(n9518)
         );
  NAND2_X1 U10674 ( .A1(n9516), .A2(n9515), .ZN(n9525) );
  INV_X1 U10675 ( .A(n9525), .ZN(n9517) );
  OR2_X1 U10676 ( .A1(n9518), .A2(n9517), .ZN(n9520) );
  AOI22_X1 U10677 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9589), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n9519) );
  OAI21_X1 U10678 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(P1_U3241) );
  INV_X1 U10679 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9540) );
  INV_X1 U10680 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9532) );
  INV_X1 U10681 ( .A(n9522), .ZN(n9524) );
  MUX2_X1 U10682 ( .A(n9524), .B(n9523), .S(n6147), .Z(n9526) );
  OAI211_X1 U10683 ( .C1(n9526), .C2(n5590), .A(P1_U4006), .B(n9525), .ZN(
        n9543) );
  XNOR2_X1 U10684 ( .A(n9528), .B(n9527), .ZN(n9530) );
  AOI22_X1 U10685 ( .A1(n9593), .A2(n9530), .B1(n9578), .B2(n9529), .ZN(n9531)
         );
  OAI211_X1 U10686 ( .C1(n9584), .C2(n9532), .A(n9543), .B(n9531), .ZN(n9533)
         );
  INV_X1 U10687 ( .A(n9533), .ZN(n9539) );
  AOI211_X1 U10688 ( .C1(n9536), .C2(n9535), .A(n9534), .B(n9553), .ZN(n9537)
         );
  INV_X1 U10689 ( .A(n9537), .ZN(n9538) );
  OAI211_X1 U10690 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9540), .A(n9539), .B(
        n9538), .ZN(P1_U3243) );
  AOI22_X1 U10691 ( .A1(n9589), .A2(P1_ADDR_REG_4__SCAN_IN), .B1(n9578), .B2(
        n9541), .ZN(n9542) );
  AND2_X1 U10692 ( .A1(n9543), .A2(n9542), .ZN(n9557) );
  INV_X1 U10693 ( .A(n9544), .ZN(n9545) );
  AOI21_X1 U10694 ( .B1(n9547), .B2(n9546), .A(n9545), .ZN(n9548) );
  OR2_X1 U10695 ( .A1(n9573), .A2(n9548), .ZN(n9555) );
  AOI21_X1 U10696 ( .B1(n9551), .B2(n9550), .A(n9549), .ZN(n9552) );
  OR2_X1 U10697 ( .A1(n9553), .A2(n9552), .ZN(n9554) );
  NAND4_X1 U10698 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(
        P1_U3245) );
  AOI22_X1 U10699 ( .A1(n9589), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9578), .B2(
        n9558), .ZN(n9569) );
  AOI21_X1 U10700 ( .B1(n9561), .B2(n9560), .A(n9559), .ZN(n9562) );
  OR2_X1 U10701 ( .A1(n9573), .A2(n9562), .ZN(n9567) );
  OAI211_X1 U10702 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9598), .ZN(n9566)
         );
  NAND4_X1 U10703 ( .A1(n9569), .A2(n9568), .A3(n9567), .A4(n9566), .ZN(
        P1_U3247) );
  AOI21_X1 U10704 ( .B1(n9572), .B2(n9571), .A(n9570), .ZN(n9574) );
  NOR2_X1 U10705 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  AOI211_X1 U10706 ( .C1(n9578), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9583)
         );
  OAI211_X1 U10707 ( .C1(n9581), .C2(n9580), .A(n9598), .B(n9579), .ZN(n9582)
         );
  OAI211_X1 U10708 ( .C1(n10129), .C2(n9584), .A(n9583), .B(n9582), .ZN(
        P1_U3250) );
  NAND3_X1 U10709 ( .A1(n9596), .A2(P1_REG1_REG_11__SCAN_IN), .A3(n9593), .ZN(
        n9588) );
  NAND3_X1 U10710 ( .A1(n9601), .A2(P1_REG2_REG_11__SCAN_IN), .A3(n9585), .ZN(
        n9586) );
  NAND3_X1 U10711 ( .A1(n9588), .A2(n9587), .A3(n9586), .ZN(n9590) );
  AOI22_X1 U10712 ( .A1(n9591), .A2(n9590), .B1(n9589), .B2(
        P1_ADDR_REG_11__SCAN_IN), .ZN(n9605) );
  INV_X1 U10713 ( .A(n9592), .ZN(n9595) );
  OAI211_X1 U10714 ( .C1(n9596), .C2(n9595), .A(n9594), .B(n9593), .ZN(n9603)
         );
  NAND2_X1 U10715 ( .A1(n9597), .A2(n10068), .ZN(n9600) );
  OAI211_X1 U10716 ( .C1(n9601), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9602)
         );
  NAND4_X1 U10717 ( .A1(n9605), .A2(n9604), .A3(n9603), .A4(n9602), .ZN(
        P1_U3252) );
  OAI21_X1 U10718 ( .B1(n9607), .B2(n6680), .A(n9606), .ZN(n9687) );
  NOR2_X1 U10719 ( .A1(n9608), .A2(n9683), .ZN(n9609) );
  OR2_X1 U10720 ( .A1(n9610), .A2(n9609), .ZN(n9684) );
  INV_X1 U10721 ( .A(n9684), .ZN(n9611) );
  AOI22_X1 U10722 ( .A1(n9687), .A2(n9613), .B1(n9612), .B2(n9611), .ZN(n9627)
         );
  XNOR2_X1 U10723 ( .A(n9615), .B(n9614), .ZN(n9621) );
  OAI22_X1 U10724 ( .A1(n6619), .A2(n9618), .B1(n9617), .B2(n9616), .ZN(n9619)
         );
  AOI21_X1 U10725 ( .B1(n9687), .B2(n9630), .A(n9619), .ZN(n9620) );
  OAI21_X1 U10726 ( .B1(n8091), .B2(n9621), .A(n9620), .ZN(n9685) );
  MUX2_X1 U10727 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9685), .S(n9646), .Z(n9625)
         );
  OAI22_X1 U10728 ( .A1(n9623), .A2(n9683), .B1(n9641), .B2(n9622), .ZN(n9624)
         );
  NOR2_X1 U10729 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  NAND2_X1 U10730 ( .A1(n9627), .A2(n9626), .ZN(P1_U3285) );
  NAND2_X1 U10731 ( .A1(n9653), .A2(n9630), .ZN(n9635) );
  AOI22_X1 U10732 ( .A1(n9633), .A2(n6488), .B1(n9632), .B2(n9631), .ZN(n9634)
         );
  OAI211_X1 U10733 ( .C1(n9636), .C2(n8091), .A(n9635), .B(n9634), .ZN(n9651)
         );
  OAI21_X1 U10734 ( .B1(n6487), .B2(n9637), .A(n9667), .ZN(n9640) );
  NOR2_X1 U10735 ( .A1(n4643), .A2(n9667), .ZN(n9638) );
  AOI211_X1 U10736 ( .C1(n9705), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9652)
         );
  INV_X1 U10737 ( .A(n9652), .ZN(n9643) );
  INV_X1 U10738 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9642) );
  OAI22_X1 U10739 ( .A1(n9643), .A2(n9710), .B1(n9642), .B2(n9641), .ZN(n9644)
         );
  AOI211_X1 U10740 ( .C1(n9645), .C2(n9653), .A(n9651), .B(n9644), .ZN(n9647)
         );
  AOI22_X1 U10741 ( .A1(n9648), .A2(n4515), .B1(n9647), .B2(n9646), .ZN(
        P1_U3290) );
  INV_X1 U10742 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U10743 ( .A1(n9649), .A2(n10093), .ZN(P1_U3292) );
  AND2_X1 U10744 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9650), .ZN(P1_U3293) );
  AND2_X1 U10745 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9650), .ZN(P1_U3294) );
  AND2_X1 U10746 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9650), .ZN(P1_U3295) );
  INV_X1 U10747 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10095) );
  NOR2_X1 U10748 ( .A1(n9649), .A2(n10095), .ZN(P1_U3296) );
  AND2_X1 U10749 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9650), .ZN(P1_U3297) );
  AND2_X1 U10750 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9650), .ZN(P1_U3298) );
  AND2_X1 U10751 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9650), .ZN(P1_U3299) );
  INV_X1 U10752 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10102) );
  NOR2_X1 U10753 ( .A1(n9649), .A2(n10102), .ZN(P1_U3300) );
  AND2_X1 U10754 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9650), .ZN(P1_U3301) );
  AND2_X1 U10755 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9650), .ZN(P1_U3302) );
  AND2_X1 U10756 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9650), .ZN(P1_U3303) );
  AND2_X1 U10757 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9650), .ZN(P1_U3304) );
  AND2_X1 U10758 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9650), .ZN(P1_U3305) );
  AND2_X1 U10759 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9650), .ZN(P1_U3306) );
  AND2_X1 U10760 ( .A1(n9650), .A2(P1_D_REG_16__SCAN_IN), .ZN(P1_U3307) );
  AND2_X1 U10761 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9650), .ZN(P1_U3308) );
  AND2_X1 U10762 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9650), .ZN(P1_U3309) );
  AND2_X1 U10763 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9650), .ZN(P1_U3310) );
  INV_X1 U10764 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9948) );
  NOR2_X1 U10765 ( .A1(n9649), .A2(n9948), .ZN(P1_U3311) );
  AND2_X1 U10766 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9650), .ZN(P1_U3312) );
  AND2_X1 U10767 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9650), .ZN(P1_U3313) );
  AND2_X1 U10768 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9650), .ZN(P1_U3314) );
  AND2_X1 U10769 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9650), .ZN(P1_U3315) );
  AND2_X1 U10770 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9650), .ZN(P1_U3316) );
  AND2_X1 U10771 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9650), .ZN(P1_U3317) );
  AND2_X1 U10772 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9650), .ZN(P1_U3318) );
  AND2_X1 U10773 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9650), .ZN(P1_U3319) );
  AND2_X1 U10774 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9650), .ZN(P1_U3320) );
  AND2_X1 U10775 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9650), .ZN(P1_U3321) );
  AOI211_X1 U10776 ( .C1(n9653), .C2(n9688), .A(n9652), .B(n9651), .ZN(n9715)
         );
  INV_X1 U10777 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U10778 ( .A1(n9714), .A2(n9715), .B1(n9654), .B2(n9712), .ZN(
        P1_U3457) );
  OAI22_X1 U10779 ( .A1(n9655), .A2(n9706), .B1(n6492), .B2(n9705), .ZN(n9657)
         );
  AOI211_X1 U10780 ( .C1(n9688), .C2(n9658), .A(n9657), .B(n9656), .ZN(n9717)
         );
  INV_X1 U10781 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U10782 ( .A1(n9714), .A2(n9717), .B1(n9659), .B2(n9712), .ZN(
        P1_U3460) );
  INV_X1 U10783 ( .A(n9660), .ZN(n9664) );
  OAI22_X1 U10784 ( .A1(n9661), .A2(n9706), .B1(n6313), .B2(n9705), .ZN(n9663)
         );
  AOI211_X1 U10785 ( .C1(n9688), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9718)
         );
  INV_X1 U10786 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9665) );
  AOI22_X1 U10787 ( .A1(n9714), .A2(n9718), .B1(n9665), .B2(n9712), .ZN(
        P1_U3463) );
  AOI22_X1 U10788 ( .A1(n9668), .A2(n9667), .B1(n9677), .B2(n9666), .ZN(n9669)
         );
  OAI211_X1 U10789 ( .C1(n9672), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9673)
         );
  INV_X1 U10790 ( .A(n9673), .ZN(n9719) );
  INV_X1 U10791 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U10792 ( .A1(n9714), .A2(n9719), .B1(n9674), .B2(n9712), .ZN(
        P1_U3466) );
  AOI21_X1 U10793 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9680) );
  NAND3_X1 U10794 ( .A1(n9317), .A2(n9678), .A3(n9710), .ZN(n9679) );
  AND3_X1 U10795 ( .A1(n9681), .A2(n9680), .A3(n9679), .ZN(n9721) );
  INV_X1 U10796 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9682) );
  AOI22_X1 U10797 ( .A1(n9714), .A2(n9721), .B1(n9682), .B2(n9712), .ZN(
        P1_U3469) );
  OAI22_X1 U10798 ( .A1(n9684), .A2(n9706), .B1(n9683), .B2(n9705), .ZN(n9686)
         );
  AOI211_X1 U10799 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9722)
         );
  INV_X1 U10800 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9689) );
  AOI22_X1 U10801 ( .A1(n9714), .A2(n9722), .B1(n9689), .B2(n9712), .ZN(
        P1_U3472) );
  OAI211_X1 U10802 ( .C1(n9692), .C2(n9705), .A(n9691), .B(n9690), .ZN(n9693)
         );
  AOI21_X1 U10803 ( .B1(n9710), .B2(n9694), .A(n9693), .ZN(n9723) );
  INV_X1 U10804 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U10805 ( .A1(n9714), .A2(n9723), .B1(n9695), .B2(n9712), .ZN(
        P1_U3475) );
  NOR2_X1 U10806 ( .A1(n9697), .A2(n9696), .ZN(n9703) );
  OAI22_X1 U10807 ( .A1(n9699), .A2(n9706), .B1(n9698), .B2(n9705), .ZN(n9701)
         );
  AOI211_X1 U10808 ( .C1(n9703), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9725)
         );
  INV_X1 U10809 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U10810 ( .A1(n9714), .A2(n9725), .B1(n9937), .B2(n9712), .ZN(
        P1_U3478) );
  OAI22_X1 U10811 ( .A1(n9707), .A2(n9706), .B1(n4606), .B2(n9705), .ZN(n9709)
         );
  AOI211_X1 U10812 ( .C1(n9711), .C2(n9710), .A(n9709), .B(n9708), .ZN(n9728)
         );
  INV_X1 U10813 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9713) );
  AOI22_X1 U10814 ( .A1(n9714), .A2(n9728), .B1(n9713), .B2(n9712), .ZN(
        P1_U3481) );
  AOI22_X1 U10815 ( .A1(n9729), .A2(n9715), .B1(n9073), .B2(n9726), .ZN(
        P1_U3524) );
  AOI22_X1 U10816 ( .A1(n9729), .A2(n9717), .B1(n9716), .B2(n9726), .ZN(
        P1_U3525) );
  AOI22_X1 U10817 ( .A1(n9729), .A2(n9718), .B1(n6137), .B2(n9726), .ZN(
        P1_U3526) );
  AOI22_X1 U10818 ( .A1(n9729), .A2(n9719), .B1(n6139), .B2(n9726), .ZN(
        P1_U3527) );
  AOI22_X1 U10819 ( .A1(n9729), .A2(n9721), .B1(n9720), .B2(n9726), .ZN(
        P1_U3528) );
  AOI22_X1 U10820 ( .A1(n9729), .A2(n9722), .B1(n6133), .B2(n9726), .ZN(
        P1_U3529) );
  AOI22_X1 U10821 ( .A1(n9729), .A2(n9723), .B1(n6144), .B2(n9726), .ZN(
        P1_U3530) );
  AOI22_X1 U10822 ( .A1(n9729), .A2(n9725), .B1(n9724), .B2(n9726), .ZN(
        P1_U3531) );
  AOI22_X1 U10823 ( .A1(n9729), .A2(n9728), .B1(n9727), .B2(n9726), .ZN(
        P1_U3532) );
  OAI211_X1 U10824 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9731), .A(n9730), .B(
        P2_IR_REG_0__SCAN_IN), .ZN(n9732) );
  AOI21_X1 U10825 ( .B1(n9733), .B2(n6254), .A(n9732), .ZN(n9742) );
  AOI22_X1 U10826 ( .A1(n9735), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9734), .ZN(n9741) );
  INV_X1 U10827 ( .A(n9736), .ZN(n9737) );
  AOI21_X1 U10828 ( .B1(n9738), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9737), .ZN(
        n9739) );
  OAI221_X1 U10829 ( .B1(n9742), .B2(n9741), .C1(n9742), .C2(n9740), .A(n9739), 
        .ZN(P2_U3245) );
  NAND2_X1 U10830 ( .A1(n9744), .A2(n9743), .ZN(n9757) );
  XNOR2_X1 U10831 ( .A(n9745), .B(n9757), .ZN(n9834) );
  XNOR2_X1 U10832 ( .A(n9746), .B(n9748), .ZN(n9747) );
  NAND2_X1 U10833 ( .A1(n9747), .A2(n9837), .ZN(n9830) );
  AOI22_X1 U10834 ( .A1(n9751), .A2(n9750), .B1(n9749), .B2(n9748), .ZN(n9752)
         );
  OAI21_X1 U10835 ( .B1(n9830), .B2(n9753), .A(n9752), .ZN(n9761) );
  NAND2_X1 U10836 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  XOR2_X1 U10837 ( .A(n9757), .B(n9756), .Z(n9760) );
  OAI21_X1 U10838 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9832) );
  AOI211_X1 U10839 ( .C1(n9762), .C2(n9834), .A(n9761), .B(n9832), .ZN(n9764)
         );
  AOI22_X1 U10840 ( .A1(n8467), .A2(n5890), .B1(n9764), .B2(n9763), .ZN(
        P2_U3291) );
  INV_X1 U10841 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9767) );
  NOR2_X1 U10842 ( .A1(n9802), .A2(n9767), .ZN(P2_U3297) );
  INV_X1 U10843 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9768) );
  NOR2_X1 U10844 ( .A1(n9802), .A2(n9768), .ZN(P2_U3298) );
  INV_X1 U10845 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9769) );
  NOR2_X1 U10846 ( .A1(n9802), .A2(n9769), .ZN(P2_U3299) );
  INV_X1 U10847 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9770) );
  NOR2_X1 U10848 ( .A1(n9802), .A2(n9770), .ZN(P2_U3300) );
  INV_X1 U10849 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9771) );
  NOR2_X1 U10850 ( .A1(n9780), .A2(n9771), .ZN(P2_U3301) );
  INV_X1 U10851 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9772) );
  NOR2_X1 U10852 ( .A1(n9780), .A2(n9772), .ZN(P2_U3302) );
  NOR2_X1 U10853 ( .A1(n9780), .A2(n10057), .ZN(P2_U3303) );
  INV_X1 U10854 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9773) );
  NOR2_X1 U10855 ( .A1(n9780), .A2(n9773), .ZN(P2_U3304) );
  INV_X1 U10856 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9774) );
  NOR2_X1 U10857 ( .A1(n9780), .A2(n9774), .ZN(P2_U3305) );
  INV_X1 U10858 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9775) );
  NOR2_X1 U10859 ( .A1(n9780), .A2(n9775), .ZN(P2_U3306) );
  INV_X1 U10860 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9776) );
  NOR2_X1 U10861 ( .A1(n9780), .A2(n9776), .ZN(P2_U3307) );
  INV_X1 U10862 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9777) );
  NOR2_X1 U10863 ( .A1(n9780), .A2(n9777), .ZN(P2_U3308) );
  INV_X1 U10864 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9778) );
  NOR2_X1 U10865 ( .A1(n9780), .A2(n9778), .ZN(P2_U3309) );
  INV_X1 U10866 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9779) );
  NOR2_X1 U10867 ( .A1(n9780), .A2(n9779), .ZN(P2_U3310) );
  NOR2_X1 U10868 ( .A1(n9802), .A2(n9781), .ZN(P2_U3311) );
  INV_X1 U10869 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9782) );
  NOR2_X1 U10870 ( .A1(n9802), .A2(n9782), .ZN(P2_U3312) );
  INV_X1 U10871 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9783) );
  NOR2_X1 U10872 ( .A1(n9802), .A2(n9783), .ZN(P2_U3313) );
  INV_X1 U10873 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9784) );
  NOR2_X1 U10874 ( .A1(n9802), .A2(n9784), .ZN(P2_U3314) );
  INV_X1 U10875 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9785) );
  NOR2_X1 U10876 ( .A1(n9802), .A2(n9785), .ZN(P2_U3315) );
  INV_X1 U10877 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9786) );
  NOR2_X1 U10878 ( .A1(n9802), .A2(n9786), .ZN(P2_U3316) );
  INV_X1 U10879 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9787) );
  NOR2_X1 U10880 ( .A1(n9802), .A2(n9787), .ZN(P2_U3317) );
  INV_X1 U10881 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9788) );
  NOR2_X1 U10882 ( .A1(n9802), .A2(n9788), .ZN(P2_U3318) );
  INV_X1 U10883 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9789) );
  NOR2_X1 U10884 ( .A1(n9802), .A2(n9789), .ZN(P2_U3319) );
  INV_X1 U10885 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9790) );
  NOR2_X1 U10886 ( .A1(n9802), .A2(n9790), .ZN(P2_U3320) );
  INV_X1 U10887 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9791) );
  NOR2_X1 U10888 ( .A1(n9802), .A2(n9791), .ZN(P2_U3321) );
  INV_X1 U10889 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9792) );
  NOR2_X1 U10890 ( .A1(n9802), .A2(n9792), .ZN(P2_U3322) );
  INV_X1 U10891 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9793) );
  NOR2_X1 U10892 ( .A1(n9802), .A2(n9793), .ZN(P2_U3323) );
  INV_X1 U10893 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9794) );
  NOR2_X1 U10894 ( .A1(n9802), .A2(n9794), .ZN(P2_U3324) );
  NOR2_X1 U10895 ( .A1(n9802), .A2(n9795), .ZN(P2_U3325) );
  NOR2_X1 U10896 ( .A1(n9802), .A2(n9796), .ZN(P2_U3326) );
  INV_X1 U10897 ( .A(n9797), .ZN(n9801) );
  OAI22_X1 U10898 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9802), .B1(n9801), .B2(
        n9798), .ZN(n9799) );
  INV_X1 U10899 ( .A(n9799), .ZN(P2_U3437) );
  OAI22_X1 U10900 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9802), .B1(n9801), .B2(
        n9800), .ZN(n9803) );
  INV_X1 U10901 ( .A(n9803), .ZN(P2_U3438) );
  AOI22_X1 U10902 ( .A1(n9806), .A2(n9885), .B1(n9805), .B2(n9804), .ZN(n9807)
         );
  AND2_X1 U10903 ( .A1(n9808), .A2(n9807), .ZN(n9890) );
  INV_X1 U10904 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9809) );
  AOI22_X1 U10905 ( .A1(n9888), .A2(n9890), .B1(n9809), .B2(n9887), .ZN(
        P2_U3451) );
  NAND3_X1 U10906 ( .A1(n9811), .A2(n9837), .A3(n9810), .ZN(n9812) );
  OAI21_X1 U10907 ( .B1(n9813), .B2(n9879), .A(n9812), .ZN(n9815) );
  AOI211_X1 U10908 ( .C1(n9885), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9891)
         );
  AOI22_X1 U10909 ( .A1(n9888), .A2(n9891), .B1(n5799), .B2(n9887), .ZN(
        P2_U3454) );
  NAND3_X1 U10910 ( .A1(n9818), .A2(n9837), .A3(n9817), .ZN(n9819) );
  OAI21_X1 U10911 ( .B1(n9820), .B2(n9879), .A(n9819), .ZN(n9822) );
  AOI211_X1 U10912 ( .C1(n9885), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9893)
         );
  AOI22_X1 U10913 ( .A1(n9888), .A2(n9893), .B1(n5815), .B2(n9887), .ZN(
        P2_U3457) );
  OAI22_X1 U10914 ( .A1(n9825), .A2(n9881), .B1(n9824), .B2(n9879), .ZN(n9828)
         );
  INV_X1 U10915 ( .A(n9826), .ZN(n9827) );
  AOI211_X1 U10916 ( .C1(n9885), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9894)
         );
  AOI22_X1 U10917 ( .A1(n9888), .A2(n9894), .B1(n5851), .B2(n9887), .ZN(
        P2_U3463) );
  OAI21_X1 U10918 ( .B1(n9831), .B2(n9879), .A(n9830), .ZN(n9833) );
  AOI211_X1 U10919 ( .C1(n9885), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9895)
         );
  AOI22_X1 U10920 ( .A1(n9888), .A2(n9895), .B1(n5891), .B2(n9887), .ZN(
        P2_U3466) );
  AOI22_X1 U10921 ( .A1(n9838), .A2(n9837), .B1(n9836), .B2(n9835), .ZN(n9841)
         );
  NAND3_X1 U10922 ( .A1(n8515), .A2(n9839), .A3(n9885), .ZN(n9840) );
  AND3_X1 U10923 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(n9897) );
  INV_X1 U10924 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U10925 ( .A1(n9888), .A2(n9897), .B1(n9843), .B2(n9887), .ZN(
        P2_U3469) );
  OAI22_X1 U10926 ( .A1(n9845), .A2(n9881), .B1(n9844), .B2(n9879), .ZN(n9847)
         );
  AOI211_X1 U10927 ( .C1(n9848), .C2(n9885), .A(n9847), .B(n9846), .ZN(n9899)
         );
  AOI22_X1 U10928 ( .A1(n9888), .A2(n9899), .B1(n5880), .B2(n9887), .ZN(
        P2_U3472) );
  INV_X1 U10929 ( .A(n9849), .ZN(n9869) );
  INV_X1 U10930 ( .A(n9850), .ZN(n9855) );
  OAI22_X1 U10931 ( .A1(n9852), .A2(n9881), .B1(n9851), .B2(n9879), .ZN(n9854)
         );
  AOI211_X1 U10932 ( .C1(n9869), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9900)
         );
  AOI22_X1 U10933 ( .A1(n9888), .A2(n9900), .B1(n5939), .B2(n9887), .ZN(
        P2_U3475) );
  INV_X1 U10934 ( .A(n9856), .ZN(n9861) );
  OAI22_X1 U10935 ( .A1(n9858), .A2(n9881), .B1(n9857), .B2(n9879), .ZN(n9860)
         );
  AOI211_X1 U10936 ( .C1(n9869), .C2(n9861), .A(n9860), .B(n9859), .ZN(n9901)
         );
  AOI22_X1 U10937 ( .A1(n9888), .A2(n9901), .B1(n5955), .B2(n9887), .ZN(
        P2_U3478) );
  INV_X1 U10938 ( .A(n9862), .ZN(n9868) );
  INV_X1 U10939 ( .A(n9863), .ZN(n9864) );
  OAI22_X1 U10940 ( .A1(n9865), .A2(n9881), .B1(n9864), .B2(n9879), .ZN(n9867)
         );
  AOI211_X1 U10941 ( .C1(n9869), .C2(n9868), .A(n9867), .B(n9866), .ZN(n9902)
         );
  INV_X1 U10942 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U10943 ( .A1(n9888), .A2(n9902), .B1(n9870), .B2(n9887), .ZN(
        P2_U3481) );
  OR2_X1 U10944 ( .A1(n9872), .A2(n9871), .ZN(n9878) );
  OAI22_X1 U10945 ( .A1(n9874), .A2(n9881), .B1(n9873), .B2(n9879), .ZN(n9875)
         );
  NOR2_X1 U10946 ( .A1(n9876), .A2(n9875), .ZN(n9877) );
  AOI22_X1 U10947 ( .A1(n9888), .A2(n9903), .B1(n5995), .B2(n9887), .ZN(
        P2_U3484) );
  OAI22_X1 U10948 ( .A1(n9882), .A2(n9881), .B1(n9880), .B2(n9879), .ZN(n9883)
         );
  AOI211_X1 U10949 ( .C1(n9886), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9905)
         );
  AOI22_X1 U10950 ( .A1(n9888), .A2(n9905), .B1(n6013), .B2(n9887), .ZN(
        P2_U3487) );
  INV_X1 U10951 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10952 ( .A1(n9906), .A2(n9890), .B1(n9889), .B2(n9904), .ZN(
        P2_U3520) );
  INV_X1 U10953 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U10954 ( .A1(n9906), .A2(n9891), .B1(n9950), .B2(n9904), .ZN(
        P2_U3521) );
  INV_X1 U10955 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U10956 ( .A1(n9906), .A2(n9893), .B1(n9892), .B2(n9904), .ZN(
        P2_U3522) );
  AOI22_X1 U10957 ( .A1(n9906), .A2(n9894), .B1(n6272), .B2(n9904), .ZN(
        P2_U3524) );
  INV_X1 U10958 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U10959 ( .A1(n9906), .A2(n9895), .B1(n9969), .B2(n9904), .ZN(
        P2_U3525) );
  INV_X1 U10960 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10961 ( .A1(n9906), .A2(n9897), .B1(n9896), .B2(n9904), .ZN(
        P2_U3526) );
  INV_X1 U10962 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U10963 ( .A1(n9906), .A2(n9899), .B1(n9898), .B2(n9904), .ZN(
        P2_U3527) );
  AOI22_X1 U10964 ( .A1(n9906), .A2(n9900), .B1(n6467), .B2(n9904), .ZN(
        P2_U3528) );
  AOI22_X1 U10965 ( .A1(n9906), .A2(n9901), .B1(n6602), .B2(n9904), .ZN(
        P2_U3529) );
  AOI22_X1 U10966 ( .A1(n9906), .A2(n9902), .B1(n6766), .B2(n9904), .ZN(
        P2_U3530) );
  AOI22_X1 U10967 ( .A1(n9906), .A2(n9903), .B1(n7025), .B2(n9904), .ZN(
        P2_U3531) );
  AOI22_X1 U10968 ( .A1(n9906), .A2(n9905), .B1(n7167), .B2(n9904), .ZN(
        P2_U3532) );
  INV_X1 U10969 ( .A(n9907), .ZN(n9908) );
  NAND2_X1 U10970 ( .A1(n9909), .A2(n9908), .ZN(n9910) );
  XOR2_X1 U10971 ( .A(n10081), .B(n9910), .Z(ADD_1071_U5) );
  XOR2_X1 U10972 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10973 ( .B1(n9913), .B2(n9912), .A(n9911), .ZN(ADD_1071_U56) );
  OAI21_X1 U10974 ( .B1(n9916), .B2(n9915), .A(n9914), .ZN(ADD_1071_U57) );
  OAI21_X1 U10975 ( .B1(n9919), .B2(n9918), .A(n9917), .ZN(ADD_1071_U58) );
  OAI21_X1 U10976 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(ADD_1071_U59) );
  OAI21_X1 U10977 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(ADD_1071_U60) );
  OAI21_X1 U10978 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(ADD_1071_U61) );
  AOI21_X1 U10979 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(ADD_1071_U62) );
  AOI21_X1 U10980 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(ADD_1071_U63) );
  AOI22_X1 U10981 ( .A1(n7292), .A2(keyinput120), .B1(keyinput98), .B2(n7602), 
        .ZN(n9935) );
  OAI221_X1 U10982 ( .B1(n7292), .B2(keyinput120), .C1(n7602), .C2(keyinput98), 
        .A(n9935), .ZN(n9944) );
  AOI22_X1 U10983 ( .A1(n10069), .A2(keyinput127), .B1(n9937), .B2(keyinput91), 
        .ZN(n9936) );
  OAI221_X1 U10984 ( .B1(n10069), .B2(keyinput127), .C1(n9937), .C2(keyinput91), .A(n9936), .ZN(n9943) );
  INV_X1 U10985 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U10986 ( .A1(n8512), .A2(keyinput65), .B1(n10100), .B2(keyinput108), 
        .ZN(n9938) );
  OAI221_X1 U10987 ( .B1(n8512), .B2(keyinput65), .C1(n10100), .C2(keyinput108), .A(n9938), .ZN(n9942) );
  XOR2_X1 U10988 ( .A(n5688), .B(keyinput70), .Z(n9940) );
  XNOR2_X1 U10989 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput126), .ZN(n9939) );
  NAND2_X1 U10990 ( .A1(n9940), .A2(n9939), .ZN(n9941) );
  NOR4_X1 U10991 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9980)
         );
  AOI22_X1 U10992 ( .A1(P2_D_REG_17__SCAN_IN), .A2(keyinput96), .B1(
        P2_IR_REG_19__SCAN_IN), .B2(keyinput67), .ZN(n9945) );
  OAI221_X1 U10993 ( .B1(P2_D_REG_17__SCAN_IN), .B2(keyinput96), .C1(
        P2_IR_REG_19__SCAN_IN), .C2(keyinput67), .A(n9945), .ZN(n9956) );
  AOI22_X1 U10994 ( .A1(n9948), .A2(keyinput110), .B1(keyinput84), .B2(n9947), 
        .ZN(n9946) );
  OAI221_X1 U10995 ( .B1(n9948), .B2(keyinput110), .C1(n9947), .C2(keyinput84), 
        .A(n9946), .ZN(n9955) );
  AOI22_X1 U10996 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(keyinput111), .B1(
        P2_D_REG_25__SCAN_IN), .B2(keyinput106), .ZN(n9949) );
  OAI221_X1 U10997 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(keyinput111), .C1(
        P2_D_REG_25__SCAN_IN), .C2(keyinput106), .A(n9949), .ZN(n9954) );
  XOR2_X1 U10998 ( .A(n9950), .B(keyinput89), .Z(n9952) );
  XNOR2_X1 U10999 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput118), .ZN(n9951) );
  NAND2_X1 U11000 ( .A1(n9952), .A2(n9951), .ZN(n9953) );
  NOR4_X1 U11001 ( .A1(n9956), .A2(n9955), .A3(n9954), .A4(n9953), .ZN(n9979)
         );
  AOI22_X1 U11002 ( .A1(n10071), .A2(keyinput104), .B1(keyinput117), .B2(n9958), .ZN(n9957) );
  OAI221_X1 U11003 ( .B1(n10071), .B2(keyinput104), .C1(n9958), .C2(
        keyinput117), .A(n9957), .ZN(n9966) );
  AOI22_X1 U11004 ( .A1(n10060), .A2(keyinput113), .B1(n10068), .B2(keyinput88), .ZN(n9959) );
  OAI221_X1 U11005 ( .B1(n10060), .B2(keyinput113), .C1(n10068), .C2(
        keyinput88), .A(n9959), .ZN(n9965) );
  AOI22_X1 U11006 ( .A1(n9961), .A2(keyinput83), .B1(keyinput125), .B2(n10103), 
        .ZN(n9960) );
  OAI221_X1 U11007 ( .B1(n9961), .B2(keyinput83), .C1(n10103), .C2(keyinput125), .A(n9960), .ZN(n9964) );
  INV_X1 U11008 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U11009 ( .A1(n10102), .A2(keyinput103), .B1(keyinput64), .B2(n10084), .ZN(n9962) );
  OAI221_X1 U11010 ( .B1(n10102), .B2(keyinput103), .C1(n10084), .C2(
        keyinput64), .A(n9962), .ZN(n9963) );
  NOR4_X1 U11011 ( .A1(n9966), .A2(n9965), .A3(n9964), .A4(n9963), .ZN(n9978)
         );
  AOI22_X1 U11012 ( .A1(n6137), .A2(keyinput97), .B1(n10093), .B2(keyinput80), 
        .ZN(n9967) );
  OAI221_X1 U11013 ( .B1(n6137), .B2(keyinput97), .C1(n10093), .C2(keyinput80), 
        .A(n9967), .ZN(n9976) );
  AOI22_X1 U11014 ( .A1(n9970), .A2(keyinput124), .B1(keyinput87), .B2(n9969), 
        .ZN(n9968) );
  OAI221_X1 U11015 ( .B1(n9970), .B2(keyinput124), .C1(n9969), .C2(keyinput87), 
        .A(n9968), .ZN(n9975) );
  AOI22_X1 U11016 ( .A1(n6013), .A2(keyinput114), .B1(n10072), .B2(keyinput105), .ZN(n9971) );
  OAI221_X1 U11017 ( .B1(n6013), .B2(keyinput114), .C1(n10072), .C2(
        keyinput105), .A(n9971), .ZN(n9974) );
  AOI22_X1 U11018 ( .A1(n7154), .A2(keyinput73), .B1(n10061), .B2(keyinput92), 
        .ZN(n9972) );
  OAI221_X1 U11019 ( .B1(n7154), .B2(keyinput73), .C1(n10061), .C2(keyinput92), 
        .A(n9972), .ZN(n9973) );
  NOR4_X1 U11020 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n9977)
         );
  AND4_X1 U11021 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(n10114)
         );
  OAI22_X1 U11022 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(keyinput79), .B1(
        keyinput115), .B2(P2_REG0_REG_11__SCAN_IN), .ZN(n9981) );
  AOI221_X1 U11023 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(keyinput79), .C1(
        P2_REG0_REG_11__SCAN_IN), .C2(keyinput115), .A(n9981), .ZN(n9988) );
  OAI22_X1 U11024 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput74), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput82), .ZN(n9982) );
  AOI221_X1 U11025 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput74), .C1(
        keyinput82), .C2(P2_REG1_REG_26__SCAN_IN), .A(n9982), .ZN(n9987) );
  OAI22_X1 U11026 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput85), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput77), .ZN(n9983) );
  AOI221_X1 U11027 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput85), .C1(
        keyinput77), .C2(P1_REG1_REG_20__SCAN_IN), .A(n9983), .ZN(n9986) );
  OAI22_X1 U11028 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(keyinput116), .B1(
        P2_REG1_REG_23__SCAN_IN), .B2(keyinput71), .ZN(n9984) );
  AOI221_X1 U11029 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(keyinput116), .C1(
        keyinput71), .C2(P2_REG1_REG_23__SCAN_IN), .A(n9984), .ZN(n9985) );
  NAND4_X1 U11030 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n10016) );
  OAI22_X1 U11031 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput119), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(keyinput76), .ZN(n9989) );
  AOI221_X1 U11032 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput119), .C1(
        keyinput76), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n9989), .ZN(n9996) );
  OAI22_X1 U11033 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput69), .B1(
        keyinput66), .B2(P2_ADDR_REG_1__SCAN_IN), .ZN(n9990) );
  AOI221_X1 U11034 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput69), .C1(
        P2_ADDR_REG_1__SCAN_IN), .C2(keyinput66), .A(n9990), .ZN(n9995) );
  OAI22_X1 U11035 ( .A1(P1_D_REG_27__SCAN_IN), .A2(keyinput107), .B1(SI_21_), 
        .B2(keyinput72), .ZN(n9991) );
  AOI221_X1 U11036 ( .B1(P1_D_REG_27__SCAN_IN), .B2(keyinput107), .C1(
        keyinput72), .C2(SI_21_), .A(n9991), .ZN(n9994) );
  OAI22_X1 U11037 ( .A1(P1_D_REG_16__SCAN_IN), .A2(keyinput122), .B1(
        keyinput99), .B2(P2_REG3_REG_13__SCAN_IN), .ZN(n9992) );
  AOI221_X1 U11038 ( .B1(P1_D_REG_16__SCAN_IN), .B2(keyinput122), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput99), .A(n9992), .ZN(n9993) );
  NAND4_X1 U11039 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n10015) );
  OAI22_X1 U11040 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput86), .B1(
        keyinput95), .B2(P2_ADDR_REG_13__SCAN_IN), .ZN(n9997) );
  AOI221_X1 U11041 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput86), .C1(
        P2_ADDR_REG_13__SCAN_IN), .C2(keyinput95), .A(n9997), .ZN(n10004) );
  OAI22_X1 U11042 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput112), .B1(
        keyinput81), .B2(P2_REG0_REG_29__SCAN_IN), .ZN(n9998) );
  AOI221_X1 U11043 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput112), .C1(
        P2_REG0_REG_29__SCAN_IN), .C2(keyinput81), .A(n9998), .ZN(n10003) );
  OAI22_X1 U11044 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput93), .B1(
        P2_IR_REG_28__SCAN_IN), .B2(keyinput94), .ZN(n9999) );
  AOI221_X1 U11045 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput93), .C1(
        keyinput94), .C2(P2_IR_REG_28__SCAN_IN), .A(n9999), .ZN(n10002) );
  OAI22_X1 U11046 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(keyinput78), .B1(
        P2_REG0_REG_1__SCAN_IN), .B2(keyinput90), .ZN(n10000) );
  AOI221_X1 U11047 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(keyinput78), .C1(
        keyinput90), .C2(P2_REG0_REG_1__SCAN_IN), .A(n10000), .ZN(n10001) );
  NAND4_X1 U11048 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(
        n10014) );
  OAI22_X1 U11049 ( .A1(P2_REG1_REG_21__SCAN_IN), .A2(keyinput102), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(keyinput109), .ZN(n10005) );
  AOI221_X1 U11050 ( .B1(P2_REG1_REG_21__SCAN_IN), .B2(keyinput102), .C1(
        keyinput109), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10005), .ZN(n10012) );
  OAI22_X1 U11051 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(keyinput75), .B1(
        keyinput121), .B2(P2_REG3_REG_8__SCAN_IN), .ZN(n10006) );
  AOI221_X1 U11052 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(keyinput75), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput121), .A(n10006), .ZN(n10011) );
  OAI22_X1 U11053 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput101), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput68), .ZN(n10007) );
  AOI221_X1 U11054 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput101), .C1(
        keyinput68), .C2(P2_DATAO_REG_17__SCAN_IN), .A(n10007), .ZN(n10010) );
  OAI22_X1 U11055 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput100), .B1(
        P1_REG2_REG_5__SCAN_IN), .B2(keyinput123), .ZN(n10008) );
  AOI221_X1 U11056 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput100), .C1(
        keyinput123), .C2(P1_REG2_REG_5__SCAN_IN), .A(n10008), .ZN(n10009) );
  NAND4_X1 U11057 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10013) );
  NOR4_X1 U11058 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10113) );
  AOI22_X1 U11059 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput6), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput36), .ZN(n10017) );
  OAI221_X1 U11060 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput6), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput36), .A(n10017), .ZN(n10024) );
  AOI22_X1 U11061 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput57), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput22), .ZN(n10018) );
  OAI221_X1 U11062 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput57), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput22), .A(n10018), .ZN(n10023) );
  AOI22_X1 U11063 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(keyinput12), .B1(
        P2_REG0_REG_11__SCAN_IN), .B2(keyinput51), .ZN(n10019) );
  OAI221_X1 U11064 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(keyinput12), .C1(
        P2_REG0_REG_11__SCAN_IN), .C2(keyinput51), .A(n10019), .ZN(n10022) );
  AOI22_X1 U11065 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(keyinput25), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput4), .ZN(n10020) );
  OAI221_X1 U11066 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(keyinput25), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput4), .A(n10020), .ZN(n10021) );
  NOR4_X1 U11067 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10052) );
  AOI22_X1 U11068 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(keyinput33), .B1(
        P1_REG2_REG_12__SCAN_IN), .B2(keyinput56), .ZN(n10025) );
  OAI221_X1 U11069 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(keyinput33), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(keyinput56), .A(n10025), .ZN(n10032) );
  AOI22_X1 U11070 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(keyinput17), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput60), .ZN(n10026) );
  OAI221_X1 U11071 ( .B1(P2_REG0_REG_29__SCAN_IN), .B2(keyinput17), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput60), .A(n10026), .ZN(n10031) );
  AOI22_X1 U11072 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(keyinput20), .B1(
        P2_REG1_REG_21__SCAN_IN), .B2(keyinput38), .ZN(n10027) );
  OAI221_X1 U11073 ( .B1(P1_DATAO_REG_29__SCAN_IN), .B2(keyinput20), .C1(
        P2_REG1_REG_21__SCAN_IN), .C2(keyinput38), .A(n10027), .ZN(n10030) );
  AOI22_X1 U11074 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(keyinput34), .B1(
        P1_REG3_REG_25__SCAN_IN), .B2(keyinput10), .ZN(n10028) );
  OAI221_X1 U11075 ( .B1(P2_REG2_REG_22__SCAN_IN), .B2(keyinput34), .C1(
        P1_REG3_REG_25__SCAN_IN), .C2(keyinput10), .A(n10028), .ZN(n10029) );
  NOR4_X1 U11076 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .ZN(
        n10051) );
  AOI22_X1 U11077 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput35), .B1(
        P1_D_REG_16__SCAN_IN), .B2(keyinput58), .ZN(n10033) );
  OAI221_X1 U11078 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput35), .C1(
        P1_D_REG_16__SCAN_IN), .C2(keyinput58), .A(n10033), .ZN(n10040) );
  AOI22_X1 U11079 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(keyinput9), .B1(
        P1_REG2_REG_5__SCAN_IN), .B2(keyinput59), .ZN(n10034) );
  OAI221_X1 U11080 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(keyinput9), .C1(
        P1_REG2_REG_5__SCAN_IN), .C2(keyinput59), .A(n10034), .ZN(n10039) );
  AOI22_X1 U11081 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput29), .B1(
        P1_REG1_REG_18__SCAN_IN), .B2(keyinput15), .ZN(n10035) );
  OAI221_X1 U11082 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput29), .C1(
        P1_REG1_REG_18__SCAN_IN), .C2(keyinput15), .A(n10035), .ZN(n10038) );
  AOI22_X1 U11083 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(keyinput47), .B1(
        P2_IR_REG_7__SCAN_IN), .B2(keyinput52), .ZN(n10036) );
  OAI221_X1 U11084 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(keyinput47), .C1(
        P2_IR_REG_7__SCAN_IN), .C2(keyinput52), .A(n10036), .ZN(n10037) );
  NOR4_X1 U11085 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(
        n10050) );
  AOI22_X1 U11086 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(keyinput18), .B1(
        P2_IR_REG_19__SCAN_IN), .B2(keyinput3), .ZN(n10041) );
  OAI221_X1 U11087 ( .B1(P2_REG1_REG_26__SCAN_IN), .B2(keyinput18), .C1(
        P2_IR_REG_19__SCAN_IN), .C2(keyinput3), .A(n10041), .ZN(n10048) );
  AOI22_X1 U11088 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(keyinput23), .B1(SI_19_), 
        .B2(keyinput53), .ZN(n10042) );
  OAI221_X1 U11089 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(keyinput23), .C1(SI_19_), 
        .C2(keyinput53), .A(n10042), .ZN(n10047) );
  AOI22_X1 U11090 ( .A1(P2_D_REG_17__SCAN_IN), .A2(keyinput32), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput46), .ZN(n10043) );
  OAI221_X1 U11091 ( .B1(P2_D_REG_17__SCAN_IN), .B2(keyinput32), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput46), .A(n10043), .ZN(n10046) );
  AOI22_X1 U11092 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(keyinput27), .B1(n5799), 
        .B2(keyinput26), .ZN(n10044) );
  OAI221_X1 U11093 ( .B1(P1_REG0_REG_8__SCAN_IN), .B2(keyinput27), .C1(n5799), 
        .C2(keyinput26), .A(n10044), .ZN(n10045) );
  NOR4_X1 U11094 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10049) );
  NAND4_X1 U11095 ( .A1(n10052), .A2(n10051), .A3(n10050), .A4(n10049), .ZN(
        n10112) );
  INV_X1 U11096 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11097 ( .A1(n10055), .A2(keyinput5), .B1(n10054), .B2(keyinput8), 
        .ZN(n10053) );
  OAI221_X1 U11098 ( .B1(n10055), .B2(keyinput5), .C1(n10054), .C2(keyinput8), 
        .A(n10053), .ZN(n10066) );
  INV_X1 U11099 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10058) );
  AOI22_X1 U11100 ( .A1(n10058), .A2(keyinput13), .B1(keyinput42), .B2(n10057), 
        .ZN(n10056) );
  OAI221_X1 U11101 ( .B1(n10058), .B2(keyinput13), .C1(n10057), .C2(keyinput42), .A(n10056), .ZN(n10065) );
  AOI22_X1 U11102 ( .A1(n10061), .A2(keyinput28), .B1(keyinput49), .B2(n10060), 
        .ZN(n10059) );
  OAI221_X1 U11103 ( .B1(n10061), .B2(keyinput28), .C1(n10060), .C2(keyinput49), .A(n10059), .ZN(n10064) );
  AOI22_X1 U11104 ( .A1(n8512), .A2(keyinput1), .B1(keyinput31), .B2(n7248), 
        .ZN(n10062) );
  OAI221_X1 U11105 ( .B1(n8512), .B2(keyinput1), .C1(n7248), .C2(keyinput31), 
        .A(n10062), .ZN(n10063) );
  NOR4_X1 U11106 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10110) );
  AOI22_X1 U11107 ( .A1(n10069), .A2(keyinput63), .B1(n10068), .B2(keyinput24), 
        .ZN(n10067) );
  OAI221_X1 U11108 ( .B1(n10069), .B2(keyinput63), .C1(n10068), .C2(keyinput24), .A(n10067), .ZN(n10079) );
  AOI22_X1 U11109 ( .A1(n10072), .A2(keyinput41), .B1(n10071), .B2(keyinput40), 
        .ZN(n10070) );
  OAI221_X1 U11110 ( .B1(n10072), .B2(keyinput41), .C1(n10071), .C2(keyinput40), .A(n10070), .ZN(n10078) );
  XOR2_X1 U11111 ( .A(n7390), .B(keyinput14), .Z(n10076) );
  XNOR2_X1 U11112 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput62), .ZN(n10075) );
  XNOR2_X1 U11113 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput11), .ZN(n10074)
         );
  XNOR2_X1 U11114 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput7), .ZN(n10073) );
  NAND4_X1 U11115 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10077) );
  NOR3_X1 U11116 ( .A1(n10079), .A2(n10078), .A3(n10077), .ZN(n10109) );
  AOI22_X1 U11117 ( .A1(n10129), .A2(keyinput45), .B1(n10081), .B2(keyinput2), 
        .ZN(n10080) );
  OAI221_X1 U11118 ( .B1(n10129), .B2(keyinput45), .C1(n10081), .C2(keyinput2), 
        .A(n10080), .ZN(n10091) );
  AOI22_X1 U11119 ( .A1(n10084), .A2(keyinput0), .B1(keyinput55), .B2(n10083), 
        .ZN(n10082) );
  OAI221_X1 U11120 ( .B1(n10084), .B2(keyinput0), .C1(n10083), .C2(keyinput55), 
        .A(n10082), .ZN(n10090) );
  XNOR2_X1 U11121 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput19), .ZN(n10088)
         );
  XNOR2_X1 U11122 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput30), .ZN(n10087) );
  XNOR2_X1 U11123 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput54), .ZN(n10086) );
  XNOR2_X1 U11124 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput37), .ZN(n10085) );
  NAND4_X1 U11125 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10089) );
  NOR3_X1 U11126 ( .A1(n10091), .A2(n10090), .A3(n10089), .ZN(n10108) );
  INV_X1 U11127 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U11128 ( .A1(n10094), .A2(keyinput21), .B1(n10093), .B2(keyinput16), 
        .ZN(n10092) );
  OAI221_X1 U11129 ( .B1(n10094), .B2(keyinput21), .C1(n10093), .C2(keyinput16), .A(n10092), .ZN(n10098) );
  XOR2_X1 U11130 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput48), .Z(n10097) );
  XNOR2_X1 U11131 ( .A(n10095), .B(keyinput43), .ZN(n10096) );
  OR3_X1 U11132 ( .A1(n10098), .A2(n10097), .A3(n10096), .ZN(n10106) );
  AOI22_X1 U11133 ( .A1(n10100), .A2(keyinput44), .B1(keyinput50), .B2(n6013), 
        .ZN(n10099) );
  OAI221_X1 U11134 ( .B1(n10100), .B2(keyinput44), .C1(n6013), .C2(keyinput50), 
        .A(n10099), .ZN(n10105) );
  AOI22_X1 U11135 ( .A1(n10103), .A2(keyinput61), .B1(n10102), .B2(keyinput39), 
        .ZN(n10101) );
  OAI221_X1 U11136 ( .B1(n10103), .B2(keyinput61), .C1(n10102), .C2(keyinput39), .A(n10101), .ZN(n10104) );
  NOR3_X1 U11137 ( .A1(n10106), .A2(n10105), .A3(n10104), .ZN(n10107) );
  NAND4_X1 U11138 ( .A1(n10110), .A2(n10109), .A3(n10108), .A4(n10107), .ZN(
        n10111) );
  AOI211_X1 U11139 ( .C1(n10114), .C2(n10113), .A(n10112), .B(n10111), .ZN(
        n10118) );
  MUX2_X1 U11140 ( .A(n10116), .B(n10115), .S(P1_U4006), .Z(n10117) );
  XNOR2_X1 U11141 ( .A(n10118), .B(n10117), .ZN(P1_U3581) );
  XOR2_X1 U11142 ( .A(n10119), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11143 ( .A1(n10121), .A2(n10120), .ZN(n10122) );
  XOR2_X1 U11144 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10122), .Z(ADD_1071_U51) );
  OAI21_X1 U11145 ( .B1(n10125), .B2(n10124), .A(n10123), .ZN(n10126) );
  XNOR2_X1 U11146 ( .A(n10126), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11147 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(ADD_1071_U47) );
  XOR2_X1 U11148 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10130), .Z(ADD_1071_U48) );
  XOR2_X1 U11149 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10131), .Z(ADD_1071_U49) );
  XOR2_X1 U11150 ( .A(n10133), .B(n10132), .Z(ADD_1071_U54) );
  XOR2_X1 U11151 ( .A(n10135), .B(n10134), .Z(ADD_1071_U53) );
  XNOR2_X1 U11152 ( .A(n10137), .B(n10136), .ZN(ADD_1071_U52) );
  INV_X1 U4829 ( .A(n5850), .ZN(n5912) );
  CLKBUF_X1 U4830 ( .A(n4935), .Z(n5666) );
  BUF_X1 U4838 ( .A(n5040), .Z(n4316) );
  CLKBUF_X1 U5003 ( .A(n5024), .Z(n8092) );
endmodule

