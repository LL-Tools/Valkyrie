

module b21_C_SARLock_k_64_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4256, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095;

  AOI21_X1 U4762 ( .B1(n9378), .B2(n9673), .A(n4611), .ZN(n4610) );
  CLKBUF_X1 U4763 ( .A(n4962), .Z(n10095) );
  INV_X2 U4764 ( .A(n5931), .ZN(n9723) );
  CLKBUF_X2 U4765 ( .A(n7275), .Z(n4260) );
  BUF_X2 U4766 ( .A(n7275), .Z(n4261) );
  INV_X1 U4767 ( .A(n10095), .ZN(n4256) );
  INV_X1 U4768 ( .A(n4256), .ZN(P1_U3084) );
  INV_X1 U4769 ( .A(n4256), .ZN(n4258) );
  CLKBUF_X2 U4770 ( .A(n5357), .Z(n7889) );
  NAND2_X1 U4771 ( .A1(n9772), .A2(n7427), .ZN(n6986) );
  CLKBUF_X3 U4772 ( .A(n5505), .Z(n7891) );
  INV_X1 U4773 ( .A(n8198), .ZN(n4643) );
  INV_X1 U4774 ( .A(n9877), .ZN(n7401) );
  AND3_X1 U4775 ( .A1(n5989), .A2(n5988), .A3(n5987), .ZN(n9844) );
  INV_X1 U4776 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U4777 ( .A1(n7674), .A2(n7673), .ZN(n8675) );
  INV_X1 U4779 ( .A(n6162), .ZN(n9668) );
  OAI211_X1 U4780 ( .C1(n7359), .C2(n5792), .A(n5791), .B(n5790), .ZN(n6012)
         );
  MUX2_X1 U4781 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5162), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5163) );
  NAND2_X1 U4782 ( .A1(n4708), .A2(n4709), .ZN(n4951) );
  NAND2_X1 U4783 ( .A1(n6610), .A2(n6609), .ZN(n9455) );
  NAND4_X1 U4784 ( .A1(n5145), .A2(n5144), .A3(n5143), .A4(n5142), .ZN(n5581)
         );
  INV_X1 U4785 ( .A(n6110), .ZN(n8760) );
  AOI211_X1 U4786 ( .C1(n9456), .C2(n9402), .A(n9401), .B(n9400), .ZN(n9403)
         );
  INV_X1 U4787 ( .A(n5139), .ZN(n7550) );
  AND2_X1 U4789 ( .A1(n7918), .A2(n5430), .ZN(n7275) );
  NAND2_X1 U4790 ( .A1(n5951), .A2(n7333), .ZN(n5535) );
  OAI211_X1 U4791 ( .C1(n8788), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8790)
         );
  OAI21_X2 U4792 ( .B1(n7877), .B2(n8655), .A(n8656), .ZN(n8549) );
  INV_X2 U4793 ( .A(n7607), .ZN(n7612) );
  XNOR2_X1 U4794 ( .A(n4904), .B(n4903), .ZN(n5348) );
  AND2_X4 U4795 ( .A1(n7918), .A2(n8541), .ZN(n6657) );
  AOI21_X2 U4796 ( .B1(n9219), .B2(n9220), .A(n9112), .ZN(n9205) );
  OAI22_X2 U4797 ( .A1(n9249), .A2(n4615), .B1(n4617), .B2(n9109), .ZN(n9219)
         );
  NAND2_X1 U4798 ( .A1(n8613), .A2(n8612), .ZN(n8611) );
  OAI21_X1 U4799 ( .B1(n4288), .B2(n10071), .A(n4806), .ZN(n4801) );
  NAND2_X1 U4800 ( .A1(n8186), .A2(n8185), .ZN(n8184) );
  AOI21_X1 U4801 ( .B1(n8164), .B2(n9771), .A(n8163), .ZN(n8426) );
  AND2_X1 U4802 ( .A1(n8675), .A2(n8592), .ZN(n4501) );
  AND2_X1 U4803 ( .A1(n9174), .A2(n4604), .ZN(n9126) );
  AOI21_X1 U4804 ( .B1(n4701), .B2(n4597), .A(n7591), .ZN(n7590) );
  OAI22_X1 U4805 ( .A1(n7999), .A2(n7998), .B1(n7571), .B2(n7570), .ZN(n8044)
         );
  AND2_X1 U4806 ( .A1(n4485), .A2(n4269), .ZN(n4484) );
  OAI22_X1 U4807 ( .A1(n8391), .A2(n8132), .B1(n8495), .B2(n8384), .ZN(n8374)
         );
  NAND2_X1 U4808 ( .A1(n6253), .A2(n6252), .ZN(n4872) );
  NAND2_X1 U4809 ( .A1(n6973), .A2(n4296), .ZN(n9789) );
  OR2_X1 U4810 ( .A1(n6287), .A2(n7514), .ZN(n6973) );
  OAI21_X1 U4811 ( .B1(n4871), .B2(n4482), .A(n6667), .ZN(n4481) );
  AOI21_X1 U4812 ( .B1(n5713), .B2(n5712), .A(n5711), .ZN(n5718) );
  NAND2_X1 U4813 ( .A1(n6037), .A2(n7396), .ZN(n6200) );
  NAND2_X1 U4814 ( .A1(n7041), .A2(n7040), .ZN(n9506) );
  NAND2_X1 U4815 ( .A1(n6907), .A2(n6906), .ZN(n8690) );
  OR2_X1 U4816 ( .A1(n8501), .A2(n7024), .ZN(n7428) );
  OR2_X1 U4817 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  XNOR2_X1 U4818 ( .A(n5291), .B(n5290), .ZN(n6739) );
  AND2_X1 U4819 ( .A1(n7405), .A2(n7406), .ZN(n6201) );
  NAND2_X1 U4820 ( .A1(n5956), .A2(n5955), .ZN(n6107) );
  NAND2_X1 U4821 ( .A1(n7371), .A2(n7375), .ZN(n4795) );
  INV_X2 U4822 ( .A(n9783), .ZN(n9813) );
  NOR2_X2 U4823 ( .A1(n7946), .A2(n7554), .ZN(n5753) );
  AND4_X1 U4824 ( .A1(n5787), .A2(n5786), .A3(n5785), .A4(n5784), .ZN(n6005)
         );
  OR2_X1 U4825 ( .A1(n8999), .A2(n9368), .ZN(n8904) );
  INV_X2 U4826 ( .A(n7359), .ZN(n7335) );
  INV_X1 U4827 ( .A(n5700), .ZN(n5505) );
  INV_X4 U4828 ( .A(n7872), .ZN(n5361) );
  AND4_X1 U4829 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n6306)
         );
  AND4_X1 U4830 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n6316)
         );
  OAI211_X1 U4831 ( .C1(n5788), .C2(n4755), .A(n5742), .B(n5741), .ZN(n8039)
         );
  NAND4_X1 U4832 ( .A1(n5455), .A2(n5454), .A3(n5453), .A4(n5452), .ZN(n8072)
         );
  AND4_X1 U4833 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n5877)
         );
  INV_X1 U4834 ( .A(n5602), .ZN(n9368) );
  AND2_X2 U4835 ( .A1(n5349), .A2(n5357), .ZN(n5377) );
  AND4_X1 U4836 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), .ZN(n7560)
         );
  AND4_X1 U4837 ( .A1(n5623), .A2(n5622), .A3(n5621), .A4(n5620), .ZN(n5931)
         );
  NAND2_X1 U4838 ( .A1(n4502), .A2(n5494), .ZN(n5700) );
  OR2_X1 U4839 ( .A1(n5348), .A2(n5586), .ZN(n5345) );
  NOR2_X1 U4840 ( .A1(n5581), .A2(n7201), .ZN(n7194) );
  AND2_X2 U4841 ( .A1(n5430), .A2(n5429), .ZN(n7328) );
  INV_X1 U4842 ( .A(n5489), .ZN(n9824) );
  NAND4_X1 U4843 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n9000)
         );
  NAND2_X1 U4844 ( .A1(n4907), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4904) );
  AND2_X1 U4845 ( .A1(n6601), .A2(n7539), .ZN(n5489) );
  AND2_X1 U4846 ( .A1(n5266), .A2(n5265), .ZN(n5269) );
  INV_X1 U4847 ( .A(n5429), .ZN(n7918) );
  INV_X1 U4848 ( .A(n7547), .ZN(n6601) );
  NAND2_X1 U4849 ( .A1(n4931), .A2(n5241), .ZN(n5494) );
  INV_X2 U4850 ( .A(n7477), .ZN(n4262) );
  MUX2_X1 U4851 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5197), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5198) );
  INV_X1 U4852 ( .A(n9256), .ZN(n5586) );
  AND2_X1 U4853 ( .A1(n5155), .A2(n5154), .ZN(n7547) );
  INV_X1 U4854 ( .A(n5138), .ZN(n7924) );
  NAND2_X2 U4855 ( .A1(n5139), .A2(n5138), .ZN(n7863) );
  NAND2_X1 U4856 ( .A1(n4929), .A2(n4923), .ZN(n7070) );
  XNOR2_X1 U4857 ( .A(n4928), .B(n4927), .ZN(n7158) );
  INV_X2 U4858 ( .A(n9481), .ZN(n7551) );
  NAND2_X1 U4859 ( .A1(n4926), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U4860 ( .A1(n4901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U4861 ( .A1(n9476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U4862 ( .A1(n5129), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5131) );
  AND2_X1 U4863 ( .A1(n4948), .A2(n4847), .ZN(n5195) );
  OR2_X1 U4864 ( .A1(n4921), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4929) );
  INV_X4 U4865 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4866 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4540) );
  NOR2_X2 U4867 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4983) );
  NOR2_X1 U4868 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4542) );
  INV_X1 U4869 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4891) );
  NOR2_X2 U4870 ( .A1(n5664), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5232) );
  NOR2_X4 U4871 ( .A1(n9284), .A2(n9430), .ZN(n9264) );
  OR2_X2 U4872 ( .A1(n9307), .A2(n9436), .ZN(n9284) );
  INV_X2 U4873 ( .A(n6283), .ZN(n5739) );
  AND2_X1 U4874 ( .A1(n5349), .A2(n5357), .ZN(n4263) );
  INV_X2 U4875 ( .A(n5700), .ZN(n4264) );
  NOR2_X1 U4876 ( .A1(n9397), .A2(n9402), .ZN(n4608) );
  INV_X1 U4877 ( .A(n8541), .ZN(n5430) );
  OR2_X1 U4878 ( .A1(n8443), .A2(n8210), .ZN(n7472) );
  AND2_X1 U4879 ( .A1(n7472), .A2(n7470), .ZN(n8228) );
  NAND2_X1 U4880 ( .A1(n4849), .A2(n5350), .ZN(n5353) );
  INV_X1 U4881 ( .A(n4399), .ZN(n4398) );
  OAI21_X1 U4882 ( .B1(n4401), .B2(n4400), .A(n8949), .ZN(n4399) );
  OAI21_X1 U4883 ( .B1(n6183), .B2(n6182), .A(n6184), .ZN(n6370) );
  NAND2_X1 U4884 ( .A1(n5181), .A2(n4885), .ZN(n5174) );
  BUF_X1 U4885 ( .A(n5788), .Z(n7359) );
  BUF_X1 U4886 ( .A(n5535), .Z(n6110) );
  AND2_X1 U4887 ( .A1(n4273), .A2(n4319), .ZN(n4531) );
  AND2_X1 U4888 ( .A1(n7428), .A2(n7477), .ZN(n4534) );
  INV_X1 U4889 ( .A(n7566), .ZN(n4699) );
  OAI21_X1 U4890 ( .B1(n7338), .B2(n8141), .A(n7368), .ZN(n7348) );
  NOR2_X1 U4891 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4543) );
  NOR2_X1 U4892 ( .A1(n8228), .A2(n4823), .ZN(n4818) );
  INV_X1 U4893 ( .A(n5156), .ZN(n4708) );
  OR2_X1 U4894 ( .A1(n9397), .A2(n9172), .ZN(n9138) );
  NOR2_X1 U4895 ( .A1(n4719), .A2(n4381), .ZN(n4380) );
  NAND2_X1 U4896 ( .A1(n4279), .A2(n4328), .ZN(n4384) );
  NAND2_X1 U4897 ( .A1(n9089), .A2(n4277), .ZN(n4387) );
  INV_X1 U4898 ( .A(n9278), .ZN(n4631) );
  AND2_X1 U4899 ( .A1(n4270), .A2(n9351), .ZN(n4716) );
  NAND2_X1 U4900 ( .A1(n4618), .A2(n4620), .ZN(n4615) );
  AOI21_X1 U4901 ( .B1(n4618), .B2(n9246), .A(n8934), .ZN(n4617) );
  XNOR2_X1 U4902 ( .A(n7352), .B(n7351), .ZN(n7350) );
  NAND2_X1 U4903 ( .A1(n7313), .A2(n7312), .ZN(n7315) );
  NAND2_X1 U4904 ( .A1(n4454), .A2(n6596), .ZN(n6689) );
  NAND2_X1 U4905 ( .A1(n6372), .A2(n4745), .ZN(n4454) );
  AOI21_X1 U4906 ( .B1(n4433), .B2(n4435), .A(n4339), .ZN(n4431) );
  INV_X1 U4907 ( .A(n4781), .ZN(n4780) );
  OAI21_X1 U4908 ( .B1(n4784), .B2(n4280), .A(n5658), .ZN(n4781) );
  NAND2_X1 U4909 ( .A1(n4457), .A2(n4455), .ZN(n5412) );
  AOI21_X1 U4910 ( .B1(n4458), .B2(n4281), .A(n4456), .ZN(n4455) );
  INV_X1 U4911 ( .A(n4884), .ZN(n4456) );
  XNOR2_X1 U4912 ( .A(n5209), .B(SI_11_), .ZN(n5208) );
  AOI21_X1 U4913 ( .B1(n4442), .B2(n4444), .A(n4440), .ZN(n4439) );
  INV_X1 U4914 ( .A(n5168), .ZN(n4440) );
  INV_X1 U4915 ( .A(n5068), .ZN(n4649) );
  OAI21_X1 U4916 ( .B1(n7333), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4367), .ZN(
        n5080) );
  NAND2_X1 U4917 ( .A1(n7333), .A2(n5701), .ZN(n4367) );
  INV_X1 U4918 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4564) );
  NOR2_X1 U4919 ( .A1(n8416), .A2(n8143), .ZN(n7531) );
  NAND2_X1 U4920 ( .A1(n7337), .A2(n7336), .ZN(n8421) );
  NAND2_X1 U4921 ( .A1(n4814), .A2(n4813), .ZN(n8203) );
  AOI21_X1 U4922 ( .B1(n4815), .B2(n4817), .A(n8207), .ZN(n4813) );
  NAND2_X1 U4923 ( .A1(n8253), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U4924 ( .A1(n8245), .A2(n4300), .ZN(n8227) );
  OR2_X1 U4925 ( .A1(n8453), .A2(n8283), .ZN(n4824) );
  AND4_X1 U4926 ( .A1(n7252), .A2(n7251), .A3(n7250), .A4(n7249), .ZN(n8267)
         );
  NAND2_X1 U4927 ( .A1(n8288), .A2(n4332), .ZN(n8274) );
  INV_X1 U4928 ( .A(n6281), .ZN(n7358) );
  INV_X1 U4929 ( .A(n4664), .ZN(n4663) );
  INV_X1 U4930 ( .A(n4660), .ZN(n4659) );
  OAI21_X1 U4931 ( .B1(n7435), .B2(n4661), .A(n7432), .ZN(n4660) );
  NAND2_X1 U4932 ( .A1(n6283), .A2(n7355), .ZN(n6281) );
  NAND2_X2 U4933 ( .A1(n7543), .A2(n7629), .ZN(n6283) );
  NAND2_X1 U4934 ( .A1(n4799), .A2(n9771), .ZN(n4798) );
  XNOR2_X1 U4935 ( .A(n5157), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7367) );
  NOR2_X1 U4936 ( .A1(n6937), .A2(n4874), .ZN(n4873) );
  INV_X1 U4937 ( .A(n6934), .ZN(n4874) );
  AOI21_X1 U4938 ( .B1(n4480), .B2(n4482), .A(n4478), .ZN(n4477) );
  INV_X1 U4939 ( .A(n6669), .ZN(n4478) );
  INV_X1 U4940 ( .A(n9097), .ZN(n9172) );
  NAND2_X1 U4941 ( .A1(n4385), .A2(n4384), .ZN(n9199) );
  NAND2_X1 U4942 ( .A1(n9227), .A2(n4378), .ZN(n4385) );
  INV_X1 U4943 ( .A(n4381), .ZN(n4378) );
  OR2_X1 U4944 ( .A1(n9430), .A2(n9250), .ZN(n9087) );
  AND2_X1 U4945 ( .A1(n4629), .A2(n4628), .ZN(n9270) );
  AND2_X1 U4946 ( .A1(n4630), .A2(n9105), .ZN(n4628) );
  NAND2_X1 U4947 ( .A1(n4711), .A2(n4276), .ZN(n4393) );
  NAND2_X1 U4948 ( .A1(n4312), .A2(n4270), .ZN(n4715) );
  AND2_X1 U4949 ( .A1(n4890), .A2(n7039), .ZN(n4741) );
  NAND2_X1 U4950 ( .A1(n6903), .A2(n6902), .ZN(n4390) );
  NOR2_X1 U4951 ( .A1(n6606), .A2(n4736), .ZN(n4735) );
  OAI21_X1 U4952 ( .B1(n6534), .B2(n4400), .A(n4398), .ZN(n6495) );
  NOR2_X1 U4953 ( .A1(n6493), .A2(n4402), .ZN(n4401) );
  INV_X1 U4954 ( .A(n6492), .ZN(n4402) );
  OR2_X1 U4955 ( .A1(n6529), .A2(n8993), .ZN(n4403) );
  INV_X1 U4956 ( .A(n8758), .ZN(n7734) );
  OR2_X1 U4957 ( .A1(n5533), .A2(n5327), .ZN(n5329) );
  OR2_X1 U4958 ( .A1(n5535), .A2(n5740), .ZN(n5328) );
  OR2_X1 U4959 ( .A1(n8888), .A2(n9016), .ZN(n9345) );
  INV_X1 U4960 ( .A(n9391), .ZN(n4633) );
  XNOR2_X1 U4961 ( .A(n6370), .B(n6369), .ZN(n7754) );
  NAND2_X1 U4962 ( .A1(n4432), .A2(n5974), .ZN(n6020) );
  NAND2_X1 U4963 ( .A1(n5691), .A2(n4436), .ZN(n4432) );
  NAND2_X1 U4964 ( .A1(n4441), .A2(n5117), .ZN(n5167) );
  NAND2_X1 U4965 ( .A1(n5116), .A2(n5115), .ZN(n4441) );
  NAND2_X1 U4966 ( .A1(n5053), .A2(n5052), .ZN(n5060) );
  INV_X1 U4967 ( .A(n5951), .ZN(n7733) );
  NAND2_X1 U4968 ( .A1(n7856), .A2(n8760), .ZN(n7859) );
  AOI21_X1 U4969 ( .B1(n8531), .B2(n8760), .A(n8759), .ZN(n9379) );
  XNOR2_X1 U4970 ( .A(n9381), .B(n9379), .ZN(n9378) );
  NOR2_X1 U4971 ( .A1(n4531), .A2(n4336), .ZN(n4530) );
  INV_X1 U4972 ( .A(n4531), .ZN(n4528) );
  NAND2_X1 U4973 ( .A1(n4273), .A2(n7521), .ZN(n4532) );
  NAND2_X1 U4974 ( .A1(n7463), .A2(n4287), .ZN(n4522) );
  AND2_X1 U4975 ( .A1(n4524), .A2(n4521), .ZN(n4520) );
  NOR2_X1 U4976 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  NAND2_X1 U4977 ( .A1(n4287), .A2(n7462), .ZN(n4521) );
  NAND2_X1 U4978 ( .A1(n8244), .A2(n4262), .ZN(n4525) );
  NAND2_X1 U4979 ( .A1(n8246), .A2(n4518), .ZN(n4517) );
  AOI21_X1 U4980 ( .B1(n4266), .B2(n4305), .A(n4519), .ZN(n4518) );
  NAND2_X1 U4981 ( .A1(n4643), .A2(n7367), .ZN(n4536) );
  OR2_X1 U4982 ( .A1(n7362), .A2(n8116), .ZN(n7497) );
  OR2_X1 U4983 ( .A1(n7011), .A2(n7010), .ZN(n7014) );
  NOR2_X1 U4984 ( .A1(n8161), .A2(n4667), .ZN(n4666) );
  INV_X1 U4985 ( .A(n4668), .ZN(n4667) );
  INV_X1 U4986 ( .A(n7487), .ZN(n4671) );
  NAND2_X1 U4987 ( .A1(n9397), .A2(n9172), .ZN(n8879) );
  INV_X1 U4988 ( .A(n4434), .ZN(n4433) );
  OAI21_X1 U4989 ( .B1(n4436), .B2(n4435), .A(n6019), .ZN(n4434) );
  NAND2_X1 U4990 ( .A1(n5216), .A2(n5215), .ZN(n5292) );
  INV_X1 U4991 ( .A(n5117), .ZN(n4444) );
  NAND2_X1 U4992 ( .A1(n4584), .A2(n7597), .ZN(n4573) );
  NAND2_X1 U4993 ( .A1(n7492), .A2(n4744), .ZN(n4743) );
  NOR2_X1 U4994 ( .A1(n7366), .A2(n7477), .ZN(n4744) );
  OR2_X1 U4995 ( .A1(n8428), .A2(n4539), .ZN(n4538) );
  NOR2_X1 U4996 ( .A1(n8458), .A2(n8463), .ZN(n4561) );
  INV_X1 U4997 ( .A(n4837), .ZN(n4833) );
  OR2_X1 U4998 ( .A1(n8490), .A2(n8483), .ZN(n4552) );
  OR2_X1 U4999 ( .A1(n7134), .A2(n5421), .ZN(n7216) );
  AND2_X1 U5000 ( .A1(n8126), .A2(n8127), .ZN(n4812) );
  OR2_X1 U5001 ( .A1(n8125), .A2(n8124), .ZN(n8128) );
  AND2_X1 U5002 ( .A1(n7019), .A2(n7435), .ZN(n8125) );
  OR2_X1 U5003 ( .A1(n8506), .A2(n6975), .ZN(n7419) );
  NAND2_X1 U5004 ( .A1(n9844), .A2(n6004), .ZN(n4556) );
  AND2_X1 U5005 ( .A1(n4943), .A2(n4942), .ZN(n4825) );
  INV_X1 U5006 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4942) );
  AND2_X1 U5007 ( .A1(n6258), .A2(n6257), .ZN(n4871) );
  AND2_X1 U5008 ( .A1(n4870), .A2(n7714), .ZN(n4869) );
  INV_X1 U5009 ( .A(n7730), .ZN(n4870) );
  INV_X1 U5010 ( .A(n4966), .ZN(n4897) );
  INV_X1 U5011 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4894) );
  NOR2_X1 U5012 ( .A1(n9566), .A2(n9567), .ZN(n9568) );
  NOR2_X1 U5013 ( .A1(n5915), .A2(n4418), .ZN(n9566) );
  AND2_X1 U5014 ( .A1(n6608), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U5015 ( .A1(n4722), .A2(n9096), .ZN(n4721) );
  INV_X1 U5016 ( .A(n4724), .ZN(n4722) );
  INV_X1 U5017 ( .A(n4384), .ZN(n4383) );
  INV_X1 U5018 ( .A(n9096), .ZN(n4720) );
  OAI21_X1 U5019 ( .B1(n7837), .B2(n4448), .A(n4446), .ZN(n8932) );
  INV_X1 U5020 ( .A(n7839), .ZN(n4448) );
  AND2_X1 U5021 ( .A1(n9173), .A2(n4447), .ZN(n4446) );
  NAND2_X1 U5022 ( .A1(n7839), .A2(n6110), .ZN(n4447) );
  NAND2_X1 U5023 ( .A1(n4328), .A2(n4277), .ZN(n4381) );
  AOI21_X1 U5024 ( .B1(n8956), .B2(n8814), .A(n8827), .ZN(n4627) );
  OR2_X1 U5025 ( .A1(n9455), .A2(n6611), .ZN(n8818) );
  INV_X1 U5026 ( .A(n4403), .ZN(n4400) );
  OR2_X1 U5027 ( .A1(n6580), .A2(n6683), .ZN(n8701) );
  NAND2_X1 U5028 ( .A1(n4621), .A2(n8905), .ZN(n8773) );
  NAND2_X1 U5029 ( .A1(n9174), .A2(n4606), .ZN(n9142) );
  AOI21_X1 U5030 ( .B1(n4775), .B2(n7329), .A(n4348), .ZN(n4774) );
  INV_X1 U5031 ( .A(n7314), .ZN(n4775) );
  INV_X1 U5032 ( .A(n7329), .ZN(n4776) );
  NAND2_X1 U5033 ( .A1(n7149), .A2(n7148), .ZN(n7313) );
  AOI21_X1 U5034 ( .B1(n4789), .B2(n4344), .A(n4788), .ZN(n4787) );
  NOR2_X1 U5035 ( .A1(n7064), .A2(n4794), .ZN(n4793) );
  INV_X1 U5036 ( .A(n6846), .ZN(n4794) );
  NAND2_X1 U5037 ( .A1(n6845), .A2(n6844), .ZN(n6847) );
  NAND2_X1 U5038 ( .A1(n6370), .A2(n6369), .ZN(n6372) );
  AOI21_X1 U5039 ( .B1(n4780), .B2(n4280), .A(n4779), .ZN(n4778) );
  INV_X1 U5040 ( .A(n5688), .ZN(n4779) );
  NOR2_X1 U5041 ( .A1(n5212), .A2(n4463), .ZN(n4462) );
  INV_X1 U5042 ( .A(n5173), .ZN(n4463) );
  INV_X1 U5043 ( .A(n5208), .ZN(n5212) );
  NAND2_X1 U5044 ( .A1(n5117), .A2(n5102), .ZN(n5112) );
  OAI21_X1 U5045 ( .B1(n7333), .B2(n4755), .A(n4754), .ZN(n5051) );
  NAND2_X1 U5046 ( .A1(n7333), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U5047 ( .A1(n9746), .A2(n4704), .ZN(n6332) );
  NOR2_X1 U5048 ( .A1(n6324), .A2(n4705), .ZN(n4704) );
  INV_X1 U5049 ( .A(n6315), .ZN(n4705) );
  AND2_X1 U5050 ( .A1(n7099), .A2(n4689), .ZN(n4688) );
  OR2_X1 U5051 ( .A1(n6865), .A2(n4690), .ZN(n4689) );
  INV_X1 U5052 ( .A(n6870), .ZN(n4690) );
  INV_X1 U5053 ( .A(n7598), .ZN(n4570) );
  INV_X1 U5054 ( .A(n4573), .ZN(n4569) );
  OR2_X1 U5055 ( .A1(n7975), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5056 ( .A1(n4681), .A2(n4679), .ZN(n5797) );
  INV_X1 U5057 ( .A(n4680), .ZN(n4679) );
  OAI21_X1 U5058 ( .B1(n9718), .B2(n4283), .A(n5802), .ZN(n4680) );
  NOR2_X1 U5059 ( .A1(n4567), .A2(n4571), .ZN(n4566) );
  AND2_X1 U5060 ( .A1(n7596), .A2(n7597), .ZN(n4571) );
  INV_X1 U5061 ( .A(n4576), .ZN(n4567) );
  NOR2_X1 U5062 ( .A1(n4579), .A2(n4582), .ZN(n4576) );
  AND2_X1 U5063 ( .A1(n7967), .A2(n4580), .ZN(n4579) );
  INV_X1 U5064 ( .A(n7966), .ZN(n4580) );
  AND2_X1 U5065 ( .A1(n4574), .A2(n4573), .ZN(n4572) );
  NAND2_X1 U5066 ( .A1(n7596), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U5067 ( .A1(n6946), .A2(n4503), .ZN(n7160) );
  OR2_X1 U5068 ( .A1(n7091), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4503) );
  NOR2_X1 U5069 ( .A1(n8093), .A2(n8092), .ZN(n8090) );
  XNOR2_X1 U5070 ( .A(n4510), .B(n7180), .ZN(n8103) );
  OR2_X1 U5071 ( .A1(n8090), .A2(n4511), .ZN(n4510) );
  AND2_X1 U5072 ( .A1(n7213), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4511) );
  NOR2_X1 U5073 ( .A1(n8176), .A2(n4669), .ZN(n4668) );
  INV_X1 U5074 ( .A(n7478), .ZN(n4669) );
  XNOR2_X1 U5075 ( .A(n8428), .B(n7625), .ZN(n8176) );
  NOR2_X1 U5076 ( .A1(n8440), .A2(n8232), .ZN(n4372) );
  AOI21_X1 U5077 ( .B1(n4818), .B2(n4816), .A(n4309), .ZN(n4815) );
  INV_X1 U5078 ( .A(n4820), .ZN(n4816) );
  INV_X1 U5079 ( .A(n4818), .ZN(n4817) );
  OR2_X1 U5080 ( .A1(n8239), .A2(n8443), .ZN(n8221) );
  NOR2_X1 U5081 ( .A1(n8246), .A2(n4821), .ZN(n4820) );
  INV_X1 U5082 ( .A(n4824), .ZN(n4821) );
  AND2_X1 U5083 ( .A1(n7369), .A2(n8229), .ZN(n8246) );
  AND2_X1 U5084 ( .A1(n8458), .A2(n8297), .ZN(n4796) );
  AND2_X1 U5085 ( .A1(n4651), .A2(n7460), .ZN(n4373) );
  NAND2_X1 U5086 ( .A1(n4274), .A2(n4653), .ZN(n4651) );
  OR2_X1 U5087 ( .A1(n8318), .A2(n8470), .ZN(n8309) );
  NOR2_X1 U5088 ( .A1(n8309), .A2(n8463), .ZN(n8290) );
  NAND2_X1 U5089 ( .A1(n8302), .A2(n4333), .ZN(n8289) );
  AOI21_X2 U5090 ( .B1(n8336), .B2(n8334), .A(n8335), .ZN(n8341) );
  OR2_X1 U5091 ( .A1(n8483), .A2(n8061), .ZN(n8334) );
  AND2_X1 U5092 ( .A1(n8483), .A2(n8385), .ZN(n4837) );
  NAND2_X1 U5093 ( .A1(n4835), .A2(n4834), .ZN(n4831) );
  INV_X1 U5094 ( .A(n8351), .ZN(n4835) );
  INV_X1 U5095 ( .A(n4831), .ZN(n8353) );
  AND4_X1 U5096 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n8403)
         );
  NOR2_X1 U5097 ( .A1(n7030), .A2(n9493), .ZN(n8392) );
  AND2_X1 U5098 ( .A1(n9807), .A2(n9854), .ZN(n9805) );
  NOR2_X1 U5099 ( .A1(n6289), .A2(n7408), .ZN(n9807) );
  NAND2_X1 U5100 ( .A1(n4839), .A2(n4838), .ZN(n6287) );
  NAND2_X1 U5101 ( .A1(n6280), .A2(n4307), .ZN(n4838) );
  INV_X1 U5102 ( .A(n4675), .ZN(n4674) );
  OAI21_X1 U5103 ( .B1(n7359), .B2(n6193), .A(n6192), .ZN(n4675) );
  NAND2_X1 U5104 ( .A1(n4844), .A2(n4845), .ZN(n6276) );
  NAND2_X1 U5105 ( .A1(n6027), .A2(n4846), .ZN(n4844) );
  NAND2_X1 U5106 ( .A1(n8155), .A2(n8161), .ZN(n8154) );
  NAND2_X1 U5107 ( .A1(n7254), .A2(n7253), .ZN(n8453) );
  XNOR2_X1 U5108 ( .A(n5194), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U5109 ( .A1(n4708), .A2(n4707), .ZN(n5192) );
  AND2_X1 U5110 ( .A1(n4709), .A2(n4316), .ZN(n4707) );
  NAND2_X1 U5111 ( .A1(n4371), .A2(n4370), .ZN(n5161) );
  INV_X1 U5112 ( .A(n4951), .ZN(n4371) );
  INV_X1 U5113 ( .A(n4476), .ZN(n4475) );
  OAI21_X1 U5114 ( .B1(n5945), .B2(n6107), .A(n6108), .ZN(n4476) );
  NAND2_X1 U5115 ( .A1(n4486), .A2(n4275), .ZN(n4857) );
  INV_X1 U5116 ( .A(n8646), .ZN(n4486) );
  INV_X1 U5117 ( .A(n7820), .ZN(n7637) );
  NAND2_X1 U5118 ( .A1(n7674), .A2(n4496), .ZN(n4492) );
  NOR2_X1 U5119 ( .A1(n4850), .A2(n8556), .ZN(n8613) );
  AND2_X1 U5120 ( .A1(n8555), .A2(n8558), .ZN(n4850) );
  AOI21_X1 U5121 ( .B1(n6178), .B2(n5357), .A(n4881), .ZN(n5358) );
  OAI21_X1 U5122 ( .B1(n8642), .B2(n8646), .A(n8565), .ZN(n8623) );
  INV_X1 U5123 ( .A(n5353), .ZN(n5352) );
  NOR2_X1 U5124 ( .A1(n7835), .A2(n4852), .ZN(n4851) );
  OR2_X1 U5125 ( .A1(n8902), .A2(n4324), .ZN(n4363) );
  NOR2_X1 U5126 ( .A1(n4429), .A2(n4428), .ZN(n4427) );
  INV_X1 U5127 ( .A(n8901), .ZN(n4429) );
  AND2_X1 U5128 ( .A1(n7805), .A2(n7804), .ZN(n9088) );
  NAND2_X1 U5129 ( .A1(n8748), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U5130 ( .A1(n5306), .A2(n5001), .ZN(n9026) );
  AND2_X1 U5131 ( .A1(n4606), .A2(n4605), .ZN(n4604) );
  AND2_X1 U5132 ( .A1(n8931), .A2(n8930), .ZN(n9118) );
  OR2_X1 U5133 ( .A1(n9094), .A2(n9173), .ZN(n9166) );
  NAND2_X1 U5134 ( .A1(n9166), .A2(n8932), .ZN(n9188) );
  INV_X1 U5135 ( .A(n9108), .ZN(n4619) );
  NAND2_X1 U5136 ( .A1(n4391), .A2(n4278), .ZN(n4739) );
  AND2_X1 U5137 ( .A1(n4739), .A2(n4737), .ZN(n9241) );
  NOR2_X1 U5138 ( .A1(n9243), .A2(n4738), .ZN(n4737) );
  INV_X1 U5139 ( .A(n9087), .ZN(n4738) );
  NAND2_X1 U5140 ( .A1(n4393), .A2(n4392), .ZN(n4391) );
  NAND2_X1 U5141 ( .A1(n9291), .A2(n9085), .ZN(n4392) );
  NAND2_X1 U5142 ( .A1(n9299), .A2(n4302), .ZN(n4629) );
  NAND2_X1 U5143 ( .A1(n4631), .A2(n9104), .ZN(n4630) );
  NAND2_X1 U5144 ( .A1(n4714), .A2(n9294), .ZN(n4713) );
  INV_X1 U5145 ( .A(n4715), .ZN(n4714) );
  NAND2_X1 U5146 ( .A1(n9350), .A2(n4295), .ZN(n4711) );
  NAND2_X1 U5147 ( .A1(n9350), .A2(n4716), .ZN(n4712) );
  NAND2_X1 U5148 ( .A1(n9325), .A2(n9102), .ZN(n9299) );
  AND2_X1 U5149 ( .A1(n9299), .A2(n9298), .ZN(n9301) );
  NAND2_X1 U5150 ( .A1(n4390), .A2(n4388), .ZN(n4742) );
  NOR2_X1 U5151 ( .A1(n4338), .A2(n4389), .ZN(n4388) );
  INV_X1 U5152 ( .A(n6904), .ZN(n4389) );
  AND2_X1 U5153 ( .A1(n9336), .A2(n9337), .ZN(n8955) );
  AOI21_X1 U5154 ( .B1(n4731), .B2(n4734), .A(n4334), .ZN(n4729) );
  NAND2_X1 U5155 ( .A1(n6498), .A2(n6497), .ZN(n6674) );
  NAND2_X1 U5156 ( .A1(n6554), .A2(n6510), .ZN(n6537) );
  NAND2_X1 U5157 ( .A1(n6552), .A2(n4304), .ZN(n6534) );
  NAND2_X1 U5158 ( .A1(n6553), .A2(n8944), .ZN(n6552) );
  INV_X1 U5159 ( .A(n9282), .ZN(n9343) );
  INV_X1 U5160 ( .A(n9345), .ZN(n9329) );
  AND2_X1 U5161 ( .A1(n9389), .A2(n9456), .ZN(n4375) );
  INV_X1 U5162 ( .A(n4361), .ZN(n4360) );
  NAND2_X1 U5163 ( .A1(n7736), .A2(n7735), .ZN(n9436) );
  NAND2_X1 U5164 ( .A1(n7698), .A2(n7697), .ZN(n9448) );
  INV_X1 U5165 ( .A(n6565), .ZN(n9682) );
  INV_X1 U5166 ( .A(n9694), .ZN(n9456) );
  INV_X1 U5167 ( .A(n7357), .ZN(n4765) );
  AND2_X1 U5168 ( .A1(n7353), .A2(n4765), .ZN(n4764) );
  OR2_X1 U5169 ( .A1(n7350), .A2(n7349), .ZN(n7354) );
  NAND2_X1 U5170 ( .A1(n4763), .A2(n7357), .ZN(n4762) );
  INV_X1 U5171 ( .A(n7353), .ZN(n4763) );
  XNOR2_X1 U5172 ( .A(n7350), .B(SI_30_), .ZN(n8744) );
  XNOR2_X1 U5173 ( .A(n7313), .B(n7312), .ZN(n7878) );
  XNOR2_X1 U5174 ( .A(n4930), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5241) );
  OAI21_X1 U5175 ( .B1(n6689), .B2(n6688), .A(n6690), .ZN(n6845) );
  OAI21_X1 U5176 ( .B1(n5412), .B2(n4280), .A(n4780), .ZN(n5689) );
  NAND2_X1 U5177 ( .A1(n4783), .A2(n5651), .ZN(n5668) );
  NAND2_X1 U5178 ( .A1(n5412), .A2(n4784), .ZN(n4783) );
  NAND2_X1 U5179 ( .A1(n5412), .A2(n5411), .ZN(n5653) );
  OAI21_X1 U5180 ( .B1(n5174), .B2(n4281), .A(n4458), .ZN(n5410) );
  OAI211_X1 U5181 ( .C1(n4645), .C2(n4588), .A(n4586), .B(n5090), .ZN(n5095)
         );
  INV_X1 U5182 ( .A(n4648), .ZN(n4647) );
  NAND2_X1 U5183 ( .A1(n4464), .A2(SI_4_), .ZN(n5068) );
  INV_X1 U5184 ( .A(n5067), .ZN(n4464) );
  XNOR2_X1 U5185 ( .A(n5080), .B(SI_5_), .ZN(n5078) );
  XNOR2_X1 U5186 ( .A(n5067), .B(SI_4_), .ZN(n5065) );
  NAND2_X1 U5187 ( .A1(n5047), .A2(n5046), .ZN(n5050) );
  NAND2_X1 U5188 ( .A1(n5055), .A2(n5054), .ZN(n5047) );
  XNOR2_X1 U5189 ( .A(n7598), .B(n7597), .ZN(n7933) );
  NAND2_X1 U5190 ( .A1(n8035), .A2(n5775), .ZN(n9719) );
  NAND2_X1 U5191 ( .A1(n5797), .A2(n5798), .ZN(n7989) );
  NAND2_X1 U5192 ( .A1(n7989), .A2(n7988), .ZN(n7987) );
  AND3_X1 U5193 ( .A1(n7270), .A2(n7269), .A3(n7268), .ZN(n8268) );
  NAND2_X1 U5194 ( .A1(n7224), .A2(n7223), .ZN(n8473) );
  OR2_X1 U5195 ( .A1(n4753), .A2(n7538), .ZN(n4751) );
  AND2_X1 U5196 ( .A1(n7540), .A2(n7539), .ZN(n4753) );
  AOI21_X1 U5197 ( .B1(n7542), .B2(n7541), .A(n7549), .ZN(n4750) );
  INV_X1 U5198 ( .A(n7548), .ZN(n4749) );
  XNOR2_X1 U5199 ( .A(n4644), .B(n4643), .ZN(n4642) );
  OAI21_X1 U5200 ( .B1(n7363), .B2(n7364), .A(n7498), .ZN(n4644) );
  OR2_X1 U5201 ( .A1(n5788), .A2(n4410), .ZN(n4693) );
  INV_X1 U5202 ( .A(n4692), .ZN(n4691) );
  OAI211_X1 U5203 ( .C1(n8154), .C2(n8141), .A(n4804), .B(n4802), .ZN(n8422)
         );
  NAND2_X1 U5204 ( .A1(n8140), .A2(n4267), .ZN(n4804) );
  NAND2_X1 U5205 ( .A1(n8154), .A2(n4803), .ZN(n4802) );
  NOR2_X1 U5206 ( .A1(n8140), .A2(n4267), .ZN(n4803) );
  INV_X1 U5207 ( .A(n4369), .ZN(n4368) );
  OAI21_X1 U5208 ( .B1(n8419), .B2(n9865), .A(n4562), .ZN(n4369) );
  NOR2_X1 U5209 ( .A1(n4808), .A2(n4797), .ZN(n4562) );
  INV_X1 U5210 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4807) );
  AOI21_X1 U5211 ( .B1(n4289), .B2(n4490), .A(n4488), .ZN(n4487) );
  NOR2_X1 U5212 ( .A1(n7075), .A2(n7074), .ZN(n4488) );
  NOR2_X1 U5213 ( .A1(n8549), .A2(n8545), .ZN(n7911) );
  NAND2_X1 U5214 ( .A1(n6935), .A2(n6934), .ZN(n6936) );
  NAND2_X1 U5215 ( .A1(n6241), .A2(n6240), .ZN(n6529) );
  NAND2_X1 U5216 ( .A1(n7757), .A2(n7756), .ZN(n9430) );
  INV_X1 U5217 ( .A(n9231), .ZN(n9420) );
  INV_X1 U5218 ( .A(n9088), .ZN(n9251) );
  NOR2_X1 U5219 ( .A1(n5034), .A2(n4351), .ZN(n5033) );
  INV_X1 U5220 ( .A(n4635), .ZN(n4634) );
  OAI21_X1 U5221 ( .B1(n9139), .B2(n9140), .A(n9348), .ZN(n4636) );
  OAI22_X1 U5222 ( .A1(n9172), .A2(n9282), .B1(n9141), .B2(n9345), .ZN(n4635)
         );
  NAND2_X1 U5223 ( .A1(n9133), .A2(n4294), .ZN(n9394) );
  OAI21_X1 U5224 ( .B1(n9199), .B2(n4724), .A(n4723), .ZN(n9165) );
  OAI21_X1 U5225 ( .B1(n9379), .B2(n9694), .A(n9382), .ZN(n4611) );
  NAND2_X1 U5226 ( .A1(n4528), .A2(n4532), .ZN(n4527) );
  INV_X1 U5227 ( .A(n7464), .ZN(n4526) );
  INV_X1 U5228 ( .A(n7466), .ZN(n4519) );
  NAND2_X1 U5229 ( .A1(n4522), .A2(n4520), .ZN(n4523) );
  NAND2_X1 U5230 ( .A1(n9137), .A2(n4453), .ZN(n4452) );
  INV_X1 U5231 ( .A(n8880), .ZN(n4453) );
  INV_X1 U5232 ( .A(n4774), .ZN(n4773) );
  NAND2_X1 U5233 ( .A1(n4776), .A2(n4770), .ZN(n4769) );
  INV_X1 U5234 ( .A(n7343), .ZN(n4770) );
  NOR2_X1 U5235 ( .A1(n4773), .A2(n7343), .ZN(n4772) );
  INV_X1 U5236 ( .A(n6201), .ZN(n7512) );
  NOR2_X1 U5237 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4895) );
  NAND2_X1 U5238 ( .A1(n4771), .A2(n4767), .ZN(n7352) );
  INV_X1 U5239 ( .A(n4768), .ZN(n4767) );
  NAND2_X1 U5240 ( .A1(n7315), .A2(n4772), .ZN(n4771) );
  OAI21_X1 U5241 ( .B1(n4773), .B2(n4769), .A(n7342), .ZN(n4768) );
  INV_X1 U5242 ( .A(n7146), .ZN(n4788) );
  NOR2_X1 U5243 ( .A1(n4747), .A2(n4746), .ZN(n4745) );
  INV_X1 U5244 ( .A(n6371), .ZN(n4746) );
  INV_X1 U5245 ( .A(n6593), .ZN(n4747) );
  INV_X1 U5246 ( .A(n5974), .ZN(n4435) );
  INV_X1 U5247 ( .A(n4443), .ZN(n4442) );
  OAI21_X1 U5248 ( .B1(n5115), .B2(n4444), .A(n4883), .ZN(n4443) );
  INV_X1 U5249 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4892) );
  NOR2_X1 U5250 ( .A1(n4283), .A2(n4683), .ZN(n4682) );
  AND2_X1 U5251 ( .A1(n7581), .A2(n7583), .ZN(n7589) );
  XNOR2_X1 U5252 ( .A(n7946), .B(n7607), .ZN(n5771) );
  NAND2_X1 U5253 ( .A1(n8188), .A2(n8216), .ZN(n4539) );
  NAND2_X1 U5254 ( .A1(n4561), .A2(n8261), .ZN(n4560) );
  INV_X1 U5255 ( .A(n8295), .ZN(n4658) );
  OR2_X1 U5256 ( .A1(n7233), .A2(n5423), .ZN(n7241) );
  OR2_X1 U5257 ( .A1(n8473), .A2(n8307), .ZN(n7457) );
  NOR2_X1 U5258 ( .A1(n8480), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U5259 ( .A1(n7009), .A2(n7428), .ZN(n4661) );
  NOR2_X1 U5260 ( .A1(n7435), .A2(n4662), .ZN(n4664) );
  OR2_X1 U5261 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  INV_X1 U5262 ( .A(n4845), .ZN(n4843) );
  NOR2_X1 U5263 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  INV_X1 U5264 ( .A(n4846), .ZN(n4841) );
  INV_X1 U5265 ( .A(n6280), .ZN(n4842) );
  OR2_X1 U5266 ( .A1(n9844), .A2(n6306), .ZN(n4846) );
  NAND2_X1 U5267 ( .A1(n9844), .A2(n6306), .ZN(n4845) );
  OR2_X1 U5268 ( .A1(n8421), .A2(n7623), .ZN(n7366) );
  NAND2_X1 U5269 ( .A1(n4665), .A2(n4670), .ZN(n7338) );
  AOI21_X1 U5270 ( .B1(n7529), .B2(n4672), .A(n4671), .ZN(n4670) );
  INV_X1 U5271 ( .A(n7481), .ZN(n4672) );
  NOR2_X1 U5272 ( .A1(n8221), .A2(n8440), .ZN(n8212) );
  NOR2_X1 U5273 ( .A1(n4945), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U5274 ( .A1(n4498), .A2(n4497), .ZN(n4496) );
  INV_X1 U5275 ( .A(n7673), .ZN(n4497) );
  NOR2_X1 U5276 ( .A1(n4498), .A2(n4495), .ZN(n4494) );
  INV_X1 U5277 ( .A(n8673), .ZN(n4495) );
  AND2_X1 U5278 ( .A1(n8605), .A2(n4499), .ZN(n4498) );
  INV_X1 U5279 ( .A(n7695), .ZN(n4499) );
  AND2_X1 U5280 ( .A1(n8605), .A2(n8592), .ZN(n4500) );
  INV_X1 U5281 ( .A(n4481), .ZN(n4480) );
  INV_X1 U5282 ( .A(n6441), .ZN(n4482) );
  INV_X1 U5283 ( .A(n8558), .ZN(n4852) );
  OR2_X1 U5284 ( .A1(n8612), .A2(n7835), .ZN(n4854) );
  NOR2_X1 U5285 ( .A1(n9568), .A2(n4345), .ZN(n9037) );
  NOR2_X1 U5286 ( .A1(n9622), .A2(n9623), .ZN(n9624) );
  INV_X1 U5287 ( .A(n5494), .ZN(n5356) );
  NOR2_X1 U5288 ( .A1(n9393), .A2(n4607), .ZN(n4606) );
  INV_X1 U5289 ( .A(n4608), .ZN(n4607) );
  OR2_X1 U5290 ( .A1(n9389), .A2(n9141), .ZN(n8931) );
  OR2_X1 U5291 ( .A1(n9393), .A2(n9157), .ZN(n8881) );
  AND2_X1 U5292 ( .A1(n9402), .A2(n9095), .ZN(n9114) );
  NAND2_X1 U5293 ( .A1(n9138), .A2(n8879), .ZN(n9116) );
  AND2_X1 U5294 ( .A1(n8932), .A2(n9184), .ZN(n9113) );
  NOR2_X1 U5295 ( .A1(n9411), .A2(n4600), .ZN(n4599) );
  INV_X1 U5296 ( .A(n4601), .ZN(n4600) );
  AND2_X1 U5297 ( .A1(n4602), .A2(n9217), .ZN(n4601) );
  NOR2_X1 U5298 ( .A1(n9420), .A2(n9426), .ZN(n4602) );
  OR2_X1 U5299 ( .A1(n7701), .A2(n7700), .ZN(n7719) );
  AND2_X1 U5300 ( .A1(n4731), .A2(n4396), .ZN(n4395) );
  NAND2_X1 U5301 ( .A1(n4398), .A2(n4400), .ZN(n4396) );
  AND2_X1 U5302 ( .A1(n6756), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U5303 ( .A1(n4733), .A2(n6605), .ZN(n4732) );
  INV_X1 U5304 ( .A(n4735), .ZN(n4733) );
  INV_X1 U5305 ( .A(n6605), .ZN(n4734) );
  INV_X1 U5306 ( .A(n7063), .ZN(n4791) );
  INV_X1 U5307 ( .A(n4790), .ZN(n4789) );
  OAI21_X1 U5308 ( .B1(n4793), .B2(n4344), .A(n7116), .ZN(n4790) );
  NOR2_X1 U5309 ( .A1(n5975), .A2(n4437), .ZN(n4436) );
  INV_X1 U5310 ( .A(n5690), .ZN(n4437) );
  INV_X1 U5311 ( .A(n5651), .ZN(n4782) );
  NOR2_X1 U5312 ( .A1(n5652), .A2(n4785), .ZN(n4784) );
  INV_X1 U5313 ( .A(n5411), .ZN(n4785) );
  AND3_X1 U5314 ( .A1(n4897), .A2(n4878), .A3(n4268), .ZN(n5297) );
  INV_X1 U5315 ( .A(n5211), .ZN(n4460) );
  INV_X1 U5316 ( .A(n4459), .ZN(n4458) );
  OAI21_X1 U5317 ( .B1(n4462), .B2(n4281), .A(n5292), .ZN(n4459) );
  NAND2_X1 U5318 ( .A1(n5100), .A2(n5099), .ZN(n5117) );
  NAND2_X1 U5319 ( .A1(n5095), .A2(n5094), .ZN(n5116) );
  AND2_X1 U5320 ( .A1(n4647), .A2(n5086), .ZN(n4585) );
  CLKBUF_X1 U5321 ( .A(n4966), .Z(n4967) );
  OAI21_X1 U5322 ( .B1(n7333), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n4362), .ZN(
        n5088) );
  NAND2_X1 U5323 ( .A1(n7333), .A2(n9976), .ZN(n4362) );
  OR2_X1 U5324 ( .A1(n7256), .A2(n5425), .ZN(n7264) );
  NAND2_X1 U5325 ( .A1(n4590), .A2(n4589), .ZN(n7956) );
  INV_X1 U5326 ( .A(n7587), .ZN(n4589) );
  OR2_X1 U5327 ( .A1(n8018), .A2(n4591), .ZN(n4590) );
  INV_X1 U5328 ( .A(n8016), .ZN(n4591) );
  NOR2_X1 U5329 ( .A1(n7582), .A2(n4702), .ZN(n4701) );
  INV_X1 U5330 ( .A(n7575), .ZN(n4702) );
  OR2_X1 U5331 ( .A1(n7954), .A2(n7589), .ZN(n7582) );
  NOR2_X1 U5332 ( .A1(n7588), .A2(n7589), .ZN(n7591) );
  AND2_X1 U5333 ( .A1(n7958), .A2(n7956), .ZN(n7588) );
  AND3_X1 U5334 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5991) );
  AOI21_X1 U5335 ( .B1(n7502), .B2(n7501), .A(n7500), .ZN(n7537) );
  AND4_X1 U5336 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n6976)
         );
  AND4_X1 U5337 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n6975)
         );
  AND2_X1 U5338 ( .A1(n6435), .A2(n4515), .ZN(n6388) );
  NAND2_X1 U5339 ( .A1(n6426), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5340 ( .A1(n6635), .A2(n4513), .ZN(n6636) );
  OR2_X1 U5341 ( .A1(n6872), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5342 ( .A1(n7163), .A2(n7162), .ZN(n8079) );
  INV_X1 U5343 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5681) );
  NOR2_X1 U5344 ( .A1(n8077), .A2(n4512), .ZN(n8093) );
  AND2_X1 U5345 ( .A1(n8082), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4512) );
  INV_X1 U5346 ( .A(n4764), .ZN(n4759) );
  AND2_X1 U5347 ( .A1(n4762), .A2(n4765), .ZN(n4761) );
  OR2_X1 U5348 ( .A1(n8146), .A2(n8421), .ZN(n8147) );
  AND2_X1 U5349 ( .A1(n4810), .A2(n4349), .ZN(n4809) );
  OR2_X1 U5350 ( .A1(n8145), .A2(n8402), .ZN(n4810) );
  NAND2_X1 U5351 ( .A1(n8168), .A2(n8139), .ZN(n8155) );
  NAND2_X1 U5352 ( .A1(n8434), .A2(n8211), .ZN(n7478) );
  NOR2_X1 U5353 ( .A1(n8221), .A2(n4539), .ZN(n8195) );
  NOR2_X1 U5354 ( .A1(n8221), .A2(n4538), .ZN(n8171) );
  NAND2_X1 U5355 ( .A1(n8184), .A2(n4357), .ZN(n8169) );
  NAND2_X1 U5356 ( .A1(n8188), .A2(n8211), .ZN(n4357) );
  OR2_X1 U5357 ( .A1(n8440), .A2(n8192), .ZN(n8138) );
  OR2_X1 U5358 ( .A1(n8453), .A2(n8060), .ZN(n8244) );
  AND2_X1 U5359 ( .A1(n8263), .A2(n8264), .ZN(n4640) );
  NOR2_X1 U5360 ( .A1(n8309), .A2(n4559), .ZN(n8275) );
  INV_X1 U5361 ( .A(n4561), .ZN(n4559) );
  AND2_X1 U5362 ( .A1(n7464), .A2(n8264), .ZN(n8281) );
  NAND2_X1 U5363 ( .A1(n8289), .A2(n8295), .ZN(n8288) );
  INV_X1 U5364 ( .A(n4657), .ZN(n4656) );
  OAI21_X1 U5365 ( .B1(n7503), .B2(n7222), .A(n7457), .ZN(n4657) );
  NAND2_X1 U5366 ( .A1(n8341), .A2(n8325), .ZN(n4655) );
  OR2_X1 U5367 ( .A1(n8393), .A2(n4550), .ZN(n8318) );
  NAND2_X1 U5368 ( .A1(n4551), .A2(n8323), .ZN(n4550) );
  NOR2_X1 U5369 ( .A1(n8393), .A2(n4549), .ZN(n8342) );
  INV_X1 U5370 ( .A(n4551), .ZN(n4549) );
  NAND2_X1 U5371 ( .A1(n4827), .A2(n4829), .ZN(n8317) );
  INV_X1 U5372 ( .A(n4830), .ZN(n4829) );
  OAI22_X1 U5373 ( .A1(n4832), .A2(n4834), .B1(n8480), .B2(n8326), .ZN(n4830)
         );
  NOR2_X1 U5374 ( .A1(n8393), .A2(n4552), .ZN(n8364) );
  NAND2_X1 U5375 ( .A1(n8128), .A2(n4303), .ZN(n8131) );
  NAND2_X1 U5376 ( .A1(n4358), .A2(n8128), .ZN(n4811) );
  NAND2_X1 U5377 ( .A1(n7023), .A2(n4664), .ZN(n7208) );
  AND4_X1 U5378 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n7024)
         );
  NAND2_X1 U5379 ( .A1(n6986), .A2(n7520), .ZN(n7023) );
  OR2_X1 U5380 ( .A1(n9766), .A2(n8501), .ZN(n7030) );
  INV_X1 U5381 ( .A(n4556), .ZN(n4555) );
  NOR2_X1 U5382 ( .A1(n4554), .A2(n5937), .ZN(n4553) );
  AND2_X1 U5383 ( .A1(n6201), .A2(n4676), .ZN(n6198) );
  NOR2_X1 U5384 ( .A1(n5937), .A2(n4556), .ZN(n6033) );
  NAND2_X1 U5385 ( .A1(n6033), .A2(n7401), .ZN(n6211) );
  NAND2_X1 U5386 ( .A1(n6007), .A2(n6006), .ZN(n6027) );
  OR2_X1 U5387 ( .A1(n5935), .A2(n9722), .ZN(n5937) );
  NOR2_X1 U5388 ( .A1(n5937), .A2(n6012), .ZN(n6000) );
  NAND2_X1 U5389 ( .A1(n7378), .A2(n7376), .ZN(n5745) );
  INV_X1 U5390 ( .A(n8402), .ZN(n9778) );
  NAND2_X1 U5391 ( .A1(n4795), .A2(n5736), .ZN(n5735) );
  INV_X1 U5392 ( .A(n9775), .ZN(n8404) );
  INV_X1 U5393 ( .A(n4809), .ZN(n4797) );
  AND2_X1 U5394 ( .A1(n8421), .A2(n9876), .ZN(n4808) );
  NAND2_X1 U5395 ( .A1(n6286), .A2(n6285), .ZN(n7408) );
  INV_X1 U5396 ( .A(n9876), .ZN(n9863) );
  NOR2_X1 U5397 ( .A1(n4848), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U5398 ( .A1(n4316), .A2(n5159), .ZN(n4848) );
  NAND2_X1 U5399 ( .A1(n4826), .A2(n4942), .ZN(n5472) );
  INV_X1 U5400 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5219) );
  INV_X1 U5401 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U5402 ( .A1(n7636), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7820) );
  INV_X1 U5403 ( .A(n7799), .ZN(n7636) );
  INV_X1 U5404 ( .A(n5355), .ZN(n4471) );
  NAND2_X1 U5405 ( .A1(n5513), .A2(n5512), .ZN(n5516) );
  AND2_X1 U5406 ( .A1(n8622), .A2(n7753), .ZN(n8565) );
  NOR2_X1 U5407 ( .A1(n5861), .A2(n5860), .ZN(n5958) );
  AND2_X1 U5408 ( .A1(n4856), .A2(n4860), .ZN(n4855) );
  INV_X1 U5409 ( .A(n8572), .ZN(n4856) );
  NAND2_X1 U5410 ( .A1(n4861), .A2(n7773), .ZN(n4860) );
  INV_X1 U5411 ( .A(n9186), .ZN(n9095) );
  NAND2_X1 U5412 ( .A1(n4872), .A2(n4871), .ZN(n6442) );
  OR2_X1 U5413 ( .A1(n7738), .A2(n7737), .ZN(n7759) );
  INV_X1 U5414 ( .A(n8622), .ZN(n4865) );
  NAND2_X1 U5415 ( .A1(n4864), .A2(n4862), .ZN(n4861) );
  INV_X1 U5416 ( .A(n8621), .ZN(n4864) );
  NAND2_X1 U5417 ( .A1(n4863), .A2(n8622), .ZN(n4862) );
  INV_X1 U5418 ( .A(n8565), .ZN(n4863) );
  OR2_X1 U5419 ( .A1(n6613), .A2(n6612), .ZN(n6764) );
  INV_X1 U5420 ( .A(n4873), .ZN(n4491) );
  AOI21_X1 U5421 ( .B1(n4873), .B2(n6676), .A(n4298), .ZN(n4490) );
  OR2_X1 U5422 ( .A1(n7797), .A2(n8635), .ZN(n7799) );
  OR2_X1 U5423 ( .A1(n6262), .A2(n10031), .ZN(n6458) );
  NAND2_X1 U5424 ( .A1(n8603), .A2(n7714), .ZN(n7731) );
  NAND2_X1 U5425 ( .A1(n4869), .A2(n4868), .ZN(n4867) );
  INV_X1 U5426 ( .A(n8605), .ZN(n4868) );
  NOR2_X1 U5427 ( .A1(n6764), .A2(n6763), .ZN(n6912) );
  NAND2_X1 U5428 ( .A1(n5280), .A2(n9015), .ZN(n5279) );
  OR2_X1 U5429 ( .A1(n5558), .A2(n5557), .ZN(n4413) );
  AND2_X1 U5430 ( .A1(n4413), .A2(n4412), .ZN(n5307) );
  NAND2_X1 U5431 ( .A1(n5018), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U5432 ( .A1(n5307), .A2(n5308), .ZN(n5306) );
  INV_X1 U5433 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10031) );
  INV_X1 U5434 ( .A(n5033), .ZN(n5004) );
  NOR2_X1 U5435 ( .A1(n5443), .A2(n4415), .ZN(n5573) );
  AND2_X1 U5436 ( .A1(n6444), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U5437 ( .A1(n5573), .A2(n5574), .ZN(n5572) );
  NAND2_X1 U5438 ( .A1(n5572), .A2(n4414), .ZN(n5446) );
  OR2_X1 U5439 ( .A1(n6496), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4414) );
  XNOR2_X1 U5440 ( .A(n9037), .B(n6905), .ZN(n5918) );
  XNOR2_X1 U5441 ( .A(n9040), .B(n9052), .ZN(n9585) );
  NOR2_X1 U5442 ( .A1(n9585), .A2(n7055), .ZN(n9584) );
  NOR2_X1 U5443 ( .A1(n9607), .A2(n4421), .ZN(n9622) );
  AND2_X1 U5444 ( .A1(n9610), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4421) );
  XNOR2_X1 U5445 ( .A(n4419), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9061) );
  OR2_X1 U5446 ( .A1(n9624), .A2(n4420), .ZN(n4419) );
  AND2_X1 U5447 ( .A1(n9627), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4420) );
  NAND2_X1 U5448 ( .A1(n8747), .A2(n8746), .ZN(n9077) );
  NAND2_X1 U5449 ( .A1(n8881), .A2(n9117), .ZN(n9134) );
  INV_X1 U5450 ( .A(n9116), .ZN(n9153) );
  OR2_X1 U5451 ( .A1(n4719), .A2(n4382), .ZN(n4379) );
  NOR2_X1 U5452 ( .A1(n4721), .A2(n4383), .ZN(n4382) );
  NAND2_X1 U5453 ( .A1(n4272), .A2(n9093), .ZN(n4724) );
  NAND2_X1 U5454 ( .A1(n4726), .A2(n4272), .ZN(n4723) );
  AND2_X1 U5455 ( .A1(n8933), .A2(n9184), .ZN(n9206) );
  NAND2_X1 U5456 ( .A1(n9264), .A2(n9260), .ZN(n9253) );
  NAND2_X1 U5457 ( .A1(n9264), .A2(n4602), .ZN(n9228) );
  NAND2_X1 U5458 ( .A1(n7635), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7779) );
  INV_X1 U5459 ( .A(n7759), .ZN(n7635) );
  OR2_X1 U5460 ( .A1(n7779), .A2(n8574), .ZN(n7797) );
  AOI21_X1 U5461 ( .B1(n4627), .B2(n8817), .A(n4625), .ZN(n4624) );
  INV_X1 U5462 ( .A(n4627), .ZN(n4626) );
  INV_X1 U5463 ( .A(n9101), .ZN(n4625) );
  OR2_X1 U5464 ( .A1(n9323), .A2(n9324), .ZN(n9325) );
  NAND2_X1 U5465 ( .A1(n4614), .A2(n4613), .ZN(n9356) );
  NOR2_X1 U5466 ( .A1(n9356), .A2(n9448), .ZN(n9318) );
  NAND2_X1 U5467 ( .A1(n7043), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7701) );
  AND2_X1 U5468 ( .A1(n6912), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U5469 ( .A1(n7042), .A2(n8814), .ZN(n9339) );
  OR2_X1 U5470 ( .A1(n6910), .A2(n8956), .ZN(n7042) );
  AND2_X1 U5471 ( .A1(n6773), .A2(n9519), .ZN(n6920) );
  OAI21_X1 U5472 ( .B1(n6761), .B2(n6760), .A(n8798), .ZN(n6908) );
  NOR2_X1 U5473 ( .A1(n6458), .A2(n6457), .ZN(n6499) );
  NOR2_X1 U5474 ( .A1(n6623), .A2(n9455), .ZN(n6773) );
  OR2_X1 U5475 ( .A1(n6575), .A2(n6674), .ZN(n6623) );
  OAI211_X1 U5476 ( .C1(n6554), .C2(n4291), .A(n8793), .B(n4622), .ZN(n6571)
         );
  NOR2_X1 U5477 ( .A1(n6542), .A2(n6529), .ZN(n6576) );
  NAND2_X1 U5478 ( .A1(n4612), .A2(n6543), .ZN(n6542) );
  OR2_X1 U5479 ( .A1(n8995), .A2(n9682), .ZN(n8785) );
  NOR2_X1 U5480 ( .A1(n6170), .A2(n6171), .ZN(n6561) );
  NAND2_X1 U5481 ( .A1(n5724), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5861) );
  AND3_X1 U5482 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5724) );
  AND2_X1 U5483 ( .A1(n4710), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U5484 ( .A1(n6165), .A2(n6167), .ZN(n6489) );
  NAND2_X1 U5485 ( .A1(n4350), .A2(n9668), .ZN(n6170) );
  NAND2_X1 U5486 ( .A1(n4598), .A2(n7201), .ZN(n7200) );
  NOR2_X1 U5487 ( .A1(n7200), .A2(n6481), .ZN(n6479) );
  INV_X1 U5488 ( .A(n8940), .ZN(n5588) );
  AND2_X1 U5489 ( .A1(n5493), .A2(n9648), .ZN(n5333) );
  XNOR2_X1 U5490 ( .A(n7344), .B(n7334), .ZN(n8681) );
  OAI21_X1 U5491 ( .B1(n7315), .B2(n4776), .A(n4774), .ZN(n7344) );
  XNOR2_X1 U5492 ( .A(n7330), .B(n7329), .ZN(n7631) );
  NAND2_X1 U5493 ( .A1(n7315), .A2(n7314), .ZN(n7330) );
  XNOR2_X1 U5494 ( .A(n7147), .B(n7146), .ZN(n7856) );
  OAI21_X1 U5495 ( .B1(n6847), .B2(n4344), .A(n4789), .ZN(n7147) );
  NAND2_X1 U5496 ( .A1(n4877), .A2(n4876), .ZN(n4921) );
  AND2_X1 U5497 ( .A1(n4920), .A2(n4317), .ZN(n4876) );
  NAND2_X1 U5498 ( .A1(n4792), .A2(n7063), .ZN(n7118) );
  NAND2_X1 U5499 ( .A1(n6372), .A2(n6371), .ZN(n6592) );
  NAND2_X1 U5500 ( .A1(n5691), .A2(n5690), .ZN(n5976) );
  NAND2_X1 U5501 ( .A1(n4461), .A2(n5211), .ZN(n5291) );
  NAND2_X1 U5502 ( .A1(n5174), .A2(n5173), .ZN(n5213) );
  XNOR2_X1 U5503 ( .A(n4359), .B(n5112), .ZN(n6282) );
  NAND2_X1 U5504 ( .A1(n5116), .A2(n5113), .ZN(n4359) );
  AOI21_X1 U5505 ( .B1(n4647), .B2(n4649), .A(n4311), .ZN(n4645) );
  XNOR2_X1 U5506 ( .A(n5061), .B(SI_3_), .ZN(n5059) );
  XNOR2_X1 U5507 ( .A(n5051), .B(n5048), .ZN(n5049) );
  OAI211_X1 U5508 ( .C1(n4637), .C2(n4410), .A(n4409), .B(n4408), .ZN(n5054)
         );
  NAND2_X1 U5509 ( .A1(n4593), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4409) );
  INV_X1 U5510 ( .A(n7333), .ZN(n7355) );
  AOI21_X1 U5511 ( .B1(n4688), .B2(n4690), .A(n4308), .ZN(n4686) );
  NAND2_X1 U5512 ( .A1(n7093), .A2(n7092), .ZN(n8495) );
  NAND2_X1 U5513 ( .A1(n7263), .A2(n7262), .ZN(n8448) );
  NOR2_X1 U5514 ( .A1(n6344), .A2(n6343), .ZN(n4879) );
  NAND2_X1 U5515 ( .A1(n6347), .A2(n6346), .ZN(n8506) );
  NAND2_X1 U5516 ( .A1(n4703), .A2(n7575), .ZN(n7955) );
  NAND2_X1 U5517 ( .A1(n7619), .A2(n9744), .ZN(n4354) );
  AND4_X1 U5518 ( .A1(n7246), .A2(n7245), .A3(n7244), .A4(n7243), .ZN(n8308)
         );
  AND3_X1 U5519 ( .A1(n7278), .A2(n7277), .A3(n7276), .ZN(n8210) );
  NAND2_X1 U5520 ( .A1(n4570), .A2(n4569), .ZN(n4583) );
  NAND2_X1 U5521 ( .A1(n7933), .A2(n7596), .ZN(n4577) );
  AND4_X1 U5522 ( .A1(n7221), .A2(n7220), .A3(n7219), .A4(n7218), .ZN(n8358)
         );
  NAND2_X1 U5523 ( .A1(n4697), .A2(n7566), .ZN(n7978) );
  NAND2_X1 U5524 ( .A1(n7976), .A2(n7975), .ZN(n4697) );
  OAI21_X1 U5525 ( .B1(n7976), .B2(n4271), .A(n4265), .ZN(n7979) );
  AND4_X1 U5526 ( .A1(n7139), .A2(n7138), .A3(n7137), .A4(n7136), .ZN(n8061)
         );
  NAND2_X1 U5527 ( .A1(n4696), .A2(n4694), .ZN(n7999) );
  AOI21_X1 U5528 ( .B1(n4265), .B2(n4271), .A(n4695), .ZN(n4694) );
  INV_X1 U5529 ( .A(n7567), .ZN(n4695) );
  NOR2_X1 U5530 ( .A1(n7598), .A2(n4575), .ZN(n8005) );
  NAND2_X1 U5531 ( .A1(n7272), .A2(n7271), .ZN(n8443) );
  AND2_X1 U5532 ( .A1(n6335), .A2(n6334), .ZN(n9854) );
  XNOR2_X1 U5533 ( .A(n7586), .B(n7585), .ZN(n8018) );
  NAND2_X1 U5534 ( .A1(n7240), .A2(n7239), .ZN(n8463) );
  NAND2_X1 U5535 ( .A1(n4687), .A2(n6870), .ZN(n7100) );
  NAND2_X1 U5536 ( .A1(n6866), .A2(n6865), .ZN(n4687) );
  NAND2_X1 U5537 ( .A1(n6874), .A2(n6873), .ZN(n9493) );
  AND2_X1 U5538 ( .A1(n8036), .A2(n8034), .ZN(n5774) );
  AND4_X1 U5539 ( .A1(n7238), .A2(n7237), .A3(n7236), .A4(n7235), .ZN(n8135)
         );
  NAND2_X1 U5540 ( .A1(n7987), .A2(n6312), .ZN(n9743) );
  NAND2_X1 U5541 ( .A1(n7601), .A2(n7966), .ZN(n4578) );
  NAND2_X1 U5542 ( .A1(n4572), .A2(n4576), .ZN(n4568) );
  NOR2_X1 U5543 ( .A1(n8051), .A2(n8052), .ZN(n8050) );
  INV_X1 U5544 ( .A(n9724), .ZN(n8021) );
  NAND2_X1 U5545 ( .A1(n7131), .A2(n7130), .ZN(n8490) );
  INV_X1 U5546 ( .A(n9734), .ZN(n9748) );
  NOR2_X1 U5547 ( .A1(n6820), .A2(n6821), .ZN(n6819) );
  NOR2_X1 U5548 ( .A1(n6783), .A2(n6782), .ZN(n6781) );
  NAND2_X1 U5549 ( .A1(n4505), .A2(n4504), .ZN(n6419) );
  NAND2_X1 U5550 ( .A1(n6085), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4504) );
  INV_X1 U5551 ( .A(n6781), .ZN(n4505) );
  NAND2_X1 U5552 ( .A1(n6419), .A2(n6420), .ZN(n6418) );
  NAND2_X1 U5553 ( .A1(n6436), .A2(n6437), .ZN(n6435) );
  OR2_X1 U5554 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  NOR2_X1 U5555 ( .A1(n6808), .A2(n6807), .ZN(n6806) );
  NOR2_X1 U5556 ( .A1(n6891), .A2(n4509), .ZN(n6808) );
  AND2_X1 U5557 ( .A1(n6896), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4509) );
  NOR2_X1 U5558 ( .A1(n6806), .A2(n4508), .ZN(n6071) );
  AND2_X1 U5559 ( .A1(n6812), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U5560 ( .A1(n6071), .A2(n6072), .ZN(n6218) );
  NAND2_X1 U5561 ( .A1(n6223), .A2(n6222), .ZN(n6635) );
  AND2_X1 U5562 ( .A1(n6374), .A2(n4514), .ZN(n6223) );
  NAND2_X1 U5563 ( .A1(n6740), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4514) );
  XNOR2_X1 U5564 ( .A(n7160), .B(n7169), .ZN(n6947) );
  NAND2_X1 U5565 ( .A1(n6947), .A2(n9966), .ZN(n7162) );
  INV_X1 U5566 ( .A(n4826), .ZN(n5977) );
  INV_X1 U5567 ( .A(n4510), .ZN(n7165) );
  NAND2_X1 U5568 ( .A1(n7346), .A2(n7345), .ZN(n8416) );
  NAND2_X1 U5569 ( .A1(n8147), .A2(n4563), .ZN(n8419) );
  OR2_X1 U5570 ( .A1(n4537), .A2(n8150), .ZN(n4563) );
  NAND2_X1 U5571 ( .A1(n4798), .A2(n4809), .ZN(n8420) );
  NAND2_X1 U5572 ( .A1(n4673), .A2(n7481), .ZN(n8162) );
  NAND2_X1 U5573 ( .A1(n8189), .A2(n4668), .ZN(n4673) );
  OAI21_X1 U5574 ( .B1(n8253), .B2(n4817), .A(n4815), .ZN(n8205) );
  NAND2_X1 U5575 ( .A1(n4819), .A2(n4822), .ZN(n8220) );
  NAND2_X1 U5576 ( .A1(n8253), .A2(n4820), .ZN(n4819) );
  NAND2_X1 U5577 ( .A1(n8253), .A2(n4824), .ZN(n8238) );
  NAND2_X1 U5578 ( .A1(n7230), .A2(n7229), .ZN(n8470) );
  NAND2_X1 U5579 ( .A1(n4831), .A2(n4828), .ZN(n8332) );
  NAND2_X1 U5580 ( .A1(n7211), .A2(n7210), .ZN(n8483) );
  NAND2_X1 U5581 ( .A1(n5488), .A2(n9788), .ZN(n9783) );
  AND2_X1 U5582 ( .A1(n5812), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9821) );
  NAND2_X1 U5583 ( .A1(n5161), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5162) );
  INV_X1 U5584 ( .A(n7367), .ZN(n7539) );
  INV_X1 U5585 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9978) );
  INV_X1 U5586 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6193) );
  INV_X1 U5587 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5792) );
  INV_X1 U5588 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U5589 ( .A1(n4507), .A2(n5224), .ZN(n4506) );
  INV_X1 U5590 ( .A(n9123), .ZN(n9157) );
  NAND2_X1 U5591 ( .A1(n7881), .A2(n7880), .ZN(n9397) );
  NAND2_X1 U5592 ( .A1(n7878), .A2(n8760), .ZN(n7881) );
  NAND2_X1 U5593 ( .A1(n6442), .A2(n6441), .ZN(n6668) );
  NAND2_X1 U5594 ( .A1(n4475), .A2(n6107), .ZN(n4473) );
  NAND2_X1 U5595 ( .A1(n4857), .A2(n4860), .ZN(n8573) );
  NAND2_X1 U5596 ( .A1(n8611), .A2(n7836), .ZN(n8582) );
  AND2_X1 U5597 ( .A1(n7861), .A2(n7842), .ZN(n9192) );
  NAND2_X1 U5598 ( .A1(n8590), .A2(n7695), .ZN(n8604) );
  NAND2_X1 U5599 ( .A1(n4405), .A2(n5536), .ZN(n5837) );
  INV_X1 U5600 ( .A(n4406), .ZN(n4405) );
  OAI22_X1 U5601 ( .A1(n5789), .A2(n6110), .B1(n5951), .B2(n9555), .ZN(n4406)
         );
  NAND2_X1 U5602 ( .A1(n4872), .A2(n6257), .ZN(n6260) );
  NOR2_X1 U5603 ( .A1(n4859), .A2(n4861), .ZN(n8625) );
  NOR3_X1 U5604 ( .A1(n8642), .A2(n8646), .A3(n4865), .ZN(n4859) );
  OAI21_X1 U5605 ( .B1(n6678), .B2(n4491), .A(n4490), .ZN(n7076) );
  NAND2_X1 U5606 ( .A1(n6678), .A2(n6677), .ZN(n6935) );
  AND2_X1 U5607 ( .A1(n5500), .A2(n5355), .ZN(n5383) );
  AND2_X1 U5608 ( .A1(n8980), .A2(n5391), .ZN(n8668) );
  OR2_X1 U5609 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  INV_X1 U5610 ( .A(n8653), .ZN(n8679) );
  NAND2_X1 U5611 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  NOR2_X1 U5612 ( .A1(n8972), .A2(n6189), .ZN(n4425) );
  NAND2_X1 U5613 ( .A1(n8975), .A2(n6189), .ZN(n4423) );
  OR2_X1 U5614 ( .A1(n7863), .A2(n5140), .ZN(n5145) );
  INV_X1 U5615 ( .A(n4413), .ZN(n5556) );
  NAND2_X1 U5616 ( .A1(n9025), .A2(n5002), .ZN(n5034) );
  NOR2_X1 U5617 ( .A1(n4417), .A2(n4416), .ZN(n5443) );
  INV_X1 U5618 ( .A(n5009), .ZN(n4416) );
  INV_X1 U5619 ( .A(n5010), .ZN(n4417) );
  NOR2_X1 U5620 ( .A1(n9584), .A2(n4411), .ZN(n9596) );
  NOR2_X1 U5621 ( .A1(n9040), .A2(n9052), .ZN(n4411) );
  OR2_X1 U5622 ( .A1(n4965), .A2(n9011), .ZN(n9632) );
  INV_X1 U5623 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5042) );
  INV_X1 U5624 ( .A(n9077), .ZN(n9384) );
  NAND2_X1 U5625 ( .A1(n4725), .A2(n9093), .ZN(n9189) );
  NAND2_X1 U5626 ( .A1(n9199), .A2(n4286), .ZN(n4725) );
  NAND2_X1 U5627 ( .A1(n4386), .A2(n4277), .ZN(n9213) );
  OR2_X1 U5628 ( .A1(n9227), .A2(n9089), .ZN(n4386) );
  NAND2_X1 U5629 ( .A1(n4616), .A2(n4618), .ZN(n9233) );
  NAND2_X1 U5630 ( .A1(n9249), .A2(n9243), .ZN(n4616) );
  AND2_X1 U5631 ( .A1(n7796), .A2(n7795), .ZN(n9231) );
  OAI21_X1 U5632 ( .B1(n9249), .B2(n9107), .A(n9243), .ZN(n9247) );
  NAND2_X1 U5633 ( .A1(n4739), .A2(n9087), .ZN(n9242) );
  INV_X1 U5634 ( .A(n4391), .ZN(n9086) );
  NAND2_X1 U5635 ( .A1(n4629), .A2(n4630), .ZN(n9277) );
  INV_X1 U5636 ( .A(n4393), .ZN(n9276) );
  NAND2_X1 U5637 ( .A1(n7717), .A2(n7716), .ZN(n9311) );
  NAND2_X1 U5638 ( .A1(n4711), .A2(n4713), .ZN(n9297) );
  NAND2_X1 U5639 ( .A1(n4712), .A2(n4715), .ZN(n9295) );
  AND2_X1 U5640 ( .A1(n4717), .A2(n4718), .ZN(n9317) );
  NAND2_X1 U5641 ( .A1(n9350), .A2(n9351), .ZN(n4717) );
  NAND2_X1 U5642 ( .A1(n4742), .A2(n7039), .ZN(n9081) );
  NAND2_X1 U5643 ( .A1(n4390), .A2(n6904), .ZN(n7038) );
  NAND2_X1 U5644 ( .A1(n6759), .A2(n6758), .ZN(n6969) );
  NAND2_X1 U5645 ( .A1(n4730), .A2(n6605), .ZN(n6757) );
  NAND2_X1 U5646 ( .A1(n6495), .A2(n4735), .ZN(n4730) );
  NAND2_X1 U5647 ( .A1(n4397), .A2(n4403), .ZN(n6570) );
  NAND2_X1 U5648 ( .A1(n6534), .A2(n4401), .ZN(n4397) );
  NAND2_X1 U5649 ( .A1(n6446), .A2(n6445), .ZN(n6580) );
  NAND2_X1 U5650 ( .A1(n6537), .A2(n8702), .ZN(n6522) );
  NAND2_X1 U5651 ( .A1(n6534), .A2(n6492), .ZN(n6521) );
  NAND2_X1 U5652 ( .A1(n6552), .A2(n6491), .ZN(n6536) );
  NAND2_X1 U5653 ( .A1(n6143), .A2(n6142), .ZN(n6164) );
  INV_X1 U5654 ( .A(n5837), .ZN(n6156) );
  NOR2_X1 U5655 ( .A1(n9388), .A2(n4375), .ZN(n4374) );
  INV_X1 U5656 ( .A(n9387), .ZN(n4376) );
  INV_X1 U5657 ( .A(n9392), .ZN(n4404) );
  NAND2_X1 U5658 ( .A1(n9393), .A2(n9456), .ZN(n4632) );
  AND2_X1 U5659 ( .A1(n5127), .A2(n5130), .ZN(n5125) );
  OAI211_X1 U5660 ( .C1(n7354), .C2(n4765), .A(n4757), .B(n4762), .ZN(n8531)
         );
  CLKBUF_X1 U5661 ( .A(n4964), .Z(n9011) );
  XNOR2_X1 U5662 ( .A(n6845), .B(n6844), .ZN(n7653) );
  INV_X1 U5663 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U5664 ( .A(n5095), .B(n5094), .ZN(n6191) );
  INV_X1 U5665 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9976) );
  INV_X1 U5666 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U5667 ( .A1(n4646), .A2(n5068), .ZN(n5079) );
  NAND2_X1 U5668 ( .A1(n5066), .A2(n5065), .ZN(n4646) );
  INV_X1 U5669 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5534) );
  INV_X1 U5670 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5502) );
  XNOR2_X1 U5671 ( .A(n4422), .B(n4980), .ZN(n5367) );
  NAND2_X1 U5672 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4422) );
  NAND2_X1 U5673 ( .A1(n9746), .A2(n6315), .ZN(n6325) );
  NAND2_X1 U5674 ( .A1(n4642), .A2(n4641), .ZN(n4752) );
  AOI21_X1 U5675 ( .B1(n4751), .B2(n4750), .A(n4749), .ZN(n4748) );
  AOI21_X1 U5676 ( .B1(n7602), .B2(n7365), .A(n7549), .ZN(n4641) );
  OR2_X1 U5677 ( .A1(n9889), .A2(n5433), .ZN(n4364) );
  OAI21_X1 U5678 ( .B1(n8422), .B2(n9829), .A(n4288), .ZN(n4366) );
  NAND2_X1 U5679 ( .A1(n10073), .A2(n9883), .ZN(n4805) );
  INV_X1 U5680 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U5681 ( .A1(n7895), .A2(n7910), .ZN(n4356) );
  INV_X1 U5682 ( .A(n4610), .ZN(n9459) );
  INV_X1 U5683 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n4609) );
  AND2_X1 U5684 ( .A1(n4700), .A2(n4698), .ZN(n4265) );
  INV_X1 U5685 ( .A(n7428), .ZN(n4662) );
  AND3_X1 U5686 ( .A1(n8264), .A2(n7465), .A3(n7477), .ZN(n4266) );
  AND2_X1 U5687 ( .A1(n8160), .A2(n8145), .ZN(n4267) );
  AND4_X1 U5688 ( .A1(n4896), .A2(n4895), .A3(n4894), .A4(n4893), .ZN(n4268)
         );
  NOR2_X1 U5689 ( .A1(n7774), .A2(n4865), .ZN(n4269) );
  OR2_X1 U5690 ( .A1(n9448), .A2(n9302), .ZN(n4270) );
  AND2_X1 U5691 ( .A1(n7975), .A2(n4699), .ZN(n4271) );
  OR2_X1 U5692 ( .A1(n9094), .A2(n9207), .ZN(n4272) );
  OAI21_X1 U5693 ( .B1(n4723), .B2(n4720), .A(n4310), .ZN(n4719) );
  AND2_X1 U5694 ( .A1(n8382), .A2(n7438), .ZN(n4273) );
  AND2_X1 U5695 ( .A1(n4658), .A2(n7454), .ZN(n4274) );
  MUX2_X1 U5696 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9483), .S(n5951), .Z(n6178) );
  NAND2_X1 U5697 ( .A1(n6112), .A2(n6111), .ZN(n6547) );
  AND2_X1 U5698 ( .A1(n4858), .A2(n4269), .ZN(n4275) );
  AND2_X1 U5699 ( .A1(n4713), .A2(n4335), .ZN(n4276) );
  NAND2_X1 U5700 ( .A1(n9038), .A2(n9039), .ZN(n9040) );
  OR2_X1 U5701 ( .A1(n7547), .A2(n4536), .ZN(n7477) );
  INV_X1 U5702 ( .A(n7597), .ZN(n4575) );
  OR2_X1 U5703 ( .A1(n9231), .A2(n9088), .ZN(n4277) );
  NOR2_X1 U5704 ( .A1(n4343), .A2(n4740), .ZN(n4278) );
  NAND2_X1 U5705 ( .A1(n9091), .A2(n4387), .ZN(n4279) );
  NAND2_X1 U5706 ( .A1(n5384), .A2(n5383), .ZN(n5501) );
  INV_X1 U5707 ( .A(n8998), .ZN(n4407) );
  AND2_X1 U5708 ( .A1(n7290), .A2(n7289), .ZN(n8188) );
  OR2_X1 U5709 ( .A1(n5667), .A2(n4782), .ZN(n4280) );
  OR2_X1 U5710 ( .A1(n5290), .A2(n4460), .ZN(n4281) );
  AND2_X1 U5711 ( .A1(n4650), .A2(n4373), .ZN(n4282) );
  NOR2_X1 U5712 ( .A1(n7834), .A2(n7833), .ZN(n7835) );
  AND2_X1 U5713 ( .A1(n5782), .A2(n5781), .ZN(n4283) );
  AND2_X1 U5714 ( .A1(n4655), .A2(n4652), .ZN(n4284) );
  NAND2_X1 U5715 ( .A1(n7075), .A2(n7074), .ZN(n4285) );
  OR2_X1 U5716 ( .A1(n9203), .A2(n9092), .ZN(n4286) );
  AND2_X1 U5717 ( .A1(n8264), .A2(n7461), .ZN(n4287) );
  AND2_X1 U5718 ( .A1(n4798), .A2(n4368), .ZN(n4288) );
  AND3_X1 U5719 ( .A1(n4875), .A2(n4891), .A3(n4983), .ZN(n4978) );
  AND2_X1 U5720 ( .A1(n4491), .A2(n4285), .ZN(n4289) );
  INV_X1 U5721 ( .A(n8945), .ZN(n6538) );
  NAND2_X1 U5722 ( .A1(n8702), .A2(n8800), .ZN(n8945) );
  NAND2_X1 U5723 ( .A1(n7670), .A2(n7665), .ZN(n4290) );
  NAND2_X1 U5724 ( .A1(n4766), .A2(n7360), .ZN(n7362) );
  INV_X1 U5725 ( .A(n5590), .ZN(n8942) );
  INV_X1 U5726 ( .A(n8700), .ZN(n4623) );
  NOR2_X1 U5727 ( .A1(n8341), .A2(n7448), .ZN(n8324) );
  INV_X1 U5728 ( .A(n7399), .ZN(n4676) );
  OAI21_X1 U5729 ( .B1(n6191), .B2(n6281), .A(n4674), .ZN(n6317) );
  NAND2_X1 U5730 ( .A1(n7280), .A2(n7279), .ZN(n8440) );
  INV_X1 U5731 ( .A(n8440), .ZN(n8216) );
  NAND2_X1 U5732 ( .A1(n4623), .A2(n8702), .ZN(n4291) );
  AND2_X1 U5733 ( .A1(n4875), .A2(n4983), .ZN(n4992) );
  INV_X1 U5734 ( .A(n9109), .ZN(n4620) );
  NOR3_X1 U5735 ( .A1(n8221), .A2(n4538), .A3(n8424), .ZN(n4537) );
  AND2_X1 U5736 ( .A1(n5075), .A2(n4941), .ZN(n5071) );
  XNOR2_X1 U5737 ( .A(n5088), .B(SI_6_), .ZN(n5086) );
  AND2_X1 U5738 ( .A1(n8935), .A2(n9108), .ZN(n9243) );
  AND3_X1 U5739 ( .A1(n7455), .A2(n7461), .A3(n7454), .ZN(n4292) );
  AND2_X1 U5740 ( .A1(n9448), .A2(n9302), .ZN(n4293) );
  OR2_X1 U5741 ( .A1(n9135), .A2(n9134), .ZN(n4294) );
  AND2_X1 U5742 ( .A1(n9294), .A2(n4716), .ZN(n4295) );
  NAND2_X1 U5743 ( .A1(n7633), .A2(n7632), .ZN(n9393) );
  AND2_X1 U5744 ( .A1(n9797), .A2(n6972), .ZN(n4296) );
  AND2_X1 U5745 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4297) );
  AND2_X1 U5746 ( .A1(n6959), .A2(n6958), .ZN(n4298) );
  NAND2_X1 U5747 ( .A1(n7215), .A2(n7214), .ZN(n8480) );
  AND2_X1 U5748 ( .A1(n8246), .A2(n8244), .ZN(n4299) );
  NAND2_X1 U5749 ( .A1(n7778), .A2(n7777), .ZN(n9426) );
  NAND2_X1 U5750 ( .A1(n4445), .A2(n7839), .ZN(n9094) );
  NAND2_X1 U5751 ( .A1(n9264), .A2(n4601), .ZN(n4603) );
  AND2_X1 U5752 ( .A1(n7248), .A2(n7247), .ZN(n8279) );
  INV_X1 U5753 ( .A(n8279), .ZN(n8458) );
  AND2_X1 U5754 ( .A1(n8228), .A2(n8229), .ZN(n4300) );
  INV_X1 U5755 ( .A(n9093), .ZN(n4727) );
  INV_X1 U5756 ( .A(n8161), .ZN(n7529) );
  NAND2_X1 U5757 ( .A1(n7487), .A2(n7486), .ZN(n8161) );
  AND2_X1 U5758 ( .A1(n4706), .A2(n6312), .ZN(n4301) );
  AND2_X1 U5759 ( .A1(n4631), .A2(n9298), .ZN(n4302) );
  NAND2_X1 U5760 ( .A1(n8130), .A2(n8129), .ZN(n4303) );
  AND2_X1 U5761 ( .A1(n8945), .A2(n6491), .ZN(n4304) );
  NAND2_X1 U5762 ( .A1(n4407), .A2(n5837), .ZN(n8905) );
  INV_X1 U5763 ( .A(n4823), .ZN(n4822) );
  NAND2_X1 U5764 ( .A1(n7464), .A2(n7460), .ZN(n4305) );
  INV_X1 U5765 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4370) );
  AND2_X1 U5766 ( .A1(n4857), .A2(n4855), .ZN(n4306) );
  INV_X1 U5767 ( .A(n4653), .ZN(n4652) );
  NAND2_X1 U5768 ( .A1(n4656), .A2(n4654), .ZN(n4653) );
  OR2_X1 U5769 ( .A1(n6275), .A2(n4843), .ZN(n4307) );
  INV_X1 U5770 ( .A(n8335), .ZN(n4836) );
  AND2_X1 U5771 ( .A1(n7103), .A2(n7102), .ZN(n4308) );
  INV_X1 U5772 ( .A(n4582), .ZN(n4581) );
  NOR2_X1 U5773 ( .A1(n7600), .A2(n7599), .ZN(n4582) );
  AOI21_X1 U5774 ( .B1(n9243), .B2(n9107), .A(n4619), .ZN(n4618) );
  OR2_X1 U5775 ( .A1(n8480), .A2(n8358), .ZN(n7222) );
  INV_X1 U5776 ( .A(n4886), .ZN(n4485) );
  NOR2_X1 U5777 ( .A1(n8443), .A2(n8248), .ZN(n4309) );
  NAND2_X1 U5778 ( .A1(n9402), .A2(n9186), .ZN(n4310) );
  AND2_X1 U5779 ( .A1(n5081), .A2(SI_5_), .ZN(n4311) );
  INV_X1 U5780 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U5781 ( .A1(n7497), .A2(n7490), .ZN(n7533) );
  INV_X1 U5782 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5073) );
  OAI21_X1 U5783 ( .B1(n4727), .B2(n4286), .A(n9188), .ZN(n4726) );
  OR2_X1 U5784 ( .A1(n8424), .A2(n8145), .ZN(n7487) );
  OR2_X1 U5785 ( .A1(n9084), .A2(n4293), .ZN(n4312) );
  AND2_X1 U5786 ( .A1(n4490), .A2(n4285), .ZN(n4313) );
  AND2_X2 U5787 ( .A1(n5342), .A2(n5494), .ZN(n5357) );
  AND2_X1 U5788 ( .A1(n5945), .A2(n6107), .ZN(n4314) );
  AND2_X1 U5789 ( .A1(n4869), .A2(n7695), .ZN(n4315) );
  AND2_X1 U5790 ( .A1(n5158), .A2(n4370), .ZN(n4316) );
  INV_X1 U5791 ( .A(n8428), .ZN(n8175) );
  NAND2_X1 U5792 ( .A1(n7301), .A2(n7300), .ZN(n8428) );
  AND2_X1 U5793 ( .A1(n4909), .A2(n4878), .ZN(n4317) );
  OR2_X1 U5794 ( .A1(n8463), .A2(n8308), .ZN(n7460) );
  AND2_X1 U5795 ( .A1(n4633), .A2(n4632), .ZN(n4318) );
  NAND2_X1 U5796 ( .A1(n8132), .A2(n7434), .ZN(n4319) );
  AND2_X1 U5797 ( .A1(n8882), .A2(n4452), .ZN(n4320) );
  OR2_X1 U5798 ( .A1(n4498), .A2(n4500), .ZN(n4321) );
  NAND2_X1 U5799 ( .A1(n4854), .A2(n8583), .ZN(n4322) );
  AND2_X1 U5800 ( .A1(n4274), .A2(n8325), .ZN(n4323) );
  OR2_X1 U5801 ( .A1(n8890), .A2(n8889), .ZN(n4324) );
  OR2_X1 U5802 ( .A1(n4855), .A2(n4886), .ZN(n4325) );
  INV_X1 U5803 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4878) );
  AND2_X1 U5804 ( .A1(n4703), .A2(n4701), .ZN(n4326) );
  OR2_X1 U5805 ( .A1(n9069), .A2(n9068), .ZN(P1_U3260) );
  INV_X1 U5806 ( .A(n5451), .ZN(n6042) );
  INV_X2 U5807 ( .A(n6042), .ZN(n7322) );
  AND2_X2 U5808 ( .A1(n5429), .A2(n8541), .ZN(n5451) );
  NAND2_X1 U5809 ( .A1(n7128), .A2(n7127), .ZN(n7976) );
  NAND2_X1 U5810 ( .A1(n8591), .A2(n4501), .ZN(n8590) );
  INV_X1 U5811 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4755) );
  INV_X1 U5812 ( .A(n5765), .ZN(n7602) );
  INV_X1 U5813 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4410) );
  NAND2_X1 U5814 ( .A1(n9415), .A2(n9234), .ZN(n4328) );
  NOR2_X1 U5815 ( .A1(n9086), .A2(n4740), .ZN(n4329) );
  NAND2_X1 U5816 ( .A1(n8684), .A2(n8683), .ZN(n9389) );
  INV_X1 U5817 ( .A(n9389), .ZN(n4605) );
  NAND2_X1 U5818 ( .A1(n7818), .A2(n7817), .ZN(n9411) );
  NOR2_X2 U5819 ( .A1(n8644), .A2(n8643), .ZN(n8642) );
  NAND2_X1 U5820 ( .A1(n4897), .A2(n4268), .ZN(n5227) );
  NOR2_X1 U5821 ( .A1(n8353), .A2(n4837), .ZN(n4330) );
  NOR3_X1 U5822 ( .A1(n8309), .A2(n8448), .A3(n4560), .ZN(n4557) );
  AND2_X1 U5823 ( .A1(n7023), .A2(n7428), .ZN(n4331) );
  OR2_X1 U5824 ( .A1(n8293), .A2(n8308), .ZN(n4332) );
  OR2_X1 U5825 ( .A1(n8136), .A2(n8135), .ZN(n4333) );
  AND2_X1 U5826 ( .A1(n9455), .A2(n8990), .ZN(n4334) );
  INV_X1 U5827 ( .A(n9402), .ZN(n9181) );
  NAND2_X1 U5828 ( .A1(n7859), .A2(n7858), .ZN(n9402) );
  NAND2_X1 U5829 ( .A1(n9311), .A2(n9330), .ZN(n4335) );
  INV_X1 U5830 ( .A(n4614), .ZN(n9355) );
  NOR2_X1 U5831 ( .A1(n7053), .A2(n9506), .ZN(n4614) );
  INV_X1 U5832 ( .A(n4558), .ZN(n8257) );
  NOR2_X1 U5833 ( .A1(n8309), .A2(n4560), .ZN(n4558) );
  OR2_X1 U5834 ( .A1(n7105), .A2(n7106), .ZN(n7128) );
  NAND2_X1 U5835 ( .A1(n4262), .A2(n7430), .ZN(n4336) );
  OR2_X1 U5836 ( .A1(n8393), .A2(n8490), .ZN(n4337) );
  NAND2_X1 U5837 ( .A1(n7317), .A2(n7316), .ZN(n8424) );
  INV_X1 U5838 ( .A(n8424), .ZN(n8160) );
  AND2_X1 U5839 ( .A1(n8690), .A2(n8988), .ZN(n4338) );
  AND2_X1 U5840 ( .A1(n7366), .A2(n7368), .ZN(n8140) );
  AND2_X1 U5841 ( .A1(n6021), .A2(SI_18_), .ZN(n4339) );
  INV_X1 U5842 ( .A(n8188), .ZN(n8434) );
  NAND2_X1 U5843 ( .A1(n7656), .A2(n7655), .ZN(n9415) );
  INV_X1 U5844 ( .A(n9415), .ZN(n9217) );
  OAI211_X1 U5845 ( .C1(n5056), .C2(n4507), .A(n5058), .B(n4506), .ZN(n6828)
         );
  NOR2_X1 U5846 ( .A1(n9301), .A2(n9104), .ZN(n4340) );
  OR2_X1 U5847 ( .A1(n7368), .A2(n4262), .ZN(n4341) );
  INV_X1 U5848 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4993) );
  AND2_X1 U5849 ( .A1(n6973), .A2(n6972), .ZN(n4342) );
  NOR2_X1 U5850 ( .A1(n9268), .A2(n9283), .ZN(n4343) );
  NAND2_X1 U5851 ( .A1(n7685), .A2(n7684), .ZN(n9360) );
  INV_X1 U5852 ( .A(n9360), .ZN(n4613) );
  OR2_X1 U5853 ( .A1(n7117), .A2(n4791), .ZN(n4344) );
  NAND2_X1 U5854 ( .A1(n7987), .A2(n4301), .ZN(n9746) );
  INV_X1 U5855 ( .A(n7204), .ZN(n4598) );
  AND2_X1 U5856 ( .A1(n9571), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4345) );
  NAND2_X1 U5857 ( .A1(n5946), .A2(n5945), .ZN(n6109) );
  AND2_X1 U5858 ( .A1(n8334), .A2(n7442), .ZN(n8356) );
  INV_X1 U5859 ( .A(n8356), .ZN(n4834) );
  AND2_X1 U5860 ( .A1(n6189), .A2(n9256), .ZN(n5347) );
  OR2_X1 U5861 ( .A1(n9704), .A2(n4609), .ZN(n4346) );
  NAND2_X1 U5862 ( .A1(n6561), .A2(n9682), .ZN(n6560) );
  INV_X1 U5863 ( .A(n6560), .ZN(n4612) );
  INV_X1 U5864 ( .A(n7009), .ZN(n7520) );
  NAND2_X1 U5865 ( .A1(n7430), .A2(n7428), .ZN(n7009) );
  NAND2_X1 U5866 ( .A1(n8335), .A2(n4833), .ZN(n4832) );
  INV_X1 U5867 ( .A(n4832), .ZN(n4828) );
  AND2_X1 U5868 ( .A1(n6935), .A2(n4873), .ZN(n4347) );
  AND2_X1 U5869 ( .A1(n7332), .A2(n7331), .ZN(n4348) );
  OR2_X1 U5870 ( .A1(n8143), .A2(n8144), .ZN(n4349) );
  INV_X1 U5871 ( .A(n9084), .ZN(n4718) );
  INV_X1 U5872 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4941) );
  INV_X1 U5873 ( .A(n9280), .ZN(n9348) );
  NOR2_X1 U5874 ( .A1(n5836), .A2(n5837), .ZN(n4350) );
  INV_X1 U5875 ( .A(n5342), .ZN(n4502) );
  NAND2_X1 U5876 ( .A1(n5382), .A2(n5403), .ZN(n5384) );
  INV_X1 U5877 ( .A(n5511), .ZN(n5517) );
  INV_X1 U5878 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4507) );
  XNOR2_X1 U5879 ( .A(n5231), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8974) );
  XOR2_X1 U5880 ( .A(n6239), .B(n6527), .Z(n4351) );
  CLKBUF_X1 U5881 ( .A(n9756), .Z(n4352) );
  NOR3_X1 U5882 ( .A1(n6058), .A2(n7629), .A3(n7543), .ZN(n9756) );
  INV_X1 U5883 ( .A(n9721), .ZN(n8046) );
  NAND2_X1 U5884 ( .A1(n9205), .A2(n9206), .ZN(n9204) );
  NOR2_X4 U5885 ( .A1(n9270), .A2(n9106), .ZN(n9249) );
  OAI21_X1 U5886 ( .B1(n6910), .B2(n4626), .A(n4624), .ZN(n9323) );
  NAND2_X1 U5887 ( .A1(n7194), .A2(n8940), .ZN(n7193) );
  AND2_X2 U5888 ( .A1(n4535), .A2(n4684), .ZN(n4826) );
  NAND2_X1 U5889 ( .A1(n8044), .A2(n8043), .ZN(n4597) );
  OAI211_X1 U5890 ( .C1(n7622), .C2(n7621), .A(n4354), .B(n4353), .ZN(n7627)
         );
  NAND2_X1 U5891 ( .A1(n7622), .A2(n7620), .ZN(n4353) );
  NOR2_X2 U5892 ( .A1(n8050), .A2(n7606), .ZN(n7927) );
  OAI211_X1 U5893 ( .C1(n7598), .C2(n4568), .A(n4578), .B(n4565), .ZN(n8051)
         );
  NAND2_X1 U5894 ( .A1(n5612), .A2(n5611), .ZN(n5610) );
  NAND2_X1 U5895 ( .A1(n4470), .A2(n4469), .ZN(n5511) );
  AOI21_X1 U5896 ( .B1(n8555), .B2(n4851), .A(n4322), .ZN(n4465) );
  NAND2_X1 U5897 ( .A1(n8581), .A2(n7855), .ZN(n8654) );
  NAND2_X1 U5898 ( .A1(n4479), .A2(n4477), .ZN(n6675) );
  NAND2_X1 U5899 ( .A1(n6678), .A2(n4313), .ZN(n4489) );
  NAND2_X1 U5900 ( .A1(n4858), .A2(n4484), .ZN(n4483) );
  NAND2_X1 U5901 ( .A1(n5845), .A2(n5844), .ZN(n5944) );
  NOR2_X1 U5902 ( .A1(n4468), .A2(n4467), .ZN(n4466) );
  OAI21_X1 U5903 ( .B1(n4483), .B2(n8646), .A(n4325), .ZN(n7811) );
  NAND3_X1 U5904 ( .A1(n4356), .A2(n4355), .A3(n7915), .ZN(P1_U3218) );
  NAND3_X1 U5905 ( .A1(n7916), .A2(n7913), .A3(n7914), .ZN(n4355) );
  NAND2_X1 U5906 ( .A1(n4489), .A2(n4487), .ZN(n7676) );
  NAND2_X1 U5907 ( .A1(n7814), .A2(n4466), .ZN(n8555) );
  NAND2_X1 U5908 ( .A1(n4853), .A2(n4465), .ZN(n8581) );
  NAND2_X1 U5909 ( .A1(n4366), .A2(n9889), .ZN(n4365) );
  INV_X1 U5910 ( .A(n8632), .ZN(n4468) );
  AND2_X1 U5911 ( .A1(n9789), .A2(n4812), .ZN(n4358) );
  NAND2_X1 U5912 ( .A1(n4636), .A2(n4634), .ZN(n9391) );
  OAI211_X1 U5913 ( .C1(n9394), .C2(n9678), .A(n4318), .B(n4404), .ZN(n9462)
         );
  OR2_X1 U5914 ( .A1(n6510), .A2(n4291), .ZN(n4622) );
  NAND2_X1 U5915 ( .A1(n9154), .A2(n9153), .ZN(n9152) );
  NOR2_X1 U5916 ( .A1(n9158), .A2(n4360), .ZN(n9396) );
  AOI21_X1 U5917 ( .B1(n9175), .B2(n9397), .A(n9696), .ZN(n4361) );
  NOR2_X2 U5918 ( .A1(n9190), .A2(n9094), .ZN(n9174) );
  NAND2_X1 U5919 ( .A1(n9318), .A2(n9442), .ZN(n9307) );
  NAND2_X1 U5920 ( .A1(n4365), .A2(n4364), .ZN(P2_U3549) );
  NAND2_X1 U5921 ( .A1(n9368), .A2(n6479), .ZN(n5836) );
  NAND2_X1 U5922 ( .A1(n8374), .A2(n8373), .ZN(n8372) );
  MUX2_X2 U5923 ( .A(n8792), .B(n8791), .S(n8884), .Z(n8804) );
  MUX2_X2 U5924 ( .A(n8854), .B(n8853), .S(n8891), .Z(n8857) );
  MUX2_X2 U5925 ( .A(n8773), .B(n8772), .S(n8884), .Z(n8782) );
  NAND2_X1 U5926 ( .A1(n4424), .A2(n4423), .ZN(n8986) );
  NAND4_X1 U5927 ( .A1(n4983), .A2(n4875), .A3(n4892), .A4(n4891), .ZN(n4966)
         );
  NAND3_X1 U5928 ( .A1(n8973), .A2(n4427), .A3(n4363), .ZN(n4426) );
  OAI21_X4 U5929 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5042), .ZN(n4639) );
  NAND2_X2 U5930 ( .A1(n8255), .A2(n8254), .ZN(n8253) );
  OAI21_X1 U5931 ( .B1(n5065), .B2(n4649), .A(n5078), .ZN(n4648) );
  NAND2_X2 U5932 ( .A1(n8190), .A2(n8191), .ZN(n8189) );
  INV_X1 U5933 ( .A(n7338), .ZN(n8142) );
  OAI21_X1 U5934 ( .B1(n6986), .B2(n4663), .A(n4659), .ZN(n8401) );
  NAND2_X2 U5935 ( .A1(n4826), .A2(n4825), .ZN(n5156) );
  AOI21_X2 U5936 ( .B1(n8208), .B2(n8207), .A(n4372), .ZN(n8190) );
  NAND2_X2 U5937 ( .A1(n8227), .A2(n7472), .ZN(n8208) );
  NAND2_X1 U5938 ( .A1(n5746), .A2(n7507), .ZN(n5881) );
  XOR2_X1 U5939 ( .A(n8142), .B(n8141), .Z(n4799) );
  NAND2_X1 U5940 ( .A1(n8773), .A2(n8774), .ZN(n6505) );
  OAI21_X1 U5941 ( .B1(n6571), .B2(n8949), .A(n8701), .ZN(n6619) );
  NAND2_X1 U5942 ( .A1(n6620), .A2(n8697), .ZN(n6761) );
  AOI21_X1 U5943 ( .B1(n9167), .B2(n9115), .A(n9114), .ZN(n9154) );
  OR2_X2 U5944 ( .A1(n9000), .A2(n9662), .ZN(n8718) );
  INV_X8 U5945 ( .A(n4596), .ZN(n7333) );
  NAND2_X1 U5946 ( .A1(n6908), .A2(n8954), .ZN(n6909) );
  NAND3_X1 U5947 ( .A1(n4376), .A2(n9390), .A3(n4374), .ZN(n9461) );
  NAND2_X1 U5948 ( .A1(n4377), .A2(n4379), .ZN(n9151) );
  NAND2_X1 U5949 ( .A1(n9227), .A2(n4380), .ZN(n4377) );
  NAND2_X1 U5950 ( .A1(n6534), .A2(n4398), .ZN(n4394) );
  NAND2_X1 U5951 ( .A1(n4394), .A2(n4395), .ZN(n4728) );
  NAND2_X2 U5952 ( .A1(n4637), .A2(n4639), .ZN(n4596) );
  NAND3_X1 U5953 ( .A1(n4639), .A2(n4637), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4408) );
  MUX2_X1 U5954 ( .A(n4981), .B(P1_REG2_REG_1__SCAN_IN), .S(n5367), .Z(n5280)
         );
  NAND3_X1 U5955 ( .A1(n8899), .A2(n8900), .A3(n5586), .ZN(n4428) );
  NAND2_X1 U5956 ( .A1(n5691), .A2(n4433), .ZN(n4430) );
  NAND2_X1 U5957 ( .A1(n4430), .A2(n4431), .ZN(n6183) );
  NAND2_X1 U5958 ( .A1(n5116), .A2(n4442), .ZN(n4438) );
  NAND2_X1 U5959 ( .A1(n4438), .A2(n4439), .ZN(n5181) );
  NAND2_X1 U5960 ( .A1(n7837), .A2(n8760), .ZN(n4445) );
  NAND2_X1 U5961 ( .A1(n4449), .A2(n4320), .ZN(n8898) );
  NAND4_X1 U5962 ( .A1(n4451), .A2(n4450), .A3(n8878), .A4(n9137), .ZN(n4449)
         );
  NAND2_X1 U5963 ( .A1(n8871), .A2(n8891), .ZN(n4450) );
  NAND2_X1 U5964 ( .A1(n8870), .A2(n8884), .ZN(n4451) );
  NAND2_X1 U5965 ( .A1(n5174), .A2(n4458), .ZN(n4457) );
  NAND2_X1 U5966 ( .A1(n5174), .A2(n4462), .ZN(n4461) );
  MUX2_X1 U5967 ( .A(n5534), .B(n5792), .S(n4596), .Z(n5067) );
  INV_X1 U5968 ( .A(n7813), .ZN(n4467) );
  NAND2_X1 U5969 ( .A1(n4471), .A2(n5500), .ZN(n4469) );
  NAND3_X1 U5970 ( .A1(n5382), .A2(n5500), .A3(n5403), .ZN(n4470) );
  NAND2_X1 U5971 ( .A1(n5297), .A2(n4910), .ZN(n4911) );
  NAND2_X1 U5972 ( .A1(n5946), .A2(n4474), .ZN(n4472) );
  NAND2_X1 U5973 ( .A1(n4472), .A2(n4473), .ZN(n6253) );
  OR2_X1 U5974 ( .A1(n4475), .A2(n4314), .ZN(n4474) );
  NAND2_X1 U5975 ( .A1(n4872), .A2(n4480), .ZN(n4479) );
  NAND2_X1 U5976 ( .A1(n8672), .A2(n4494), .ZN(n4493) );
  NAND2_X1 U5977 ( .A1(n8672), .A2(n8673), .ZN(n8591) );
  NAND3_X1 U5978 ( .A1(n4493), .A2(n4492), .A3(n4321), .ZN(n8603) );
  MUX2_X1 U5979 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6061), .S(n6828), .Z(n6820)
         );
  NAND2_X1 U5980 ( .A1(n4523), .A2(n4516), .ZN(n7467) );
  AOI21_X1 U5981 ( .B1(n4292), .B2(n4266), .A(n4517), .ZN(n4516) );
  NAND2_X1 U5982 ( .A1(n7431), .A2(n4530), .ZN(n4529) );
  OAI211_X1 U5983 ( .C1(n4533), .C2(n4531), .A(n4529), .B(n4527), .ZN(n7441)
         );
  NAND2_X1 U5984 ( .A1(n7426), .A2(n4534), .ZN(n4533) );
  AND2_X2 U5985 ( .A1(n5075), .A2(n4540), .ZN(n4535) );
  INV_X1 U5986 ( .A(n4537), .ZN(n8146) );
  NOR2_X1 U5987 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4547) );
  NOR2_X1 U5988 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4546) );
  NOR2_X1 U5989 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4545) );
  AND2_X2 U5990 ( .A1(n5057), .A2(n4940), .ZN(n5075) );
  NOR2_X2 U5991 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5057) );
  NOR2_X2 U5992 ( .A1(n4544), .A2(n4541), .ZN(n4684) );
  NAND3_X1 U5993 ( .A1(n4543), .A2(n4542), .A3(n5104), .ZN(n4541) );
  NAND4_X1 U5994 ( .A1(n4548), .A2(n4547), .A3(n4546), .A4(n4545), .ZN(n4544)
         );
  NOR2_X1 U5995 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4548) );
  NAND2_X1 U5996 ( .A1(n7401), .A2(n9848), .ZN(n4554) );
  NAND2_X1 U5997 ( .A1(n4555), .A2(n4553), .ZN(n6289) );
  INV_X1 U5998 ( .A(n4557), .ZN(n8239) );
  NAND2_X1 U5999 ( .A1(n4564), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U6000 ( .A1(n7598), .A2(n4566), .ZN(n4565) );
  NAND3_X1 U6001 ( .A1(n4577), .A2(n4583), .A3(n4581), .ZN(n7969) );
  OR2_X1 U6002 ( .A1(n8008), .A2(n8007), .ZN(n4584) );
  NAND2_X1 U6003 ( .A1(n5066), .A2(n4585), .ZN(n4586) );
  NAND2_X1 U6004 ( .A1(n4587), .A2(n4645), .ZN(n5087) );
  NAND2_X1 U6005 ( .A1(n5066), .A2(n4647), .ZN(n4587) );
  INV_X1 U6006 ( .A(n5086), .ZN(n4588) );
  INV_X1 U6007 ( .A(n4639), .ZN(n4593) );
  INV_X1 U6008 ( .A(n4637), .ZN(n4595) );
  NAND3_X1 U6009 ( .A1(n5260), .A2(n4594), .A3(n4592), .ZN(n5045) );
  NAND2_X1 U6010 ( .A1(n4593), .A2(n4297), .ZN(n4592) );
  NAND2_X1 U6011 ( .A1(n4595), .A2(n4297), .ZN(n4594) );
  NAND3_X1 U6012 ( .A1(n4639), .A2(n4637), .A3(n5043), .ZN(n5260) );
  NAND2_X1 U6013 ( .A1(n9264), .A2(n4599), .ZN(n9190) );
  INV_X1 U6014 ( .A(n4603), .ZN(n9215) );
  AND2_X1 U6015 ( .A1(n9174), .A2(n4608), .ZN(n9158) );
  NAND2_X1 U6016 ( .A1(n9174), .A2(n9181), .ZN(n9175) );
  OAI21_X1 U6017 ( .B1(n4610), .B2(n9702), .A(n4346), .ZN(P1_U3522) );
  INV_X1 U6018 ( .A(n8771), .ZN(n4621) );
  NAND2_X2 U6019 ( .A1(n5831), .A2(n8904), .ZN(n8771) );
  NAND2_X2 U6020 ( .A1(n8911), .A2(n5591), .ZN(n5831) );
  NAND2_X2 U6021 ( .A1(n6473), .A2(n8718), .ZN(n8911) );
  INV_X1 U6022 ( .A(n5587), .ZN(n5591) );
  XNOR2_X2 U6023 ( .A(n7204), .B(n9002), .ZN(n8940) );
  NAND2_X2 U6024 ( .A1(n5371), .A2(n5370), .ZN(n7204) );
  NAND3_X1 U6025 ( .A1(n9152), .A2(n9137), .A3(n9138), .ZN(n9136) );
  NAND2_X1 U6026 ( .A1(n6909), .A2(n8691), .ZN(n6910) );
  NAND2_X2 U6027 ( .A1(n8942), .A2(n8722), .ZN(n6473) );
  NAND2_X1 U6028 ( .A1(n7193), .A2(n5589), .ZN(n8722) );
  NAND2_X1 U6029 ( .A1(n9204), .A2(n9113), .ZN(n9167) );
  NAND2_X2 U6030 ( .A1(n4638), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4637) );
  NAND2_X2 U6031 ( .A1(n8262), .A2(n4299), .ZN(n8245) );
  NAND2_X2 U6032 ( .A1(n8280), .A2(n4640), .ZN(n8262) );
  NAND2_X1 U6033 ( .A1(n4323), .A2(n8341), .ZN(n4650) );
  NAND2_X1 U6034 ( .A1(n4655), .A2(n4656), .ZN(n8304) );
  INV_X1 U6035 ( .A(n8305), .ZN(n4654) );
  NAND2_X1 U6036 ( .A1(n8189), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U6037 ( .A1(n8189), .A2(n7478), .ZN(n8177) );
  OAI21_X1 U6038 ( .B1(n8035), .B2(n4678), .A(n4677), .ZN(n5800) );
  AOI21_X1 U6039 ( .B1(n9718), .B2(n4683), .A(n4283), .ZN(n4677) );
  INV_X1 U6040 ( .A(n9718), .ZN(n4678) );
  NAND2_X1 U6041 ( .A1(n8035), .A2(n4682), .ZN(n4681) );
  INV_X1 U6042 ( .A(n5775), .ZN(n4683) );
  NAND2_X1 U6043 ( .A1(n9719), .A2(n9718), .ZN(n9717) );
  NAND3_X1 U6044 ( .A1(n4684), .A2(n5075), .A3(n4941), .ZN(n5696) );
  NAND2_X1 U6045 ( .A1(n6866), .A2(n4688), .ZN(n4685) );
  NAND2_X1 U6046 ( .A1(n4685), .A2(n4686), .ZN(n7105) );
  NAND2_X2 U6047 ( .A1(n4693), .A2(n4691), .ZN(n7946) );
  OAI22_X1 U6048 ( .A1(n6281), .A2(n5618), .B1(n6283), .B2(n6828), .ZN(n4692)
         );
  NAND2_X1 U6049 ( .A1(n7976), .A2(n4265), .ZN(n4696) );
  INV_X1 U6050 ( .A(n7982), .ZN(n4700) );
  NAND2_X1 U6051 ( .A1(n8044), .A2(n8043), .ZN(n4703) );
  INV_X1 U6052 ( .A(n9742), .ZN(n4706) );
  NOR2_X2 U6053 ( .A1(n5156), .A2(n4945), .ZN(n4948) );
  NAND3_X1 U6054 ( .A1(n6143), .A2(n6161), .A3(n6142), .ZN(n4710) );
  NAND2_X1 U6055 ( .A1(n4728), .A2(n4729), .ZN(n6903) );
  NAND2_X1 U6056 ( .A1(n6495), .A2(n6494), .ZN(n6607) );
  INV_X1 U6057 ( .A(n6494), .ZN(n4736) );
  AND2_X1 U6058 ( .A1(n9436), .A2(n9303), .ZN(n4740) );
  NAND2_X1 U6059 ( .A1(n4742), .A2(n4741), .ZN(n9083) );
  AND3_X2 U6060 ( .A1(n4897), .A2(n4317), .A3(n4268), .ZN(n5413) );
  OR2_X2 U6061 ( .A1(n5128), .A2(n4993), .ZN(n4939) );
  AND2_X2 U6062 ( .A1(n5413), .A2(n4935), .ZN(n5128) );
  NAND3_X1 U6063 ( .A1(n7494), .A2(n4341), .A3(n4743), .ZN(n7502) );
  NAND2_X1 U6064 ( .A1(n4752), .A2(n4748), .ZN(P2_U3244) );
  INV_X1 U6065 ( .A(n7354), .ZN(n4756) );
  NAND2_X1 U6066 ( .A1(n7354), .A2(n4764), .ZN(n4757) );
  NAND2_X1 U6067 ( .A1(n4761), .A2(n4756), .ZN(n4760) );
  NAND3_X1 U6068 ( .A1(n4760), .A2(n7358), .A3(n4758), .ZN(n4766) );
  NAND3_X1 U6069 ( .A1(n7354), .A2(n4762), .A3(n4759), .ZN(n4758) );
  NAND2_X1 U6070 ( .A1(n5412), .A2(n4780), .ZN(n4777) );
  NAND2_X1 U6071 ( .A1(n4777), .A2(n4778), .ZN(n5691) );
  NAND2_X1 U6072 ( .A1(n6847), .A2(n4789), .ZN(n4786) );
  NAND2_X1 U6073 ( .A1(n4786), .A2(n4787), .ZN(n7149) );
  NAND2_X1 U6074 ( .A1(n6847), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U6075 ( .A1(n6847), .A2(n6846), .ZN(n7065) );
  NOR2_X1 U6076 ( .A1(n4795), .A2(n7506), .ZN(n7508) );
  OAI21_X1 U6077 ( .B1(n5736), .B2(n4795), .A(n5735), .ZN(n9834) );
  XNOR2_X1 U6078 ( .A(n4795), .B(n5743), .ZN(n5619) );
  AOI21_X2 U6079 ( .B1(n8274), .B2(n8137), .A(n4796), .ZN(n8255) );
  OAI21_X1 U6080 ( .B1(n8422), .B2(n4805), .A(n4800), .ZN(P2_U3517) );
  OR2_X1 U6081 ( .A1(n10073), .A2(n4807), .ZN(n4806) );
  NAND2_X1 U6082 ( .A1(n4811), .A2(n8131), .ZN(n8391) );
  NOR2_X1 U6083 ( .A1(n8243), .A2(n8268), .ZN(n4823) );
  NAND2_X1 U6084 ( .A1(n8351), .A2(n4828), .ZN(n4827) );
  NAND2_X1 U6085 ( .A1(n6027), .A2(n4840), .ZN(n4839) );
  NAND2_X1 U6086 ( .A1(n5366), .A2(n5610), .ZN(n5381) );
  NAND2_X1 U6087 ( .A1(n4264), .A2(n6481), .ZN(n4849) );
  NAND2_X1 U6088 ( .A1(n8556), .A2(n7836), .ZN(n4853) );
  INV_X1 U6089 ( .A(n8642), .ZN(n4858) );
  NAND3_X1 U6090 ( .A1(n5719), .A2(n5721), .A3(n5844), .ZN(n5845) );
  NAND2_X1 U6091 ( .A1(n5719), .A2(n5844), .ZN(n5720) );
  NAND2_X1 U6092 ( .A1(n8590), .A2(n4315), .ZN(n4866) );
  NAND2_X1 U6093 ( .A1(n4866), .A2(n4867), .ZN(n8644) );
  NOR2_X2 U6094 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4875) );
  INV_X1 U6095 ( .A(n5227), .ZN(n4877) );
  AND2_X2 U6096 ( .A1(n6292), .A2(n7405), .ZN(n4887) );
  OAI21_X1 U6097 ( .B1(n7361), .B2(n7531), .A(n7492), .ZN(n7363) );
  XNOR2_X1 U6098 ( .A(n7118), .B(n7117), .ZN(n7837) );
  NAND2_X1 U6099 ( .A1(n5583), .A2(n5590), .ZN(n6472) );
  AND2_X1 U6100 ( .A1(n9789), .A2(n8127), .ZN(n6992) );
  NAND2_X1 U6101 ( .A1(n5192), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5160) );
  OR2_X1 U6102 ( .A1(n5535), .A2(n5618), .ZN(n5370) );
  NAND2_X1 U6103 ( .A1(n4907), .A2(n4906), .ZN(n5262) );
  OR2_X1 U6104 ( .A1(n5337), .A2(n5264), .ZN(n5265) );
  OR2_X1 U6105 ( .A1(n5337), .A2(n5141), .ZN(n5142) );
  NAND2_X1 U6106 ( .A1(n5198), .A2(n8535), .ZN(n8541) );
  NAND2_X1 U6107 ( .A1(n8535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6108 ( .A1(n5195), .A2(n5193), .ZN(n8535) );
  AOI21_X2 U6109 ( .B1(n6200), .B2(n6199), .A(n6198), .ZN(n6292) );
  AOI21_X1 U6110 ( .B1(n6400), .B2(n6345), .A(n4879), .ZN(n6649) );
  AND4_X1 U6111 ( .A1(n5669), .A2(n4914), .A3(n4913), .A4(n4909), .ZN(n4880)
         );
  AND2_X1 U6112 ( .A1(n5356), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4881) );
  INV_X1 U6113 ( .A(n9207), .ZN(n9173) );
  AND4_X1 U6114 ( .A1(n4916), .A2(n4908), .A3(n4915), .A4(n5980), .ZN(n4882)
         );
  AND2_X1 U6115 ( .A1(n5168), .A2(n5122), .ZN(n4883) );
  AND2_X1 U6116 ( .A1(n5411), .A2(n5296), .ZN(n4884) );
  AND2_X1 U6117 ( .A1(n5173), .A2(n5172), .ZN(n4885) );
  AND2_X1 U6118 ( .A1(n7792), .A2(n7791), .ZN(n4886) );
  NOR2_X1 U6119 ( .A1(n6172), .A2(n6189), .ZN(n4888) );
  AND2_X1 U6120 ( .A1(n7311), .A2(n7310), .ZN(n7625) );
  NOR2_X1 U6121 ( .A1(n8126), .A2(n7418), .ZN(n4889) );
  OR2_X1 U6122 ( .A1(n9506), .A2(n9342), .ZN(n4890) );
  INV_X1 U6123 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4893) );
  INV_X1 U6124 ( .A(n7372), .ZN(n5746) );
  INV_X1 U6125 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4940) );
  AND2_X1 U6126 ( .A1(n4882), .A2(n4880), .ZN(n4910) );
  INV_X1 U6127 ( .A(n5112), .ZN(n5114) );
  OAI21_X1 U6128 ( .B1(n8008), .B2(n8248), .A(n8006), .ZN(n7595) );
  INV_X1 U6129 ( .A(n7496), .ZN(n7501) );
  OR2_X1 U6130 ( .A1(n7281), .A2(n10013), .ZN(n7292) );
  OR2_X1 U6131 ( .A1(n6744), .A2(n6743), .ZN(n6876) );
  NAND2_X1 U6132 ( .A1(n5881), .A2(n7376), .ZN(n5930) );
  NOR2_X1 U6133 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4943) );
  INV_X1 U6134 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5104) );
  INV_X1 U6135 ( .A(n7861), .ZN(n7638) );
  INV_X1 U6136 ( .A(n7719), .ZN(n7634) );
  INV_X1 U6137 ( .A(n9134), .ZN(n9137) );
  AND2_X1 U6138 ( .A1(n8738), .A2(n9166), .ZN(n9115) );
  OR2_X1 U6139 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4933) );
  AND2_X1 U6140 ( .A1(n5114), .A2(n5113), .ZN(n5115) );
  INV_X1 U6141 ( .A(n7595), .ZN(n7596) );
  OR2_X1 U6142 ( .A1(n7273), .A2(n8011), .ZN(n7281) );
  INV_X1 U6143 ( .A(n8140), .ZN(n8141) );
  INV_X1 U6144 ( .A(n5745), .ZN(n7507) );
  XNOR2_X1 U6145 ( .A(n7851), .B(n5361), .ZN(n7854) );
  INV_X1 U6146 ( .A(n6261), .ZN(n6258) );
  INV_X1 U6147 ( .A(n5723), .ZN(n5721) );
  OR2_X1 U6148 ( .A1(n7882), .A2(n7641), .ZN(n7896) );
  NAND2_X1 U6149 ( .A1(n7638), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U6150 ( .A1(n7637), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U6151 ( .A1(n7634), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7738) );
  OR2_X1 U6152 ( .A1(n6119), .A2(n10056), .ZN(n6262) );
  OR2_X1 U6153 ( .A1(n9554), .A2(n5015), .ZN(n9556) );
  NAND2_X1 U6154 ( .A1(n5128), .A2(n5125), .ZN(n9476) );
  INV_X1 U6155 ( .A(n5232), .ZN(n5693) );
  NAND2_X1 U6156 ( .A1(n5120), .A2(n5119), .ZN(n5168) );
  XNOR2_X1 U6157 ( .A(n8443), .B(n7607), .ZN(n8008) );
  NAND2_X1 U6158 ( .A1(n7480), .A2(n7478), .ZN(n8185) );
  OR2_X1 U6159 ( .A1(n9764), .A2(n9765), .ZN(n9766) );
  OR2_X1 U6160 ( .A1(n6295), .A2(n6294), .ZN(n6348) );
  NAND2_X1 U6161 ( .A1(n9723), .A2(n5874), .ZN(n7378) );
  INV_X1 U6162 ( .A(n7016), .ZN(n9773) );
  OAI21_X1 U6163 ( .B1(n5876), .B2(n7507), .A(n5875), .ZN(n5926) );
  OR2_X1 U6164 ( .A1(n7841), .A2(n7840), .ZN(n7861) );
  XNOR2_X1 U6165 ( .A(n5539), .B(n5361), .ZN(n5710) );
  AND2_X1 U6166 ( .A1(n7731), .A2(n7730), .ZN(n8646) );
  AND2_X1 U6167 ( .A1(n7642), .A2(n7896), .ZN(n9145) );
  INV_X1 U6168 ( .A(n7783), .ZN(n7898) );
  INV_X1 U6169 ( .A(n9393), .ZN(n9148) );
  AND2_X1 U6170 ( .A1(n8807), .A2(n8691), .ZN(n8954) );
  AND2_X1 U6171 ( .A1(n5593), .A2(n5592), .ZN(n9280) );
  OR2_X1 U6172 ( .A1(n6172), .A2(n8974), .ZN(n9696) );
  AND2_X1 U6173 ( .A1(n5690), .A2(n5663), .ZN(n5688) );
  AND2_X1 U6174 ( .A1(n7321), .A2(n7320), .ZN(n8158) );
  OR2_X1 U6175 ( .A1(n7553), .A2(n9863), .ZN(n9734) );
  AND2_X1 U6176 ( .A1(n7288), .A2(n7287), .ZN(n8232) );
  AND4_X1 U6177 ( .A1(n7110), .A2(n7109), .A3(n7108), .A4(n7107), .ZN(n8405)
         );
  INV_X1 U6178 ( .A(n4352), .ZN(n8091) );
  INV_X1 U6179 ( .A(n8132), .ZN(n8400) );
  INV_X1 U6180 ( .A(n8369), .ZN(n9809) );
  AND2_X1 U6181 ( .A1(n9790), .A2(n8511), .ZN(n9829) );
  AND2_X1 U6182 ( .A1(n5459), .A2(n5458), .ZN(n9814) );
  AND2_X1 U6183 ( .A1(n5091), .A2(n5085), .ZN(n6079) );
  INV_X1 U6184 ( .A(n4259), .ZN(n8983) );
  OR2_X1 U6185 ( .A1(n9177), .A2(n7863), .ZN(n7869) );
  AND2_X1 U6186 ( .A1(n9541), .A2(n9011), .ZN(n9628) );
  AND2_X1 U6187 ( .A1(n9111), .A2(n8863), .ZN(n9220) );
  OR2_X1 U6189 ( .A1(n9696), .A2(n6131), .ZN(n9367) );
  INV_X1 U6190 ( .A(n9369), .ZN(n9361) );
  OR2_X1 U6191 ( .A1(n6172), .A2(n5347), .ZN(n9694) );
  OR2_X1 U6192 ( .A1(n9441), .A2(n9678), .ZN(n9447) );
  INV_X1 U6193 ( .A(n9700), .ZN(n9678) );
  XNOR2_X1 U6194 ( .A(n5096), .B(SI_7_), .ZN(n5094) );
  OR2_X1 U6195 ( .A1(n4958), .A2(n6849), .ZN(n6053) );
  INV_X2 U6196 ( .A(n7560), .ZN(n8070) );
  INV_X1 U6197 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7190) );
  AND2_X1 U6198 ( .A1(n8362), .A2(n8361), .ZN(n8488) );
  INV_X1 U6199 ( .A(n9889), .ZN(n9887) );
  INV_X1 U6200 ( .A(n10073), .ZN(n10071) );
  INV_X1 U6201 ( .A(n9816), .ZN(n9819) );
  INV_X1 U6202 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10041) );
  AND2_X1 U6203 ( .A1(n5499), .A2(n5498), .ZN(n8671) );
  NAND2_X1 U6204 ( .A1(n7869), .A2(n7868), .ZN(n9186) );
  OR2_X1 U6205 ( .A1(P1_U3083), .A2(n5029), .ZN(n9641) );
  OR2_X1 U6206 ( .A1(n5257), .A2(n5275), .ZN(n9713) );
  OR2_X1 U6207 ( .A1(n6141), .A2(n5275), .ZN(n9702) );
  AND2_X1 U6208 ( .A1(n5494), .A2(n5237), .ZN(n9648) );
  NOR2_X1 U6209 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4896) );
  INV_X1 U6210 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4909) );
  NOR2_X1 U6211 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4898) );
  NAND2_X1 U6212 ( .A1(n5413), .A2(n4898), .ZN(n5664) );
  NOR2_X1 U6213 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5233) );
  INV_X1 U6214 ( .A(n5233), .ZN(n4899) );
  NOR2_X1 U6215 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(n4899), .ZN(n4900) );
  NAND2_X1 U6216 ( .A1(n5232), .A2(n4900), .ZN(n4901) );
  INV_X1 U6217 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4913) );
  AOI21_X1 U6218 ( .B1(n5231), .B2(n4913), .A(n4993), .ZN(n4905) );
  INV_X1 U6219 ( .A(n4905), .ZN(n4902) );
  INV_X1 U6220 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6221 ( .A1(n4902), .A2(n4914), .ZN(n4907) );
  INV_X1 U6222 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U6223 ( .A1(n4905), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4906) );
  INV_X1 U6224 ( .A(n5262), .ZN(n8968) );
  NAND2_X1 U6225 ( .A1(n8983), .A2(n8968), .ZN(n8888) );
  NOR2_X1 U6226 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4916) );
  NOR2_X1 U6227 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4908) );
  INV_X1 U6228 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4915) );
  INV_X1 U6229 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5980) );
  INV_X1 U6230 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U6231 ( .A1(n4911), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4925) );
  INV_X1 U6232 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4924) );
  XNOR2_X1 U6233 ( .A(n4925), .B(n4924), .ZN(n6730) );
  INV_X1 U6234 ( .A(n6730), .ZN(n4912) );
  OR2_X1 U6235 ( .A1(n8888), .A2(n4912), .ZN(n4932) );
  AND4_X1 U6236 ( .A1(n5669), .A2(n4914), .A3(n5980), .A4(n4913), .ZN(n4919)
         );
  INV_X1 U6237 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5235) );
  AND3_X1 U6238 ( .A1(n5235), .A2(n4915), .A3(n4924), .ZN(n4918) );
  NOR2_X1 U6239 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4917) );
  NAND4_X1 U6240 ( .A1(n4919), .A2(n4918), .A3(n4917), .A4(n4916), .ZN(n4934)
         );
  INV_X1 U6241 ( .A(n4934), .ZN(n4920) );
  NAND2_X1 U6242 ( .A1(n4921), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4922) );
  MUX2_X1 U6243 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4922), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n4923) );
  NAND2_X1 U6244 ( .A1(n4925), .A2(n4924), .ZN(n4926) );
  INV_X1 U6245 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4927) );
  NOR2_X1 U6246 ( .A1(n7070), .A2(n7158), .ZN(n4931) );
  NAND2_X1 U6247 ( .A1(n4929), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4930) );
  NAND2_X1 U6248 ( .A1(n5356), .A2(n6730), .ZN(n5028) );
  NAND2_X1 U6249 ( .A1(n4932), .A2(n5028), .ZN(n4963) );
  NOR2_X1 U6250 ( .A1(n4934), .A2(n4933), .ZN(n4935) );
  NAND2_X1 U6251 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4936) );
  NAND2_X1 U6252 ( .A1(n4939), .A2(n4936), .ZN(n4937) );
  XNOR2_X2 U6253 ( .A(n4937), .B(P1_IR_REG_28__SCAN_IN), .ZN(n4964) );
  INV_X1 U6254 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4938) );
  XNOR2_X2 U6255 ( .A(n4939), .B(n4938), .ZN(n9071) );
  NAND2_X4 U6256 ( .A1(n4964), .A2(n9071), .ZN(n5951) );
  OAI21_X1 U6257 ( .B1(n4963), .B2(n7733), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  INV_X1 U6258 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n4962) );
  OR2_X2 U6259 ( .A1(n5028), .A2(P1_U3084), .ZN(n9001) );
  INV_X1 U6260 ( .A(n9001), .ZN(P1_U4006) );
  INV_X1 U6261 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4954) );
  INV_X1 U6262 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4944) );
  INV_X1 U6263 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4959) );
  INV_X1 U6264 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4956) );
  NAND4_X1 U6265 ( .A1(n4954), .A2(n4944), .A3(n4959), .A4(n4956), .ZN(n4945)
         );
  NOR2_X1 U6266 ( .A1(n4948), .A2(n5224), .ZN(n4946) );
  MUX2_X1 U6267 ( .A(n5224), .B(n4946), .S(P2_IR_REG_25__SCAN_IN), .Z(n4947)
         );
  INV_X1 U6268 ( .A(n4947), .ZN(n4949) );
  NAND2_X1 U6269 ( .A1(n4949), .A2(n4951), .ZN(n7071) );
  INV_X1 U6270 ( .A(n7071), .ZN(n4953) );
  NAND2_X1 U6271 ( .A1(n4951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4950) );
  MUX2_X1 U6272 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4950), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n4952) );
  NAND2_X1 U6273 ( .A1(n4952), .A2(n5161), .ZN(n7126) );
  INV_X1 U6274 ( .A(n7126), .ZN(n5458) );
  NAND2_X1 U6275 ( .A1(n4953), .A2(n5458), .ZN(n4958) );
  NOR2_X1 U6276 ( .A1(n5156), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6277 ( .A1(n5151), .A2(n4954), .ZN(n5154) );
  NAND2_X1 U6278 ( .A1(n5154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4960) );
  NAND2_X1 U6279 ( .A1(n4960), .A2(n4959), .ZN(n4955) );
  NAND2_X1 U6280 ( .A1(n4955), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4957) );
  XNOR2_X1 U6281 ( .A(n4957), .B(n4956), .ZN(n6849) );
  XNOR2_X1 U6282 ( .A(n4960), .B(n4959), .ZN(n5812) );
  INV_X1 U6283 ( .A(n9821), .ZN(n4961) );
  NOR2_X2 U6284 ( .A1(n6053), .A2(n4961), .ZN(P2_U3966) );
  NOR2_X1 U6285 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10031), .ZN(n6465) );
  NOR2_X1 U6286 ( .A1(n4963), .A2(n4962), .ZN(n5026) );
  INV_X1 U6287 ( .A(n9071), .ZN(n9013) );
  AND2_X1 U6288 ( .A1(n5026), .A2(n9013), .ZN(n9541) );
  INV_X1 U6289 ( .A(n9541), .ZN(n4965) );
  OR2_X1 U6290 ( .A1(n4967), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4976) );
  NOR2_X1 U6291 ( .A1(n4976), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n4970) );
  INV_X1 U6292 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U6293 ( .A1(n4970), .A2(n4968), .ZN(n5005) );
  NAND2_X1 U6294 ( .A1(n5005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4969) );
  XNOR2_X1 U6295 ( .A(n4969), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6239) );
  INV_X1 U6296 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6527) );
  OR2_X1 U6297 ( .A1(n4970), .A2(n4993), .ZN(n4971) );
  XNOR2_X1 U6298 ( .A(n4971), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9028) );
  OR2_X1 U6299 ( .A1(n9028), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5002) );
  NOR2_X1 U6300 ( .A1(n9028), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4972) );
  AOI21_X1 U6301 ( .B1(n9028), .B2(P1_REG2_REG_8__SCAN_IN), .A(n4972), .ZN(
        n9027) );
  NAND2_X1 U6302 ( .A1(n4976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4973) );
  XNOR2_X1 U6303 ( .A(n4973), .B(P1_IR_REG_7__SCAN_IN), .ZN(n5312) );
  OR2_X1 U6304 ( .A1(n5312), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5001) );
  NOR2_X1 U6305 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n5312), .ZN(n4974) );
  AOI21_X1 U6306 ( .B1(n5312), .B2(P1_REG2_REG_7__SCAN_IN), .A(n4974), .ZN(
        n5308) );
  NAND2_X1 U6307 ( .A1(n4967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4975) );
  MUX2_X1 U6308 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4975), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n4977) );
  AND2_X1 U6309 ( .A1(n4977), .A2(n4976), .ZN(n5018) );
  OR2_X1 U6310 ( .A1(n4978), .A2(n4993), .ZN(n4979) );
  XNOR2_X1 U6311 ( .A(n4979), .B(P1_IR_REG_5__SCAN_IN), .ZN(n5069) );
  INV_X1 U6312 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4981) );
  INV_X1 U6313 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4980) );
  AND2_X1 U6314 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9015) );
  INV_X1 U6315 ( .A(n5367), .ZN(n5288) );
  NAND2_X1 U6316 ( .A1(n5288), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U6317 ( .A1(n5279), .A2(n4982), .ZN(n9020) );
  OR2_X1 U6318 ( .A1(n4983), .A2(n4993), .ZN(n4985) );
  INV_X1 U6319 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6320 ( .A1(n4985), .A2(n4984), .ZN(n4987) );
  OAI21_X1 U6321 ( .B1(n4985), .B2(n4984), .A(n4987), .ZN(n5330) );
  XNOR2_X1 U6322 ( .A(n5330), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U6323 ( .A1(n9020), .A2(n9021), .ZN(n9019) );
  INV_X1 U6324 ( .A(n5330), .ZN(n9010) );
  NAND2_X1 U6325 ( .A1(n9010), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6326 ( .A1(n9019), .A2(n4986), .ZN(n5635) );
  INV_X1 U6327 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U6328 ( .A1(n4987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4989) );
  INV_X1 U6329 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4988) );
  XNOR2_X1 U6330 ( .A(n4989), .B(n4988), .ZN(n5647) );
  MUX2_X1 U6331 ( .A(n4990), .B(P1_REG2_REG_3__SCAN_IN), .S(n5647), .Z(n5636)
         );
  NAND2_X1 U6332 ( .A1(n5635), .A2(n5636), .ZN(n5634) );
  OR2_X1 U6333 ( .A1(n5647), .A2(n4990), .ZN(n4991) );
  NAND2_X1 U6334 ( .A1(n5634), .A2(n4991), .ZN(n9550) );
  NOR2_X1 U6335 ( .A1(n4992), .A2(n4993), .ZN(n4994) );
  MUX2_X1 U6336 ( .A(n4993), .B(n4994), .S(P1_IR_REG_4__SCAN_IN), .Z(n4995) );
  INV_X1 U6337 ( .A(n4995), .ZN(n4997) );
  INV_X1 U6338 ( .A(n4978), .ZN(n4996) );
  NAND2_X1 U6339 ( .A1(n4997), .A2(n4996), .ZN(n9555) );
  INV_X1 U6340 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5522) );
  XNOR2_X1 U6341 ( .A(n9555), .B(n5522), .ZN(n9549) );
  INV_X1 U6342 ( .A(n9555), .ZN(n9551) );
  OAI22_X1 U6343 ( .A1(n9550), .A2(n9549), .B1(n9551), .B2(
        P1_REG2_REG_4__SCAN_IN), .ZN(n5317) );
  NOR2_X1 U6344 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n5069), .ZN(n4998) );
  AOI21_X1 U6345 ( .B1(n5069), .B2(P1_REG2_REG_5__SCAN_IN), .A(n4998), .ZN(
        n5318) );
  NAND2_X1 U6346 ( .A1(n5317), .A2(n5318), .ZN(n5316) );
  OAI21_X1 U6347 ( .B1(n5069), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5316), .ZN(
        n5558) );
  INV_X1 U6348 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4999) );
  MUX2_X1 U6349 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n4999), .S(n5018), .Z(n5000)
         );
  INV_X1 U6350 ( .A(n5000), .ZN(n5557) );
  NAND2_X1 U6351 ( .A1(n9027), .A2(n9026), .ZN(n9025) );
  NAND2_X1 U6352 ( .A1(n6239), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6353 ( .A1(n5004), .A2(n5003), .ZN(n5010) );
  OR2_X1 U6354 ( .A1(n5005), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6355 ( .A1(n5006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5187) );
  XNOR2_X1 U6356 ( .A(n5187), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6444) );
  OR2_X1 U6357 ( .A1(n6444), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6358 ( .A1(n6444), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5007) );
  AND2_X1 U6359 ( .A1(n5008), .A2(n5007), .ZN(n5009) );
  NOR2_X1 U6360 ( .A1(n5010), .A2(n5009), .ZN(n5011) );
  NOR3_X1 U6361 ( .A1(n9632), .A2(n5443), .A3(n5011), .ZN(n5032) );
  NOR2_X1 U6362 ( .A1(n6239), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6363 ( .A1(n9028), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5021) );
  INV_X1 U6364 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5960) );
  MUX2_X1 U6365 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n5960), .S(n9028), .Z(n9032)
         );
  NOR2_X1 U6366 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n5312), .ZN(n5020) );
  NAND2_X1 U6367 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n5069), .ZN(n5017) );
  INV_X1 U6368 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5545) );
  MUX2_X1 U6369 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5545), .S(n5069), .Z(n5323)
         );
  INV_X1 U6370 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5521) );
  INV_X1 U6371 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5264) );
  MUX2_X1 U6372 ( .A(n5264), .B(P1_REG1_REG_1__SCAN_IN), .S(n5367), .Z(n5283)
         );
  AND2_X1 U6373 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n5284) );
  NAND2_X1 U6374 ( .A1(n5283), .A2(n5284), .ZN(n9007) );
  OR2_X1 U6375 ( .A1(n5367), .A2(n5264), .ZN(n9003) );
  NAND2_X1 U6376 ( .A1(n9007), .A2(n9003), .ZN(n5012) );
  MUX2_X1 U6377 ( .A(n9706), .B(P1_REG1_REG_2__SCAN_IN), .S(n5330), .Z(n9005)
         );
  AND2_X1 U6378 ( .A1(n5012), .A2(n9005), .ZN(n9006) );
  NOR2_X1 U6379 ( .A1(n5330), .A2(n9706), .ZN(n5640) );
  INV_X1 U6380 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5394) );
  MUX2_X1 U6381 ( .A(n5394), .B(P1_REG1_REG_3__SCAN_IN), .S(n5647), .Z(n5013)
         );
  OAI21_X1 U6382 ( .B1(n9006), .B2(n5640), .A(n5013), .ZN(n5643) );
  OR2_X1 U6383 ( .A1(n5647), .A2(n5394), .ZN(n5014) );
  NAND2_X1 U6384 ( .A1(n5643), .A2(n5014), .ZN(n9554) );
  MUX2_X1 U6385 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n5521), .S(n9555), .Z(n5015)
         );
  INV_X1 U6386 ( .A(n9556), .ZN(n5016) );
  AOI21_X1 U6387 ( .B1(n9555), .B2(n5521), .A(n5016), .ZN(n5324) );
  NAND2_X1 U6388 ( .A1(n5323), .A2(n5324), .ZN(n5322) );
  NAND2_X1 U6389 ( .A1(n5017), .A2(n5322), .ZN(n5561) );
  INV_X1 U6390 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9709) );
  INV_X1 U6391 ( .A(n5018), .ZN(n5848) );
  AOI22_X1 U6392 ( .A1(n5018), .A2(n9709), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n5848), .ZN(n5560) );
  NOR2_X1 U6393 ( .A1(n5561), .A2(n5560), .ZN(n5559) );
  NOR2_X1 U6394 ( .A1(n5018), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5019) );
  NOR2_X1 U6395 ( .A1(n5559), .A2(n5019), .ZN(n5305) );
  INV_X1 U6396 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5859) );
  MUX2_X1 U6397 ( .A(n5859), .B(P1_REG1_REG_7__SCAN_IN), .S(n5312), .Z(n5304)
         );
  NOR2_X1 U6398 ( .A1(n5305), .A2(n5304), .ZN(n5303) );
  NOR2_X1 U6399 ( .A1(n5020), .A2(n5303), .ZN(n9033) );
  NAND2_X1 U6400 ( .A1(n9032), .A2(n9033), .ZN(n9031) );
  NAND2_X1 U6401 ( .A1(n5021), .A2(n9031), .ZN(n5037) );
  INV_X1 U6402 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9714) );
  INV_X1 U6403 ( .A(n6239), .ZN(n5148) );
  INV_X1 U6404 ( .A(n5023), .ZN(n5022) );
  OAI21_X1 U6405 ( .B1(n9714), .B2(n5148), .A(n5022), .ZN(n5036) );
  NOR2_X1 U6406 ( .A1(n5037), .A2(n5036), .ZN(n5035) );
  NOR2_X1 U6407 ( .A1(n5023), .A2(n5035), .ZN(n5025) );
  INV_X1 U6408 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9491) );
  INV_X1 U6409 ( .A(n6444), .ZN(n5437) );
  AOI22_X1 U6410 ( .A1(n6444), .A2(n9491), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n5437), .ZN(n5024) );
  NOR2_X1 U6411 ( .A1(n5025), .A2(n5024), .ZN(n5436) );
  AOI21_X1 U6412 ( .B1(n5025), .B2(n5024), .A(n5436), .ZN(n5027) );
  INV_X1 U6413 ( .A(n9011), .ZN(n9016) );
  AND2_X1 U6414 ( .A1(n5026), .A2(n9016), .ZN(n9542) );
  AND2_X1 U6415 ( .A1(n9542), .A2(n9071), .ZN(n9616) );
  INV_X1 U6416 ( .A(n9616), .ZN(n9638) );
  NOR2_X1 U6417 ( .A1(n5027), .A2(n9638), .ZN(n5031) );
  INV_X1 U6418 ( .A(n9628), .ZN(n5920) );
  INV_X1 U6419 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9965) );
  INV_X1 U6420 ( .A(n5028), .ZN(n5029) );
  OAI22_X1 U6421 ( .A1(n5920), .A2(n5437), .B1(n9965), .B2(n9641), .ZN(n5030)
         );
  OR4_X1 U6422 ( .A1(n6465), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(P1_U3251)
         );
  INV_X1 U6423 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U6424 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10056), .ZN(n6269) );
  AOI211_X1 U6425 ( .C1(n4351), .C2(n5034), .A(n5033), .B(n9632), .ZN(n5041)
         );
  AOI21_X1 U6426 ( .B1(n5037), .B2(n5036), .A(n5035), .ZN(n5038) );
  NOR2_X1 U6427 ( .A1(n9638), .A2(n5038), .ZN(n5040) );
  INV_X1 U6428 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10090) );
  OAI22_X1 U6429 ( .A1(n5920), .A2(n5148), .B1(n10090), .B2(n9641), .ZN(n5039)
         );
  OR4_X1 U6430 ( .A1(n6269), .A2(n5041), .A3(n5040), .A4(n5039), .ZN(P1_U3250)
         );
  NAND2_X1 U6431 ( .A1(n7355), .A2(n4258), .ZN(n9478) );
  INV_X1 U6432 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5327) );
  NOR2_X1 U6433 ( .A1(n7355), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9481) );
  AND2_X1 U6434 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5043) );
  INV_X1 U6435 ( .A(SI_1_), .ZN(n5044) );
  XNOR2_X1 U6436 ( .A(n5045), .B(n5044), .ZN(n5055) );
  NAND2_X1 U6437 ( .A1(n5045), .A2(SI_1_), .ZN(n5046) );
  INV_X1 U6438 ( .A(SI_2_), .ZN(n5048) );
  XNOR2_X1 U6439 ( .A(n5050), .B(n5049), .ZN(n5740) );
  OAI222_X1 U6440 ( .A1(n9478), .A2(n5327), .B1(n7551), .B2(n5740), .C1(
        P1_U3084), .C2(n5330), .ZN(P1_U3351) );
  NAND2_X1 U6441 ( .A1(n5050), .A2(n5049), .ZN(n5053) );
  NAND2_X1 U6442 ( .A1(n5051), .A2(SI_2_), .ZN(n5052) );
  MUX2_X1 U6443 ( .A(n5779), .B(n5502), .S(n7333), .Z(n5061) );
  XNOR2_X1 U6444 ( .A(n5060), .B(n5059), .ZN(n5776) );
  OAI222_X1 U6445 ( .A1(n9478), .A2(n5502), .B1(n7551), .B2(n5776), .C1(n4258), 
        .C2(n5647), .ZN(P1_U3350) );
  NAND2_X1 U6446 ( .A1(n7333), .A2(P2_U3152), .ZN(n8539) );
  AND2_X1 U6447 ( .A1(n7355), .A2(P2_U3152), .ZN(n8537) );
  INV_X1 U6448 ( .A(n8537), .ZN(n7920) );
  XNOR2_X1 U6449 ( .A(n5055), .B(n5054), .ZN(n5618) );
  NAND2_X1 U6450 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5056) );
  INV_X1 U6451 ( .A(n5057), .ZN(n5058) );
  OAI222_X1 U6452 ( .A1(n8539), .A2(n4410), .B1(n7920), .B2(n5618), .C1(
        P2_U3152), .C2(n6828), .ZN(P2_U3357) );
  INV_X1 U6453 ( .A(n9478), .ZN(n5694) );
  INV_X1 U6454 ( .A(n5694), .ZN(n7154) );
  INV_X1 U6455 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5368) );
  OAI222_X1 U6456 ( .A1(n7154), .A2(n5368), .B1(n7551), .B2(n5618), .C1(
        P1_U3084), .C2(n5367), .ZN(P1_U3352) );
  NAND2_X1 U6457 ( .A1(n5060), .A2(n5059), .ZN(n5064) );
  INV_X1 U6458 ( .A(n5061), .ZN(n5062) );
  NAND2_X1 U6459 ( .A1(n5062), .A2(SI_3_), .ZN(n5063) );
  NAND2_X2 U6460 ( .A1(n5064), .A2(n5063), .ZN(n5066) );
  XNOR2_X1 U6461 ( .A(n5066), .B(n5065), .ZN(n5789) );
  OAI222_X1 U6462 ( .A1(n9478), .A2(n5534), .B1(n7551), .B2(n5789), .C1(n4258), 
        .C2(n9555), .ZN(P1_U3349) );
  XNOR2_X1 U6463 ( .A(n5079), .B(n5078), .ZN(n5986) );
  INV_X1 U6464 ( .A(n5069), .ZN(n5704) );
  OAI222_X1 U6465 ( .A1(n9478), .A2(n5701), .B1(n7551), .B2(n5986), .C1(
        P1_U3084), .C2(n5704), .ZN(P1_U3348) );
  INV_X1 U6466 ( .A(n8539), .ZN(n6696) );
  INV_X1 U6467 ( .A(n6696), .ZN(n8533) );
  INV_X1 U6468 ( .A(n8537), .ZN(n8543) );
  OR2_X1 U6469 ( .A1(n5057), .A2(n5224), .ZN(n5070) );
  XNOR2_X1 U6470 ( .A(n5070), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6085) );
  INV_X1 U6471 ( .A(n6085), .ZN(n6790) );
  OAI222_X1 U6472 ( .A1(n8533), .A2(n4755), .B1(n8543), .B2(n5740), .C1(
        P2_U3152), .C2(n6790), .ZN(P2_U3356) );
  INV_X1 U6473 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6474 ( .A1(n5071), .A2(n5072), .ZN(n5108) );
  NAND2_X1 U6475 ( .A1(n5108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U6476 ( .A(n5082), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6089) );
  INV_X1 U6477 ( .A(n6089), .ZN(n6399) );
  OAI222_X1 U6478 ( .A1(n8533), .A2(n5073), .B1(n7920), .B2(n5986), .C1(
        P2_U3152), .C2(n6399), .ZN(P2_U3353) );
  OR2_X1 U6479 ( .A1(n5071), .A2(n5224), .ZN(n5074) );
  XNOR2_X1 U6480 ( .A(n5074), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6426) );
  INV_X1 U6481 ( .A(n6426), .ZN(n6440) );
  OAI222_X1 U6482 ( .A1(n8533), .A2(n5792), .B1(n7920), .B2(n5789), .C1(
        P2_U3152), .C2(n6440), .ZN(P2_U3354) );
  NOR2_X1 U6483 ( .A1(n5075), .A2(n5224), .ZN(n5076) );
  MUX2_X1 U6484 ( .A(n5224), .B(n5076), .S(P2_IR_REG_3__SCAN_IN), .Z(n5077) );
  NOR2_X1 U6485 ( .A1(n5077), .A2(n5071), .ZN(n6086) );
  INV_X1 U6486 ( .A(n6086), .ZN(n6423) );
  OAI222_X1 U6487 ( .A1(n8533), .A2(n5779), .B1(n8543), .B2(n5776), .C1(
        P2_U3152), .C2(n6423), .ZN(P2_U3355) );
  INV_X1 U6488 ( .A(n5080), .ZN(n5081) );
  XNOR2_X1 U6489 ( .A(n5087), .B(n5086), .ZN(n6028) );
  INV_X1 U6490 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6491 ( .A1(n5082), .A2(n5105), .ZN(n5083) );
  NAND2_X1 U6492 ( .A1(n5083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5084) );
  INV_X1 U6493 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6494 ( .A1(n5084), .A2(n5106), .ZN(n5091) );
  OR2_X1 U6495 ( .A1(n5084), .A2(n5106), .ZN(n5085) );
  INV_X1 U6496 ( .A(n6079), .ZN(n6803) );
  OAI222_X1 U6497 ( .A1(n8533), .A2(n6031), .B1(n7920), .B2(n6028), .C1(
        P2_U3152), .C2(n6803), .ZN(P2_U3352) );
  OAI222_X1 U6498 ( .A1(n9478), .A2(n9976), .B1(n7551), .B2(n6028), .C1(n4258), 
        .C2(n5848), .ZN(P1_U3347) );
  INV_X1 U6499 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6500 ( .A1(n5089), .A2(SI_6_), .ZN(n5090) );
  MUX2_X1 U6501 ( .A(n6193), .B(n5947), .S(n7333), .Z(n5096) );
  NAND2_X1 U6502 ( .A1(n5091), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U6503 ( .A(n5092), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6837) );
  INV_X1 U6504 ( .A(n6837), .ZN(n5093) );
  OAI222_X1 U6505 ( .A1(n8533), .A2(n6193), .B1(n8543), .B2(n6191), .C1(
        P2_U3152), .C2(n5093), .ZN(P2_U3351) );
  INV_X1 U6506 ( .A(n5312), .ZN(n5950) );
  OAI222_X1 U6507 ( .A1(n9478), .A2(n5947), .B1(n7551), .B2(n6191), .C1(
        P1_U3084), .C2(n5950), .ZN(P1_U3346) );
  INV_X1 U6508 ( .A(n5096), .ZN(n5097) );
  NAND2_X1 U6509 ( .A1(n5097), .A2(SI_7_), .ZN(n5113) );
  INV_X1 U6510 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5098) );
  MUX2_X1 U6511 ( .A(n9978), .B(n5098), .S(n7333), .Z(n5100) );
  INV_X1 U6512 ( .A(SI_8_), .ZN(n5099) );
  INV_X1 U6513 ( .A(n5100), .ZN(n5101) );
  NAND2_X1 U6514 ( .A1(n5101), .A2(SI_8_), .ZN(n5102) );
  INV_X1 U6515 ( .A(n6282), .ZN(n5111) );
  AOI22_X1 U6516 ( .A1(n9028), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n5694), .ZN(n5103) );
  OAI21_X1 U6517 ( .B1(n5111), .B2(n7551), .A(n5103), .ZN(P1_U3345) );
  NAND3_X1 U6518 ( .A1(n5106), .A2(n5105), .A3(n5104), .ZN(n5107) );
  OR2_X1 U6519 ( .A1(n5108), .A2(n5107), .ZN(n5123) );
  NAND2_X1 U6520 ( .A1(n5123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5110) );
  INV_X1 U6521 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5109) );
  XNOR2_X1 U6522 ( .A(n5110), .B(n5109), .ZN(n6861) );
  OAI222_X1 U6523 ( .A1(n8533), .A2(n9978), .B1(n8543), .B2(n5111), .C1(
        P2_U3152), .C2(n6861), .ZN(P2_U3350) );
  INV_X1 U6524 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5118) );
  INV_X1 U6525 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5150) );
  MUX2_X1 U6526 ( .A(n5118), .B(n5150), .S(n7333), .Z(n5120) );
  INV_X1 U6527 ( .A(SI_9_), .ZN(n5119) );
  INV_X1 U6528 ( .A(n5120), .ZN(n5121) );
  NAND2_X1 U6529 ( .A1(n5121), .A2(SI_9_), .ZN(n5122) );
  XNOR2_X1 U6530 ( .A(n5167), .B(n4883), .ZN(n6333) );
  INV_X1 U6531 ( .A(n6333), .ZN(n5149) );
  NOR2_X1 U6532 ( .A1(n5123), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5223) );
  OR2_X1 U6533 ( .A1(n5223), .A2(n5224), .ZN(n5176) );
  XNOR2_X1 U6534 ( .A(n5176), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U6535 ( .A1(n6896), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n6696), .ZN(n5124) );
  OAI21_X1 U6536 ( .B1(n5149), .B2(n7920), .A(n5124), .ZN(P2_U3349) );
  INV_X1 U6537 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5137) );
  NOR2_X1 U6538 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5127) );
  INV_X1 U6539 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5130) );
  INV_X1 U6540 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9477) );
  XNOR2_X2 U6541 ( .A(n5126), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6542 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  XNOR2_X2 U6543 ( .A(n5131), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6544 ( .A1(n7550), .A2(n5138), .ZN(n5337) );
  INV_X1 U6545 ( .A(n5337), .ZN(n5393) );
  INV_X2 U6546 ( .A(n5393), .ZN(n8753) );
  INV_X1 U6547 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5135) );
  AND2_X4 U6548 ( .A1(n7550), .A2(n7924), .ZN(n8748) );
  NAND2_X1 U6549 ( .A1(n8748), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6550 ( .A1(n7924), .A2(n5139), .ZN(n5336) );
  CLKBUF_X3 U6551 ( .A(n5336), .Z(n7783) );
  INV_X1 U6552 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5132) );
  OR2_X1 U6553 ( .A1(n7783), .A2(n5132), .ZN(n5133) );
  OAI211_X1 U6554 ( .C1(n8753), .C2(n5135), .A(n5134), .B(n5133), .ZN(n9073)
         );
  NAND2_X1 U6555 ( .A1(n9073), .A2(P1_U4006), .ZN(n5136) );
  OAI21_X1 U6556 ( .B1(P1_U4006), .B2(n5137), .A(n5136), .ZN(P1_U3586) );
  INV_X1 U6557 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5147) );
  INV_X1 U6558 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5140) );
  INV_X1 U6559 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9012) );
  OR2_X1 U6560 ( .A1(n5336), .A2(n9012), .ZN(n5144) );
  INV_X1 U6561 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6562 ( .A1(n5581), .A2(P1_U4006), .ZN(n5146) );
  OAI21_X1 U6563 ( .B1(P1_U4006), .B2(n5147), .A(n5146), .ZN(P1_U3555) );
  OAI222_X1 U6564 ( .A1(n7154), .A2(n5150), .B1(n7551), .B2(n5149), .C1(n5148), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  NAND2_X1 U6565 ( .A1(n6053), .A2(n9821), .ZN(n9815) );
  INV_X1 U6566 ( .A(n9815), .ZN(n7545) );
  INV_X1 U6567 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6568 ( .A1(n5152), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5153) );
  MUX2_X1 U6569 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5153), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5155) );
  NAND2_X1 U6570 ( .A1(n5156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6571 ( .A1(n7547), .A2(n7367), .ZN(n5478) );
  INV_X1 U6572 ( .A(n5478), .ZN(n6056) );
  NAND2_X1 U6573 ( .A1(n7545), .A2(n6056), .ZN(n5166) );
  OR2_X1 U6574 ( .A1(n5812), .A2(P2_U3152), .ZN(n7549) );
  NAND2_X1 U6575 ( .A1(n9815), .A2(n7549), .ZN(n5164) );
  INV_X1 U6576 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5158) );
  INV_X1 U6577 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5159) );
  XNOR2_X2 U6578 ( .A(n5160), .B(n5159), .ZN(n7629) );
  NAND2_X2 U6579 ( .A1(n5163), .A2(n5192), .ZN(n7543) );
  NAND2_X1 U6580 ( .A1(n5164), .A2(n5739), .ZN(n5165) );
  AND2_X1 U6581 ( .A1(n5166), .A2(n5165), .ZN(n8106) );
  INV_X1 U6582 ( .A(n8106), .ZN(n9754) );
  NOR2_X1 U6583 ( .A1(n9754), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U6584 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5185) );
  MUX2_X1 U6585 ( .A(n10041), .B(n5185), .S(n7333), .Z(n5170) );
  INV_X1 U6586 ( .A(SI_10_), .ZN(n5169) );
  NAND2_X1 U6587 ( .A1(n5170), .A2(n5169), .ZN(n5173) );
  INV_X1 U6588 ( .A(n5170), .ZN(n5171) );
  NAND2_X1 U6589 ( .A1(n5171), .A2(SI_10_), .ZN(n5172) );
  INV_X1 U6590 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5175) );
  INV_X1 U6591 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5191) );
  MUX2_X1 U6592 ( .A(n5175), .B(n5191), .S(n7333), .Z(n5209) );
  XNOR2_X1 U6593 ( .A(n5213), .B(n5208), .ZN(n6650) );
  INV_X1 U6594 ( .A(n6650), .ZN(n5190) );
  INV_X1 U6595 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6596 ( .A1(n5176), .A2(n5221), .ZN(n5177) );
  NAND2_X1 U6597 ( .A1(n5177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5182) );
  INV_X1 U6598 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6599 ( .A1(n5182), .A2(n5220), .ZN(n5178) );
  NAND2_X1 U6600 ( .A1(n5178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5179) );
  XNOR2_X1 U6601 ( .A(n5179), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6651) );
  AOI22_X1 U6602 ( .A1(n6651), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6696), .ZN(n5180) );
  OAI21_X1 U6603 ( .B1(n5190), .B2(n8543), .A(n5180), .ZN(P2_U3347) );
  XNOR2_X1 U6604 ( .A(n5181), .B(n4885), .ZN(n6443) );
  INV_X1 U6605 ( .A(n6443), .ZN(n5184) );
  XNOR2_X1 U6606 ( .A(n5182), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6812) );
  INV_X1 U6607 ( .A(n6812), .ZN(n5183) );
  OAI222_X1 U6608 ( .A1(n8533), .A2(n10041), .B1(n7920), .B2(n5184), .C1(n5183), .C2(P2_U3152), .ZN(P2_U3348) );
  OAI222_X1 U6609 ( .A1(n7154), .A2(n5185), .B1(n7551), .B2(n5184), .C1(n5437), 
        .C2(n4258), .ZN(P1_U3343) );
  INV_X1 U6610 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6611 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6612 ( .A1(n5188), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6613 ( .A(n5189), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6496) );
  INV_X1 U6614 ( .A(n6496), .ZN(n5576) );
  OAI222_X1 U6615 ( .A1(n7154), .A2(n5191), .B1(n7551), .B2(n5190), .C1(n5576), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U6616 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5193) );
  INV_X1 U6617 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6618 ( .A1(n5196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6619 ( .A1(n4260), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6620 ( .A1(n6657), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6621 ( .A1(n7322), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5199) );
  AND3_X1 U6622 ( .A1(n5201), .A2(n5200), .A3(n5199), .ZN(n8143) );
  INV_X2 U6623 ( .A(P2_U3966), .ZN(n8071) );
  NAND2_X1 U6624 ( .A1(n8071), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5202) );
  OAI21_X1 U6625 ( .B1(n8143), .B2(n8071), .A(n5202), .ZN(P2_U3582) );
  INV_X1 U6626 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10022) );
  NAND2_X1 U6627 ( .A1(n4261), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6628 ( .A1(n6657), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6629 ( .A1(n5451), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5203) );
  AND3_X1 U6630 ( .A1(n5205), .A2(n5204), .A3(n5203), .ZN(n8116) );
  INV_X1 U6631 ( .A(n8116), .ZN(n5206) );
  NAND2_X1 U6632 ( .A1(n5206), .A2(P2_U3966), .ZN(n5207) );
  OAI21_X1 U6633 ( .B1(P2_U3966), .B2(n10022), .A(n5207), .ZN(P2_U3583) );
  INV_X1 U6634 ( .A(n5209), .ZN(n5210) );
  NAND2_X1 U6635 ( .A1(n5210), .A2(SI_11_), .ZN(n5211) );
  INV_X1 U6636 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5214) );
  INV_X1 U6637 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5230) );
  MUX2_X1 U6638 ( .A(n5214), .B(n5230), .S(n7333), .Z(n5216) );
  INV_X1 U6639 ( .A(SI_12_), .ZN(n5215) );
  INV_X1 U6640 ( .A(n5216), .ZN(n5217) );
  NAND2_X1 U6641 ( .A1(n5217), .A2(SI_12_), .ZN(n5218) );
  NAND2_X1 U6642 ( .A1(n5292), .A2(n5218), .ZN(n5290) );
  INV_X1 U6643 ( .A(n6739), .ZN(n5229) );
  AND3_X1 U6644 ( .A1(n5221), .A2(n5220), .A3(n5219), .ZN(n5222) );
  AND2_X1 U6645 ( .A1(n5223), .A2(n5222), .ZN(n5301) );
  OR2_X1 U6646 ( .A1(n5301), .A2(n5224), .ZN(n5225) );
  XNOR2_X1 U6647 ( .A(n5225), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6740) );
  AOI22_X1 U6648 ( .A1(n6740), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n6696), .ZN(n5226) );
  OAI21_X1 U6649 ( .B1(n5229), .B2(n8543), .A(n5226), .ZN(P2_U3346) );
  NAND2_X1 U6650 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  XNOR2_X1 U6651 ( .A(n5228), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6608) );
  INV_X1 U6652 ( .A(n6608), .ZN(n5439) );
  OAI222_X1 U6653 ( .A1(n7154), .A2(n5230), .B1(n7551), .B2(n5229), .C1(n4258), 
        .C2(n5439), .ZN(P1_U3341) );
  INV_X1 U6654 ( .A(n8974), .ZN(n6189) );
  NAND2_X1 U6655 ( .A1(n5232), .A2(n5233), .ZN(n5234) );
  NAND2_X1 U6656 ( .A1(n5234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5236) );
  XNOR2_X2 U6657 ( .A(n5236), .B(n5235), .ZN(n9256) );
  OR2_X1 U6658 ( .A1(n8888), .A2(n5347), .ZN(n5493) );
  AND2_X1 U6659 ( .A1(n6730), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6660 ( .A1(n7070), .A2(P1_B_REG_SCAN_IN), .ZN(n5239) );
  INV_X1 U6661 ( .A(n7158), .ZN(n5238) );
  MUX2_X1 U6662 ( .A(n5239), .B(P1_B_REG_SCAN_IN), .S(n5238), .Z(n5240) );
  NAND2_X1 U6663 ( .A1(n5240), .A2(n5241), .ZN(n9643) );
  NOR2_X1 U6664 ( .A1(n9643), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5243) );
  INV_X1 U6665 ( .A(n5241), .ZN(n7123) );
  AND2_X1 U6666 ( .A1(n7158), .A2(n7123), .ZN(n5242) );
  NOR2_X1 U6667 ( .A1(n5243), .A2(n5242), .ZN(n9646) );
  NAND2_X1 U6668 ( .A1(n5333), .A2(n9646), .ZN(n5257) );
  NAND2_X1 U6669 ( .A1(n4259), .A2(n5262), .ZN(n6172) );
  NAND2_X1 U6670 ( .A1(n7123), .A2(n7070), .ZN(n5244) );
  OAI21_X1 U6671 ( .B1(n9643), .B2(P1_D_REG_1__SCAN_IN), .A(n5244), .ZN(n5332)
         );
  INV_X1 U6672 ( .A(n5332), .ZN(n9475) );
  NOR4_X1 U6673 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5248) );
  NOR4_X1 U6674 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5247) );
  NOR4_X1 U6675 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5246) );
  NOR4_X1 U6676 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5245) );
  NAND4_X1 U6677 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n5254)
         );
  NOR2_X1 U6678 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n5252) );
  NOR4_X1 U6679 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5251) );
  NOR4_X1 U6680 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5250) );
  NOR4_X1 U6681 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5249) );
  NAND4_X1 U6682 ( .A1(n5252), .A2(n5251), .A3(n5250), .A4(n5249), .ZN(n5253)
         );
  NOR2_X1 U6683 ( .A1(n5254), .A2(n5253), .ZN(n5255) );
  NOR2_X1 U6684 ( .A1(n9643), .A2(n5255), .ZN(n5331) );
  NOR2_X1 U6685 ( .A1(n9475), .A2(n5331), .ZN(n5256) );
  OAI21_X1 U6686 ( .B1(n9696), .B2(n9256), .A(n5256), .ZN(n5275) );
  INV_X2 U6687 ( .A(n9713), .ZN(n9716) );
  INV_X1 U6688 ( .A(SI_0_), .ZN(n5259) );
  INV_X1 U6689 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5258) );
  OAI21_X1 U6690 ( .B1(n7355), .B2(n5259), .A(n5258), .ZN(n5261) );
  AND2_X1 U6691 ( .A1(n5261), .A2(n5260), .ZN(n9483) );
  INV_X1 U6692 ( .A(n6178), .ZN(n7201) );
  AND2_X1 U6693 ( .A1(n5581), .A2(n7201), .ZN(n8715) );
  NOR2_X1 U6694 ( .A1(n7194), .A2(n8715), .ZN(n8941) );
  OR2_X2 U6695 ( .A1(n5262), .A2(n8974), .ZN(n5342) );
  OR2_X1 U6696 ( .A1(n5345), .A2(n5342), .ZN(n5390) );
  INV_X1 U6697 ( .A(n5390), .ZN(n6144) );
  INV_X1 U6698 ( .A(n6172), .ZN(n5263) );
  OR3_X1 U6699 ( .A1(n8941), .A2(n6144), .A3(n5263), .ZN(n5271) );
  OR2_X1 U6700 ( .A1(n5336), .A2(n4981), .ZN(n5266) );
  INV_X1 U6701 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7202) );
  OR2_X1 U6702 ( .A1(n7863), .A2(n7202), .ZN(n5268) );
  NAND2_X1 U6703 ( .A1(n8748), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5267) );
  NAND3_X2 U6704 ( .A1(n5269), .A2(n5268), .A3(n5267), .ZN(n9002) );
  NAND2_X1 U6705 ( .A1(n9329), .A2(n9002), .ZN(n5270) );
  NAND2_X1 U6706 ( .A1(n5271), .A2(n5270), .ZN(n6179) );
  INV_X1 U6707 ( .A(n6179), .ZN(n5272) );
  OAI21_X1 U6708 ( .B1(n7201), .B2(n6172), .A(n5272), .ZN(n5276) );
  NAND2_X1 U6709 ( .A1(n5276), .A2(n9716), .ZN(n5273) );
  OAI21_X1 U6710 ( .B1(n9716), .B2(n5141), .A(n5273), .ZN(P1_U3523) );
  INV_X1 U6711 ( .A(n9646), .ZN(n5274) );
  NAND2_X1 U6712 ( .A1(n5333), .A2(n5274), .ZN(n6141) );
  INV_X2 U6713 ( .A(n9702), .ZN(n9704) );
  INV_X1 U6714 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6715 ( .A1(n5276), .A2(n9704), .ZN(n5277) );
  OAI21_X1 U6716 ( .B1(n9704), .B2(n5278), .A(n5277), .ZN(P1_U3454) );
  OAI21_X1 U6717 ( .B1(n5280), .B2(n9015), .A(n5279), .ZN(n5282) );
  INV_X1 U6718 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n5281) );
  OAI22_X1 U6719 ( .A1(n9632), .A2(n5282), .B1(n9641), .B2(n5281), .ZN(n5287)
         );
  OAI211_X1 U6720 ( .C1(n5284), .C2(n5283), .A(n9616), .B(n9007), .ZN(n5285)
         );
  OAI21_X1 U6721 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7202), .A(n5285), .ZN(n5286) );
  AOI211_X1 U6722 ( .C1(n9628), .C2(n5288), .A(n5287), .B(n5286), .ZN(n5289)
         );
  INV_X1 U6723 ( .A(n5289), .ZN(P1_U3242) );
  INV_X1 U6724 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5299) );
  INV_X1 U6725 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9992) );
  MUX2_X1 U6726 ( .A(n9992), .B(n5299), .S(n7333), .Z(n5294) );
  INV_X1 U6727 ( .A(SI_13_), .ZN(n5293) );
  NAND2_X1 U6728 ( .A1(n5294), .A2(n5293), .ZN(n5411) );
  INV_X1 U6729 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6730 ( .A1(n5295), .A2(SI_13_), .ZN(n5296) );
  XNOR2_X1 U6731 ( .A(n5410), .B(n4884), .ZN(n6871) );
  INV_X1 U6732 ( .A(n6871), .ZN(n5302) );
  OR2_X1 U6733 ( .A1(n5297), .A2(n4993), .ZN(n5298) );
  XNOR2_X1 U6734 ( .A(n5298), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9571) );
  INV_X1 U6735 ( .A(n9571), .ZN(n5912) );
  OAI222_X1 U6736 ( .A1(n7154), .A2(n5299), .B1(n7551), .B2(n5302), .C1(n5912), 
        .C2(n4258), .ZN(P1_U3340) );
  INV_X1 U6737 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6738 ( .A1(n5301), .A2(n5300), .ZN(n5683) );
  NAND2_X1 U6739 ( .A1(n5683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5415) );
  XNOR2_X1 U6740 ( .A(n5415), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6872) );
  INV_X1 U6741 ( .A(n6872), .ZN(n6631) );
  OAI222_X1 U6742 ( .A1(n8533), .A2(n9992), .B1(n7920), .B2(n5302), .C1(n6631), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  AOI21_X1 U6743 ( .B1(n5305), .B2(n5304), .A(n5303), .ZN(n5315) );
  INV_X1 U6744 ( .A(n9632), .ZN(n9553) );
  OAI21_X1 U6745 ( .B1(n5308), .B2(n5307), .A(n5306), .ZN(n5311) );
  AND2_X1 U6746 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5966) );
  INV_X1 U6747 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n5309) );
  NOR2_X1 U6748 ( .A1(n9641), .A2(n5309), .ZN(n5310) );
  AOI211_X1 U6749 ( .C1(n9553), .C2(n5311), .A(n5966), .B(n5310), .ZN(n5314)
         );
  NAND2_X1 U6750 ( .A1(n9628), .A2(n5312), .ZN(n5313) );
  OAI211_X1 U6751 ( .C1(n5315), .C2(n9638), .A(n5314), .B(n5313), .ZN(P1_U3248) );
  OAI21_X1 U6752 ( .B1(n5318), .B2(n5317), .A(n5316), .ZN(n5321) );
  AND2_X1 U6753 ( .A1(n4258), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5730) );
  INV_X1 U6754 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n5319) );
  NOR2_X1 U6755 ( .A1(n9641), .A2(n5319), .ZN(n5320) );
  AOI211_X1 U6756 ( .C1(n9553), .C2(n5321), .A(n5730), .B(n5320), .ZN(n5326)
         );
  OAI211_X1 U6757 ( .C1(n5324), .C2(n5323), .A(n9616), .B(n5322), .ZN(n5325)
         );
  OAI211_X1 U6758 ( .C1(n5920), .C2(n5704), .A(n5326), .B(n5325), .ZN(P1_U3246) );
  NAND2_X2 U6759 ( .A1(n5951), .A2(n7355), .ZN(n5533) );
  OAI211_X2 U6760 ( .C1(n5951), .C2(n5330), .A(n5329), .B(n5328), .ZN(n6481)
         );
  INV_X2 U6761 ( .A(n6481), .ZN(n9662) );
  NOR2_X1 U6762 ( .A1(n5332), .A2(n5331), .ZN(n6139) );
  AND2_X1 U6763 ( .A1(n6139), .A2(n9646), .ZN(n5391) );
  INV_X1 U6764 ( .A(n5391), .ZN(n5387) );
  NAND3_X1 U6765 ( .A1(n4888), .A2(n9648), .A3(n5387), .ZN(n5498) );
  AND2_X1 U6766 ( .A1(n5498), .A2(n5333), .ZN(n8580) );
  NAND2_X1 U6767 ( .A1(n8580), .A2(n9456), .ZN(n8653) );
  NAND2_X1 U6768 ( .A1(n6481), .A2(n5357), .ZN(n5344) );
  NAND2_X1 U6769 ( .A1(n8748), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5341) );
  INV_X1 U6770 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5334) );
  OR2_X1 U6771 ( .A1(n7863), .A2(n5334), .ZN(n5340) );
  INV_X1 U6772 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5335) );
  OR2_X1 U6773 ( .A1(n5336), .A2(n5335), .ZN(n5339) );
  OR2_X1 U6774 ( .A1(n5337), .A2(n9706), .ZN(n5338) );
  NAND2_X1 U6775 ( .A1(n9000), .A2(n5505), .ZN(n5343) );
  NAND2_X1 U6776 ( .A1(n5344), .A2(n5343), .ZN(n5346) );
  AND2_X4 U6777 ( .A1(n5345), .A2(n5342), .ZN(n7872) );
  XNOR2_X1 U6778 ( .A(n5346), .B(n7872), .ZN(n5351) );
  NAND2_X1 U6779 ( .A1(n4259), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6780 ( .A1(n5377), .A2(n9000), .ZN(n5350) );
  NAND2_X1 U6781 ( .A1(n5351), .A2(n5352), .ZN(n5500) );
  INV_X1 U6782 ( .A(n5351), .ZN(n5354) );
  NAND2_X1 U6783 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6784 ( .A1(n5581), .A2(n5505), .ZN(n5359) );
  NAND2_X1 U6785 ( .A1(n5359), .A2(n5358), .ZN(n5611) );
  INV_X1 U6786 ( .A(n5611), .ZN(n5360) );
  NAND2_X1 U6787 ( .A1(n5361), .A2(n5360), .ZN(n5366) );
  NAND2_X1 U6788 ( .A1(n4263), .A2(n5581), .ZN(n5365) );
  INV_X1 U6789 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5362) );
  NOR2_X1 U6790 ( .A1(n5494), .A2(n5362), .ZN(n5363) );
  AOI21_X1 U6791 ( .B1(n5505), .B2(n6178), .A(n5363), .ZN(n5364) );
  AND2_X1 U6792 ( .A1(n5365), .A2(n5364), .ZN(n5612) );
  INV_X1 U6793 ( .A(n5381), .ZN(n5376) );
  OAI22_X1 U6794 ( .A1(n5533), .A2(n5368), .B1(n5951), .B2(n5367), .ZN(n5369)
         );
  INV_X1 U6795 ( .A(n5369), .ZN(n5371) );
  NAND2_X1 U6796 ( .A1(n7204), .A2(n5357), .ZN(n5373) );
  NAND2_X1 U6797 ( .A1(n9002), .A2(n5505), .ZN(n5372) );
  NAND2_X1 U6798 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  XNOR2_X1 U6799 ( .A(n5374), .B(n7872), .ZN(n5380) );
  INV_X1 U6800 ( .A(n5380), .ZN(n5375) );
  NAND2_X1 U6801 ( .A1(n5376), .A2(n5375), .ZN(n5402) );
  NAND2_X1 U6802 ( .A1(n5377), .A2(n9002), .ZN(n5379) );
  NAND2_X1 U6803 ( .A1(n4264), .A2(n7204), .ZN(n5378) );
  AND2_X1 U6804 ( .A1(n5379), .A2(n5378), .ZN(n5405) );
  NAND2_X1 U6805 ( .A1(n5402), .A2(n5405), .ZN(n5382) );
  NAND2_X1 U6806 ( .A1(n5381), .A2(n5380), .ZN(n5403) );
  OAI21_X1 U6807 ( .B1(n5383), .B2(n5384), .A(n5501), .ZN(n5386) );
  AND2_X1 U6808 ( .A1(n8888), .A2(n9648), .ZN(n5385) );
  NAND3_X1 U6809 ( .A1(n5385), .A2(n9694), .A3(n5391), .ZN(n8664) );
  INV_X1 U6810 ( .A(n8664), .ZN(n8647) );
  NAND2_X1 U6811 ( .A1(n5386), .A2(n8647), .ZN(n5401) );
  NAND2_X1 U6812 ( .A1(n9694), .A2(n5387), .ZN(n5495) );
  NAND2_X1 U6813 ( .A1(n8580), .A2(n5495), .ZN(n5616) );
  NAND2_X1 U6814 ( .A1(n9648), .A2(n9016), .ZN(n5388) );
  NOR2_X1 U6815 ( .A1(n5390), .A2(n5388), .ZN(n8980) );
  INV_X1 U6816 ( .A(n8668), .ZN(n8598) );
  INV_X1 U6817 ( .A(n9002), .ZN(n5614) );
  NAND2_X1 U6818 ( .A1(n9648), .A2(n9011), .ZN(n5389) );
  NOR2_X1 U6819 ( .A1(n5390), .A2(n5389), .ZN(n5392) );
  AND2_X1 U6820 ( .A1(n5392), .A2(n5391), .ZN(n8659) );
  INV_X1 U6821 ( .A(n8659), .ZN(n8666) );
  NAND2_X1 U6822 ( .A1(n8748), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5398) );
  OR2_X1 U6823 ( .A1(n7863), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5397) );
  OR2_X1 U6824 ( .A1(n7783), .A2(n4990), .ZN(n5396) );
  OR2_X1 U6825 ( .A1(n5337), .A2(n5394), .ZN(n5395) );
  NAND4_X1 U6826 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n8999)
         );
  INV_X1 U6827 ( .A(n8999), .ZN(n5830) );
  OAI22_X1 U6828 ( .A1(n8598), .A2(n5614), .B1(n8666), .B2(n5830), .ZN(n5399)
         );
  AOI21_X1 U6829 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n5616), .A(n5399), .ZN(
        n5400) );
  OAI211_X1 U6830 ( .C1(n9662), .C2(n8653), .A(n5401), .B(n5400), .ZN(P1_U3235) );
  NAND2_X1 U6831 ( .A1(n5402), .A2(n5403), .ZN(n5404) );
  XNOR2_X1 U6832 ( .A(n5405), .B(n5404), .ZN(n5409) );
  NOR2_X1 U6833 ( .A1(n9694), .A2(n4598), .ZN(n9650) );
  INV_X1 U6834 ( .A(n5581), .ZN(n7196) );
  INV_X1 U6835 ( .A(n9000), .ZN(n7195) );
  OAI22_X1 U6836 ( .A1(n8598), .A2(n7196), .B1(n8666), .B2(n7195), .ZN(n5406)
         );
  AOI21_X1 U6837 ( .B1(n8580), .B2(n9650), .A(n5406), .ZN(n5408) );
  NAND2_X1 U6838 ( .A1(n5616), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5407) );
  OAI211_X1 U6839 ( .C1(n5409), .C2(n8664), .A(n5408), .B(n5407), .ZN(P1_U3220) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5414) );
  INV_X1 U6841 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5418) );
  MUX2_X1 U6842 ( .A(n5418), .B(n5414), .S(n7333), .Z(n5649) );
  XNOR2_X1 U6843 ( .A(n5649), .B(SI_14_), .ZN(n5648) );
  XNOR2_X1 U6844 ( .A(n5653), .B(n5648), .ZN(n7090) );
  INV_X1 U6845 ( .A(n7090), .ZN(n5417) );
  OR2_X1 U6846 ( .A1(n5413), .A2(n4993), .ZN(n5670) );
  XNOR2_X1 U6847 ( .A(n5670), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6905) );
  INV_X1 U6848 ( .A(n6905), .ZN(n9049) );
  OAI222_X1 U6849 ( .A1(n7154), .A2(n5414), .B1(n7551), .B2(n5417), .C1(n9049), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U6850 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6851 ( .A1(n5415), .A2(n5679), .ZN(n5416) );
  NAND2_X1 U6852 ( .A1(n5416), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5674) );
  XNOR2_X1 U6853 ( .A(n5674), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7091) );
  INV_X1 U6854 ( .A(n7091), .ZN(n6950) );
  OAI222_X1 U6855 ( .A1(n8539), .A2(n5418), .B1(n7920), .B2(n5417), .C1(n6950), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U6856 ( .A1(n5991), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6040) );
  INV_X1 U6857 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6039) );
  NOR2_X1 U6858 ( .A1(n6040), .A2(n6039), .ZN(n6203) );
  NAND2_X1 U6859 ( .A1(n6203), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6295) );
  INV_X1 U6860 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6294) );
  INV_X1 U6861 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6364) );
  NOR2_X1 U6862 ( .A1(n6348), .A2(n6364), .ZN(n6355) );
  NAND2_X1 U6863 ( .A1(n6355), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6655) );
  INV_X1 U6864 ( .A(n6655), .ZN(n5419) );
  NAND2_X1 U6865 ( .A1(n5419), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6744) );
  INV_X1 U6866 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6743) );
  INV_X1 U6867 ( .A(n6876), .ZN(n5420) );
  NAND2_X1 U6868 ( .A1(n5420), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U6869 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5421) );
  INV_X1 U6870 ( .A(n7216), .ZN(n5422) );
  NAND2_X1 U6871 ( .A1(n5422), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U6872 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5423) );
  INV_X1 U6873 ( .A(n7241), .ZN(n5424) );
  NAND2_X1 U6874 ( .A1(n5424), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U6875 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5425) );
  INV_X1 U6876 ( .A(n7264), .ZN(n5426) );
  NAND2_X1 U6877 ( .A1(n5426), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7273) );
  INV_X1 U6878 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8011) );
  INV_X1 U6879 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10013) );
  INV_X1 U6880 ( .A(n7292), .ZN(n5427) );
  NAND2_X1 U6881 ( .A1(n5427), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7303) );
  INV_X1 U6882 ( .A(n7303), .ZN(n5428) );
  NAND2_X1 U6883 ( .A1(n5428), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7319) );
  INV_X1 U6884 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7318) );
  OR2_X1 U6885 ( .A1(n7319), .A2(n7318), .ZN(n7321) );
  INV_X1 U6886 ( .A(n7321), .ZN(n8148) );
  INV_X1 U6887 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5433) );
  INV_X1 U6888 ( .A(n4260), .ZN(n7325) );
  NAND2_X1 U6889 ( .A1(n5451), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6890 ( .A1(n6657), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5431) );
  OAI211_X1 U6891 ( .C1(n5433), .C2(n7325), .A(n5432), .B(n5431), .ZN(n5434)
         );
  AOI21_X1 U6892 ( .B1(n8148), .B2(n7328), .A(n5434), .ZN(n7623) );
  NAND2_X1 U6893 ( .A1(n8071), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5435) );
  OAI21_X1 U6894 ( .B1(n7623), .B2(n8071), .A(n5435), .ZN(P2_U3581) );
  INV_X1 U6895 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9531) );
  AOI21_X1 U6896 ( .B1(n5437), .B2(n9491), .A(n5436), .ZN(n5571) );
  AOI22_X1 U6897 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n5576), .B1(n6496), .B2(
        n9531), .ZN(n5570) );
  NOR2_X1 U6898 ( .A1(n5571), .A2(n5570), .ZN(n5569) );
  AOI21_X1 U6899 ( .B1(n9531), .B2(n5576), .A(n5569), .ZN(n5441) );
  INV_X1 U6900 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5438) );
  AOI22_X1 U6901 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n5439), .B1(n6608), .B2(
        n5438), .ZN(n5440) );
  NOR2_X1 U6902 ( .A1(n5441), .A2(n5440), .ZN(n5909) );
  AOI21_X1 U6903 ( .B1(n5441), .B2(n5440), .A(n5909), .ZN(n5450) );
  INV_X1 U6904 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6905 ( .A1(n4258), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6938) );
  OAI21_X1 U6906 ( .B1(n9641), .B2(n5442), .A(n6938), .ZN(n5448) );
  INV_X1 U6907 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U6908 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6496), .B1(n5576), .B2(
        n6514), .ZN(n5574) );
  NAND2_X1 U6909 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6608), .ZN(n5444) );
  OAI21_X1 U6910 ( .B1(n6608), .B2(P1_REG2_REG_12__SCAN_IN), .A(n5444), .ZN(
        n5445) );
  NOR2_X1 U6911 ( .A1(n5445), .A2(n5446), .ZN(n5915) );
  AOI211_X1 U6912 ( .C1(n5446), .C2(n5445), .A(n5915), .B(n9632), .ZN(n5447)
         );
  AOI211_X1 U6913 ( .C1(n9628), .C2(n6608), .A(n5448), .B(n5447), .ZN(n5449)
         );
  OAI21_X1 U6914 ( .B1(n5450), .B2(n9638), .A(n5449), .ZN(P1_U3253) );
  NAND2_X1 U6915 ( .A1(n7328), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6916 ( .A1(n7275), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6917 ( .A1(n5451), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6918 ( .A1(n6657), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5452) );
  INV_X1 U6919 ( .A(n8072), .ZN(n7555) );
  NAND2_X1 U6920 ( .A1(n7355), .A2(SI_0_), .ZN(n5456) );
  XNOR2_X1 U6921 ( .A(n5456), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8544) );
  MUX2_X1 U6922 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8544), .S(n6283), .Z(n7554) );
  NAND2_X1 U6923 ( .A1(n7555), .A2(n7554), .ZN(n5743) );
  INV_X1 U6924 ( .A(n7554), .ZN(n9823) );
  NAND2_X1 U6925 ( .A1(n8072), .A2(n9823), .ZN(n7370) );
  NAND2_X1 U6926 ( .A1(n5743), .A2(n7370), .ZN(n7504) );
  INV_X1 U6927 ( .A(n7504), .ZN(n9825) );
  XNOR2_X1 U6928 ( .A(n6849), .B(P2_B_REG_SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6929 ( .A1(n5457), .A2(n7071), .ZN(n5459) );
  INV_X1 U6930 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9817) );
  AND2_X1 U6931 ( .A1(n6849), .A2(n7126), .ZN(n9818) );
  AOI21_X1 U6932 ( .B1(n9814), .B2(n9817), .A(n9818), .ZN(n5904) );
  INV_X1 U6933 ( .A(n5904), .ZN(n5896) );
  INV_X1 U6934 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U6935 ( .A1(n9814), .A2(n9820), .ZN(n5461) );
  AND2_X1 U6936 ( .A1(n7071), .A2(n7126), .ZN(n9822) );
  INV_X1 U6937 ( .A(n9822), .ZN(n5460) );
  NAND2_X1 U6938 ( .A1(n5461), .A2(n5460), .ZN(n5894) );
  INV_X1 U6939 ( .A(n5894), .ZN(n5805) );
  NOR4_X1 U6940 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5465) );
  NOR4_X1 U6941 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5464) );
  NOR4_X1 U6942 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5463) );
  NOR4_X1 U6943 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5462) );
  NAND4_X1 U6944 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n5471)
         );
  NOR2_X1 U6945 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n5469) );
  NOR4_X1 U6946 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5468) );
  NOR4_X1 U6947 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5467) );
  NOR4_X1 U6948 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5466) );
  NAND4_X1 U6949 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n5470)
         );
  OAI21_X1 U6950 ( .B1(n5471), .B2(n5470), .A(n9814), .ZN(n5804) );
  NAND2_X1 U6951 ( .A1(n5472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5477) );
  INV_X1 U6952 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6953 ( .A1(n5477), .A2(n5476), .ZN(n5473) );
  NAND2_X1 U6954 ( .A1(n5473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5475) );
  INV_X1 U6955 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U6956 ( .A(n5475), .B(n5474), .ZN(n7506) );
  XNOR2_X1 U6957 ( .A(n5477), .B(n5476), .ZN(n8198) );
  AND2_X1 U6958 ( .A1(n7506), .A2(n8198), .ZN(n7544) );
  NOR2_X1 U6959 ( .A1(n5478), .A2(n7544), .ZN(n7552) );
  NOR2_X1 U6960 ( .A1(n9815), .A2(n7552), .ZN(n5479) );
  AND2_X1 U6961 ( .A1(n5804), .A2(n5479), .ZN(n5895) );
  NAND3_X1 U6962 ( .A1(n5896), .A2(n5805), .A3(n5895), .ZN(n5488) );
  AND2_X2 U6963 ( .A1(n5489), .A2(n7506), .ZN(n9878) );
  NAND2_X1 U6964 ( .A1(n9878), .A2(n4643), .ZN(n5893) );
  INV_X1 U6965 ( .A(n5893), .ZN(n5480) );
  NAND2_X1 U6966 ( .A1(n7545), .A2(n5480), .ZN(n9788) );
  AND2_X1 U6967 ( .A1(n7506), .A2(n7367), .ZN(n5761) );
  XNOR2_X1 U6968 ( .A(n6601), .B(n5761), .ZN(n5481) );
  NAND2_X1 U6969 ( .A1(n5481), .A2(n8198), .ZN(n9790) );
  NAND2_X1 U6970 ( .A1(n5761), .A2(n4643), .ZN(n5927) );
  NAND2_X1 U6971 ( .A1(n9790), .A2(n5927), .ZN(n9770) );
  NAND2_X1 U6972 ( .A1(n9783), .A2(n9770), .ZN(n8412) );
  NAND2_X1 U6973 ( .A1(n7547), .A2(n4643), .ZN(n7536) );
  INV_X1 U6974 ( .A(n7506), .ZN(n7535) );
  NAND2_X1 U6975 ( .A1(n7535), .A2(n7367), .ZN(n7365) );
  AND2_X1 U6976 ( .A1(n7536), .A2(n7365), .ZN(n9795) );
  NAND2_X1 U6977 ( .A1(n4261), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6978 ( .A1(n7328), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6979 ( .A1(n6657), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6980 ( .A1(n5451), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5482) );
  AND2_X1 U6981 ( .A1(n7629), .A2(n6056), .ZN(n9775) );
  OAI22_X1 U6982 ( .A1(n9825), .A2(n9795), .B1(n7560), .B2(n8404), .ZN(n9827)
         );
  INV_X1 U6983 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9755) );
  INV_X1 U6984 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5486) );
  OAI22_X1 U6985 ( .A1(n9783), .A2(n9755), .B1(n5486), .B2(n9788), .ZN(n5487)
         );
  AOI21_X1 U6986 ( .B1(n9827), .B2(n9783), .A(n5487), .ZN(n5492) );
  OR2_X1 U6987 ( .A1(n5488), .A2(n4643), .ZN(n6001) );
  INV_X1 U6988 ( .A(n6001), .ZN(n8344) );
  NAND2_X1 U6989 ( .A1(n8344), .A2(n9878), .ZN(n8369) );
  OR2_X1 U6990 ( .A1(n9824), .A2(n7506), .ZN(n9782) );
  INV_X1 U6991 ( .A(n9782), .ZN(n5490) );
  NAND2_X1 U6992 ( .A1(n9783), .A2(n5490), .ZN(n8398) );
  INV_X1 U6993 ( .A(n8398), .ZN(n9803) );
  OAI21_X1 U6994 ( .B1(n9809), .B2(n9803), .A(n7554), .ZN(n5491) );
  OAI211_X1 U6995 ( .C1(n9825), .C2(n8412), .A(n5492), .B(n5491), .ZN(P2_U3296) );
  AND3_X1 U6996 ( .A1(n5494), .A2(n6730), .A3(n5493), .ZN(n5496) );
  NAND2_X1 U6997 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  NAND2_X1 U6998 ( .A1(n5497), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6999 ( .A1(n5377), .A2(n8999), .ZN(n5507) );
  OR2_X1 U7000 ( .A1(n5533), .A2(n5502), .ZN(n5504) );
  OR2_X1 U7001 ( .A1(n5535), .A2(n5776), .ZN(n5503) );
  OAI211_X1 U7002 ( .C1(n5951), .C2(n5647), .A(n5504), .B(n5503), .ZN(n5602)
         );
  NAND2_X1 U7003 ( .A1(n7891), .A2(n5602), .ZN(n5506) );
  AND2_X1 U7004 ( .A1(n5507), .A2(n5506), .ZN(n5513) );
  NAND2_X1 U7005 ( .A1(n8999), .A2(n4264), .ZN(n5509) );
  NAND2_X1 U7006 ( .A1(n5602), .A2(n7889), .ZN(n5508) );
  NAND2_X1 U7007 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  XNOR2_X1 U7008 ( .A(n5510), .B(n7872), .ZN(n5512) );
  NAND2_X1 U7009 ( .A1(n5511), .A2(n5516), .ZN(n5532) );
  INV_X1 U7010 ( .A(n5512), .ZN(n5515) );
  INV_X1 U7011 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U7012 ( .A1(n5515), .A2(n5514), .ZN(n5531) );
  INV_X1 U7013 ( .A(n5531), .ZN(n5520) );
  INV_X1 U7014 ( .A(n5516), .ZN(n5518) );
  OAI21_X1 U7015 ( .B1(n5520), .B2(n5518), .A(n5517), .ZN(n5519) );
  OAI211_X1 U7016 ( .C1(n5532), .C2(n5520), .A(n8647), .B(n5519), .ZN(n5530)
         );
  NAND2_X1 U7017 ( .A1(n8748), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5526) );
  OR2_X1 U7018 ( .A1(n8753), .A2(n5521), .ZN(n5525) );
  XNOR2_X1 U7019 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6152) );
  OR2_X1 U7020 ( .A1(n7863), .A2(n6152), .ZN(n5524) );
  OR2_X1 U7021 ( .A1(n7783), .A2(n5522), .ZN(n5523) );
  NAND4_X1 U7022 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n8998)
         );
  AND2_X1 U7023 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5639) );
  AOI21_X1 U7024 ( .B1(n8659), .B2(n8998), .A(n5639), .ZN(n5527) );
  OAI21_X1 U7025 ( .B1(n8598), .B2(n7195), .A(n5527), .ZN(n5528) );
  AOI21_X1 U7026 ( .B1(n8679), .B2(n5602), .A(n5528), .ZN(n5529) );
  OAI211_X1 U7027 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8671), .A(n5530), .B(
        n5529), .ZN(P1_U3216) );
  NAND2_X1 U7028 ( .A1(n5532), .A2(n5531), .ZN(n5713) );
  NAND2_X1 U7029 ( .A1(n8998), .A2(n7891), .ZN(n5538) );
  OR2_X1 U7030 ( .A1(n8758), .A2(n5534), .ZN(n5536) );
  NAND2_X1 U7031 ( .A1(n5837), .A2(n7889), .ZN(n5537) );
  NAND2_X1 U7032 ( .A1(n5538), .A2(n5537), .ZN(n5539) );
  NAND2_X1 U7033 ( .A1(n5377), .A2(n8998), .ZN(n5541) );
  NAND2_X1 U7034 ( .A1(n7891), .A2(n5837), .ZN(n5540) );
  NAND2_X1 U7035 ( .A1(n5541), .A2(n5540), .ZN(n5709) );
  INV_X1 U7036 ( .A(n5709), .ZN(n5707) );
  XNOR2_X1 U7037 ( .A(n5710), .B(n5707), .ZN(n5542) );
  XNOR2_X1 U7038 ( .A(n5713), .B(n5542), .ZN(n5555) );
  INV_X1 U7039 ( .A(n7863), .ZN(n7897) );
  AOI21_X1 U7040 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5543) );
  NOR2_X1 U7041 ( .A1(n5543), .A2(n5724), .ZN(n6132) );
  NAND2_X1 U7042 ( .A1(n7897), .A2(n6132), .ZN(n5550) );
  INV_X1 U7043 ( .A(n8748), .ZN(n7824) );
  INV_X1 U7044 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5544) );
  OR2_X1 U7045 ( .A1(n7824), .A2(n5544), .ZN(n5549) );
  OR2_X1 U7046 ( .A1(n8753), .A2(n5545), .ZN(n5548) );
  INV_X1 U7047 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5546) );
  OR2_X1 U7048 ( .A1(n7783), .A2(n5546), .ZN(n5547) );
  NAND4_X1 U7049 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n8997)
         );
  AND2_X1 U7050 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9559) );
  AOI21_X1 U7051 ( .B1(n8659), .B2(n8997), .A(n9559), .ZN(n5551) );
  OAI21_X1 U7052 ( .B1(n8598), .B2(n5830), .A(n5551), .ZN(n5553) );
  NOR2_X1 U7053 ( .A1(n8671), .A2(n6152), .ZN(n5552) );
  AOI211_X1 U7054 ( .C1(n8679), .C2(n5837), .A(n5553), .B(n5552), .ZN(n5554)
         );
  OAI21_X1 U7055 ( .B1(n5555), .B2(n8664), .A(n5554), .ZN(P1_U3228) );
  AOI211_X1 U7056 ( .C1(n5558), .C2(n5557), .A(n5556), .B(n9632), .ZN(n5568)
         );
  AOI21_X1 U7057 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(n5562) );
  OAI22_X1 U7058 ( .A1(n5848), .A2(n5920), .B1(n9638), .B2(n5562), .ZN(n5567)
         );
  INV_X1 U7059 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n5565) );
  INV_X1 U7060 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5563) );
  NOR2_X1 U7061 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5563), .ZN(n5867) );
  INV_X1 U7062 ( .A(n5867), .ZN(n5564) );
  OAI21_X1 U7063 ( .B1(n9641), .B2(n5565), .A(n5564), .ZN(n5566) );
  OR3_X1 U7064 ( .A1(n5568), .A2(n5567), .A3(n5566), .ZN(P1_U3247) );
  AOI21_X1 U7065 ( .B1(n5571), .B2(n5570), .A(n5569), .ZN(n5580) );
  OAI21_X1 U7066 ( .B1(n5574), .B2(n5573), .A(n5572), .ZN(n5578) );
  INV_X1 U7067 ( .A(n9641), .ZN(n9544) );
  AND2_X1 U7068 ( .A1(n4258), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6681) );
  AOI21_X1 U7069 ( .B1(n9544), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6681), .ZN(
        n5575) );
  OAI21_X1 U7070 ( .B1(n5920), .B2(n5576), .A(n5575), .ZN(n5577) );
  AOI21_X1 U7071 ( .B1(n5578), .B2(n9553), .A(n5577), .ZN(n5579) );
  OAI21_X1 U7072 ( .B1(n5580), .B2(n9638), .A(n5579), .ZN(P1_U3252) );
  INV_X1 U7073 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5607) );
  AND2_X1 U7074 ( .A1(n5581), .A2(n6178), .ZN(n7192) );
  NAND2_X1 U7075 ( .A1(n5588), .A2(n7192), .ZN(n7191) );
  NAND2_X1 U7076 ( .A1(n9002), .A2(n7204), .ZN(n5582) );
  NAND2_X1 U7077 ( .A1(n7191), .A2(n5582), .ZN(n6470) );
  INV_X1 U7078 ( .A(n6470), .ZN(n5583) );
  NAND2_X1 U7079 ( .A1(n9000), .A2(n9662), .ZN(n8720) );
  NAND2_X2 U7080 ( .A1(n8718), .A2(n8720), .ZN(n5590) );
  NAND2_X1 U7081 ( .A1(n7195), .A2(n9662), .ZN(n5584) );
  NAND2_X1 U7082 ( .A1(n6472), .A2(n5584), .ZN(n5585) );
  NAND2_X1 U7083 ( .A1(n8999), .A2(n9368), .ZN(n8724) );
  NAND2_X1 U7084 ( .A1(n8904), .A2(n8724), .ZN(n5587) );
  NAND2_X1 U7085 ( .A1(n5585), .A2(n5587), .ZN(n5827) );
  OAI21_X1 U7086 ( .B1(n5585), .B2(n5587), .A(n5827), .ZN(n9374) );
  INV_X1 U7087 ( .A(n9374), .ZN(n5605) );
  NAND2_X1 U7088 ( .A1(n4259), .A2(n5586), .ZN(n8884) );
  OR2_X1 U7089 ( .A1(n8884), .A2(n8974), .ZN(n9653) );
  NAND2_X1 U7090 ( .A1(n5614), .A2(n7204), .ZN(n5589) );
  OAI21_X1 U7091 ( .B1(n5591), .B2(n8911), .A(n5831), .ZN(n5596) );
  OR2_X1 U7092 ( .A1(n4259), .A2(n9256), .ZN(n5593) );
  OR2_X1 U7093 ( .A1(n6189), .A2(n5262), .ZN(n5592) );
  OR2_X1 U7094 ( .A1(n8888), .A2(n9011), .ZN(n9282) );
  NAND2_X1 U7095 ( .A1(n9343), .A2(n9000), .ZN(n5594) );
  OAI21_X1 U7096 ( .B1(n4407), .B2(n9345), .A(n5594), .ZN(n5595) );
  AOI21_X1 U7097 ( .B1(n5596), .B2(n9348), .A(n5595), .ZN(n5600) );
  OR2_X1 U7098 ( .A1(n4502), .A2(n5345), .ZN(n5598) );
  NAND3_X1 U7099 ( .A1(n4259), .A2(n8968), .A3(n5347), .ZN(n5597) );
  AND2_X1 U7100 ( .A1(n5598), .A2(n5597), .ZN(n9385) );
  INV_X1 U7101 ( .A(n9385), .ZN(n7052) );
  NAND2_X1 U7102 ( .A1(n9374), .A2(n7052), .ZN(n5599) );
  NAND2_X1 U7103 ( .A1(n5600), .A2(n5599), .ZN(n9365) );
  INV_X1 U7104 ( .A(n9365), .ZN(n5604) );
  OR2_X1 U7105 ( .A1(n6479), .A2(n9368), .ZN(n5601) );
  AND2_X1 U7106 ( .A1(n5836), .A2(n5601), .ZN(n9371) );
  INV_X1 U7107 ( .A(n9696), .ZN(n9673) );
  AOI22_X1 U7108 ( .A1(n9371), .A2(n9673), .B1(n9456), .B2(n5602), .ZN(n5603)
         );
  OAI211_X1 U7109 ( .C1(n5605), .C2(n9653), .A(n5604), .B(n5603), .ZN(n5608)
         );
  NAND2_X1 U7110 ( .A1(n5608), .A2(n9704), .ZN(n5606) );
  OAI21_X1 U7111 ( .B1(n9704), .B2(n5607), .A(n5606), .ZN(P1_U3463) );
  NAND2_X1 U7112 ( .A1(n5608), .A2(n9716), .ZN(n5609) );
  OAI21_X1 U7113 ( .B1(n9716), .B2(n5394), .A(n5609), .ZN(P1_U3526) );
  OAI21_X1 U7114 ( .B1(n5612), .B2(n5611), .A(n5610), .ZN(n5613) );
  INV_X1 U7115 ( .A(n5613), .ZN(n9014) );
  OAI22_X1 U7116 ( .A1(n9014), .A2(n8664), .B1(n5614), .B2(n8666), .ZN(n5615)
         );
  AOI21_X1 U7117 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n5616), .A(n5615), .ZN(
        n5617) );
  OAI21_X1 U7118 ( .B1(n7201), .B2(n8653), .A(n5617), .ZN(P1_U3230) );
  NAND2_X1 U7119 ( .A1(n6283), .A2(n7333), .ZN(n5788) );
  INV_X1 U7120 ( .A(n6828), .ZN(n6082) );
  NAND2_X1 U7121 ( .A1(n7560), .A2(n7946), .ZN(n7375) );
  INV_X1 U7122 ( .A(n7946), .ZN(n9831) );
  NAND2_X1 U7123 ( .A1(n8070), .A2(n9831), .ZN(n7371) );
  INV_X1 U7124 ( .A(n9795), .ZN(n9771) );
  NAND2_X1 U7125 ( .A1(n5619), .A2(n9771), .ZN(n5626) );
  NAND2_X1 U7126 ( .A1(n6657), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7127 ( .A1(n7275), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7128 ( .A1(n5451), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7129 ( .A1(n7328), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5620) );
  INV_X1 U7130 ( .A(n7629), .ZN(n5624) );
  NAND2_X1 U7131 ( .A1(n5624), .A2(n6056), .ZN(n8402) );
  AOI22_X1 U7132 ( .A1(n9723), .A2(n9775), .B1(n9778), .B2(n8072), .ZN(n5625)
         );
  NAND2_X1 U7133 ( .A1(n5626), .A2(n5625), .ZN(n9832) );
  INV_X1 U7134 ( .A(n9832), .ZN(n5633) );
  INV_X1 U7135 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7136 ( .A1(n7946), .A2(n7554), .ZN(n5627) );
  NAND2_X1 U7137 ( .A1(n5627), .A2(n9878), .ZN(n5628) );
  OR2_X1 U7138 ( .A1(n5628), .A2(n5753), .ZN(n9830) );
  INV_X1 U7139 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5629) );
  OAI22_X1 U7140 ( .A1(n6001), .A2(n9830), .B1(n5629), .B2(n9788), .ZN(n5630)
         );
  AOI21_X1 U7141 ( .B1(n9813), .B2(P2_REG2_REG_1__SCAN_IN), .A(n5630), .ZN(
        n5632) );
  NAND2_X1 U7142 ( .A1(n8072), .A2(n7554), .ZN(n5736) );
  INV_X1 U7143 ( .A(n8412), .ZN(n6195) );
  AOI22_X1 U7144 ( .A1(n9834), .A2(n6195), .B1(n9803), .B2(n7946), .ZN(n5631)
         );
  OAI211_X1 U7145 ( .C1(n5633), .C2(n9813), .A(n5632), .B(n5631), .ZN(P2_U3295) );
  OAI211_X1 U7146 ( .C1(n5636), .C2(n5635), .A(n9553), .B(n5634), .ZN(n5637)
         );
  INV_X1 U7147 ( .A(n5637), .ZN(n5638) );
  AOI211_X1 U7148 ( .C1(n9544), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n5639), .B(
        n5638), .ZN(n5646) );
  MUX2_X1 U7149 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n5394), .S(n5647), .Z(n5642)
         );
  INV_X1 U7150 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7151 ( .A1(n5642), .A2(n5641), .ZN(n5644) );
  OAI211_X1 U7152 ( .C1(n9006), .C2(n5644), .A(n9616), .B(n5643), .ZN(n5645)
         );
  OAI211_X1 U7153 ( .C1(n5920), .C2(n5647), .A(n5646), .B(n5645), .ZN(P1_U3244) );
  INV_X1 U7154 ( .A(n5648), .ZN(n5652) );
  INV_X1 U7155 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7156 ( .A1(n5650), .A2(SI_14_), .ZN(n5651) );
  INV_X1 U7157 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5678) );
  INV_X1 U7158 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5673) );
  MUX2_X1 U7159 ( .A(n5678), .B(n5673), .S(n7333), .Z(n5655) );
  INV_X1 U7160 ( .A(SI_15_), .ZN(n5654) );
  NAND2_X1 U7161 ( .A1(n5655), .A2(n5654), .ZN(n5658) );
  INV_X1 U7162 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7163 ( .A1(n5656), .A2(SI_15_), .ZN(n5657) );
  NAND2_X1 U7164 ( .A1(n5658), .A2(n5657), .ZN(n5667) );
  INV_X1 U7165 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5686) );
  INV_X1 U7166 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5659) );
  MUX2_X1 U7167 ( .A(n5686), .B(n5659), .S(n7333), .Z(n5661) );
  INV_X1 U7168 ( .A(SI_16_), .ZN(n5660) );
  NAND2_X1 U7169 ( .A1(n5661), .A2(n5660), .ZN(n5690) );
  INV_X1 U7170 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7171 ( .A1(n5662), .A2(SI_16_), .ZN(n5663) );
  XNOR2_X1 U7172 ( .A(n5689), .B(n5688), .ZN(n7683) );
  INV_X1 U7173 ( .A(n7683), .ZN(n5687) );
  NAND2_X1 U7174 ( .A1(n5664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5665) );
  XNOR2_X1 U7175 ( .A(n5665), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9599) );
  AOI22_X1 U7176 ( .A1(n9599), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n5694), .ZN(n5666) );
  OAI21_X1 U7177 ( .B1(n5687), .B2(n7551), .A(n5666), .ZN(P1_U3337) );
  XNOR2_X1 U7178 ( .A(n5668), .B(n5667), .ZN(n7129) );
  INV_X1 U7179 ( .A(n7129), .ZN(n5677) );
  NAND2_X1 U7180 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  NAND2_X1 U7181 ( .A1(n5671), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  XNOR2_X1 U7182 ( .A(n5672), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9588) );
  INV_X1 U7183 ( .A(n9588), .ZN(n9052) );
  OAI222_X1 U7184 ( .A1(n7154), .A2(n5673), .B1(n7551), .B2(n5677), .C1(
        P1_U3084), .C2(n9052), .ZN(P1_U3338) );
  NAND2_X1 U7185 ( .A1(n5674), .A2(n5681), .ZN(n5675) );
  NAND2_X1 U7186 ( .A1(n5675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U7187 ( .A(n5676), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7169) );
  INV_X1 U7188 ( .A(n7169), .ZN(n7161) );
  OAI222_X1 U7189 ( .A1(n8533), .A2(n5678), .B1(n7920), .B2(n5677), .C1(
        P2_U3152), .C2(n7161), .ZN(P2_U3343) );
  INV_X1 U7190 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5680) );
  NAND3_X1 U7191 ( .A1(n5681), .A2(n5680), .A3(n5679), .ZN(n5682) );
  OAI21_X1 U7192 ( .B1(n5683), .B2(n5682), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5684) );
  MUX2_X1 U7193 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5684), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5685) );
  AND2_X1 U7194 ( .A1(n5685), .A2(n5696), .ZN(n8082) );
  INV_X1 U7195 ( .A(n8082), .ZN(n7173) );
  OAI222_X1 U7196 ( .A1(P2_U3152), .A2(n7173), .B1(n7920), .B2(n5687), .C1(
        n5686), .C2(n8533), .ZN(P2_U3342) );
  INV_X1 U7197 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5699) );
  INV_X1 U7198 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5692) );
  MUX2_X1 U7199 ( .A(n5699), .B(n5692), .S(n7333), .Z(n5972) );
  XNOR2_X1 U7200 ( .A(n5972), .B(SI_17_), .ZN(n5971) );
  XNOR2_X1 U7201 ( .A(n5976), .B(n5971), .ZN(n7696) );
  INV_X1 U7202 ( .A(n7696), .ZN(n5698) );
  NAND2_X1 U7203 ( .A1(n5693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7204 ( .A(n5981), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9610) );
  AOI22_X1 U7205 ( .A1(n9610), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n5694), .ZN(n5695) );
  OAI21_X1 U7206 ( .B1(n5698), .B2(n7551), .A(n5695), .ZN(P1_U3336) );
  NAND2_X1 U7207 ( .A1(n5696), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5697) );
  XNOR2_X1 U7208 ( .A(n5697), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7213) );
  INV_X1 U7209 ( .A(n7213), .ZN(n8089) );
  OAI222_X1 U7210 ( .A1(n8539), .A2(n5699), .B1(n7920), .B2(n5698), .C1(n8089), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U7211 ( .A1(n5377), .A2(n8997), .ZN(n5706) );
  OR2_X1 U7212 ( .A1(n6110), .A2(n5986), .ZN(n5703) );
  OR2_X1 U7213 ( .A1(n8758), .A2(n5701), .ZN(n5702) );
  OAI211_X1 U7214 ( .C1(n5951), .C2(n5704), .A(n5703), .B(n5702), .ZN(n6162)
         );
  NAND2_X1 U7215 ( .A1(n4264), .A2(n6162), .ZN(n5705) );
  NAND2_X1 U7216 ( .A1(n5706), .A2(n5705), .ZN(n5723) );
  INV_X1 U7217 ( .A(n5710), .ZN(n5708) );
  NAND2_X1 U7218 ( .A1(n5708), .A2(n5707), .ZN(n5712) );
  AND2_X1 U7219 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  NAND2_X1 U7220 ( .A1(n8997), .A2(n7891), .ZN(n5715) );
  NAND2_X1 U7221 ( .A1(n6162), .A2(n7889), .ZN(n5714) );
  NAND2_X1 U7222 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  XNOR2_X1 U7223 ( .A(n5716), .B(n7872), .ZN(n5717) );
  OR2_X1 U7224 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  NAND2_X1 U7225 ( .A1(n5718), .A2(n5717), .ZN(n5844) );
  INV_X1 U7226 ( .A(n5845), .ZN(n5722) );
  AOI21_X1 U7227 ( .B1(n5723), .B2(n5720), .A(n5722), .ZN(n5734) );
  INV_X1 U7228 ( .A(n8671), .ZN(n8618) );
  NAND2_X1 U7229 ( .A1(n8748), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5728) );
  OR2_X1 U7230 ( .A1(n8753), .A2(n9709), .ZN(n5727) );
  OAI21_X1 U7231 ( .B1(n5724), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5861), .ZN(
        n6174) );
  OR2_X1 U7232 ( .A1(n7863), .A2(n6174), .ZN(n5726) );
  OR2_X1 U7233 ( .A1(n7783), .A2(n4999), .ZN(n5725) );
  NAND4_X1 U7234 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n5725), .ZN(n8996)
         );
  INV_X1 U7235 ( .A(n8996), .ZN(n6559) );
  NOR2_X1 U7236 ( .A1(n8666), .A2(n6559), .ZN(n5729) );
  AOI211_X1 U7237 ( .C1(n8668), .C2(n8998), .A(n5730), .B(n5729), .ZN(n5731)
         );
  OAI21_X1 U7238 ( .B1(n9668), .B2(n8653), .A(n5731), .ZN(n5732) );
  AOI21_X1 U7239 ( .B1(n6132), .B2(n8618), .A(n5732), .ZN(n5733) );
  OAI21_X1 U7240 ( .B1(n5734), .B2(n8664), .A(n5733), .ZN(P1_U3225) );
  NAND2_X1 U7241 ( .A1(n5735), .A2(n7946), .ZN(n5738) );
  INV_X1 U7242 ( .A(n5736), .ZN(n5760) );
  NAND2_X1 U7243 ( .A1(n5760), .A2(n8070), .ZN(n5737) );
  NAND2_X1 U7244 ( .A1(n5738), .A2(n5737), .ZN(n5876) );
  NAND2_X1 U7245 ( .A1(n5739), .A2(n6085), .ZN(n5742) );
  OR2_X1 U7246 ( .A1(n6281), .A2(n5740), .ZN(n5741) );
  INV_X1 U7247 ( .A(n8039), .ZN(n5874) );
  NAND2_X1 U7248 ( .A1(n5931), .A2(n8039), .ZN(n7376) );
  XNOR2_X1 U7249 ( .A(n5745), .B(n5876), .ZN(n5901) );
  NAND2_X1 U7250 ( .A1(n7375), .A2(n5743), .ZN(n5744) );
  NAND2_X1 U7251 ( .A1(n5744), .A2(n7371), .ZN(n7372) );
  OAI21_X1 U7252 ( .B1(n5746), .B2(n7507), .A(n5881), .ZN(n5752) );
  INV_X1 U7253 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7254 ( .A1(n7328), .A2(n5747), .ZN(n5751) );
  NAND2_X1 U7255 ( .A1(n4260), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7256 ( .A1(n5451), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7257 ( .A1(n6657), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5748) );
  INV_X1 U7258 ( .A(n5877), .ZN(n8069) );
  AOI222_X1 U7259 ( .A1(n9771), .A2(n5752), .B1(n8070), .B2(n9778), .C1(n8069), 
        .C2(n9775), .ZN(n5900) );
  INV_X1 U7260 ( .A(n5900), .ZN(n5758) );
  OR2_X1 U7261 ( .A1(n5874), .A2(n5753), .ZN(n5754) );
  NAND2_X1 U7262 ( .A1(n5753), .A2(n5874), .ZN(n5935) );
  AND2_X1 U7263 ( .A1(n5754), .A2(n5935), .ZN(n5898) );
  NAND2_X1 U7264 ( .A1(n9809), .A2(n5898), .ZN(n5756) );
  INV_X1 U7265 ( .A(n9788), .ZN(n9802) );
  AOI22_X1 U7266 ( .A1(n9813), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n9802), .ZN(n5755) );
  OAI211_X1 U7267 ( .C1(n5874), .C2(n8398), .A(n5756), .B(n5755), .ZN(n5757)
         );
  AOI21_X1 U7268 ( .B1(n5758), .B2(n9783), .A(n5757), .ZN(n5759) );
  OAI21_X1 U7269 ( .B1(n8412), .B2(n5901), .A(n5759), .ZN(P2_U3294) );
  AND2_X2 U7270 ( .A1(n9878), .A2(n8198), .ZN(n5765) );
  NAND2_X1 U7271 ( .A1(n5760), .A2(n7602), .ZN(n7557) );
  NAND3_X1 U7272 ( .A1(n9824), .A2(n7539), .A3(n7536), .ZN(n5763) );
  INV_X1 U7273 ( .A(n5761), .ZN(n5762) );
  NAND2_X2 U7274 ( .A1(n5763), .A2(n5762), .ZN(n7607) );
  NAND2_X1 U7275 ( .A1(n9823), .A2(n7612), .ZN(n5764) );
  AND2_X1 U7276 ( .A1(n7557), .A2(n5764), .ZN(n7949) );
  OR2_X1 U7277 ( .A1(n7560), .A2(n5765), .ZN(n5773) );
  XNOR2_X1 U7278 ( .A(n5773), .B(n5771), .ZN(n7948) );
  NAND2_X1 U7279 ( .A1(n7949), .A2(n7948), .ZN(n7947) );
  NOR2_X1 U7280 ( .A1(n5931), .A2(n5765), .ZN(n5766) );
  XNOR2_X1 U7281 ( .A(n8039), .B(n7607), .ZN(n5767) );
  NAND2_X1 U7282 ( .A1(n5766), .A2(n5767), .ZN(n5775) );
  INV_X1 U7283 ( .A(n5766), .ZN(n5769) );
  INV_X1 U7284 ( .A(n5767), .ZN(n5768) );
  NAND2_X1 U7285 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  AND2_X1 U7286 ( .A1(n5775), .A2(n5770), .ZN(n8036) );
  INV_X1 U7287 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7288 ( .A1(n5773), .A2(n5772), .ZN(n8034) );
  NAND2_X1 U7289 ( .A1(n7947), .A2(n5774), .ZN(n8035) );
  OR2_X1 U7290 ( .A1(n5877), .A2(n5765), .ZN(n5780) );
  NAND2_X1 U7291 ( .A1(n5739), .A2(n6086), .ZN(n5778) );
  OR2_X1 U7292 ( .A1(n6281), .A2(n5776), .ZN(n5777) );
  OAI211_X1 U7293 ( .C1(n5788), .C2(n5779), .A(n5778), .B(n5777), .ZN(n9722)
         );
  XNOR2_X1 U7294 ( .A(n9722), .B(n7607), .ZN(n5781) );
  XNOR2_X1 U7295 ( .A(n5780), .B(n5781), .ZN(n9718) );
  INV_X1 U7296 ( .A(n5780), .ZN(n5782) );
  INV_X1 U7297 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5783) );
  XNOR2_X1 U7298 ( .A(n5783), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7299 ( .A1(n7328), .A2(n5888), .ZN(n5787) );
  NAND2_X1 U7300 ( .A1(n4260), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7301 ( .A1(n6657), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7302 ( .A1(n7322), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5784) );
  OR2_X1 U7303 ( .A1(n6005), .A2(n5765), .ZN(n5793) );
  NAND2_X1 U7304 ( .A1(n5739), .A2(n6426), .ZN(n5791) );
  OR2_X1 U7305 ( .A1(n6281), .A2(n5789), .ZN(n5790) );
  XNOR2_X1 U7306 ( .A(n6012), .B(n7612), .ZN(n5794) );
  NAND2_X1 U7307 ( .A1(n5793), .A2(n5794), .ZN(n5802) );
  INV_X1 U7308 ( .A(n5793), .ZN(n5796) );
  INV_X1 U7309 ( .A(n5794), .ZN(n5795) );
  NAND2_X1 U7310 ( .A1(n5796), .A2(n5795), .ZN(n5798) );
  INV_X1 U7311 ( .A(n7989), .ZN(n5803) );
  INV_X1 U7312 ( .A(n5797), .ZN(n5799) );
  NAND2_X1 U7313 ( .A1(n5799), .A2(n5798), .ZN(n5801) );
  AOI22_X1 U7314 ( .A1(n5803), .A2(n5802), .B1(n5801), .B2(n5800), .ZN(n5825)
         );
  NAND3_X1 U7315 ( .A1(n5805), .A2(n5904), .A3(n5804), .ZN(n5811) );
  OR2_X1 U7316 ( .A1(n5811), .A2(n9815), .ZN(n5810) );
  INV_X1 U7317 ( .A(n5810), .ZN(n5808) );
  OR2_X1 U7318 ( .A1(n9824), .A2(n8198), .ZN(n5806) );
  NAND2_X2 U7319 ( .A1(n9782), .A2(n5806), .ZN(n9876) );
  NOR2_X1 U7320 ( .A1(n9876), .A2(n6056), .ZN(n5807) );
  NAND2_X1 U7321 ( .A1(n5808), .A2(n5807), .ZN(n9744) );
  INV_X1 U7322 ( .A(n7544), .ZN(n5809) );
  NOR2_X1 U7323 ( .A1(n5810), .A2(n5809), .ZN(n9741) );
  INV_X1 U7324 ( .A(n9741), .ZN(n5816) );
  NOR2_X2 U7325 ( .A1(n5816), .A2(n8402), .ZN(n9724) );
  NAND2_X1 U7326 ( .A1(n5811), .A2(n5893), .ZN(n5814) );
  AND2_X1 U7327 ( .A1(n6053), .A2(n5812), .ZN(n5813) );
  NAND2_X1 U7328 ( .A1(n5814), .A2(n5813), .ZN(n7617) );
  OR2_X1 U7329 ( .A1(n7617), .A2(n7552), .ZN(n5815) );
  NAND2_X1 U7330 ( .A1(n5815), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9752) );
  INV_X1 U7331 ( .A(n9752), .ZN(n8054) );
  AOI22_X1 U7332 ( .A1(n9724), .A2(n8069), .B1(n8054), .B2(n5888), .ZN(n5824)
         );
  OR2_X1 U7333 ( .A1(n7617), .A2(P2_U3152), .ZN(n7553) );
  NOR2_X1 U7334 ( .A1(n5816), .A2(n8404), .ZN(n9721) );
  NAND2_X1 U7335 ( .A1(n6657), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5821) );
  AOI21_X1 U7336 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5817) );
  NOR2_X1 U7337 ( .A1(n5817), .A2(n5991), .ZN(n7990) );
  NAND2_X1 U7338 ( .A1(n7328), .A2(n7990), .ZN(n5820) );
  NAND2_X1 U7339 ( .A1(n4261), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7340 ( .A1(n7322), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7341 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6424) );
  OAI21_X1 U7342 ( .B1(n8046), .B2(n6306), .A(n6424), .ZN(n5822) );
  AOI21_X1 U7343 ( .B1(n9748), .B2(n6012), .A(n5822), .ZN(n5823) );
  OAI211_X1 U7344 ( .C1(n5825), .C2(n9744), .A(n5824), .B(n5823), .ZN(P2_U3232) );
  NAND2_X1 U7345 ( .A1(n5830), .A2(n9368), .ZN(n5826) );
  NAND2_X1 U7346 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  NAND2_X1 U7347 ( .A1(n8998), .A2(n6156), .ZN(n8774) );
  NAND2_X1 U7348 ( .A1(n8905), .A2(n8774), .ZN(n5832) );
  NAND2_X1 U7349 ( .A1(n5828), .A2(n5832), .ZN(n6143) );
  OAI21_X1 U7350 ( .B1(n5828), .B2(n5832), .A(n6143), .ZN(n6158) );
  INV_X1 U7351 ( .A(n6158), .ZN(n5839) );
  INV_X1 U7352 ( .A(n8997), .ZN(n5829) );
  OAI22_X1 U7353 ( .A1(n5830), .A2(n9282), .B1(n5829), .B2(n9345), .ZN(n5835)
         );
  XNOR2_X1 U7354 ( .A(n8771), .B(n5832), .ZN(n5833) );
  NOR2_X1 U7355 ( .A1(n5833), .A2(n9280), .ZN(n5834) );
  AOI211_X1 U7356 ( .C1(n7052), .C2(n6158), .A(n5835), .B(n5834), .ZN(n6160)
         );
  AOI211_X1 U7357 ( .C1(n5837), .C2(n5836), .A(n9696), .B(n4350), .ZN(n6151)
         );
  AOI21_X1 U7358 ( .B1(n9456), .B2(n5837), .A(n6151), .ZN(n5838) );
  OAI211_X1 U7359 ( .C1(n5839), .C2(n9653), .A(n6160), .B(n5838), .ZN(n5841)
         );
  NAND2_X1 U7360 ( .A1(n5841), .A2(n9716), .ZN(n5840) );
  OAI21_X1 U7361 ( .B1(n9716), .B2(n5521), .A(n5840), .ZN(P1_U3527) );
  INV_X1 U7362 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7363 ( .A1(n5841), .A2(n9704), .ZN(n5842) );
  OAI21_X1 U7364 ( .B1(n9704), .B2(n5843), .A(n5842), .ZN(P1_U3466) );
  NAND2_X1 U7365 ( .A1(n8996), .A2(n7891), .ZN(n5850) );
  OR2_X1 U7366 ( .A1(n6110), .A2(n6028), .ZN(n5847) );
  OR2_X1 U7367 ( .A1(n8758), .A2(n9976), .ZN(n5846) );
  OAI211_X1 U7368 ( .C1(n5951), .C2(n5848), .A(n5847), .B(n5846), .ZN(n6171)
         );
  NAND2_X1 U7369 ( .A1(n6171), .A2(n7889), .ZN(n5849) );
  NAND2_X1 U7370 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  XNOR2_X1 U7371 ( .A(n5851), .B(n5361), .ZN(n5854) );
  NAND2_X1 U7372 ( .A1(n5377), .A2(n8996), .ZN(n5853) );
  NAND2_X1 U7373 ( .A1(n7891), .A2(n6171), .ZN(n5852) );
  NAND2_X1 U7374 ( .A1(n5853), .A2(n5852), .ZN(n5855) );
  NAND2_X1 U7375 ( .A1(n5854), .A2(n5855), .ZN(n5943) );
  INV_X1 U7376 ( .A(n5854), .ZN(n5857) );
  INV_X1 U7377 ( .A(n5855), .ZN(n5856) );
  NAND2_X1 U7378 ( .A1(n5857), .A2(n5856), .ZN(n5945) );
  NAND2_X1 U7379 ( .A1(n5943), .A2(n5945), .ZN(n5858) );
  XNOR2_X1 U7380 ( .A(n5944), .B(n5858), .ZN(n5873) );
  INV_X1 U7381 ( .A(n6171), .ZN(n6487) );
  NOR2_X1 U7382 ( .A1(n9694), .A2(n6487), .ZN(n9672) );
  NAND2_X1 U7383 ( .A1(n8748), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5866) );
  OR2_X1 U7384 ( .A1(n8753), .A2(n5859), .ZN(n5865) );
  AND2_X1 U7385 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  OR2_X1 U7386 ( .A1(n5862), .A2(n5958), .ZN(n6562) );
  OR2_X1 U7387 ( .A1(n7863), .A2(n6562), .ZN(n5864) );
  INV_X1 U7388 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6563) );
  OR2_X1 U7389 ( .A1(n7783), .A2(n6563), .ZN(n5863) );
  NAND4_X1 U7390 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n8995)
         );
  AOI21_X1 U7391 ( .B1(n8659), .B2(n8995), .A(n5867), .ZN(n5869) );
  NAND2_X1 U7392 ( .A1(n8668), .A2(n8997), .ZN(n5868) );
  NAND2_X1 U7393 ( .A1(n5869), .A2(n5868), .ZN(n5871) );
  NOR2_X1 U7394 ( .A1(n8671), .A2(n6174), .ZN(n5870) );
  AOI211_X1 U7395 ( .C1(n8580), .C2(n9672), .A(n5871), .B(n5870), .ZN(n5872)
         );
  OAI21_X1 U7396 ( .B1(n5873), .B2(n8664), .A(n5872), .ZN(P1_U3237) );
  NAND2_X1 U7397 ( .A1(n5931), .A2(n5874), .ZN(n5875) );
  NAND2_X1 U7398 ( .A1(n5877), .A2(n9722), .ZN(n5884) );
  INV_X1 U7399 ( .A(n9722), .ZN(n9836) );
  NAND2_X1 U7400 ( .A1(n8069), .A2(n9836), .ZN(n7395) );
  NAND2_X1 U7401 ( .A1(n5884), .A2(n7395), .ZN(n7385) );
  NAND2_X1 U7402 ( .A1(n5926), .A2(n7385), .ZN(n5925) );
  NAND2_X1 U7403 ( .A1(n5877), .A2(n9836), .ZN(n5878) );
  NAND2_X1 U7404 ( .A1(n5925), .A2(n5878), .ZN(n5879) );
  NAND2_X1 U7405 ( .A1(n6005), .A2(n6012), .ZN(n7387) );
  INV_X1 U7406 ( .A(n6005), .ZN(n9720) );
  INV_X1 U7407 ( .A(n6012), .ZN(n6004) );
  NAND2_X1 U7408 ( .A1(n9720), .A2(n6004), .ZN(n6036) );
  NAND2_X1 U7409 ( .A1(n7387), .A2(n6036), .ZN(n7505) );
  NAND2_X1 U7410 ( .A1(n5879), .A2(n7505), .ZN(n6007) );
  OAI21_X1 U7411 ( .B1(n5879), .B2(n7505), .A(n6007), .ZN(n5880) );
  INV_X1 U7412 ( .A(n5880), .ZN(n6014) );
  INV_X1 U7413 ( .A(n7385), .ZN(n7509) );
  NAND2_X1 U7414 ( .A1(n5930), .A2(n7509), .ZN(n5929) );
  INV_X1 U7415 ( .A(n5884), .ZN(n7389) );
  NOR2_X1 U7416 ( .A1(n7505), .A2(n7389), .ZN(n5882) );
  NAND2_X2 U7417 ( .A1(n5929), .A2(n5882), .ZN(n6037) );
  NAND2_X1 U7418 ( .A1(n6037), .A2(n9771), .ZN(n5887) );
  INV_X1 U7419 ( .A(n7505), .ZN(n5883) );
  AOI21_X1 U7420 ( .B1(n5929), .B2(n5884), .A(n5883), .ZN(n5886) );
  INV_X1 U7421 ( .A(n6306), .ZN(n8068) );
  AOI22_X1 U7422 ( .A1(n9775), .A2(n8068), .B1(n8069), .B2(n9778), .ZN(n5885)
         );
  OAI21_X1 U7423 ( .B1(n5887), .B2(n5886), .A(n5885), .ZN(n6010) );
  INV_X1 U7424 ( .A(n9878), .ZN(n9865) );
  AOI211_X1 U7425 ( .C1(n6012), .C2(n5937), .A(n9865), .B(n6000), .ZN(n6011)
         );
  NAND2_X1 U7426 ( .A1(n6011), .A2(n8344), .ZN(n5890) );
  AOI22_X1 U7427 ( .A1(n9813), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n5888), .B2(
        n9802), .ZN(n5889) );
  OAI211_X1 U7428 ( .C1(n6004), .C2(n8398), .A(n5890), .B(n5889), .ZN(n5891)
         );
  AOI21_X1 U7429 ( .B1(n9783), .B2(n6010), .A(n5891), .ZN(n5892) );
  OAI21_X1 U7430 ( .B1(n6014), .B2(n8412), .A(n5892), .ZN(P2_U3292) );
  AND3_X1 U7431 ( .A1(n5895), .A2(n5894), .A3(n5893), .ZN(n5905) );
  AND2_X2 U7432 ( .A1(n5905), .A2(n5896), .ZN(n10073) );
  INV_X1 U7433 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5903) );
  AND2_X1 U7434 ( .A1(n7506), .A2(n4643), .ZN(n5897) );
  NAND2_X1 U7435 ( .A1(n6601), .A2(n5897), .ZN(n8511) );
  AOI22_X1 U7436 ( .A1(n5898), .A2(n9878), .B1(n8039), .B2(n9876), .ZN(n5899)
         );
  OAI211_X1 U7437 ( .C1(n9829), .C2(n5901), .A(n5900), .B(n5899), .ZN(n5906)
         );
  NAND2_X1 U7438 ( .A1(n5906), .A2(n10073), .ZN(n5902) );
  OAI21_X1 U7439 ( .B1(n10073), .B2(n5903), .A(n5902), .ZN(P2_U3457) );
  AND2_X2 U7440 ( .A1(n5905), .A2(n5904), .ZN(n9889) );
  INV_X1 U7441 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7442 ( .A1(n5906), .A2(n9889), .ZN(n5907) );
  OAI21_X1 U7443 ( .B1(n9889), .B2(n6083), .A(n5907), .ZN(P2_U3522) );
  INV_X1 U7444 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9525) );
  NOR2_X1 U7445 ( .A1(n6608), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5908) );
  NOR2_X1 U7446 ( .A1(n5909), .A2(n5908), .ZN(n9579) );
  OR2_X1 U7447 ( .A1(n9571), .A2(n9525), .ZN(n5911) );
  NAND2_X1 U7448 ( .A1(n9571), .A2(n9525), .ZN(n5910) );
  AND2_X1 U7449 ( .A1(n5911), .A2(n5910), .ZN(n9578) );
  NOR2_X1 U7450 ( .A1(n9579), .A2(n9578), .ZN(n9577) );
  AOI21_X1 U7451 ( .B1(n9525), .B2(n5912), .A(n9577), .ZN(n5914) );
  INV_X1 U7452 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9518) );
  AOI22_X1 U7453 ( .A1(n6905), .A2(n9518), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9049), .ZN(n5913) );
  NOR2_X1 U7454 ( .A1(n5914), .A2(n5913), .ZN(n9048) );
  AOI21_X1 U7455 ( .B1(n5914), .B2(n5913), .A(n9048), .ZN(n5924) );
  OR2_X1 U7456 ( .A1(n9571), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7457 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9571), .ZN(n5916) );
  NAND2_X1 U7458 ( .A1(n5917), .A2(n5916), .ZN(n9567) );
  INV_X1 U7459 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U7460 ( .A1(n5918), .A2(n9953), .ZN(n9038) );
  OAI21_X1 U7461 ( .B1(n5918), .B2(n9953), .A(n9038), .ZN(n5922) );
  INV_X1 U7462 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6763) );
  NOR2_X1 U7463 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6763), .ZN(n7084) );
  AOI21_X1 U7464 ( .B1(n9544), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7084), .ZN(
        n5919) );
  OAI21_X1 U7465 ( .B1(n5920), .B2(n9049), .A(n5919), .ZN(n5921) );
  AOI21_X1 U7466 ( .B1(n5922), .B2(n9553), .A(n5921), .ZN(n5923) );
  OAI21_X1 U7467 ( .B1(n5924), .B2(n9638), .A(n5923), .ZN(P1_U3255) );
  OAI21_X1 U7468 ( .B1(n5926), .B2(n7385), .A(n5925), .ZN(n9840) );
  INV_X1 U7469 ( .A(n9840), .ZN(n5942) );
  INV_X1 U7470 ( .A(n5927), .ZN(n5928) );
  NAND2_X1 U7471 ( .A1(n9783), .A2(n5928), .ZN(n7029) );
  OAI21_X1 U7472 ( .B1(n7509), .B2(n5930), .A(n5929), .ZN(n5933) );
  OAI22_X1 U7473 ( .A1(n6005), .A2(n8404), .B1(n5931), .B2(n8402), .ZN(n5932)
         );
  AOI21_X1 U7474 ( .B1(n5933), .B2(n9771), .A(n5932), .ZN(n5934) );
  OAI21_X1 U7475 ( .B1(n5942), .B2(n9790), .A(n5934), .ZN(n9838) );
  NAND2_X1 U7476 ( .A1(n9838), .A2(n9783), .ZN(n5941) );
  INV_X1 U7477 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6062) );
  OAI22_X1 U7478 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n9788), .B1(n9783), .B2(
        n6062), .ZN(n5939) );
  NAND2_X1 U7479 ( .A1(n5935), .A2(n9722), .ZN(n5936) );
  NAND2_X1 U7480 ( .A1(n5937), .A2(n5936), .ZN(n9837) );
  NOR2_X1 U7481 ( .A1(n8369), .A2(n9837), .ZN(n5938) );
  AOI211_X1 U7482 ( .C1(n9803), .C2(n9722), .A(n5939), .B(n5938), .ZN(n5940)
         );
  OAI211_X1 U7483 ( .C1(n5942), .C2(n7029), .A(n5941), .B(n5940), .ZN(P2_U3293) );
  NAND2_X1 U7484 ( .A1(n5944), .A2(n5943), .ZN(n5946) );
  NAND2_X1 U7485 ( .A1(n8995), .A2(n7891), .ZN(n5953) );
  OR2_X1 U7486 ( .A1(n6191), .A2(n6110), .ZN(n5949) );
  OR2_X1 U7487 ( .A1(n8758), .A2(n5947), .ZN(n5948) );
  OAI211_X1 U7488 ( .C1(n5951), .C2(n5950), .A(n5949), .B(n5948), .ZN(n6565)
         );
  NAND2_X1 U7489 ( .A1(n6565), .A2(n7889), .ZN(n5952) );
  NAND2_X1 U7490 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  XNOR2_X1 U7491 ( .A(n5954), .B(n5361), .ZN(n6108) );
  NAND2_X1 U7492 ( .A1(n5377), .A2(n8995), .ZN(n5956) );
  NAND2_X1 U7493 ( .A1(n6565), .A2(n7891), .ZN(n5955) );
  XNOR2_X1 U7494 ( .A(n6108), .B(n6107), .ZN(n5957) );
  XNOR2_X1 U7495 ( .A(n6109), .B(n5957), .ZN(n5970) );
  NAND2_X1 U7496 ( .A1(n8748), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5964) );
  INV_X1 U7497 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6545) );
  OR2_X1 U7498 ( .A1(n7783), .A2(n6545), .ZN(n5963) );
  NAND2_X1 U7499 ( .A1(n5958), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6119) );
  OR2_X1 U7500 ( .A1(n5958), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7501 ( .A1(n6119), .A2(n5959), .ZN(n6544) );
  OR2_X1 U7502 ( .A1(n7863), .A2(n6544), .ZN(n5962) );
  OR2_X1 U7503 ( .A1(n8753), .A2(n5960), .ZN(n5961) );
  NAND4_X1 U7504 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(n8994)
         );
  INV_X1 U7505 ( .A(n8994), .ZN(n6558) );
  NOR2_X1 U7506 ( .A1(n8666), .A2(n6558), .ZN(n5965) );
  AOI211_X1 U7507 ( .C1(n8668), .C2(n8996), .A(n5966), .B(n5965), .ZN(n5967)
         );
  OAI21_X1 U7508 ( .B1(n8671), .B2(n6562), .A(n5967), .ZN(n5968) );
  AOI21_X1 U7509 ( .B1(n8679), .B2(n6565), .A(n5968), .ZN(n5969) );
  OAI21_X1 U7510 ( .B1(n5970), .B2(n8664), .A(n5969), .ZN(P1_U3211) );
  INV_X1 U7511 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5979) );
  INV_X1 U7512 ( .A(n5971), .ZN(n5975) );
  INV_X1 U7513 ( .A(n5972), .ZN(n5973) );
  NAND2_X1 U7514 ( .A1(n5973), .A2(SI_17_), .ZN(n5974) );
  MUX2_X1 U7515 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7333), .Z(n6021) );
  XNOR2_X1 U7516 ( .A(n6021), .B(SI_18_), .ZN(n6018) );
  XNOR2_X1 U7517 ( .A(n6020), .B(n6018), .ZN(n7715) );
  INV_X1 U7518 ( .A(n7715), .ZN(n5984) );
  NAND2_X1 U7519 ( .A1(n5977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  XNOR2_X1 U7520 ( .A(n5978), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8108) );
  INV_X1 U7521 ( .A(n8108), .ZN(n7180) );
  OAI222_X1 U7522 ( .A1(n8539), .A2(n5979), .B1(n7920), .B2(n5984), .C1(
        P2_U3152), .C2(n7180), .ZN(P2_U3340) );
  INV_X1 U7523 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7524 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  NAND2_X1 U7525 ( .A1(n5982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7526 ( .A(n5983), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9627) );
  INV_X1 U7527 ( .A(n9627), .ZN(n9058) );
  OAI222_X1 U7528 ( .A1(n7154), .A2(n5985), .B1(n7551), .B2(n5984), .C1(n4258), 
        .C2(n9058), .ZN(P1_U3335) );
  NAND2_X1 U7529 ( .A1(n6037), .A2(n6036), .ZN(n5990) );
  NAND2_X1 U7530 ( .A1(n7335), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7531 ( .A1(n6281), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7532 ( .A1(n5739), .A2(n6089), .ZN(n5987) );
  INV_X1 U7533 ( .A(n9844), .ZN(n7994) );
  NAND2_X1 U7534 ( .A1(n6306), .A2(n7994), .ZN(n7382) );
  NAND2_X1 U7535 ( .A1(n8068), .A2(n9844), .ZN(n7397) );
  NAND2_X1 U7536 ( .A1(n7382), .A2(n7397), .ZN(n7511) );
  XNOR2_X1 U7537 ( .A(n5990), .B(n7511), .ZN(n5997) );
  OAI21_X1 U7538 ( .B1(n5991), .B2(P2_REG3_REG_6__SCAN_IN), .A(n6040), .ZN(
        n9751) );
  INV_X1 U7539 ( .A(n9751), .ZN(n5992) );
  NAND2_X1 U7540 ( .A1(n7328), .A2(n5992), .ZN(n5996) );
  NAND2_X1 U7541 ( .A1(n4260), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7542 ( .A1(n6657), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7543 ( .A1(n7322), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5993) );
  NAND4_X1 U7544 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n8067)
         );
  AOI222_X1 U7545 ( .A1(n9771), .A2(n5997), .B1(n8067), .B2(n9775), .C1(n9720), 
        .C2(n9778), .ZN(n9843) );
  INV_X1 U7546 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10025) );
  INV_X1 U7547 ( .A(n7990), .ZN(n5998) );
  OAI22_X1 U7548 ( .A1(n9783), .A2(n10025), .B1(n5998), .B2(n9788), .ZN(n6003)
         );
  INV_X1 U7549 ( .A(n6033), .ZN(n5999) );
  OAI211_X1 U7550 ( .C1(n9844), .C2(n6000), .A(n5999), .B(n9878), .ZN(n9842)
         );
  NOR2_X1 U7551 ( .A1(n9842), .A2(n6001), .ZN(n6002) );
  AOI211_X1 U7552 ( .C1(n9803), .C2(n7994), .A(n6003), .B(n6002), .ZN(n6009)
         );
  NAND2_X1 U7553 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  XNOR2_X1 U7554 ( .A(n6027), .B(n7511), .ZN(n9846) );
  NAND2_X1 U7555 ( .A1(n9846), .A2(n6195), .ZN(n6008) );
  OAI211_X1 U7556 ( .C1(n9843), .C2(n9813), .A(n6009), .B(n6008), .ZN(P2_U3291) );
  INV_X1 U7557 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9980) );
  AOI211_X1 U7558 ( .C1(n6012), .C2(n9876), .A(n6011), .B(n6010), .ZN(n6013)
         );
  OAI21_X1 U7559 ( .B1(n9829), .B2(n6014), .A(n6013), .ZN(n6016) );
  NAND2_X1 U7560 ( .A1(n6016), .A2(n10073), .ZN(n6015) );
  OAI21_X1 U7561 ( .B1(n10073), .B2(n9980), .A(n6015), .ZN(P2_U3463) );
  NAND2_X1 U7562 ( .A1(n6016), .A2(n9889), .ZN(n6017) );
  OAI21_X1 U7563 ( .B1(n9889), .B2(n6427), .A(n6017), .ZN(P2_U3524) );
  INV_X1 U7564 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6026) );
  INV_X1 U7565 ( .A(n6018), .ZN(n6019) );
  INV_X1 U7566 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10055) );
  MUX2_X1 U7567 ( .A(n6026), .B(n10055), .S(n7333), .Z(n6023) );
  INV_X1 U7568 ( .A(SI_19_), .ZN(n6022) );
  NAND2_X1 U7569 ( .A1(n6023), .A2(n6022), .ZN(n6184) );
  INV_X1 U7570 ( .A(n6023), .ZN(n6024) );
  NAND2_X1 U7571 ( .A1(n6024), .A2(SI_19_), .ZN(n6025) );
  NAND2_X1 U7572 ( .A1(n6184), .A2(n6025), .ZN(n6182) );
  XNOR2_X1 U7573 ( .A(n6183), .B(n6182), .ZN(n7732) );
  INV_X1 U7574 ( .A(n7732), .ZN(n7159) );
  OAI222_X1 U7575 ( .A1(n8539), .A2(n6026), .B1(n7920), .B2(n7159), .C1(n8198), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U7576 ( .A1(n5739), .A2(n6079), .ZN(n6030) );
  OR2_X1 U7577 ( .A1(n6281), .A2(n6028), .ZN(n6029) );
  OAI211_X1 U7578 ( .C1(n7359), .C2(n6031), .A(n6030), .B(n6029), .ZN(n9877)
         );
  XNOR2_X1 U7579 ( .A(n8067), .B(n9877), .ZN(n7515) );
  INV_X1 U7580 ( .A(n7515), .ZN(n6032) );
  XNOR2_X1 U7581 ( .A(n6276), .B(n6032), .ZN(n9884) );
  INV_X1 U7582 ( .A(n9884), .ZN(n6052) );
  OR2_X1 U7583 ( .A1(n6033), .A2(n7401), .ZN(n6034) );
  AND2_X1 U7584 ( .A1(n6211), .A2(n6034), .ZN(n9879) );
  OAI22_X1 U7585 ( .A1(n8398), .A2(n7401), .B1(n9788), .B2(n9751), .ZN(n6035)
         );
  AOI21_X1 U7586 ( .B1(n9879), .B2(n9809), .A(n6035), .ZN(n6051) );
  INV_X1 U7587 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6049) );
  AND2_X1 U7588 ( .A1(n6036), .A2(n7397), .ZN(n7396) );
  NAND2_X1 U7589 ( .A1(n6200), .A2(n7382), .ZN(n6038) );
  XNOR2_X1 U7590 ( .A(n6038), .B(n7515), .ZN(n6048) );
  AND2_X1 U7591 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  NOR2_X1 U7592 ( .A1(n6203), .A2(n6041), .ZN(n6326) );
  NAND2_X1 U7593 ( .A1(n7328), .A2(n6326), .ZN(n6046) );
  NAND2_X1 U7594 ( .A1(n4261), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7595 ( .A1(n6657), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7596 ( .A1(n7322), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6043) );
  OR2_X1 U7597 ( .A1(n6316), .A2(n8404), .ZN(n6047) );
  OAI21_X1 U7598 ( .B1(n6306), .B2(n8402), .A(n6047), .ZN(n9740) );
  AOI21_X1 U7599 ( .B1(n6048), .B2(n9771), .A(n9740), .ZN(n9881) );
  MUX2_X1 U7600 ( .A(n6049), .B(n9881), .S(n9783), .Z(n6050) );
  OAI211_X1 U7601 ( .C1(n6052), .C2(n8412), .A(n6051), .B(n6050), .ZN(P2_U3290) );
  OAI21_X1 U7602 ( .B1(n6053), .B2(P2_U3152), .A(n7549), .ZN(n6054) );
  INV_X1 U7603 ( .A(n6054), .ZN(n6055) );
  OAI21_X1 U7604 ( .B1(n9815), .B2(n6056), .A(n6055), .ZN(n6074) );
  NAND2_X1 U7605 ( .A1(n6074), .A2(n6283), .ZN(n6057) );
  NAND2_X1 U7606 ( .A1(n6057), .A2(n8071), .ZN(n6100) );
  INV_X1 U7607 ( .A(n6100), .ZN(n6058) );
  INV_X1 U7608 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6059) );
  MUX2_X1 U7609 ( .A(n6059), .B(P2_REG2_REG_11__SCAN_IN), .S(n6651), .Z(n6060)
         );
  INV_X1 U7610 ( .A(n6060), .ZN(n6072) );
  INV_X1 U7611 ( .A(n6861), .ZN(n6067) );
  NAND2_X1 U7612 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n6821) );
  AOI21_X1 U7613 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n6082), .A(n6819), .ZN(
        n6783) );
  XNOR2_X1 U7614 ( .A(n6085), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6782) );
  MUX2_X1 U7615 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6062), .S(n6086), .Z(n6420)
         );
  OAI21_X1 U7616 ( .B1(n6423), .B2(n6062), .A(n6418), .ZN(n6436) );
  XOR2_X1 U7617 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6426), .Z(n6437) );
  NAND2_X1 U7618 ( .A1(n6089), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6063) );
  OAI21_X1 U7619 ( .B1(n6089), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6063), .ZN(
        n6387) );
  INV_X1 U7620 ( .A(n6389), .ZN(n6064) );
  AOI21_X1 U7621 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6089), .A(n6064), .ZN(
        n6795) );
  MUX2_X1 U7622 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6049), .S(n6079), .Z(n6065)
         );
  INV_X1 U7623 ( .A(n6065), .ZN(n6794) );
  NOR2_X1 U7624 ( .A1(n6795), .A2(n6794), .ZN(n6793) );
  AOI21_X1 U7625 ( .B1(n6079), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6793), .ZN(
        n6833) );
  NAND2_X1 U7626 ( .A1(n6837), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6066) );
  OAI21_X1 U7627 ( .B1(n6837), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6066), .ZN(
        n6832) );
  NOR2_X1 U7628 ( .A1(n6833), .A2(n6832), .ZN(n6831) );
  AOI21_X1 U7629 ( .B1(n6837), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6831), .ZN(
        n6852) );
  XOR2_X1 U7630 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6861), .Z(n6851) );
  NOR2_X1 U7631 ( .A1(n6852), .A2(n6851), .ZN(n6850) );
  AOI21_X1 U7632 ( .B1(n6067), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6850), .ZN(
        n6893) );
  OR2_X1 U7633 ( .A1(n6896), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7634 ( .A1(n6896), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7635 ( .A1(n6069), .A2(n6068), .ZN(n6892) );
  NOR2_X1 U7636 ( .A1(n6893), .A2(n6892), .ZN(n6891) );
  NAND2_X1 U7637 ( .A1(n6812), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6070) );
  OAI21_X1 U7638 ( .B1(n6812), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6070), .ZN(
        n6807) );
  OAI21_X1 U7639 ( .B1(n6072), .B2(n6071), .A(n6218), .ZN(n6105) );
  AND2_X1 U7640 ( .A1(n6283), .A2(n7543), .ZN(n6073) );
  NAND2_X1 U7641 ( .A1(n6074), .A2(n6073), .ZN(n9759) );
  INV_X1 U7642 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6075) );
  MUX2_X1 U7643 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6075), .S(n6651), .Z(n6099)
         );
  INV_X1 U7644 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7645 ( .A1(n6812), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6097) );
  MUX2_X1 U7646 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6076), .S(n6812), .Z(n6811)
         );
  NAND2_X1 U7647 ( .A1(n6896), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6096) );
  INV_X1 U7648 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6077) );
  MUX2_X1 U7649 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6077), .S(n6896), .Z(n6898)
         );
  INV_X1 U7650 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7651 ( .A1(n6837), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6093) );
  INV_X1 U7652 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6078) );
  MUX2_X1 U7653 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6078), .S(n6837), .Z(n6836)
         );
  NAND2_X1 U7654 ( .A1(n6079), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6092) );
  INV_X1 U7655 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6080) );
  MUX2_X1 U7656 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6080), .S(n6079), .Z(n6799)
         );
  NAND2_X1 U7657 ( .A1(n6089), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6091) );
  INV_X1 U7658 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6081) );
  MUX2_X1 U7659 ( .A(n6081), .B(P2_REG1_REG_1__SCAN_IN), .S(n6828), .Z(n6824)
         );
  NAND3_X1 U7660 ( .A1(n6824), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U7661 ( .A1(n6082), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6785) );
  MUX2_X1 U7662 ( .A(n6083), .B(P2_REG1_REG_2__SCAN_IN), .S(n6085), .Z(n6784)
         );
  AOI21_X1 U7663 ( .B1(n6823), .B2(n6785), .A(n6784), .ZN(n6084) );
  INV_X1 U7664 ( .A(n6084), .ZN(n6787) );
  NAND2_X1 U7665 ( .A1(n6085), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6414) );
  INV_X1 U7666 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U7667 ( .A(n10016), .B(P2_REG1_REG_3__SCAN_IN), .S(n6086), .Z(n6413)
         );
  AOI21_X1 U7668 ( .B1(n6787), .B2(n6414), .A(n6413), .ZN(n6430) );
  INV_X1 U7669 ( .A(n6430), .ZN(n6088) );
  NAND2_X1 U7670 ( .A1(n6086), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6425) );
  MUX2_X1 U7671 ( .A(n6427), .B(P2_REG1_REG_4__SCAN_IN), .S(n6426), .Z(n6087)
         );
  AOI21_X1 U7672 ( .B1(n6088), .B2(n6425), .A(n6087), .ZN(n6432) );
  AOI21_X1 U7673 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6426), .A(n6432), .ZN(
        n6393) );
  INV_X1 U7674 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9874) );
  MUX2_X1 U7675 ( .A(n9874), .B(P2_REG1_REG_5__SCAN_IN), .S(n6089), .Z(n6392)
         );
  OR2_X1 U7676 ( .A1(n6393), .A2(n6392), .ZN(n6090) );
  NAND2_X1 U7677 ( .A1(n6091), .A2(n6090), .ZN(n6800) );
  NAND2_X1 U7678 ( .A1(n6799), .A2(n6800), .ZN(n6798) );
  NAND2_X1 U7679 ( .A1(n6092), .A2(n6798), .ZN(n6835) );
  NAND2_X1 U7680 ( .A1(n6836), .A2(n6835), .ZN(n6834) );
  NAND2_X1 U7681 ( .A1(n6093), .A2(n6834), .ZN(n6853) );
  MUX2_X1 U7682 ( .A(n6095), .B(P2_REG1_REG_8__SCAN_IN), .S(n6861), .Z(n6094)
         );
  NAND2_X1 U7683 ( .A1(n6853), .A2(n6094), .ZN(n6854) );
  OAI21_X1 U7684 ( .B1(n6861), .B2(n6095), .A(n6854), .ZN(n6899) );
  NAND2_X1 U7685 ( .A1(n6898), .A2(n6899), .ZN(n6897) );
  NAND2_X1 U7686 ( .A1(n6096), .A2(n6897), .ZN(n6810) );
  NAND2_X1 U7687 ( .A1(n6811), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U7688 ( .A1(n6097), .A2(n6809), .ZN(n6098) );
  NAND2_X1 U7689 ( .A1(n6099), .A2(n6098), .ZN(n6224) );
  OAI21_X1 U7690 ( .B1(n6099), .B2(n6098), .A(n6224), .ZN(n6103) );
  NAND2_X1 U7691 ( .A1(n6100), .A2(n7629), .ZN(n9757) );
  INV_X1 U7692 ( .A(n9757), .ZN(n8109) );
  NAND2_X1 U7693 ( .A1(n8109), .A2(n6651), .ZN(n6102) );
  AND2_X1 U7694 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6663) );
  AOI21_X1 U7695 ( .B1(n9754), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6663), .ZN(
        n6101) );
  OAI211_X1 U7696 ( .C1(n9759), .C2(n6103), .A(n6102), .B(n6101), .ZN(n6104)
         );
  AOI21_X1 U7697 ( .B1(n4352), .B2(n6105), .A(n6104), .ZN(n6106) );
  INV_X1 U7698 ( .A(n6106), .ZN(P2_U3256) );
  NAND2_X1 U7699 ( .A1(n6282), .A2(n8760), .ZN(n6112) );
  AOI22_X1 U7700 ( .A1(n7734), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7733), .B2(
        n9028), .ZN(n6111) );
  NAND2_X1 U7701 ( .A1(n6547), .A2(n7889), .ZN(n6114) );
  NAND2_X1 U7702 ( .A1(n8994), .A2(n7891), .ZN(n6113) );
  NAND2_X1 U7703 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  XNOR2_X1 U7704 ( .A(n6115), .B(n7872), .ZN(n6254) );
  NAND2_X1 U7705 ( .A1(n6547), .A2(n7891), .ZN(n6117) );
  NAND2_X1 U7706 ( .A1(n5377), .A2(n8994), .ZN(n6116) );
  AND2_X1 U7707 ( .A1(n6117), .A2(n6116), .ZN(n6251) );
  INV_X1 U7708 ( .A(n6251), .ZN(n6255) );
  XNOR2_X1 U7709 ( .A(n6254), .B(n6255), .ZN(n6118) );
  XNOR2_X1 U7710 ( .A(n6253), .B(n6118), .ZN(n6130) );
  AND2_X1 U7711 ( .A1(n9456), .A2(n6547), .ZN(n9687) );
  NAND2_X1 U7712 ( .A1(n8748), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7713 ( .A1(n6119), .A2(n10056), .ZN(n6120) );
  NAND2_X1 U7714 ( .A1(n6262), .A2(n6120), .ZN(n6526) );
  OR2_X1 U7715 ( .A1(n7863), .A2(n6526), .ZN(n6123) );
  OR2_X1 U7716 ( .A1(n7783), .A2(n6527), .ZN(n6122) );
  OR2_X1 U7717 ( .A1(n8753), .A2(n9714), .ZN(n6121) );
  NAND4_X1 U7718 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(n8993)
         );
  INV_X1 U7719 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6125) );
  NOR2_X1 U7720 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6125), .ZN(n9030) );
  AOI21_X1 U7721 ( .B1(n8659), .B2(n8993), .A(n9030), .ZN(n6127) );
  NAND2_X1 U7722 ( .A1(n8668), .A2(n8995), .ZN(n6126) );
  OAI211_X1 U7723 ( .C1(n8671), .C2(n6544), .A(n6127), .B(n6126), .ZN(n6128)
         );
  AOI21_X1 U7724 ( .B1(n8580), .B2(n9687), .A(n6128), .ZN(n6129) );
  OAI21_X1 U7725 ( .B1(n6130), .B2(n8664), .A(n6129), .ZN(P1_U3219) );
  OAI211_X1 U7726 ( .C1(n4350), .C2(n9668), .A(n9673), .B(n6170), .ZN(n9667)
         );
  INV_X1 U7727 ( .A(n9667), .ZN(n6138) );
  NAND2_X1 U7728 ( .A1(n9648), .A2(n5586), .ZN(n6131) );
  INV_X1 U7729 ( .A(n6132), .ZN(n6133) );
  NAND2_X1 U7730 ( .A1(n9329), .A2(n8996), .ZN(n9666) );
  OAI21_X1 U7731 ( .B1(n9367), .B2(n6133), .A(n9666), .ZN(n6137) );
  OR2_X1 U7732 ( .A1(n8997), .A2(n9668), .ZN(n8781) );
  NAND2_X1 U7733 ( .A1(n8997), .A2(n9668), .ZN(n8783) );
  NAND2_X1 U7734 ( .A1(n8781), .A2(n8783), .ZN(n6161) );
  XNOR2_X1 U7735 ( .A(n6505), .B(n6161), .ZN(n6134) );
  NAND2_X1 U7736 ( .A1(n6134), .A2(n9348), .ZN(n6136) );
  NAND2_X1 U7737 ( .A1(n9343), .A2(n8998), .ZN(n6135) );
  NAND2_X1 U7738 ( .A1(n6136), .A2(n6135), .ZN(n9669) );
  AOI211_X1 U7739 ( .C1(n6138), .C2(n9256), .A(n6137), .B(n9669), .ZN(n6148)
         );
  INV_X1 U7740 ( .A(n6139), .ZN(n6140) );
  OR2_X1 U7741 ( .A1(n6141), .A2(n6140), .ZN(n6150) );
  AND2_X2 U7742 ( .A1(n6150), .A2(n9367), .ZN(n9364) );
  NAND2_X1 U7743 ( .A1(n4407), .A2(n6156), .ZN(n6142) );
  XNOR2_X1 U7744 ( .A(n6164), .B(n6161), .ZN(n9671) );
  NOR2_X1 U7745 ( .A1(n6144), .A2(n7872), .ZN(n6145) );
  NAND2_X1 U7746 ( .A1(n6776), .A2(n6145), .ZN(n9335) );
  INV_X1 U7747 ( .A(n9335), .ZN(n9352) );
  NAND2_X1 U7748 ( .A1(n6776), .A2(n4888), .ZN(n9369) );
  OAI22_X1 U7749 ( .A1(n6776), .A2(n5546), .B1(n9369), .B2(n9668), .ZN(n6146)
         );
  AOI21_X1 U7750 ( .B1(n9671), .B2(n9352), .A(n6146), .ZN(n6147) );
  OAI21_X1 U7751 ( .B1(n6148), .B2(n9364), .A(n6147), .ZN(P1_U3286) );
  NAND2_X1 U7752 ( .A1(n4502), .A2(n5586), .ZN(n6149) );
  NOR2_X1 U7753 ( .A1(n9364), .A2(n6149), .ZN(n9373) );
  OR2_X1 U7754 ( .A1(n6150), .A2(n5586), .ZN(n9357) );
  INV_X1 U7755 ( .A(n9357), .ZN(n9211) );
  NAND2_X1 U7756 ( .A1(n6151), .A2(n9211), .ZN(n6155) );
  NOR2_X1 U7757 ( .A1(n9367), .A2(n6152), .ZN(n6153) );
  AOI21_X1 U7758 ( .B1(n9364), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6153), .ZN(
        n6154) );
  OAI211_X1 U7759 ( .C1(n6156), .C2(n9369), .A(n6155), .B(n6154), .ZN(n6157)
         );
  AOI21_X1 U7760 ( .B1(n9373), .B2(n6158), .A(n6157), .ZN(n6159) );
  OAI21_X1 U7761 ( .B1(n6160), .B2(n9364), .A(n6159), .ZN(P1_U3287) );
  NAND2_X1 U7762 ( .A1(n8997), .A2(n6162), .ZN(n6163) );
  OR2_X1 U7763 ( .A1(n8996), .A2(n6487), .ZN(n8786) );
  NAND2_X1 U7764 ( .A1(n8996), .A2(n6487), .ZN(n8908) );
  NAND2_X1 U7765 ( .A1(n8786), .A2(n8908), .ZN(n6167) );
  OAI21_X1 U7766 ( .B1(n6165), .B2(n6167), .A(n6489), .ZN(n6166) );
  INV_X1 U7767 ( .A(n6166), .ZN(n9677) );
  INV_X1 U7768 ( .A(n8783), .ZN(n6506) );
  OAI21_X1 U7769 ( .B1(n6505), .B2(n6506), .A(n8781), .ZN(n6168) );
  INV_X1 U7770 ( .A(n6167), .ZN(n8778) );
  XNOR2_X1 U7771 ( .A(n6168), .B(n8778), .ZN(n6169) );
  AOI222_X1 U7772 ( .A1(n9348), .A2(n6169), .B1(n8997), .B2(n9343), .C1(n8995), 
        .C2(n9329), .ZN(n9676) );
  MUX2_X1 U7773 ( .A(n4999), .B(n9676), .S(n6776), .Z(n6177) );
  AOI21_X1 U7774 ( .B1(n6171), .B2(n6170), .A(n6561), .ZN(n9674) );
  INV_X1 U7775 ( .A(n5347), .ZN(n8978) );
  OR2_X1 U7776 ( .A1(n6172), .A2(n8978), .ZN(n6173) );
  NOR2_X1 U7777 ( .A1(n9364), .A2(n6173), .ZN(n9372) );
  OAI22_X1 U7778 ( .A1(n9369), .A2(n6487), .B1(n6174), .B2(n9367), .ZN(n6175)
         );
  AOI21_X1 U7779 ( .B1(n9674), .B2(n9372), .A(n6175), .ZN(n6176) );
  OAI211_X1 U7780 ( .C1(n9335), .C2(n9677), .A(n6177), .B(n6176), .ZN(P1_U3285) );
  OAI21_X1 U7781 ( .B1(n9372), .B2(n9361), .A(n6178), .ZN(n6181) );
  INV_X1 U7782 ( .A(n9367), .ZN(n9287) );
  AOI22_X1 U7783 ( .A1(n6179), .A2(n6776), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9287), .ZN(n6180) );
  OAI211_X1 U7784 ( .C1(n6776), .C2(n9012), .A(n6181), .B(n6180), .ZN(P1_U3291) );
  INV_X1 U7785 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6238) );
  INV_X1 U7786 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7755) );
  MUX2_X1 U7787 ( .A(n6238), .B(n7755), .S(n7333), .Z(n6186) );
  INV_X1 U7788 ( .A(SI_20_), .ZN(n6185) );
  NAND2_X1 U7789 ( .A1(n6186), .A2(n6185), .ZN(n6371) );
  INV_X1 U7790 ( .A(n6186), .ZN(n6187) );
  NAND2_X1 U7791 ( .A1(n6187), .A2(SI_20_), .ZN(n6188) );
  AND2_X1 U7792 ( .A1(n6371), .A2(n6188), .ZN(n6369) );
  INV_X1 U7793 ( .A(n7754), .ZN(n6237) );
  OAI222_X1 U7794 ( .A1(P1_U3084), .A2(n6189), .B1(n7551), .B2(n6237), .C1(
        n7755), .C2(n7154), .ZN(P1_U3333) );
  NOR2_X1 U7795 ( .A1(n8067), .A2(n9877), .ZN(n6274) );
  OR2_X1 U7796 ( .A1(n6276), .A2(n6274), .ZN(n6190) );
  NAND2_X1 U7797 ( .A1(n8067), .A2(n9877), .ZN(n6277) );
  NAND2_X1 U7798 ( .A1(n6190), .A2(n6277), .ZN(n6194) );
  NAND2_X1 U7799 ( .A1(n5739), .A2(n6837), .ZN(n6192) );
  NAND2_X1 U7800 ( .A1(n6316), .A2(n6317), .ZN(n7406) );
  INV_X1 U7801 ( .A(n6316), .ZN(n8066) );
  INV_X1 U7802 ( .A(n6317), .ZN(n9848) );
  NAND2_X1 U7803 ( .A1(n8066), .A2(n9848), .ZN(n7405) );
  XNOR2_X1 U7804 ( .A(n6194), .B(n6201), .ZN(n9852) );
  INV_X1 U7805 ( .A(n9852), .ZN(n6217) );
  INV_X1 U7806 ( .A(n8067), .ZN(n7992) );
  NAND2_X1 U7807 ( .A1(n7992), .A2(n9877), .ZN(n6196) );
  AND2_X1 U7808 ( .A1(n7382), .A2(n6196), .ZN(n7391) );
  NAND2_X1 U7809 ( .A1(n6200), .A2(n7391), .ZN(n6197) );
  NAND2_X1 U7810 ( .A1(n8067), .A2(n7401), .ZN(n7399) );
  NAND2_X1 U7811 ( .A1(n6197), .A2(n7399), .ZN(n6202) );
  AND2_X1 U7812 ( .A1(n7391), .A2(n6201), .ZN(n6199) );
  OAI211_X1 U7813 ( .C1(n6202), .C2(n6201), .A(n6292), .B(n9771), .ZN(n6210)
         );
  OR2_X1 U7814 ( .A1(n6203), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7815 ( .A1(n6295), .A2(n6204), .ZN(n9739) );
  INV_X1 U7816 ( .A(n9739), .ZN(n6290) );
  NAND2_X1 U7817 ( .A1(n7328), .A2(n6290), .ZN(n6208) );
  NAND2_X1 U7818 ( .A1(n4260), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7819 ( .A1(n6657), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7820 ( .A1(n5451), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6205) );
  NAND4_X1 U7821 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .ZN(n8065)
         );
  AOI22_X1 U7822 ( .A1(n9775), .A2(n8065), .B1(n8067), .B2(n9778), .ZN(n6209)
         );
  NAND2_X1 U7823 ( .A1(n6210), .A2(n6209), .ZN(n9851) );
  INV_X1 U7824 ( .A(n6211), .ZN(n6212) );
  OAI21_X1 U7825 ( .B1(n6212), .B2(n9848), .A(n6289), .ZN(n9849) );
  AOI22_X1 U7826 ( .A1(n9813), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n6326), .B2(
        n9802), .ZN(n6214) );
  NAND2_X1 U7827 ( .A1(n9803), .A2(n6317), .ZN(n6213) );
  OAI211_X1 U7828 ( .C1(n9849), .C2(n8369), .A(n6214), .B(n6213), .ZN(n6215)
         );
  AOI21_X1 U7829 ( .B1(n9851), .B2(n9783), .A(n6215), .ZN(n6216) );
  OAI21_X1 U7830 ( .B1(n6217), .B2(n8412), .A(n6216), .ZN(P2_U3289) );
  INV_X1 U7831 ( .A(n6651), .ZN(n6220) );
  INV_X1 U7832 ( .A(n6218), .ZN(n6219) );
  AOI21_X1 U7833 ( .B1(n6220), .B2(n6059), .A(n6219), .ZN(n6375) );
  XOR2_X1 U7834 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6740), .Z(n6376) );
  NAND2_X1 U7835 ( .A1(n6375), .A2(n6376), .ZN(n6374) );
  NOR2_X1 U7836 ( .A1(n6872), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6221) );
  AOI21_X1 U7837 ( .B1(n6872), .B2(P2_REG2_REG_13__SCAN_IN), .A(n6221), .ZN(
        n6222) );
  OAI21_X1 U7838 ( .B1(n6223), .B2(n6222), .A(n6635), .ZN(n6235) );
  INV_X1 U7839 ( .A(n6224), .ZN(n6225) );
  AOI21_X1 U7840 ( .B1(n6651), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6225), .ZN(
        n6379) );
  INV_X1 U7841 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6226) );
  MUX2_X1 U7842 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6226), .S(n6740), .Z(n6378)
         );
  NAND2_X1 U7843 ( .A1(n6379), .A2(n6378), .ZN(n6377) );
  INV_X1 U7844 ( .A(n6740), .ZN(n6386) );
  NAND2_X1 U7845 ( .A1(n6386), .A2(n6226), .ZN(n6227) );
  NAND2_X1 U7846 ( .A1(n6377), .A2(n6227), .ZN(n6229) );
  INV_X1 U7847 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9499) );
  MUX2_X1 U7848 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9499), .S(n6872), .Z(n6228)
         );
  AND2_X1 U7849 ( .A1(n6229), .A2(n6228), .ZN(n6630) );
  NOR2_X1 U7850 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  NOR2_X1 U7851 ( .A1(n6630), .A2(n6230), .ZN(n6233) );
  NAND2_X1 U7852 ( .A1(n8109), .A2(n6872), .ZN(n6232) );
  AND2_X1 U7853 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6884) );
  AOI21_X1 U7854 ( .B1(n9754), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6884), .ZN(
        n6231) );
  OAI211_X1 U7855 ( .C1(n6233), .C2(n9759), .A(n6232), .B(n6231), .ZN(n6234)
         );
  AOI21_X1 U7856 ( .B1(n4352), .B2(n6235), .A(n6234), .ZN(n6236) );
  INV_X1 U7857 ( .A(n6236), .ZN(P2_U3258) );
  OAI222_X1 U7858 ( .A1(n8539), .A2(n6238), .B1(P2_U3152), .B2(n7506), .C1(
        n8543), .C2(n6237), .ZN(P2_U3338) );
  NAND2_X1 U7859 ( .A1(n6333), .A2(n8760), .ZN(n6241) );
  AOI22_X1 U7860 ( .A1(n7734), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7733), .B2(
        n6239), .ZN(n6240) );
  NAND2_X1 U7861 ( .A1(n6529), .A2(n7889), .ZN(n6243) );
  NAND2_X1 U7862 ( .A1(n8993), .A2(n7891), .ZN(n6242) );
  NAND2_X1 U7863 ( .A1(n6243), .A2(n6242), .ZN(n6244) );
  XNOR2_X1 U7864 ( .A(n6244), .B(n7872), .ZN(n6246) );
  AND2_X1 U7865 ( .A1(n5377), .A2(n8993), .ZN(n6245) );
  AOI21_X1 U7866 ( .B1(n6529), .B2(n7891), .A(n6245), .ZN(n6247) );
  NAND2_X1 U7867 ( .A1(n6246), .A2(n6247), .ZN(n6441) );
  INV_X1 U7868 ( .A(n6246), .ZN(n6249) );
  INV_X1 U7869 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U7870 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND2_X1 U7871 ( .A1(n6441), .A2(n6250), .ZN(n6261) );
  NAND2_X1 U7872 ( .A1(n6254), .A2(n6251), .ZN(n6252) );
  INV_X1 U7873 ( .A(n6254), .ZN(n6256) );
  NAND2_X1 U7874 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  INV_X1 U7875 ( .A(n6442), .ZN(n6259) );
  AOI21_X1 U7876 ( .B1(n6261), .B2(n6260), .A(n6259), .ZN(n6273) );
  NAND2_X1 U7877 ( .A1(n8748), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6267) );
  OR2_X1 U7878 ( .A1(n8753), .A2(n9491), .ZN(n6266) );
  NAND2_X1 U7879 ( .A1(n6262), .A2(n10031), .ZN(n6263) );
  NAND2_X1 U7880 ( .A1(n6458), .A2(n6263), .ZN(n6577) );
  OR2_X1 U7881 ( .A1(n7863), .A2(n6577), .ZN(n6265) );
  INV_X1 U7882 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6578) );
  OR2_X1 U7883 ( .A1(n7783), .A2(n6578), .ZN(n6264) );
  NAND4_X1 U7884 ( .A1(n6267), .A2(n6266), .A3(n6265), .A4(n6264), .ZN(n8992)
         );
  INV_X1 U7885 ( .A(n8992), .ZN(n6683) );
  NOR2_X1 U7886 ( .A1(n8666), .A2(n6683), .ZN(n6268) );
  AOI211_X1 U7887 ( .C1(n8668), .C2(n8994), .A(n6269), .B(n6268), .ZN(n6270)
         );
  OAI21_X1 U7888 ( .B1(n8671), .B2(n6526), .A(n6270), .ZN(n6271) );
  AOI21_X1 U7889 ( .B1(n8679), .B2(n6529), .A(n6271), .ZN(n6272) );
  OAI21_X1 U7890 ( .B1(n6273), .B2(n8664), .A(n6272), .ZN(P1_U3229) );
  AND2_X1 U7891 ( .A1(n6316), .A2(n9848), .ZN(n6279) );
  OR2_X1 U7892 ( .A1(n6274), .A2(n6279), .ZN(n6275) );
  AND2_X1 U7893 ( .A1(n7512), .A2(n6277), .ZN(n6278) );
  INV_X1 U7894 ( .A(n6287), .ZN(n6288) );
  NAND2_X1 U7895 ( .A1(n6282), .A2(n7358), .ZN(n6286) );
  OAI22_X1 U7896 ( .A1(n7359), .A2(n9978), .B1(n6283), .B2(n6861), .ZN(n6284)
         );
  INV_X1 U7897 ( .A(n6284), .ZN(n6285) );
  XNOR2_X1 U7898 ( .A(n8065), .B(n7408), .ZN(n7514) );
  INV_X1 U7899 ( .A(n7514), .ZN(n6293) );
  OAI21_X1 U7900 ( .B1(n6288), .B2(n6293), .A(n6973), .ZN(n6587) );
  AOI21_X1 U7901 ( .B1(n7408), .B2(n6289), .A(n9807), .ZN(n6584) );
  INV_X1 U7902 ( .A(n7408), .ZN(n9735) );
  AOI22_X1 U7903 ( .A1(n9813), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n6290), .B2(
        n9802), .ZN(n6291) );
  OAI21_X1 U7904 ( .B1(n9735), .B2(n8398), .A(n6291), .ZN(n6304) );
  NAND2_X2 U7905 ( .A1(n4887), .A2(n7514), .ZN(n9792) );
  OAI21_X1 U7906 ( .B1(n4887), .B2(n7514), .A(n9792), .ZN(n6302) );
  NAND2_X1 U7907 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  AND2_X1 U7908 ( .A1(n6348), .A2(n6296), .ZN(n9801) );
  NAND2_X1 U7909 ( .A1(n7328), .A2(n9801), .ZN(n6300) );
  NAND2_X1 U7910 ( .A1(n4261), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7911 ( .A1(n6657), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7912 ( .A1(n7322), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6297) );
  NAND4_X1 U7913 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n8064)
         );
  NAND2_X1 U7914 ( .A1(n8064), .A2(n9775), .ZN(n6301) );
  OAI21_X1 U7915 ( .B1(n6316), .B2(n8402), .A(n6301), .ZN(n9729) );
  AOI21_X1 U7916 ( .B1(n6302), .B2(n9771), .A(n9729), .ZN(n6586) );
  NOR2_X1 U7917 ( .A1(n6586), .A2(n9813), .ZN(n6303) );
  AOI211_X1 U7918 ( .C1(n6584), .C2(n9809), .A(n6304), .B(n6303), .ZN(n6305)
         );
  OAI21_X1 U7919 ( .B1(n8412), .B2(n6587), .A(n6305), .ZN(P2_U3288) );
  NOR2_X1 U7920 ( .A1(n6306), .A2(n5765), .ZN(n6307) );
  XNOR2_X1 U7921 ( .A(n9844), .B(n7612), .ZN(n6308) );
  NAND2_X1 U7922 ( .A1(n6307), .A2(n6308), .ZN(n6312) );
  INV_X1 U7923 ( .A(n6307), .ZN(n6310) );
  INV_X1 U7924 ( .A(n6308), .ZN(n6309) );
  NAND2_X1 U7925 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  AND2_X1 U7926 ( .A1(n6312), .A2(n6311), .ZN(n7988) );
  NAND2_X1 U7927 ( .A1(n8067), .A2(n7602), .ZN(n6314) );
  XNOR2_X1 U7928 ( .A(n9877), .B(n7612), .ZN(n6313) );
  XNOR2_X1 U7929 ( .A(n6314), .B(n6313), .ZN(n9742) );
  NAND2_X1 U7930 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  NOR2_X1 U7931 ( .A1(n6316), .A2(n5765), .ZN(n6318) );
  XNOR2_X1 U7932 ( .A(n6317), .B(n7607), .ZN(n6319) );
  NAND2_X1 U7933 ( .A1(n6318), .A2(n6319), .ZN(n6331) );
  INV_X1 U7934 ( .A(n6318), .ZN(n6321) );
  INV_X1 U7935 ( .A(n6319), .ZN(n6320) );
  NAND2_X1 U7936 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  NAND2_X1 U7937 ( .A1(n6331), .A2(n6322), .ZN(n6324) );
  INV_X1 U7938 ( .A(n6332), .ZN(n6323) );
  AOI211_X1 U7939 ( .C1(n6325), .C2(n6324), .A(n9744), .B(n6323), .ZN(n6330)
         );
  AOI22_X1 U7940 ( .A1(n9724), .A2(n8067), .B1(n6326), .B2(n8054), .ZN(n6328)
         );
  AND2_X1 U7941 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6838) );
  AOI21_X1 U7942 ( .B1(n9721), .B2(n8065), .A(n6838), .ZN(n6327) );
  OAI211_X1 U7943 ( .C1(n9848), .C2(n9734), .A(n6328), .B(n6327), .ZN(n6329)
         );
  OR2_X1 U7944 ( .A1(n6330), .A2(n6329), .ZN(P2_U3215) );
  NAND2_X1 U7945 ( .A1(n6332), .A2(n6331), .ZN(n6400) );
  XNOR2_X1 U7946 ( .A(n7408), .B(n7607), .ZN(n6341) );
  NAND2_X1 U7947 ( .A1(n8065), .A2(n7602), .ZN(n6340) );
  XNOR2_X1 U7948 ( .A(n6341), .B(n6340), .ZN(n9732) );
  NAND2_X1 U7949 ( .A1(n6333), .A2(n7358), .ZN(n6335) );
  AOI22_X1 U7950 ( .A1(n7335), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5739), .B2(
        n6896), .ZN(n6334) );
  XNOR2_X1 U7951 ( .A(n9854), .B(n7612), .ZN(n6339) );
  INV_X1 U7952 ( .A(n6339), .ZN(n6337) );
  AND2_X1 U7953 ( .A1(n8064), .A2(n7602), .ZN(n6338) );
  INV_X1 U7954 ( .A(n6338), .ZN(n6336) );
  NAND2_X1 U7955 ( .A1(n6337), .A2(n6336), .ZN(n6402) );
  AND2_X1 U7956 ( .A1(n9732), .A2(n6402), .ZN(n6345) );
  INV_X1 U7957 ( .A(n6402), .ZN(n6344) );
  NAND2_X1 U7958 ( .A1(n6339), .A2(n6338), .ZN(n6403) );
  INV_X1 U7959 ( .A(n6340), .ZN(n6342) );
  NAND2_X1 U7960 ( .A1(n6342), .A2(n6341), .ZN(n6401) );
  AND2_X1 U7961 ( .A1(n6403), .A2(n6401), .ZN(n6343) );
  NAND2_X1 U7962 ( .A1(n6443), .A2(n7358), .ZN(n6347) );
  AOI22_X1 U7963 ( .A1(n7335), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5739), .B2(
        n6812), .ZN(n6346) );
  XNOR2_X1 U7964 ( .A(n8506), .B(n7607), .ZN(n6644) );
  NAND2_X1 U7965 ( .A1(n4260), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6354) );
  AND2_X1 U7966 ( .A1(n6348), .A2(n6364), .ZN(n6349) );
  OR2_X1 U7967 ( .A1(n6355), .A2(n6349), .ZN(n6999) );
  INV_X1 U7968 ( .A(n6999), .ZN(n6350) );
  NAND2_X1 U7969 ( .A1(n7328), .A2(n6350), .ZN(n6353) );
  NAND2_X1 U7970 ( .A1(n5451), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U7971 ( .A1(n6657), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6351) );
  NOR2_X1 U7972 ( .A1(n6975), .A2(n5765), .ZN(n6645) );
  XNOR2_X1 U7973 ( .A(n6644), .B(n6645), .ZN(n6648) );
  XNOR2_X1 U7974 ( .A(n6649), .B(n6648), .ZN(n6368) );
  INV_X1 U7975 ( .A(n6355), .ZN(n6357) );
  INV_X1 U7976 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U7977 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  NAND2_X1 U7978 ( .A1(n6655), .A2(n6358), .ZN(n9787) );
  INV_X1 U7979 ( .A(n9787), .ZN(n6359) );
  NAND2_X1 U7980 ( .A1(n7328), .A2(n6359), .ZN(n6363) );
  NAND2_X1 U7981 ( .A1(n4261), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U7982 ( .A1(n7322), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U7983 ( .A1(n6657), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6360) );
  INV_X1 U7984 ( .A(n6976), .ZN(n8063) );
  NOR2_X1 U7985 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6364), .ZN(n6813) );
  INV_X1 U7986 ( .A(n8064), .ZN(n6974) );
  OAI22_X1 U7987 ( .A1(n8021), .A2(n6974), .B1(n6999), .B2(n9752), .ZN(n6365)
         );
  AOI211_X1 U7988 ( .C1(n9721), .C2(n8063), .A(n6813), .B(n6365), .ZN(n6367)
         );
  NAND2_X1 U7989 ( .A1(n9748), .A2(n8506), .ZN(n6366) );
  OAI211_X1 U7990 ( .C1(n6368), .C2(n9744), .A(n6367), .B(n6366), .ZN(P2_U3219) );
  INV_X1 U7991 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6373) );
  INV_X1 U7992 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7776) );
  MUX2_X1 U7993 ( .A(n6373), .B(n7776), .S(n7333), .Z(n6594) );
  XNOR2_X1 U7994 ( .A(n6594), .B(SI_21_), .ZN(n6593) );
  XNOR2_X1 U7995 ( .A(n6592), .B(n6593), .ZN(n7775) );
  INV_X1 U7996 ( .A(n7775), .ZN(n6604) );
  OAI222_X1 U7997 ( .A1(n8539), .A2(n6373), .B1(P2_U3152), .B2(n7539), .C1(
        n8543), .C2(n6604), .ZN(P2_U3337) );
  OAI211_X1 U7998 ( .C1(n6376), .C2(n6375), .A(n4352), .B(n6374), .ZN(n6385)
         );
  INV_X1 U7999 ( .A(n9759), .ZN(n9753) );
  OAI21_X1 U8000 ( .B1(n6379), .B2(n6378), .A(n6377), .ZN(n6383) );
  INV_X1 U8001 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6654) );
  NOR2_X1 U8002 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6654), .ZN(n6382) );
  INV_X1 U8003 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U8004 ( .A1(n8106), .A2(n6380), .ZN(n6381) );
  AOI211_X1 U8005 ( .C1(n9753), .C2(n6383), .A(n6382), .B(n6381), .ZN(n6384)
         );
  OAI211_X1 U8006 ( .C1(n9757), .C2(n6386), .A(n6385), .B(n6384), .ZN(P2_U3257) );
  INV_X1 U8007 ( .A(n6387), .ZN(n6391) );
  INV_X1 U8008 ( .A(n6388), .ZN(n6390) );
  OAI211_X1 U8009 ( .C1(n6391), .C2(n6390), .A(n4352), .B(n6389), .ZN(n6398)
         );
  INV_X1 U8010 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7991) );
  NOR2_X1 U8011 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7991), .ZN(n6396) );
  XNOR2_X1 U8012 ( .A(n6393), .B(n6392), .ZN(n6394) );
  NOR2_X1 U8013 ( .A1(n9759), .A2(n6394), .ZN(n6395) );
  AOI211_X1 U8014 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9754), .A(n6396), .B(
        n6395), .ZN(n6397) );
  OAI211_X1 U8015 ( .C1(n9757), .C2(n6399), .A(n6398), .B(n6397), .ZN(P2_U3250) );
  NAND2_X1 U8016 ( .A1(n6400), .A2(n9732), .ZN(n9731) );
  NAND2_X1 U8017 ( .A1(n9731), .A2(n6401), .ZN(n6405) );
  NAND2_X1 U8018 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  XNOR2_X1 U8019 ( .A(n6405), .B(n6404), .ZN(n6411) );
  INV_X1 U8020 ( .A(n9744), .ZN(n9730) );
  NAND2_X1 U8021 ( .A1(n8065), .A2(n9778), .ZN(n6406) );
  OAI21_X1 U8022 ( .B1(n6975), .B2(n8404), .A(n6406), .ZN(n9799) );
  AND2_X1 U8023 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6888) );
  AOI21_X1 U8024 ( .B1(n9741), .B2(n9799), .A(n6888), .ZN(n6409) );
  INV_X1 U8025 ( .A(n9801), .ZN(n6407) );
  OR2_X1 U8026 ( .A1(n9752), .A2(n6407), .ZN(n6408) );
  OAI211_X1 U8027 ( .C1(n9734), .C2(n9854), .A(n6409), .B(n6408), .ZN(n6410)
         );
  AOI21_X1 U8028 ( .B1(n6411), .B2(n9730), .A(n6410), .ZN(n6412) );
  INV_X1 U8029 ( .A(n6412), .ZN(P2_U3233) );
  NOR2_X1 U8030 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5747), .ZN(n6417) );
  AND3_X1 U8031 ( .A1(n6787), .A2(n6414), .A3(n6413), .ZN(n6415) );
  NOR3_X1 U8032 ( .A1(n9759), .A2(n6430), .A3(n6415), .ZN(n6416) );
  AOI211_X1 U8033 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9754), .A(n6417), .B(
        n6416), .ZN(n6422) );
  OAI211_X1 U8034 ( .C1(n6420), .C2(n6419), .A(n4352), .B(n6418), .ZN(n6421)
         );
  OAI211_X1 U8035 ( .C1(n9757), .C2(n6423), .A(n6422), .B(n6421), .ZN(P2_U3248) );
  INV_X1 U8036 ( .A(n6424), .ZN(n6434) );
  INV_X1 U8037 ( .A(n6425), .ZN(n6429) );
  INV_X1 U8038 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6427) );
  MUX2_X1 U8039 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6427), .S(n6426), .Z(n6428)
         );
  NOR3_X1 U8040 ( .A1(n6430), .A2(n6429), .A3(n6428), .ZN(n6431) );
  NOR3_X1 U8041 ( .A1(n9759), .A2(n6432), .A3(n6431), .ZN(n6433) );
  AOI211_X1 U8042 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9754), .A(n6434), .B(
        n6433), .ZN(n6439) );
  OAI211_X1 U8043 ( .C1(n6437), .C2(n6436), .A(n4352), .B(n6435), .ZN(n6438)
         );
  OAI211_X1 U8044 ( .C1(n9757), .C2(n6440), .A(n6439), .B(n6438), .ZN(P2_U3249) );
  NAND2_X1 U8045 ( .A1(n6443), .A2(n8760), .ZN(n6446) );
  AOI22_X1 U8046 ( .A1(n7734), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7733), .B2(
        n6444), .ZN(n6445) );
  NAND2_X1 U8047 ( .A1(n6580), .A2(n7889), .ZN(n6448) );
  NAND2_X1 U8048 ( .A1(n8992), .A2(n4264), .ZN(n6447) );
  NAND2_X1 U8049 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  XNOR2_X1 U8050 ( .A(n6449), .B(n5361), .ZN(n6452) );
  NAND2_X1 U8051 ( .A1(n6580), .A2(n7891), .ZN(n6451) );
  NAND2_X1 U8052 ( .A1(n5377), .A2(n8992), .ZN(n6450) );
  NAND2_X1 U8053 ( .A1(n6451), .A2(n6450), .ZN(n6453) );
  NAND2_X1 U8054 ( .A1(n6452), .A2(n6453), .ZN(n6667) );
  INV_X1 U8055 ( .A(n6452), .ZN(n6455) );
  INV_X1 U8056 ( .A(n6453), .ZN(n6454) );
  NAND2_X1 U8057 ( .A1(n6455), .A2(n6454), .ZN(n6669) );
  NAND2_X1 U8058 ( .A1(n6667), .A2(n6669), .ZN(n6456) );
  XNOR2_X1 U8059 ( .A(n6668), .B(n6456), .ZN(n6469) );
  NAND2_X1 U8060 ( .A1(n8748), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6463) );
  OR2_X1 U8061 ( .A1(n8753), .A2(n9531), .ZN(n6462) );
  INV_X1 U8062 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6457) );
  AND2_X1 U8063 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  OR2_X1 U8064 ( .A1(n6459), .A2(n6499), .ZN(n6680) );
  OR2_X1 U8065 ( .A1(n7863), .A2(n6680), .ZN(n6461) );
  OR2_X1 U8066 ( .A1(n7783), .A2(n6514), .ZN(n6460) );
  NAND4_X1 U8067 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n8991)
         );
  INV_X1 U8068 ( .A(n8991), .ZN(n6622) );
  NOR2_X1 U8069 ( .A1(n8666), .A2(n6622), .ZN(n6464) );
  AOI211_X1 U8070 ( .C1(n8668), .C2(n8993), .A(n6465), .B(n6464), .ZN(n6466)
         );
  OAI21_X1 U8071 ( .B1(n8671), .B2(n6577), .A(n6466), .ZN(n6467) );
  AOI21_X1 U8072 ( .B1(n8679), .B2(n6580), .A(n6467), .ZN(n6468) );
  OAI21_X1 U8073 ( .B1(n6469), .B2(n8664), .A(n6468), .ZN(P1_U3215) );
  NAND2_X1 U8074 ( .A1(n6470), .A2(n8942), .ZN(n6471) );
  NAND2_X1 U8075 ( .A1(n6472), .A2(n6471), .ZN(n9659) );
  NAND2_X1 U8076 ( .A1(n9659), .A2(n7052), .ZN(n6477) );
  OAI21_X1 U8077 ( .B1(n8942), .B2(n8722), .A(n6473), .ZN(n6474) );
  NAND2_X1 U8078 ( .A1(n6474), .A2(n9348), .ZN(n6476) );
  AOI22_X1 U8079 ( .A1(n9343), .A2(n9002), .B1(n9329), .B2(n8999), .ZN(n6475)
         );
  NAND3_X1 U8080 ( .A1(n6477), .A2(n6476), .A3(n6475), .ZN(n9664) );
  INV_X1 U8081 ( .A(n9664), .ZN(n6486) );
  NAND2_X1 U8082 ( .A1(n7200), .A2(n6481), .ZN(n6478) );
  NAND2_X1 U8083 ( .A1(n9673), .A2(n6478), .ZN(n6480) );
  OR2_X1 U8084 ( .A1(n6480), .A2(n6479), .ZN(n9660) );
  AOI22_X1 U8085 ( .A1(n9364), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9287), .ZN(n6483) );
  NAND2_X1 U8086 ( .A1(n9361), .A2(n6481), .ZN(n6482) );
  OAI211_X1 U8087 ( .C1(n9357), .C2(n9660), .A(n6483), .B(n6482), .ZN(n6484)
         );
  AOI21_X1 U8088 ( .B1(n9373), .B2(n9659), .A(n6484), .ZN(n6485) );
  OAI21_X1 U8089 ( .B1(n9364), .B2(n6486), .A(n6485), .ZN(P1_U3289) );
  NAND2_X1 U8090 ( .A1(n6559), .A2(n6487), .ZN(n6488) );
  NAND2_X1 U8091 ( .A1(n6489), .A2(n6488), .ZN(n6553) );
  NAND2_X1 U8092 ( .A1(n9682), .A2(n8995), .ZN(n8789) );
  NAND2_X1 U8093 ( .A1(n8785), .A2(n8789), .ZN(n8944) );
  INV_X1 U8094 ( .A(n8995), .ZN(n6490) );
  NAND2_X1 U8095 ( .A1(n6490), .A2(n9682), .ZN(n6491) );
  INV_X1 U8096 ( .A(n6547), .ZN(n6543) );
  NAND2_X1 U8097 ( .A1(n6543), .A2(n8994), .ZN(n8702) );
  NAND2_X1 U8098 ( .A1(n6558), .A2(n6547), .ZN(n8800) );
  NAND2_X1 U8099 ( .A1(n6547), .A2(n8994), .ZN(n6492) );
  AND2_X1 U8100 ( .A1(n6529), .A2(n8993), .ZN(n6493) );
  NAND2_X1 U8101 ( .A1(n6580), .A2(n6683), .ZN(n8794) );
  NAND2_X1 U8102 ( .A1(n8701), .A2(n8794), .ZN(n8949) );
  OR2_X1 U8103 ( .A1(n6580), .A2(n8992), .ZN(n6494) );
  NAND2_X1 U8104 ( .A1(n6650), .A2(n8760), .ZN(n6498) );
  AOI22_X1 U8105 ( .A1(n7734), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7733), .B2(
        n6496), .ZN(n6497) );
  OR2_X1 U8106 ( .A1(n6674), .A2(n6622), .ZN(n8697) );
  NAND2_X1 U8107 ( .A1(n6674), .A2(n6622), .ZN(n8692) );
  NAND2_X1 U8108 ( .A1(n8697), .A2(n8692), .ZN(n8950) );
  XNOR2_X1 U8109 ( .A(n6607), .B(n8950), .ZN(n9530) );
  INV_X1 U8110 ( .A(n9530), .ZN(n6519) );
  NAND2_X1 U8111 ( .A1(n8748), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6504) );
  INV_X1 U8112 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6625) );
  OR2_X1 U8113 ( .A1(n7783), .A2(n6625), .ZN(n6503) );
  NAND2_X1 U8114 ( .A1(n6499), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6613) );
  OR2_X1 U8115 ( .A1(n6499), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8116 ( .A1(n6613), .A2(n6500), .ZN(n6942) );
  OR2_X1 U8117 ( .A1(n7863), .A2(n6942), .ZN(n6502) );
  OR2_X1 U8118 ( .A1(n8753), .A2(n5438), .ZN(n6501) );
  NAND4_X1 U8119 ( .A1(n6504), .A2(n6503), .A3(n6502), .A4(n6501), .ZN(n8990)
         );
  INV_X1 U8120 ( .A(n8990), .ZN(n6611) );
  NAND2_X1 U8121 ( .A1(n8786), .A2(n8781), .ZN(n8906) );
  INV_X1 U8122 ( .A(n8906), .ZN(n8726) );
  NAND2_X1 U8123 ( .A1(n6505), .A2(n8726), .ZN(n6508) );
  NAND2_X1 U8124 ( .A1(n8786), .A2(n6506), .ZN(n6507) );
  AND2_X1 U8125 ( .A1(n6507), .A2(n8908), .ZN(n8728) );
  NAND2_X1 U8126 ( .A1(n6508), .A2(n8728), .ZN(n6556) );
  OR2_X2 U8127 ( .A1(n6556), .A2(n8944), .ZN(n6554) );
  INV_X1 U8128 ( .A(n8785), .ZN(n6509) );
  NOR2_X1 U8129 ( .A1(n8945), .A2(n6509), .ZN(n6510) );
  INV_X1 U8130 ( .A(n8993), .ZN(n6511) );
  NOR2_X1 U8131 ( .A1(n6529), .A2(n6511), .ZN(n8700) );
  NAND2_X1 U8132 ( .A1(n6529), .A2(n6511), .ZN(n8793) );
  INV_X1 U8133 ( .A(n8950), .ZN(n8810) );
  XNOR2_X1 U8134 ( .A(n6619), .B(n8810), .ZN(n6512) );
  OAI222_X1 U8135 ( .A1(n9345), .A2(n6611), .B1(n9282), .B2(n6683), .C1(n9280), 
        .C2(n6512), .ZN(n9528) );
  INV_X1 U8137 ( .A(n6580), .ZN(n9485) );
  NAND2_X1 U8138 ( .A1(n6576), .A2(n9485), .ZN(n6575) );
  INV_X1 U8139 ( .A(n6575), .ZN(n6513) );
  INV_X1 U8140 ( .A(n6674), .ZN(n9526) );
  OAI21_X1 U8141 ( .B1(n6513), .B2(n9526), .A(n6623), .ZN(n9527) );
  INV_X1 U8142 ( .A(n9372), .ZN(n9313) );
  OAI22_X1 U8143 ( .A1(n6776), .A2(n6514), .B1(n6680), .B2(n9367), .ZN(n6515)
         );
  AOI21_X1 U8144 ( .B1(n9361), .B2(n6674), .A(n6515), .ZN(n6516) );
  OAI21_X1 U8145 ( .B1(n9527), .B2(n9313), .A(n6516), .ZN(n6517) );
  AOI21_X1 U8146 ( .B1(n9528), .B2(n6776), .A(n6517), .ZN(n6518) );
  OAI21_X1 U8147 ( .B1(n6519), .B2(n9335), .A(n6518), .ZN(P1_U3280) );
  INV_X1 U8148 ( .A(n8793), .ZN(n6520) );
  OR2_X1 U8149 ( .A1(n6520), .A2(n8700), .ZN(n8948) );
  XOR2_X1 U8150 ( .A(n8948), .B(n6521), .Z(n9701) );
  INV_X1 U8151 ( .A(n9701), .ZN(n6533) );
  XOR2_X1 U8152 ( .A(n8948), .B(n6522), .Z(n6523) );
  OAI222_X1 U8153 ( .A1(n9282), .A2(n6558), .B1(n9345), .B2(n6683), .C1(n9280), 
        .C2(n6523), .ZN(n9698) );
  INV_X1 U8154 ( .A(n6529), .ZN(n9695) );
  INV_X1 U8155 ( .A(n6542), .ZN(n6525) );
  INV_X1 U8156 ( .A(n6576), .ZN(n6524) );
  OAI21_X1 U8157 ( .B1(n9695), .B2(n6525), .A(n6524), .ZN(n9697) );
  OAI22_X1 U8158 ( .A1(n6776), .A2(n6527), .B1(n6526), .B2(n9367), .ZN(n6528)
         );
  AOI21_X1 U8159 ( .B1(n9361), .B2(n6529), .A(n6528), .ZN(n6530) );
  OAI21_X1 U8160 ( .B1(n9697), .B2(n9313), .A(n6530), .ZN(n6531) );
  AOI21_X1 U8161 ( .B1(n9698), .B2(n6776), .A(n6531), .ZN(n6532) );
  OAI21_X1 U8162 ( .B1(n6533), .B2(n9335), .A(n6532), .ZN(P1_U3282) );
  INV_X1 U8163 ( .A(n6534), .ZN(n6535) );
  AOI21_X1 U8164 ( .B1(n6538), .B2(n6536), .A(n6535), .ZN(n9692) );
  INV_X1 U8165 ( .A(n9692), .ZN(n6551) );
  NAND2_X1 U8166 ( .A1(n6537), .A2(n9348), .ZN(n6541) );
  AOI21_X1 U8167 ( .B1(n6554), .B2(n8785), .A(n6538), .ZN(n6540) );
  AOI22_X1 U8168 ( .A1(n9329), .A2(n8993), .B1(n9343), .B2(n8995), .ZN(n6539)
         );
  OAI21_X1 U8169 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(n9691) );
  OAI21_X1 U8170 ( .B1(n4612), .B2(n6543), .A(n6542), .ZN(n9689) );
  OAI22_X1 U8171 ( .A1(n6776), .A2(n6545), .B1(n6544), .B2(n9367), .ZN(n6546)
         );
  AOI21_X1 U8172 ( .B1(n9361), .B2(n6547), .A(n6546), .ZN(n6548) );
  OAI21_X1 U8173 ( .B1(n9689), .B2(n9313), .A(n6548), .ZN(n6549) );
  AOI21_X1 U8174 ( .B1(n9691), .B2(n6776), .A(n6549), .ZN(n6550) );
  OAI21_X1 U8175 ( .B1(n6551), .B2(n9335), .A(n6550), .ZN(P1_U3283) );
  OAI21_X1 U8176 ( .B1(n6553), .B2(n8944), .A(n6552), .ZN(n9685) );
  INV_X1 U8177 ( .A(n9685), .ZN(n6569) );
  INV_X1 U8178 ( .A(n6554), .ZN(n6555) );
  AOI21_X1 U8179 ( .B1(n8944), .B2(n6556), .A(n6555), .ZN(n6557) );
  OAI222_X1 U8180 ( .A1(n9282), .A2(n6559), .B1(n9345), .B2(n6558), .C1(n9280), 
        .C2(n6557), .ZN(n9683) );
  OAI211_X1 U8181 ( .C1(n6561), .C2(n9682), .A(n6560), .B(n9673), .ZN(n9681)
         );
  OAI22_X1 U8182 ( .A1(n6776), .A2(n6563), .B1(n6562), .B2(n9367), .ZN(n6564)
         );
  AOI21_X1 U8183 ( .B1(n9361), .B2(n6565), .A(n6564), .ZN(n6566) );
  OAI21_X1 U8184 ( .B1(n9681), .B2(n9357), .A(n6566), .ZN(n6567) );
  AOI21_X1 U8185 ( .B1(n9683), .B2(n6776), .A(n6567), .ZN(n6568) );
  OAI21_X1 U8186 ( .B1(n6569), .B2(n9335), .A(n6568), .ZN(P1_U3284) );
  XNOR2_X1 U8187 ( .A(n6570), .B(n8949), .ZN(n9487) );
  XNOR2_X1 U8188 ( .A(n6571), .B(n8949), .ZN(n6573) );
  AOI22_X1 U8189 ( .A1(n9343), .A2(n8993), .B1(n9329), .B2(n8991), .ZN(n6572)
         );
  OAI21_X1 U8190 ( .B1(n6573), .B2(n9280), .A(n6572), .ZN(n6574) );
  AOI21_X1 U8191 ( .B1(n9487), .B2(n7052), .A(n6574), .ZN(n9489) );
  OAI211_X1 U8192 ( .C1(n6576), .C2(n9485), .A(n9673), .B(n6575), .ZN(n9484)
         );
  OAI22_X1 U8193 ( .A1(n6776), .A2(n6578), .B1(n6577), .B2(n9367), .ZN(n6579)
         );
  AOI21_X1 U8194 ( .B1(n9361), .B2(n6580), .A(n6579), .ZN(n6581) );
  OAI21_X1 U8195 ( .B1(n9484), .B2(n9357), .A(n6581), .ZN(n6582) );
  AOI21_X1 U8196 ( .B1(n9487), .B2(n9373), .A(n6582), .ZN(n6583) );
  OAI21_X1 U8197 ( .B1(n9489), .B2(n9364), .A(n6583), .ZN(P1_U3281) );
  INV_X1 U8198 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6589) );
  AOI22_X1 U8199 ( .A1(n6584), .A2(n9878), .B1(n7408), .B2(n9876), .ZN(n6585)
         );
  OAI211_X1 U8200 ( .C1(n6587), .C2(n9829), .A(n6586), .B(n6585), .ZN(n6590)
         );
  NAND2_X1 U8201 ( .A1(n6590), .A2(n10073), .ZN(n6588) );
  OAI21_X1 U8202 ( .B1(n10073), .B2(n6589), .A(n6588), .ZN(P2_U3475) );
  NAND2_X1 U8203 ( .A1(n6590), .A2(n9889), .ZN(n6591) );
  OAI21_X1 U8204 ( .B1(n9889), .B2(n6095), .A(n6591), .ZN(P2_U3528) );
  INV_X1 U8205 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7794) );
  INV_X1 U8206 ( .A(n6594), .ZN(n6595) );
  NAND2_X1 U8207 ( .A1(n6595), .A2(SI_21_), .ZN(n6596) );
  INV_X1 U8208 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6603) );
  MUX2_X1 U8209 ( .A(n6603), .B(n7794), .S(n7333), .Z(n6598) );
  INV_X1 U8210 ( .A(SI_22_), .ZN(n6597) );
  NAND2_X1 U8211 ( .A1(n6598), .A2(n6597), .ZN(n6690) );
  INV_X1 U8212 ( .A(n6598), .ZN(n6599) );
  NAND2_X1 U8213 ( .A1(n6599), .A2(SI_22_), .ZN(n6600) );
  NAND2_X1 U8214 ( .A1(n6690), .A2(n6600), .ZN(n6688) );
  XNOR2_X1 U8215 ( .A(n6689), .B(n6688), .ZN(n7793) );
  INV_X1 U8216 ( .A(n7793), .ZN(n6602) );
  OAI222_X1 U8217 ( .A1(n9478), .A2(n7794), .B1(n7551), .B2(n6602), .C1(
        P1_U3084), .C2(n4259), .ZN(P1_U3331) );
  OAI222_X1 U8218 ( .A1(n8539), .A2(n6603), .B1(n7920), .B2(n6602), .C1(n6601), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  OAI222_X1 U8219 ( .A1(n4258), .A2(n5262), .B1(n7551), .B2(n6604), .C1(n7776), 
        .C2(n7154), .ZN(P1_U3332) );
  NOR2_X1 U8220 ( .A1(n6674), .A2(n8991), .ZN(n6606) );
  NAND2_X1 U8221 ( .A1(n6674), .A2(n8991), .ZN(n6605) );
  NAND2_X1 U8222 ( .A1(n6739), .A2(n8760), .ZN(n6610) );
  AOI22_X1 U8223 ( .A1(n7734), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7733), .B2(
        n6608), .ZN(n6609) );
  NAND2_X1 U8224 ( .A1(n9455), .A2(n6611), .ZN(n8798) );
  NAND2_X1 U8225 ( .A1(n8818), .A2(n8798), .ZN(n6756) );
  XNOR2_X1 U8226 ( .A(n6757), .B(n6756), .ZN(n9458) );
  NAND2_X1 U8227 ( .A1(n8748), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6618) );
  INV_X1 U8228 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6775) );
  OR2_X1 U8229 ( .A1(n7783), .A2(n6775), .ZN(n6617) );
  INV_X1 U8230 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U8231 ( .A1(n6613), .A2(n6612), .ZN(n6614) );
  NAND2_X1 U8232 ( .A1(n6764), .A2(n6614), .ZN(n6967) );
  OR2_X1 U8233 ( .A1(n7863), .A2(n6967), .ZN(n6616) );
  OR2_X1 U8234 ( .A1(n8753), .A2(n9525), .ZN(n6615) );
  NAND4_X1 U8235 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n8989)
         );
  INV_X1 U8236 ( .A(n8989), .ZN(n6939) );
  NAND2_X1 U8237 ( .A1(n6619), .A2(n8692), .ZN(n6620) );
  INV_X1 U8238 ( .A(n6756), .ZN(n8953) );
  XNOR2_X1 U8239 ( .A(n6761), .B(n8953), .ZN(n6621) );
  OAI222_X1 U8240 ( .A1(n9282), .A2(n6622), .B1(n9345), .B2(n6939), .C1(n9280), 
        .C2(n6621), .ZN(n9453) );
  NAND2_X1 U8241 ( .A1(n9453), .A2(n6776), .ZN(n6629) );
  AOI211_X1 U8242 ( .C1(n9455), .C2(n6623), .A(n9696), .B(n6773), .ZN(n9454)
         );
  INV_X1 U8243 ( .A(n9455), .ZN(n6624) );
  NOR2_X1 U8244 ( .A1(n6624), .A2(n9369), .ZN(n6627) );
  OAI22_X1 U8245 ( .A1(n6776), .A2(n6625), .B1(n6942), .B2(n9367), .ZN(n6626)
         );
  AOI211_X1 U8246 ( .C1(n9454), .C2(n9211), .A(n6627), .B(n6626), .ZN(n6628)
         );
  OAI211_X1 U8247 ( .C1(n9458), .C2(n9335), .A(n6629), .B(n6628), .ZN(P1_U3279) );
  AOI21_X1 U8248 ( .B1(n6631), .B2(n9499), .A(n6630), .ZN(n6633) );
  INV_X1 U8249 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6949) );
  AOI22_X1 U8250 ( .A1(n7091), .A2(n6949), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n6950), .ZN(n6632) );
  NOR2_X1 U8251 ( .A1(n6633), .A2(n6632), .ZN(n6948) );
  AOI21_X1 U8252 ( .B1(n6633), .B2(n6632), .A(n6948), .ZN(n6643) );
  INV_X1 U8253 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6634) );
  AOI22_X1 U8254 ( .A1(n7091), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n6634), .B2(
        n6950), .ZN(n6637) );
  NAND2_X1 U8255 ( .A1(n6637), .A2(n6636), .ZN(n6946) );
  OAI21_X1 U8256 ( .B1(n6637), .B2(n6636), .A(n6946), .ZN(n6641) );
  NOR2_X1 U8257 ( .A1(n9757), .A2(n6950), .ZN(n6640) );
  INV_X1 U8258 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U8259 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7111) );
  OAI21_X1 U8260 ( .B1(n8106), .B2(n6638), .A(n7111), .ZN(n6639) );
  AOI211_X1 U8261 ( .C1(n6641), .C2(n4352), .A(n6640), .B(n6639), .ZN(n6642)
         );
  OAI21_X1 U8262 ( .B1(n6643), .B2(n9759), .A(n6642), .ZN(P2_U3259) );
  INV_X1 U8263 ( .A(n6644), .ZN(n6647) );
  INV_X1 U8264 ( .A(n6645), .ZN(n6646) );
  OAI22_X1 U8265 ( .A1(n6649), .A2(n6648), .B1(n6647), .B2(n6646), .ZN(n6733)
         );
  NAND2_X1 U8266 ( .A1(n6650), .A2(n7358), .ZN(n6653) );
  AOI22_X1 U8267 ( .A1(n7335), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5739), .B2(
        n6651), .ZN(n6652) );
  NAND2_X1 U8268 ( .A1(n6653), .A2(n6652), .ZN(n9765) );
  XNOR2_X1 U8269 ( .A(n9765), .B(n7612), .ZN(n6734) );
  NOR2_X1 U8270 ( .A1(n6976), .A2(n5765), .ZN(n6735) );
  XNOR2_X1 U8271 ( .A(n6734), .B(n6735), .ZN(n6732) );
  XNOR2_X1 U8272 ( .A(n6733), .B(n6732), .ZN(n6666) );
  NAND2_X1 U8273 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  AND2_X1 U8274 ( .A1(n6744), .A2(n6656), .ZN(n6980) );
  NAND2_X1 U8275 ( .A1(n7328), .A2(n6980), .ZN(n6661) );
  NAND2_X1 U8276 ( .A1(n4261), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8277 ( .A1(n7322), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U8278 ( .A1(n6657), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6658) );
  INV_X1 U8279 ( .A(n7024), .ZN(n9776) );
  OAI22_X1 U8280 ( .A1(n8021), .A2(n6975), .B1(n9787), .B2(n9752), .ZN(n6662)
         );
  AOI211_X1 U8281 ( .C1(n9721), .C2(n9776), .A(n6663), .B(n6662), .ZN(n6665)
         );
  NAND2_X1 U8282 ( .A1(n9748), .A2(n9765), .ZN(n6664) );
  OAI211_X1 U8283 ( .C1(n6666), .C2(n9744), .A(n6665), .B(n6664), .ZN(P2_U3238) );
  NAND2_X1 U8284 ( .A1(n6674), .A2(n7889), .ZN(n6671) );
  NAND2_X1 U8285 ( .A1(n8991), .A2(n7891), .ZN(n6670) );
  NAND2_X1 U8286 ( .A1(n6671), .A2(n6670), .ZN(n6672) );
  XNOR2_X1 U8287 ( .A(n6672), .B(n7872), .ZN(n6930) );
  AND2_X1 U8288 ( .A1(n5377), .A2(n8991), .ZN(n6673) );
  AOI21_X1 U8289 ( .B1(n6674), .B2(n4264), .A(n6673), .ZN(n6931) );
  XNOR2_X1 U8290 ( .A(n6930), .B(n6931), .ZN(n6676) );
  AOI21_X1 U8291 ( .B1(n6675), .B2(n6676), .A(n8664), .ZN(n6679) );
  INV_X1 U8292 ( .A(n6675), .ZN(n6678) );
  INV_X1 U8293 ( .A(n6676), .ZN(n6677) );
  NAND2_X1 U8294 ( .A1(n6679), .A2(n6935), .ZN(n6687) );
  INV_X1 U8295 ( .A(n6680), .ZN(n6685) );
  AOI21_X1 U8296 ( .B1(n8659), .B2(n8990), .A(n6681), .ZN(n6682) );
  OAI21_X1 U8297 ( .B1(n8598), .B2(n6683), .A(n6682), .ZN(n6684) );
  AOI21_X1 U8298 ( .B1(n6685), .B2(n8618), .A(n6684), .ZN(n6686) );
  OAI211_X1 U8299 ( .C1(n9526), .C2(n8653), .A(n6687), .B(n6686), .ZN(P1_U3234) );
  INV_X1 U8300 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6691) );
  INV_X1 U8301 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7654) );
  MUX2_X1 U8302 ( .A(n6691), .B(n7654), .S(n7333), .Z(n6693) );
  INV_X1 U8303 ( .A(SI_23_), .ZN(n6692) );
  NAND2_X1 U8304 ( .A1(n6693), .A2(n6692), .ZN(n6846) );
  INV_X1 U8305 ( .A(n6693), .ZN(n6694) );
  NAND2_X1 U8306 ( .A1(n6694), .A2(SI_23_), .ZN(n6695) );
  AND2_X1 U8307 ( .A1(n6846), .A2(n6695), .ZN(n6844) );
  INV_X1 U8308 ( .A(n7653), .ZN(n6698) );
  NAND2_X1 U8309 ( .A1(n6696), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6697) );
  OAI211_X1 U8310 ( .C1(n6698), .C2(n7920), .A(n7549), .B(n6697), .ZN(P2_U3335) );
  INV_X1 U8311 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10084) );
  NOR2_X1 U8312 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6699) );
  AOI21_X1 U8313 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6699), .ZN(n9897) );
  NOR2_X1 U8314 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6700) );
  AOI21_X1 U8315 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6700), .ZN(n9900) );
  NOR2_X1 U8316 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6701) );
  AOI21_X1 U8317 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6701), .ZN(n9903) );
  NOR2_X1 U8318 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6702) );
  AOI21_X1 U8319 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6702), .ZN(n9906) );
  NOR2_X1 U8320 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6703) );
  AOI21_X1 U8321 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6703), .ZN(n9909) );
  NOR2_X1 U8322 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6710) );
  XNOR2_X1 U8323 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10094) );
  NAND2_X1 U8324 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6708) );
  XOR2_X1 U8325 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10092) );
  NAND2_X1 U8326 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6706) );
  XOR2_X1 U8327 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10087) );
  AOI21_X1 U8328 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9890) );
  INV_X1 U8329 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6704) );
  NAND3_X1 U8330 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9892) );
  OAI21_X1 U8331 ( .B1(n9890), .B2(n6704), .A(n9892), .ZN(n10086) );
  NAND2_X1 U8332 ( .A1(n10087), .A2(n10086), .ZN(n6705) );
  NAND2_X1 U8333 ( .A1(n6706), .A2(n6705), .ZN(n10091) );
  NAND2_X1 U8334 ( .A1(n10092), .A2(n10091), .ZN(n6707) );
  NAND2_X1 U8335 ( .A1(n6708), .A2(n6707), .ZN(n10093) );
  NOR2_X1 U8336 ( .A1(n10094), .A2(n10093), .ZN(n6709) );
  NOR2_X1 U8337 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  NOR2_X1 U8338 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6711), .ZN(n10079) );
  AND2_X1 U8339 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6711), .ZN(n10078) );
  NOR2_X1 U8340 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10078), .ZN(n6712) );
  NOR2_X1 U8341 ( .A1(n10079), .A2(n6712), .ZN(n6713) );
  NAND2_X1 U8342 ( .A1(n6713), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6715) );
  XOR2_X1 U8343 ( .A(n6713), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10076) );
  NAND2_X1 U8344 ( .A1(n10076), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U8345 ( .A1(n6715), .A2(n6714), .ZN(n6716) );
  NAND2_X1 U8346 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n6716), .ZN(n6718) );
  XOR2_X1 U8347 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n6716), .Z(n10077) );
  NAND2_X1 U8348 ( .A1(n10077), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U8349 ( .A1(n6718), .A2(n6717), .ZN(n6719) );
  NAND2_X1 U8350 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n6719), .ZN(n6721) );
  XOR2_X1 U8351 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n6719), .Z(n10081) );
  NAND2_X1 U8352 ( .A1(n10081), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U8353 ( .A1(n6721), .A2(n6720), .ZN(n6722) );
  AND2_X1 U8354 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6722), .ZN(n6723) );
  XNOR2_X1 U8355 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n6722), .ZN(n10089) );
  NOR2_X1 U8356 ( .A1(n10090), .A2(n10089), .ZN(n10088) );
  NOR2_X1 U8357 ( .A1(n6723), .A2(n10088), .ZN(n9918) );
  NAND2_X1 U8358 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n6724) );
  OAI21_X1 U8359 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6724), .ZN(n9917) );
  NOR2_X1 U8360 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  AOI21_X1 U8361 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9916), .ZN(n9915) );
  NAND2_X1 U8362 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n6725) );
  OAI21_X1 U8363 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6725), .ZN(n9914) );
  NOR2_X1 U8364 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  AOI21_X1 U8365 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9913), .ZN(n9912) );
  NOR2_X1 U8366 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6726) );
  AOI21_X1 U8367 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6726), .ZN(n9911) );
  NAND2_X1 U8368 ( .A1(n9912), .A2(n9911), .ZN(n9910) );
  OAI21_X1 U8369 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9910), .ZN(n9908) );
  NAND2_X1 U8370 ( .A1(n9909), .A2(n9908), .ZN(n9907) );
  OAI21_X1 U8371 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9907), .ZN(n9905) );
  NAND2_X1 U8372 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  OAI21_X1 U8373 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9904), .ZN(n9902) );
  NAND2_X1 U8374 ( .A1(n9903), .A2(n9902), .ZN(n9901) );
  OAI21_X1 U8375 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9901), .ZN(n9899) );
  NAND2_X1 U8376 ( .A1(n9900), .A2(n9899), .ZN(n9898) );
  OAI21_X1 U8377 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9898), .ZN(n9896) );
  NAND2_X1 U8378 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  OAI21_X1 U8379 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9895), .ZN(n10083) );
  NOR2_X1 U8380 ( .A1(n10084), .A2(n10083), .ZN(n6727) );
  NAND2_X1 U8381 ( .A1(n10084), .A2(n10083), .ZN(n10082) );
  OAI21_X1 U8382 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n6727), .A(n10082), .ZN(
        n6729) );
  XNOR2_X1 U8383 ( .A(n7190), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6728) );
  XNOR2_X1 U8384 ( .A(n6729), .B(n6728), .ZN(ADD_1071_U4) );
  NAND2_X1 U8385 ( .A1(n7653), .A2(n9481), .ZN(n6731) );
  NOR2_X1 U8386 ( .A1(n6730), .A2(n4258), .ZN(n8977) );
  INV_X1 U8387 ( .A(n8977), .ZN(n8982) );
  OAI211_X1 U8388 ( .C1(n7654), .C2(n9478), .A(n6731), .B(n8982), .ZN(P1_U3330) );
  NAND2_X1 U8389 ( .A1(n6733), .A2(n6732), .ZN(n6738) );
  INV_X1 U8390 ( .A(n6734), .ZN(n6736) );
  NAND2_X1 U8391 ( .A1(n6736), .A2(n6735), .ZN(n6737) );
  NAND2_X1 U8392 ( .A1(n6738), .A2(n6737), .ZN(n6866) );
  NAND2_X1 U8393 ( .A1(n6739), .A2(n7358), .ZN(n6742) );
  AOI22_X1 U8394 ( .A1(n7335), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5739), .B2(
        n6740), .ZN(n6741) );
  NAND2_X2 U8395 ( .A1(n6742), .A2(n6741), .ZN(n8501) );
  XNOR2_X1 U8396 ( .A(n8501), .B(n7612), .ZN(n6867) );
  NOR2_X1 U8397 ( .A1(n7024), .A2(n5765), .ZN(n6868) );
  XNOR2_X1 U8398 ( .A(n6867), .B(n6868), .ZN(n6865) );
  XNOR2_X1 U8399 ( .A(n6866), .B(n6865), .ZN(n6755) );
  INV_X1 U8400 ( .A(n6980), .ZN(n6752) );
  NAND2_X1 U8401 ( .A1(n6744), .A2(n6743), .ZN(n6745) );
  AND2_X1 U8402 ( .A1(n6876), .A2(n6745), .ZN(n7032) );
  NAND2_X1 U8403 ( .A1(n7328), .A2(n7032), .ZN(n6749) );
  NAND2_X1 U8404 ( .A1(n4261), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U8405 ( .A1(n7322), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U8406 ( .A1(n6657), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6746) );
  OR2_X1 U8407 ( .A1(n6976), .A2(n8402), .ZN(n6750) );
  OAI21_X1 U8408 ( .B1(n8403), .B2(n8404), .A(n6750), .ZN(n6987) );
  AOI22_X1 U8409 ( .A1(n9741), .A2(n6987), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n6751) );
  OAI21_X1 U8410 ( .B1(n6752), .B2(n9752), .A(n6751), .ZN(n6753) );
  AOI21_X1 U8411 ( .B1(n9748), .B2(n8501), .A(n6753), .ZN(n6754) );
  OAI21_X1 U8412 ( .B1(n6755), .B2(n9744), .A(n6754), .ZN(P2_U3226) );
  NAND2_X1 U8413 ( .A1(n6871), .A2(n8760), .ZN(n6759) );
  AOI22_X1 U8414 ( .A1(n7734), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7733), .B2(
        n9571), .ZN(n6758) );
  OR2_X1 U8415 ( .A1(n6969), .A2(n6939), .ZN(n8807) );
  NAND2_X1 U8416 ( .A1(n6969), .A2(n6939), .ZN(n8691) );
  XNOR2_X1 U8417 ( .A(n6903), .B(n8954), .ZN(n9522) );
  INV_X1 U8418 ( .A(n8818), .ZN(n6760) );
  INV_X1 U8419 ( .A(n8954), .ZN(n6762) );
  XNOR2_X1 U8420 ( .A(n6908), .B(n6762), .ZN(n6771) );
  NAND2_X1 U8421 ( .A1(n8748), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6769) );
  OR2_X1 U8422 ( .A1(n8753), .A2(n9518), .ZN(n6768) );
  AND2_X1 U8423 ( .A1(n6764), .A2(n6763), .ZN(n6765) );
  OR2_X1 U8424 ( .A1(n6765), .A2(n6912), .ZN(n7086) );
  OR2_X1 U8425 ( .A1(n7863), .A2(n7086), .ZN(n6767) );
  OR2_X1 U8426 ( .A1(n7783), .A2(n9953), .ZN(n6766) );
  NAND4_X1 U8427 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n8988)
         );
  AOI22_X1 U8428 ( .A1(n9343), .A2(n8990), .B1(n9329), .B2(n8988), .ZN(n6770)
         );
  OAI21_X1 U8429 ( .B1(n6771), .B2(n9280), .A(n6770), .ZN(n6772) );
  AOI21_X1 U8430 ( .B1(n9522), .B2(n7052), .A(n6772), .ZN(n9524) );
  INV_X1 U8431 ( .A(n6969), .ZN(n9519) );
  NOR2_X1 U8432 ( .A1(n6773), .A2(n9519), .ZN(n6774) );
  OR2_X1 U8433 ( .A1(n6920), .A2(n6774), .ZN(n9520) );
  OAI22_X1 U8434 ( .A1(n6776), .A2(n6775), .B1(n6967), .B2(n9367), .ZN(n6777)
         );
  AOI21_X1 U8435 ( .B1(n6969), .B2(n9361), .A(n6777), .ZN(n6778) );
  OAI21_X1 U8436 ( .B1(n9520), .B2(n9313), .A(n6778), .ZN(n6779) );
  AOI21_X1 U8437 ( .B1(n9522), .B2(n9373), .A(n6779), .ZN(n6780) );
  OAI21_X1 U8438 ( .B1(n9524), .B2(n9364), .A(n6780), .ZN(P1_U3278) );
  AOI211_X1 U8439 ( .C1(n6783), .C2(n6782), .A(n6781), .B(n8091), .ZN(n6792)
         );
  AOI22_X1 U8440 ( .A1(n9754), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n6789) );
  NAND3_X1 U8441 ( .A1(n6823), .A2(n6785), .A3(n6784), .ZN(n6786) );
  NAND3_X1 U8442 ( .A1(n9753), .A2(n6787), .A3(n6786), .ZN(n6788) );
  OAI211_X1 U8443 ( .C1(n9757), .C2(n6790), .A(n6789), .B(n6788), .ZN(n6791)
         );
  OR2_X1 U8444 ( .A1(n6792), .A2(n6791), .ZN(P2_U3247) );
  AOI211_X1 U8445 ( .C1(n6795), .C2(n6794), .A(n6793), .B(n8091), .ZN(n6805)
         );
  INV_X1 U8446 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6796) );
  NOR2_X1 U8447 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6796), .ZN(n6797) );
  AOI21_X1 U8448 ( .B1(n9754), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6797), .ZN(
        n6802) );
  OAI211_X1 U8449 ( .C1(n6800), .C2(n6799), .A(n9753), .B(n6798), .ZN(n6801)
         );
  OAI211_X1 U8450 ( .C1(n9757), .C2(n6803), .A(n6802), .B(n6801), .ZN(n6804)
         );
  OR2_X1 U8451 ( .A1(n6805), .A2(n6804), .ZN(P2_U3251) );
  AOI211_X1 U8452 ( .C1(n6808), .C2(n6807), .A(n6806), .B(n8091), .ZN(n6818)
         );
  OAI21_X1 U8453 ( .B1(n6811), .B2(n6810), .A(n6809), .ZN(n6816) );
  NAND2_X1 U8454 ( .A1(n8109), .A2(n6812), .ZN(n6815) );
  AOI21_X1 U8455 ( .B1(n9754), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6813), .ZN(
        n6814) );
  OAI211_X1 U8456 ( .C1(n9759), .C2(n6816), .A(n6815), .B(n6814), .ZN(n6817)
         );
  OR2_X1 U8457 ( .A1(n6818), .A2(n6817), .ZN(P2_U3255) );
  AOI211_X1 U8458 ( .C1(n6821), .C2(n6820), .A(n6819), .B(n8091), .ZN(n6830)
         );
  AOI22_X1 U8459 ( .A1(n9754), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n6827) );
  INV_X1 U8460 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6822) );
  INV_X1 U8461 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U8462 ( .A1(n6822), .A2(n9870), .ZN(n6825) );
  OAI211_X1 U8463 ( .C1(n6825), .C2(n6824), .A(n9753), .B(n6823), .ZN(n6826)
         );
  OAI211_X1 U8464 ( .C1(n9757), .C2(n6828), .A(n6827), .B(n6826), .ZN(n6829)
         );
  OR2_X1 U8465 ( .A1(n6830), .A2(n6829), .ZN(P2_U3246) );
  AOI211_X1 U8466 ( .C1(n6833), .C2(n6832), .A(n6831), .B(n8091), .ZN(n6843)
         );
  OAI21_X1 U8467 ( .B1(n6836), .B2(n6835), .A(n6834), .ZN(n6841) );
  NAND2_X1 U8468 ( .A1(n8109), .A2(n6837), .ZN(n6840) );
  AOI21_X1 U8469 ( .B1(n9754), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6838), .ZN(
        n6839) );
  OAI211_X1 U8470 ( .C1(n9759), .C2(n6841), .A(n6840), .B(n6839), .ZN(n6842)
         );
  OR2_X1 U8471 ( .A1(n6843), .A2(n6842), .ZN(P2_U3252) );
  INV_X1 U8472 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n6848) );
  INV_X1 U8473 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7816) );
  MUX2_X1 U8474 ( .A(n6848), .B(n7816), .S(n7333), .Z(n7061) );
  XNOR2_X1 U8475 ( .A(n7061), .B(SI_24_), .ZN(n7060) );
  XNOR2_X1 U8476 ( .A(n7065), .B(n7060), .ZN(n7815) );
  INV_X1 U8477 ( .A(n7815), .ZN(n7157) );
  OAI222_X1 U8478 ( .A1(P2_U3152), .A2(n6849), .B1(n7920), .B2(n7157), .C1(
        n6848), .C2(n8539), .ZN(P2_U3334) );
  AOI211_X1 U8479 ( .C1(n6852), .C2(n6851), .A(n6850), .B(n8091), .ZN(n6864)
         );
  INV_X1 U8480 ( .A(n6853), .ZN(n6857) );
  MUX2_X1 U8481 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6095), .S(n6861), .Z(n6856)
         );
  INV_X1 U8482 ( .A(n6854), .ZN(n6855) );
  AOI211_X1 U8483 ( .C1(n6857), .C2(n6856), .A(n9759), .B(n6855), .ZN(n6863)
         );
  INV_X1 U8484 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6858) );
  NOR2_X1 U8485 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6858), .ZN(n6859) );
  AOI21_X1 U8486 ( .B1(n9754), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6859), .ZN(
        n6860) );
  OAI21_X1 U8487 ( .B1(n9757), .B2(n6861), .A(n6860), .ZN(n6862) );
  OR3_X1 U8488 ( .A1(n6864), .A2(n6863), .A3(n6862), .ZN(P2_U3253) );
  INV_X1 U8489 ( .A(n6867), .ZN(n6869) );
  NAND2_X1 U8490 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  NAND2_X1 U8491 ( .A1(n6871), .A2(n7358), .ZN(n6874) );
  AOI22_X1 U8492 ( .A1(n7335), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5739), .B2(
        n6872), .ZN(n6873) );
  XNOR2_X1 U8493 ( .A(n9493), .B(n7612), .ZN(n7101) );
  NOR2_X1 U8494 ( .A1(n8403), .A2(n5765), .ZN(n7102) );
  XNOR2_X1 U8495 ( .A(n7101), .B(n7102), .ZN(n7099) );
  XNOR2_X1 U8496 ( .A(n7100), .B(n7099), .ZN(n6887) );
  NAND2_X1 U8497 ( .A1(n4261), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6881) );
  INV_X1 U8498 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8499 ( .A1(n6876), .A2(n6875), .ZN(n6877) );
  AND2_X1 U8500 ( .A1(n7134), .A2(n6877), .ZN(n8396) );
  NAND2_X1 U8501 ( .A1(n7328), .A2(n8396), .ZN(n6880) );
  NAND2_X1 U8502 ( .A1(n7322), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U8503 ( .A1(n6657), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6878) );
  NAND4_X1 U8504 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n8384)
         );
  INV_X1 U8505 ( .A(n7032), .ZN(n6882) );
  OAI22_X1 U8506 ( .A1(n8021), .A2(n7024), .B1(n6882), .B2(n9752), .ZN(n6883)
         );
  AOI211_X1 U8507 ( .C1(n9721), .C2(n8384), .A(n6884), .B(n6883), .ZN(n6886)
         );
  NAND2_X1 U8508 ( .A1(n9493), .A2(n9748), .ZN(n6885) );
  OAI211_X1 U8509 ( .C1(n6887), .C2(n9744), .A(n6886), .B(n6885), .ZN(P2_U3236) );
  INV_X1 U8510 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6890) );
  INV_X1 U8511 ( .A(n6888), .ZN(n6889) );
  OAI21_X1 U8512 ( .B1(n8106), .B2(n6890), .A(n6889), .ZN(n6895) );
  AOI211_X1 U8513 ( .C1(n6893), .C2(n6892), .A(n6891), .B(n8091), .ZN(n6894)
         );
  AOI211_X1 U8514 ( .C1(n8109), .C2(n6896), .A(n6895), .B(n6894), .ZN(n6901)
         );
  OAI211_X1 U8515 ( .C1(n6899), .C2(n6898), .A(n9753), .B(n6897), .ZN(n6900)
         );
  NAND2_X1 U8516 ( .A1(n6901), .A2(n6900), .ZN(P2_U3254) );
  OR2_X1 U8517 ( .A1(n6969), .A2(n8989), .ZN(n6902) );
  NAND2_X1 U8518 ( .A1(n6969), .A2(n8989), .ZN(n6904) );
  NAND2_X1 U8519 ( .A1(n7090), .A2(n8760), .ZN(n6907) );
  AOI22_X1 U8520 ( .A1(n7734), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7733), .B2(
        n6905), .ZN(n6906) );
  INV_X1 U8521 ( .A(n8988), .ZN(n8689) );
  XNOR2_X1 U8522 ( .A(n8690), .B(n8689), .ZN(n8956) );
  XOR2_X1 U8523 ( .A(n7038), .B(n8956), .Z(n9517) );
  INV_X1 U8524 ( .A(n9517), .ZN(n6925) );
  NAND2_X1 U8525 ( .A1(n6910), .A2(n8956), .ZN(n6911) );
  NAND3_X1 U8526 ( .A1(n7042), .A2(n9348), .A3(n6911), .ZN(n6919) );
  NAND2_X1 U8527 ( .A1(n8748), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6917) );
  INV_X1 U8528 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9053) );
  OR2_X1 U8529 ( .A1(n8753), .A2(n9053), .ZN(n6916) );
  NOR2_X1 U8530 ( .A1(n6912), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6913) );
  OR2_X1 U8531 ( .A1(n7043), .A2(n6913), .ZN(n8670) );
  OR2_X1 U8532 ( .A1(n7863), .A2(n8670), .ZN(n6915) );
  INV_X1 U8533 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7055) );
  OR2_X1 U8534 ( .A1(n7783), .A2(n7055), .ZN(n6914) );
  NAND4_X1 U8535 ( .A1(n6917), .A2(n6916), .A3(n6915), .A4(n6914), .ZN(n9342)
         );
  AOI22_X1 U8536 ( .A1(n9343), .A2(n8989), .B1(n9329), .B2(n9342), .ZN(n6918)
         );
  NAND2_X1 U8537 ( .A1(n6919), .A2(n6918), .ZN(n9516) );
  INV_X1 U8538 ( .A(n8690), .ZN(n9514) );
  NAND2_X1 U8539 ( .A1(n6920), .A2(n9514), .ZN(n7053) );
  OAI211_X1 U8540 ( .C1(n6920), .C2(n9514), .A(n9673), .B(n7053), .ZN(n9513)
         );
  OAI22_X1 U8541 ( .A1(n6776), .A2(n9953), .B1(n7086), .B2(n9367), .ZN(n6921)
         );
  AOI21_X1 U8542 ( .B1(n8690), .B2(n9361), .A(n6921), .ZN(n6922) );
  OAI21_X1 U8543 ( .B1(n9513), .B2(n9357), .A(n6922), .ZN(n6923) );
  AOI21_X1 U8544 ( .B1(n9516), .B2(n6776), .A(n6923), .ZN(n6924) );
  OAI21_X1 U8545 ( .B1(n6925), .B2(n9335), .A(n6924), .ZN(P1_U3277) );
  NAND2_X1 U8546 ( .A1(n9455), .A2(n7889), .ZN(n6927) );
  NAND2_X1 U8547 ( .A1(n8990), .A2(n4264), .ZN(n6926) );
  NAND2_X1 U8548 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  XNOR2_X1 U8549 ( .A(n6928), .B(n7872), .ZN(n6959) );
  AND2_X1 U8550 ( .A1(n5377), .A2(n8990), .ZN(n6929) );
  AOI21_X1 U8551 ( .B1(n9455), .B2(n7891), .A(n6929), .ZN(n6958) );
  XNOR2_X1 U8552 ( .A(n6959), .B(n6958), .ZN(n6937) );
  INV_X1 U8553 ( .A(n6930), .ZN(n6933) );
  INV_X1 U8554 ( .A(n6931), .ZN(n6932) );
  NAND2_X1 U8555 ( .A1(n6933), .A2(n6932), .ZN(n6934) );
  AOI21_X1 U8556 ( .B1(n6937), .B2(n6936), .A(n4347), .ZN(n6945) );
  OAI21_X1 U8557 ( .B1(n8666), .B2(n6939), .A(n6938), .ZN(n6940) );
  AOI21_X1 U8558 ( .B1(n8668), .B2(n8991), .A(n6940), .ZN(n6941) );
  OAI21_X1 U8559 ( .B1(n8671), .B2(n6942), .A(n6941), .ZN(n6943) );
  AOI21_X1 U8560 ( .B1(n8679), .B2(n9455), .A(n6943), .ZN(n6944) );
  OAI21_X1 U8561 ( .B1(n6945), .B2(n8664), .A(n6944), .ZN(P1_U3222) );
  INV_X1 U8562 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9966) );
  OAI21_X1 U8563 ( .B1(n6947), .B2(n9966), .A(n7162), .ZN(n6956) );
  AOI21_X1 U8564 ( .B1(n6950), .B2(n6949), .A(n6948), .ZN(n7168) );
  XNOR2_X1 U8565 ( .A(n7168), .B(n7161), .ZN(n6951) );
  NAND2_X1 U8566 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n6951), .ZN(n7170) );
  OAI211_X1 U8567 ( .C1(n6951), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9753), .B(
        n7170), .ZN(n6954) );
  AND2_X1 U8568 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6952) );
  AOI21_X1 U8569 ( .B1(n9754), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n6952), .ZN(
        n6953) );
  OAI211_X1 U8570 ( .C1(n9757), .C2(n7161), .A(n6954), .B(n6953), .ZN(n6955)
         );
  AOI21_X1 U8571 ( .B1(n4352), .B2(n6956), .A(n6955), .ZN(n6957) );
  INV_X1 U8572 ( .A(n6957), .ZN(P2_U3260) );
  NAND2_X1 U8573 ( .A1(n6969), .A2(n7889), .ZN(n6961) );
  NAND2_X1 U8574 ( .A1(n8989), .A2(n4264), .ZN(n6960) );
  NAND2_X1 U8575 ( .A1(n6961), .A2(n6960), .ZN(n6962) );
  XNOR2_X1 U8576 ( .A(n6962), .B(n7872), .ZN(n7075) );
  AND2_X1 U8577 ( .A1(n5377), .A2(n8989), .ZN(n6963) );
  AOI21_X1 U8578 ( .B1(n6969), .B2(n7891), .A(n6963), .ZN(n7074) );
  XNOR2_X1 U8579 ( .A(n7075), .B(n7074), .ZN(n6964) );
  XNOR2_X1 U8580 ( .A(n7076), .B(n6964), .ZN(n6971) );
  NOR2_X1 U8581 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6612), .ZN(n9572) );
  NOR2_X1 U8582 ( .A1(n8666), .A2(n8689), .ZN(n6965) );
  AOI211_X1 U8583 ( .C1(n8668), .C2(n8990), .A(n9572), .B(n6965), .ZN(n6966)
         );
  OAI21_X1 U8584 ( .B1(n8671), .B2(n6967), .A(n6966), .ZN(n6968) );
  AOI21_X1 U8585 ( .B1(n8679), .B2(n6969), .A(n6968), .ZN(n6970) );
  OAI21_X1 U8586 ( .B1(n6971), .B2(n8664), .A(n6970), .ZN(P1_U3232) );
  NAND2_X1 U8587 ( .A1(n8501), .A2(n7024), .ZN(n7430) );
  NAND2_X1 U8588 ( .A1(n8065), .A2(n7408), .ZN(n6972) );
  NAND2_X1 U8589 ( .A1(n9854), .A2(n8064), .ZN(n7418) );
  INV_X1 U8590 ( .A(n9854), .ZN(n9804) );
  NAND2_X1 U8591 ( .A1(n6974), .A2(n9804), .ZN(n7415) );
  NAND2_X1 U8592 ( .A1(n7418), .A2(n7415), .ZN(n9797) );
  NAND2_X1 U8593 ( .A1(n9854), .A2(n6974), .ZN(n8127) );
  NAND2_X1 U8594 ( .A1(n8506), .A2(n6975), .ZN(n7421) );
  NAND2_X1 U8595 ( .A1(n7419), .A2(n7421), .ZN(n8126) );
  NAND2_X1 U8596 ( .A1(n6992), .A2(n8126), .ZN(n7013) );
  INV_X1 U8597 ( .A(n6975), .ZN(n9777) );
  NAND2_X1 U8598 ( .A1(n8506), .A2(n9777), .ZN(n7012) );
  NAND2_X1 U8599 ( .A1(n7013), .A2(n7012), .ZN(n9769) );
  OR2_X1 U8600 ( .A1(n9765), .A2(n6976), .ZN(n7427) );
  NAND2_X1 U8601 ( .A1(n9765), .A2(n6976), .ZN(n7425) );
  NAND2_X1 U8602 ( .A1(n7427), .A2(n7425), .ZN(n7016) );
  NAND2_X1 U8603 ( .A1(n9769), .A2(n7016), .ZN(n6977) );
  NAND2_X1 U8604 ( .A1(n9765), .A2(n8063), .ZN(n7008) );
  NAND2_X1 U8605 ( .A1(n6977), .A2(n7008), .ZN(n6978) );
  XOR2_X1 U8606 ( .A(n7520), .B(n6978), .Z(n8504) );
  INV_X1 U8607 ( .A(n8506), .ZN(n7002) );
  NAND2_X1 U8608 ( .A1(n9805), .A2(n7002), .ZN(n9764) );
  INV_X1 U8609 ( .A(n7030), .ZN(n6979) );
  AOI211_X1 U8610 ( .C1(n8501), .C2(n9766), .A(n9865), .B(n6979), .ZN(n8500)
         );
  INV_X1 U8611 ( .A(n8501), .ZN(n6982) );
  AOI22_X1 U8612 ( .A1(n9813), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n6980), .B2(
        n9802), .ZN(n6981) );
  OAI21_X1 U8613 ( .B1(n6982), .B2(n8398), .A(n6981), .ZN(n6990) );
  INV_X1 U8614 ( .A(n9797), .ZN(n7516) );
  INV_X1 U8615 ( .A(n8065), .ZN(n6983) );
  NAND2_X1 U8616 ( .A1(n6983), .A2(n7408), .ZN(n9791) );
  AND2_X1 U8617 ( .A1(n7516), .A2(n9791), .ZN(n6993) );
  INV_X1 U8618 ( .A(n8126), .ZN(n6996) );
  AND2_X1 U8619 ( .A1(n6993), .A2(n6996), .ZN(n6984) );
  AOI21_X2 U8620 ( .B1(n9792), .B2(n6984), .A(n4889), .ZN(n6994) );
  NAND2_X1 U8621 ( .A1(n6994), .A2(n7419), .ZN(n9774) );
  NAND2_X1 U8622 ( .A1(n9774), .A2(n9773), .ZN(n9772) );
  INV_X1 U8623 ( .A(n6986), .ZN(n6985) );
  AOI21_X1 U8624 ( .B1(n6985), .B2(n7009), .A(n9795), .ZN(n6988) );
  AOI21_X1 U8625 ( .B1(n6988), .B2(n7023), .A(n6987), .ZN(n8503) );
  NOR2_X1 U8626 ( .A1(n8503), .A2(n9813), .ZN(n6989) );
  AOI211_X1 U8627 ( .C1(n8500), .C2(n8344), .A(n6990), .B(n6989), .ZN(n6991)
         );
  OAI21_X1 U8628 ( .B1(n8504), .B2(n8412), .A(n6991), .ZN(P2_U3284) );
  OAI21_X1 U8629 ( .B1(n6992), .B2(n8126), .A(n7013), .ZN(n8510) );
  AOI22_X1 U8630 ( .A1(n8063), .A2(n9775), .B1(n8064), .B2(n9778), .ZN(n6998)
         );
  NAND2_X1 U8631 ( .A1(n9792), .A2(n6993), .ZN(n9793) );
  NAND2_X1 U8632 ( .A1(n9793), .A2(n7418), .ZN(n6995) );
  OAI211_X1 U8633 ( .C1(n6996), .C2(n6995), .A(n6994), .B(n9771), .ZN(n6997)
         );
  OAI211_X1 U8634 ( .C1(n8510), .C2(n9790), .A(n6998), .B(n6997), .ZN(n8505)
         );
  INV_X1 U8635 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7000) );
  OAI22_X1 U8636 ( .A1(n9783), .A2(n7000), .B1(n6999), .B2(n9788), .ZN(n7001)
         );
  AOI21_X1 U8637 ( .B1(n9803), .B2(n8506), .A(n7001), .ZN(n7005) );
  OR2_X1 U8638 ( .A1(n9805), .A2(n7002), .ZN(n7003) );
  AND2_X1 U8639 ( .A1(n9764), .A2(n7003), .ZN(n8507) );
  NAND2_X1 U8640 ( .A1(n8507), .A2(n9809), .ZN(n7004) );
  OAI211_X1 U8641 ( .C1(n8510), .C2(n7029), .A(n7005), .B(n7004), .ZN(n7006)
         );
  AOI21_X1 U8642 ( .B1(n8505), .B2(n9783), .A(n7006), .ZN(n7007) );
  INV_X1 U8643 ( .A(n7007), .ZN(P2_U3286) );
  OR2_X1 U8644 ( .A1(n8501), .A2(n9776), .ZN(n7015) );
  INV_X1 U8645 ( .A(n7015), .ZN(n7011) );
  AND2_X1 U8646 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  AND2_X1 U8647 ( .A1(n7012), .A2(n7014), .ZN(n8130) );
  NAND2_X1 U8648 ( .A1(n7013), .A2(n8130), .ZN(n7020) );
  INV_X1 U8649 ( .A(n7014), .ZN(n7018) );
  AND2_X1 U8650 ( .A1(n7016), .A2(n7015), .ZN(n7017) );
  AND2_X1 U8651 ( .A1(n7019), .A2(n7020), .ZN(n7022) );
  OR2_X1 U8652 ( .A1(n9493), .A2(n8403), .ZN(n7433) );
  NAND2_X1 U8653 ( .A1(n9493), .A2(n8403), .ZN(n7432) );
  NAND2_X1 U8654 ( .A1(n7433), .A2(n7432), .ZN(n7435) );
  NAND2_X1 U8655 ( .A1(n7020), .A2(n8125), .ZN(n7021) );
  OAI21_X1 U8656 ( .B1(n7022), .B2(n7435), .A(n7021), .ZN(n7028) );
  INV_X1 U8657 ( .A(n7435), .ZN(n7521) );
  OAI21_X1 U8658 ( .B1(n4331), .B2(n7521), .A(n7208), .ZN(n7026) );
  INV_X1 U8659 ( .A(n8384), .ZN(n7436) );
  OAI22_X1 U8660 ( .A1(n7436), .A2(n8404), .B1(n7024), .B2(n8402), .ZN(n7025)
         );
  AOI21_X1 U8661 ( .B1(n7026), .B2(n9771), .A(n7025), .ZN(n7027) );
  OAI21_X1 U8662 ( .B1(n7028), .B2(n9790), .A(n7027), .ZN(n9496) );
  INV_X1 U8663 ( .A(n9496), .ZN(n7037) );
  INV_X1 U8664 ( .A(n7028), .ZN(n9498) );
  INV_X1 U8665 ( .A(n7029), .ZN(n9810) );
  AND2_X1 U8666 ( .A1(n7030), .A2(n9493), .ZN(n7031) );
  OR2_X1 U8667 ( .A1(n7031), .A2(n8392), .ZN(n9495) );
  AOI22_X1 U8668 ( .A1(n9813), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7032), .B2(
        n9802), .ZN(n7034) );
  NAND2_X1 U8669 ( .A1(n9493), .A2(n9803), .ZN(n7033) );
  OAI211_X1 U8670 ( .C1(n9495), .C2(n8369), .A(n7034), .B(n7033), .ZN(n7035)
         );
  AOI21_X1 U8671 ( .B1(n9498), .B2(n9810), .A(n7035), .ZN(n7036) );
  OAI21_X1 U8672 ( .B1(n7037), .B2(n9813), .A(n7036), .ZN(P2_U3283) );
  OR2_X1 U8673 ( .A1(n8690), .A2(n8988), .ZN(n7039) );
  NAND2_X1 U8674 ( .A1(n7129), .A2(n8760), .ZN(n7041) );
  AOI22_X1 U8675 ( .A1(n7734), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7733), .B2(
        n9588), .ZN(n7040) );
  INV_X1 U8676 ( .A(n9342), .ZN(n8597) );
  OR2_X1 U8677 ( .A1(n9506), .A2(n8597), .ZN(n9336) );
  NAND2_X1 U8678 ( .A1(n9506), .A2(n8597), .ZN(n9337) );
  INV_X1 U8679 ( .A(n8955), .ZN(n8823) );
  XNOR2_X1 U8680 ( .A(n9081), .B(n8823), .ZN(n9510) );
  OR2_X1 U8681 ( .A1(n8690), .A2(n8689), .ZN(n8814) );
  XNOR2_X1 U8682 ( .A(n9339), .B(n8955), .ZN(n7050) );
  NAND2_X1 U8683 ( .A1(n8748), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7048) );
  INV_X1 U8684 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9354) );
  OR2_X1 U8685 ( .A1(n7783), .A2(n9354), .ZN(n7047) );
  OR2_X1 U8686 ( .A1(n7043), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7044) );
  NAND2_X1 U8687 ( .A1(n7701), .A2(n7044), .ZN(n9353) );
  OR2_X1 U8688 ( .A1(n7863), .A2(n9353), .ZN(n7046) );
  INV_X1 U8689 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9047) );
  OR2_X1 U8690 ( .A1(n8753), .A2(n9047), .ZN(n7045) );
  NAND4_X1 U8691 ( .A1(n7048), .A2(n7047), .A3(n7046), .A4(n7045), .ZN(n9328)
         );
  AOI22_X1 U8692 ( .A1(n9343), .A2(n8988), .B1(n9329), .B2(n9328), .ZN(n7049)
         );
  OAI21_X1 U8693 ( .B1(n7050), .B2(n9280), .A(n7049), .ZN(n7051) );
  AOI21_X1 U8694 ( .B1(n9510), .B2(n7052), .A(n7051), .ZN(n9512) );
  NAND2_X1 U8695 ( .A1(n7053), .A2(n9506), .ZN(n7054) );
  NAND2_X1 U8696 ( .A1(n9355), .A2(n7054), .ZN(n9508) );
  OAI22_X1 U8697 ( .A1(n6776), .A2(n7055), .B1(n8670), .B2(n9367), .ZN(n7056)
         );
  AOI21_X1 U8698 ( .B1(n9506), .B2(n9361), .A(n7056), .ZN(n7057) );
  OAI21_X1 U8699 ( .B1(n9508), .B2(n9313), .A(n7057), .ZN(n7058) );
  AOI21_X1 U8700 ( .B1(n9510), .B2(n9373), .A(n7058), .ZN(n7059) );
  OAI21_X1 U8701 ( .B1(n9512), .B2(n9364), .A(n7059), .ZN(P1_U3276) );
  INV_X1 U8702 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7838) );
  INV_X1 U8703 ( .A(n7060), .ZN(n7064) );
  INV_X1 U8704 ( .A(n7061), .ZN(n7062) );
  NAND2_X1 U8705 ( .A1(n7062), .A2(SI_24_), .ZN(n7063) );
  INV_X1 U8706 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7073) );
  MUX2_X1 U8707 ( .A(n7073), .B(n7838), .S(n7333), .Z(n7067) );
  INV_X1 U8708 ( .A(SI_25_), .ZN(n7066) );
  NAND2_X1 U8709 ( .A1(n7067), .A2(n7066), .ZN(n7116) );
  INV_X1 U8710 ( .A(n7067), .ZN(n7068) );
  NAND2_X1 U8711 ( .A1(n7068), .A2(SI_25_), .ZN(n7069) );
  NAND2_X1 U8712 ( .A1(n7116), .A2(n7069), .ZN(n7117) );
  INV_X1 U8713 ( .A(n7837), .ZN(n7072) );
  OAI222_X1 U8714 ( .A1(n9478), .A2(n7838), .B1(n7551), .B2(n7072), .C1(n7070), 
        .C2(n4258), .ZN(P1_U3328) );
  OAI222_X1 U8715 ( .A1(n8539), .A2(n7073), .B1(n7920), .B2(n7072), .C1(
        P2_U3152), .C2(n7071), .ZN(P2_U3333) );
  NAND2_X1 U8716 ( .A1(n8690), .A2(n7889), .ZN(n7078) );
  NAND2_X1 U8717 ( .A1(n8988), .A2(n4264), .ZN(n7077) );
  NAND2_X1 U8718 ( .A1(n7078), .A2(n7077), .ZN(n7079) );
  XNOR2_X1 U8719 ( .A(n7079), .B(n5361), .ZN(n7670) );
  NAND2_X1 U8720 ( .A1(n8690), .A2(n4264), .ZN(n7081) );
  NAND2_X1 U8721 ( .A1(n5377), .A2(n8988), .ZN(n7080) );
  NAND2_X1 U8722 ( .A1(n7081), .A2(n7080), .ZN(n7665) );
  INV_X1 U8723 ( .A(n7665), .ZN(n7671) );
  XNOR2_X1 U8724 ( .A(n7670), .B(n7671), .ZN(n7082) );
  XNOR2_X1 U8725 ( .A(n7676), .B(n7082), .ZN(n7089) );
  NOR2_X1 U8726 ( .A1(n8666), .A2(n8597), .ZN(n7083) );
  AOI211_X1 U8727 ( .C1(n8668), .C2(n8989), .A(n7084), .B(n7083), .ZN(n7085)
         );
  OAI21_X1 U8728 ( .B1(n8671), .B2(n7086), .A(n7085), .ZN(n7087) );
  AOI21_X1 U8729 ( .B1(n8690), .B2(n8679), .A(n7087), .ZN(n7088) );
  OAI21_X1 U8730 ( .B1(n7089), .B2(n8664), .A(n7088), .ZN(P1_U3213) );
  NAND2_X1 U8731 ( .A1(n7090), .A2(n7358), .ZN(n7093) );
  AOI22_X1 U8732 ( .A1(n7335), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5739), .B2(
        n7091), .ZN(n7092) );
  XNOR2_X1 U8733 ( .A(n8495), .B(n7612), .ZN(n7094) );
  NAND2_X1 U8734 ( .A1(n8384), .A2(n7602), .ZN(n7095) );
  NAND2_X1 U8735 ( .A1(n7094), .A2(n7095), .ZN(n7127) );
  INV_X1 U8736 ( .A(n7094), .ZN(n7097) );
  INV_X1 U8737 ( .A(n7095), .ZN(n7096) );
  NAND2_X1 U8738 ( .A1(n7097), .A2(n7096), .ZN(n7098) );
  NAND2_X1 U8739 ( .A1(n7127), .A2(n7098), .ZN(n7106) );
  INV_X1 U8740 ( .A(n7101), .ZN(n7103) );
  INV_X1 U8741 ( .A(n7128), .ZN(n7104) );
  AOI21_X1 U8742 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7115) );
  NAND2_X1 U8743 ( .A1(n6657), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7110) );
  XNOR2_X1 U8744 ( .A(n7134), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U8745 ( .A1(n7328), .A2(n8377), .ZN(n7109) );
  NAND2_X1 U8746 ( .A1(n4260), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U8747 ( .A1(n7322), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7107) );
  INV_X1 U8748 ( .A(n8403), .ZN(n8123) );
  AOI22_X1 U8749 ( .A1(n9724), .A2(n8123), .B1(n8396), .B2(n8054), .ZN(n7112)
         );
  OAI211_X1 U8750 ( .C1(n8046), .C2(n8405), .A(n7112), .B(n7111), .ZN(n7113)
         );
  AOI21_X1 U8751 ( .B1(n9748), .B2(n8495), .A(n7113), .ZN(n7114) );
  OAI21_X1 U8752 ( .B1(n7115), .B2(n9744), .A(n7114), .ZN(P2_U3217) );
  INV_X1 U8753 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7124) );
  INV_X1 U8754 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7857) );
  MUX2_X1 U8755 ( .A(n7124), .B(n7857), .S(n7333), .Z(n7120) );
  INV_X1 U8756 ( .A(SI_26_), .ZN(n7119) );
  NAND2_X1 U8757 ( .A1(n7120), .A2(n7119), .ZN(n7148) );
  INV_X1 U8758 ( .A(n7120), .ZN(n7121) );
  NAND2_X1 U8759 ( .A1(n7121), .A2(SI_26_), .ZN(n7122) );
  AND2_X1 U8760 ( .A1(n7148), .A2(n7122), .ZN(n7146) );
  INV_X1 U8761 ( .A(n7856), .ZN(n7125) );
  OAI222_X1 U8762 ( .A1(n7123), .A2(P1_U3084), .B1(n7551), .B2(n7125), .C1(
        n7857), .C2(n7154), .ZN(P1_U3327) );
  OAI222_X1 U8763 ( .A1(P2_U3152), .A2(n7126), .B1(n8543), .B2(n7125), .C1(
        n7124), .C2(n8533), .ZN(P2_U3332) );
  NOR2_X1 U8764 ( .A1(n8405), .A2(n5765), .ZN(n7566) );
  NAND2_X1 U8765 ( .A1(n7129), .A2(n7358), .ZN(n7131) );
  AOI22_X1 U8766 ( .A1(n7335), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5739), .B2(
        n7169), .ZN(n7130) );
  XNOR2_X1 U8767 ( .A(n8490), .B(n7612), .ZN(n7975) );
  XOR2_X1 U8768 ( .A(n7566), .B(n7975), .Z(n7132) );
  XNOR2_X1 U8769 ( .A(n7976), .B(n7132), .ZN(n7145) );
  NAND2_X1 U8770 ( .A1(n6657), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7139) );
  INV_X1 U8771 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7140) );
  INV_X1 U8772 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7133) );
  OAI21_X1 U8773 ( .B1(n7134), .B2(n7140), .A(n7133), .ZN(n7135) );
  AND2_X1 U8774 ( .A1(n7135), .A2(n7216), .ZN(n8366) );
  NAND2_X1 U8775 ( .A1(n7328), .A2(n8366), .ZN(n7138) );
  NAND2_X1 U8776 ( .A1(n4261), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8777 ( .A1(n7322), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7136) );
  OAI22_X1 U8778 ( .A1(n8046), .A2(n8061), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7140), .ZN(n7143) );
  INV_X1 U8779 ( .A(n8377), .ZN(n7141) );
  OAI22_X1 U8780 ( .A1(n8021), .A2(n7436), .B1(n9752), .B2(n7141), .ZN(n7142)
         );
  AOI211_X1 U8781 ( .C1(n8490), .C2(n9748), .A(n7143), .B(n7142), .ZN(n7144)
         );
  OAI21_X1 U8782 ( .B1(n7145), .B2(n9744), .A(n7144), .ZN(P2_U3243) );
  INV_X1 U8783 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7879) );
  INV_X1 U8784 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7156) );
  MUX2_X1 U8785 ( .A(n7156), .B(n7879), .S(n7333), .Z(n7151) );
  INV_X1 U8786 ( .A(SI_27_), .ZN(n7150) );
  NAND2_X1 U8787 ( .A1(n7151), .A2(n7150), .ZN(n7314) );
  INV_X1 U8788 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U8789 ( .A1(n7152), .A2(SI_27_), .ZN(n7153) );
  AND2_X1 U8790 ( .A1(n7314), .A2(n7153), .ZN(n7312) );
  INV_X1 U8791 ( .A(n7878), .ZN(n7155) );
  OAI222_X1 U8792 ( .A1(n7154), .A2(n7879), .B1(n7551), .B2(n7155), .C1(n9071), 
        .C2(P1_U3084), .ZN(P1_U3326) );
  OAI222_X1 U8793 ( .A1(n8539), .A2(n7156), .B1(n7920), .B2(n7155), .C1(n7543), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  OAI222_X1 U8794 ( .A1(n7158), .A2(n4258), .B1(n7551), .B2(n7157), .C1(n7816), 
        .C2(n9478), .ZN(P1_U3329) );
  OAI222_X1 U8795 ( .A1(n9478), .A2(n10055), .B1(n7551), .B2(n7159), .C1(n4258), .C2(n9256), .ZN(P1_U3334) );
  NAND2_X1 U8796 ( .A1(n7161), .A2(n7160), .ZN(n7163) );
  XNOR2_X1 U8797 ( .A(n8082), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8078) );
  NOR2_X1 U8798 ( .A1(n8079), .A2(n8078), .ZN(n8077) );
  NAND2_X1 U8799 ( .A1(n7213), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7164) );
  OAI21_X1 U8800 ( .B1(n7213), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7164), .ZN(
        n8092) );
  INV_X1 U8801 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U8802 ( .A1(n8103), .A2(n8102), .ZN(n8101) );
  NAND2_X1 U8803 ( .A1(n7165), .A2(n7180), .ZN(n7166) );
  NAND2_X1 U8804 ( .A1(n8101), .A2(n7166), .ZN(n7167) );
  XNOR2_X1 U8805 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n7167), .ZN(n7186) );
  INV_X1 U8806 ( .A(n7186), .ZN(n7184) );
  INV_X1 U8807 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7182) );
  INV_X1 U8808 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7179) );
  INV_X1 U8809 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7178) );
  NAND2_X1 U8810 ( .A1(n7169), .A2(n7168), .ZN(n7171) );
  NAND2_X1 U8811 ( .A1(n7171), .A2(n7170), .ZN(n8075) );
  INV_X1 U8812 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7172) );
  NAND2_X1 U8813 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  OAI21_X1 U8814 ( .B1(n7173), .B2(n7172), .A(n7174), .ZN(n8074) );
  NOR2_X1 U8815 ( .A1(n8075), .A2(n8074), .ZN(n8073) );
  INV_X1 U8816 ( .A(n7174), .ZN(n7175) );
  NOR2_X1 U8817 ( .A1(n8073), .A2(n7175), .ZN(n8086) );
  XNOR2_X1 U8818 ( .A(n7213), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8085) );
  INV_X1 U8819 ( .A(n8085), .ZN(n7176) );
  NAND2_X1 U8820 ( .A1(n8086), .A2(n7176), .ZN(n7177) );
  OAI21_X1 U8821 ( .B1(n7178), .B2(n8089), .A(n7177), .ZN(n8100) );
  AOI22_X1 U8822 ( .A1(n8108), .A2(n7179), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n7180), .ZN(n8099) );
  NOR2_X1 U8823 ( .A1(n8100), .A2(n8099), .ZN(n8098) );
  AOI21_X1 U8824 ( .B1(n7180), .B2(n7179), .A(n8098), .ZN(n7181) );
  XNOR2_X1 U8825 ( .A(n7182), .B(n7181), .ZN(n7185) );
  OAI21_X1 U8826 ( .B1(n7185), .B2(n9759), .A(n9757), .ZN(n7183) );
  AOI21_X1 U8827 ( .B1(n7184), .B2(n4352), .A(n7183), .ZN(n7188) );
  AOI22_X1 U8828 ( .A1(n7186), .A2(n4352), .B1(n9753), .B2(n7185), .ZN(n7187)
         );
  MUX2_X1 U8829 ( .A(n7188), .B(n7187), .S(n8198), .Z(n7189) );
  NAND2_X1 U8830 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7941) );
  OAI211_X1 U8831 ( .C1(n8106), .C2(n7190), .A(n7189), .B(n7941), .ZN(P2_U3264) );
  OAI21_X1 U8832 ( .B1(n5588), .B2(n7192), .A(n7191), .ZN(n9654) );
  INV_X1 U8833 ( .A(n9373), .ZN(n7207) );
  OAI21_X1 U8834 ( .B1(n8940), .B2(n7194), .A(n7193), .ZN(n7198) );
  OAI22_X1 U8835 ( .A1(n7196), .A2(n9282), .B1(n7195), .B2(n9345), .ZN(n7197)
         );
  AOI21_X1 U8836 ( .B1(n7198), .B2(n9348), .A(n7197), .ZN(n7199) );
  OAI21_X1 U8837 ( .B1(n9385), .B2(n9654), .A(n7199), .ZN(n9656) );
  OAI211_X1 U8838 ( .C1(n4598), .C2(n7201), .A(n9673), .B(n7200), .ZN(n9651)
         );
  OAI22_X1 U8839 ( .A1(n9651), .A2(n5586), .B1(n9367), .B2(n7202), .ZN(n7203)
         );
  OAI21_X1 U8840 ( .B1(n9656), .B2(n7203), .A(n6776), .ZN(n7206) );
  AOI22_X1 U8841 ( .A1(n9361), .A2(n7204), .B1(n9364), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7205) );
  OAI211_X1 U8842 ( .C1(n9654), .C2(n7207), .A(n7206), .B(n7205), .ZN(P1_U3290) );
  XNOR2_X1 U8843 ( .A(n8495), .B(n8384), .ZN(n8132) );
  OR2_X2 U8844 ( .A1(n8401), .A2(n8400), .ZN(n8407) );
  OR2_X1 U8845 ( .A1(n8495), .A2(n7436), .ZN(n8380) );
  OR2_X1 U8846 ( .A1(n8490), .A2(n8405), .ZN(n7439) );
  AND2_X1 U8847 ( .A1(n8380), .A2(n7439), .ZN(n7209) );
  NAND2_X1 U8848 ( .A1(n8407), .A2(n7209), .ZN(n8355) );
  NAND2_X1 U8849 ( .A1(n7683), .A2(n7358), .ZN(n7211) );
  AOI22_X1 U8850 ( .A1(n7335), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5739), .B2(
        n8082), .ZN(n7210) );
  NAND2_X1 U8851 ( .A1(n8483), .A2(n8061), .ZN(n7442) );
  NAND2_X1 U8852 ( .A1(n8490), .A2(n8405), .ZN(n8354) );
  AND2_X1 U8853 ( .A1(n7442), .A2(n8354), .ZN(n7212) );
  NAND2_X1 U8854 ( .A1(n8355), .A2(n7212), .ZN(n8336) );
  NAND2_X1 U8855 ( .A1(n7696), .A2(n7358), .ZN(n7215) );
  AOI22_X1 U8856 ( .A1(n7335), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5739), .B2(
        n7213), .ZN(n7214) );
  NAND2_X1 U8857 ( .A1(n5451), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U8858 ( .A1(n4260), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7220) );
  INV_X1 U8859 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U8860 ( .A1(n7216), .A2(n9989), .ZN(n7217) );
  AND2_X1 U8861 ( .A1(n7233), .A2(n7217), .ZN(n8345) );
  NAND2_X1 U8862 ( .A1(n7328), .A2(n8345), .ZN(n7219) );
  NAND2_X1 U8863 ( .A1(n6657), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U8864 ( .A1(n8480), .A2(n8358), .ZN(n7446) );
  NAND2_X1 U8865 ( .A1(n7222), .A2(n7446), .ZN(n8335) );
  INV_X1 U8866 ( .A(n7222), .ZN(n7448) );
  NAND2_X1 U8867 ( .A1(n7715), .A2(n7358), .ZN(n7224) );
  AOI22_X1 U8868 ( .A1(n7335), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5739), .B2(
        n8108), .ZN(n7223) );
  XNOR2_X1 U8869 ( .A(n7233), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U8870 ( .A1(n7328), .A2(n8321), .ZN(n7228) );
  NAND2_X1 U8871 ( .A1(n4260), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8872 ( .A1(n6657), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7226) );
  NAND2_X1 U8873 ( .A1(n7322), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7225) );
  NAND4_X1 U8874 ( .A1(n7228), .A2(n7227), .A3(n7226), .A4(n7225), .ZN(n8338)
         );
  INV_X1 U8875 ( .A(n8338), .ZN(n8307) );
  NAND2_X1 U8876 ( .A1(n8473), .A2(n8307), .ZN(n7452) );
  NAND2_X1 U8877 ( .A1(n7457), .A2(n7452), .ZN(n7503) );
  NAND2_X1 U8878 ( .A1(n7732), .A2(n7358), .ZN(n7230) );
  AOI22_X1 U8879 ( .A1(n7335), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5739), .B2(
        n4643), .ZN(n7229) );
  INV_X1 U8880 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7232) );
  INV_X1 U8881 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7231) );
  OAI21_X1 U8882 ( .B1(n7233), .B2(n7232), .A(n7231), .ZN(n7234) );
  AND2_X1 U8883 ( .A1(n7234), .A2(n7241), .ZN(n8311) );
  NAND2_X1 U8884 ( .A1(n7328), .A2(n8311), .ZN(n7238) );
  NAND2_X1 U8885 ( .A1(n4260), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U8886 ( .A1(n6657), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U8887 ( .A1(n5451), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7235) );
  OR2_X1 U8888 ( .A1(n8470), .A2(n8135), .ZN(n7459) );
  NAND2_X1 U8889 ( .A1(n8470), .A2(n8135), .ZN(n7454) );
  NAND2_X1 U8890 ( .A1(n7459), .A2(n7454), .ZN(n8305) );
  INV_X1 U8891 ( .A(n7454), .ZN(n8294) );
  NAND2_X1 U8892 ( .A1(n7754), .A2(n7358), .ZN(n7240) );
  NAND2_X1 U8893 ( .A1(n7335), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8894 ( .A1(n6657), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7246) );
  INV_X1 U8895 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10010) );
  NAND2_X1 U8896 ( .A1(n7241), .A2(n10010), .ZN(n7242) );
  AND2_X1 U8897 ( .A1(n7256), .A2(n7242), .ZN(n8291) );
  NAND2_X1 U8898 ( .A1(n7328), .A2(n8291), .ZN(n7245) );
  NAND2_X1 U8899 ( .A1(n4261), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7244) );
  NAND2_X1 U8900 ( .A1(n7322), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7243) );
  NAND2_X1 U8901 ( .A1(n8463), .A2(n8308), .ZN(n7461) );
  NAND2_X1 U8902 ( .A1(n7460), .A2(n7461), .ZN(n8295) );
  NAND2_X1 U8903 ( .A1(n7775), .A2(n7358), .ZN(n7248) );
  NAND2_X1 U8904 ( .A1(n7335), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7247) );
  NAND2_X1 U8905 ( .A1(n4261), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7252) );
  XNOR2_X1 U8906 ( .A(n7256), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U8907 ( .A1(n7328), .A2(n8277), .ZN(n7251) );
  NAND2_X1 U8908 ( .A1(n5451), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7250) );
  NAND2_X1 U8909 ( .A1(n6657), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7249) );
  OR2_X1 U8910 ( .A1(n8458), .A2(n8267), .ZN(n7464) );
  NAND2_X1 U8911 ( .A1(n8458), .A2(n8267), .ZN(n8264) );
  NAND2_X2 U8912 ( .A1(n4282), .A2(n8281), .ZN(n8280) );
  NAND2_X1 U8913 ( .A1(n7793), .A2(n7358), .ZN(n7254) );
  NAND2_X1 U8914 ( .A1(n7335), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7253) );
  INV_X1 U8915 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7960) );
  INV_X1 U8916 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7255) );
  OAI21_X1 U8917 ( .B1(n7256), .B2(n7960), .A(n7255), .ZN(n7257) );
  AND2_X1 U8918 ( .A1(n7257), .A2(n7264), .ZN(n8259) );
  NAND2_X1 U8919 ( .A1(n8259), .A2(n7328), .ZN(n7261) );
  NAND2_X1 U8920 ( .A1(n6657), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U8921 ( .A1(n7322), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7259) );
  NAND2_X1 U8922 ( .A1(n4261), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7258) );
  AND4_X1 U8923 ( .A1(n7261), .A2(n7260), .A3(n7259), .A4(n7258), .ZN(n8060)
         );
  NAND2_X1 U8924 ( .A1(n8453), .A2(n8060), .ZN(n7465) );
  NAND2_X1 U8925 ( .A1(n8244), .A2(n7465), .ZN(n8254) );
  INV_X1 U8926 ( .A(n8254), .ZN(n8263) );
  NAND2_X1 U8927 ( .A1(n7653), .A2(n7358), .ZN(n7263) );
  NAND2_X1 U8928 ( .A1(n7335), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7262) );
  INV_X1 U8929 ( .A(n7328), .ZN(n7305) );
  INV_X1 U8930 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U8931 ( .A1(n7264), .A2(n7934), .ZN(n7265) );
  NAND2_X1 U8932 ( .A1(n7273), .A2(n7265), .ZN(n8240) );
  OR2_X1 U8933 ( .A1(n7305), .A2(n8240), .ZN(n7270) );
  NAND2_X1 U8934 ( .A1(n4261), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7267) );
  NAND2_X1 U8935 ( .A1(n5451), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7266) );
  AND2_X1 U8936 ( .A1(n7267), .A2(n7266), .ZN(n7269) );
  NAND2_X1 U8937 ( .A1(n6657), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7268) );
  OR2_X1 U8938 ( .A1(n8448), .A2(n8268), .ZN(n7369) );
  NAND2_X1 U8939 ( .A1(n8448), .A2(n8268), .ZN(n8229) );
  NAND2_X1 U8940 ( .A1(n7815), .A2(n7358), .ZN(n7272) );
  NAND2_X1 U8941 ( .A1(n7335), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U8942 ( .A1(n7273), .A2(n8011), .ZN(n7274) );
  NAND2_X1 U8943 ( .A1(n7281), .A2(n7274), .ZN(n8223) );
  OR2_X1 U8944 ( .A1(n8223), .A2(n7305), .ZN(n7278) );
  AOI22_X1 U8945 ( .A1(n4260), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n7322), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U8946 ( .A1(n6657), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7276) );
  NAND2_X1 U8947 ( .A1(n8443), .A2(n8210), .ZN(n7470) );
  NAND2_X1 U8948 ( .A1(n7837), .A2(n7358), .ZN(n7280) );
  NAND2_X1 U8949 ( .A1(n7335), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U8950 ( .A1(n7281), .A2(n10013), .ZN(n7282) );
  AND2_X1 U8951 ( .A1(n7292), .A2(n7282), .ZN(n8213) );
  NAND2_X1 U8952 ( .A1(n8213), .A2(n7328), .ZN(n7288) );
  INV_X1 U8953 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n7285) );
  NAND2_X1 U8954 ( .A1(n6657), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7284) );
  NAND2_X1 U8955 ( .A1(n7322), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7283) );
  OAI211_X1 U8956 ( .C1(n7285), .C2(n7325), .A(n7284), .B(n7283), .ZN(n7286)
         );
  INV_X1 U8957 ( .A(n7286), .ZN(n7287) );
  XNOR2_X1 U8958 ( .A(n8440), .B(n8232), .ZN(n8204) );
  INV_X1 U8959 ( .A(n8204), .ZN(n8207) );
  INV_X1 U8960 ( .A(n8232), .ZN(n8192) );
  NAND2_X1 U8961 ( .A1(n7856), .A2(n7358), .ZN(n7290) );
  NAND2_X1 U8962 ( .A1(n7335), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7289) );
  INV_X1 U8963 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7291) );
  NAND2_X1 U8964 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  NAND2_X1 U8965 ( .A1(n7303), .A2(n7293), .ZN(n8053) );
  OR2_X1 U8966 ( .A1(n8053), .A2(n7305), .ZN(n7299) );
  INV_X1 U8967 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7296) );
  NAND2_X1 U8968 ( .A1(n6657), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7295) );
  NAND2_X1 U8969 ( .A1(n7322), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7294) );
  OAI211_X1 U8970 ( .C1(n7296), .C2(n7325), .A(n7295), .B(n7294), .ZN(n7297)
         );
  INV_X1 U8971 ( .A(n7297), .ZN(n7298) );
  NAND2_X1 U8972 ( .A1(n7299), .A2(n7298), .ZN(n8179) );
  NAND2_X1 U8973 ( .A1(n8188), .A2(n8179), .ZN(n7480) );
  INV_X1 U8974 ( .A(n8179), .ZN(n8211) );
  INV_X1 U8975 ( .A(n8185), .ZN(n8191) );
  NAND2_X1 U8976 ( .A1(n7878), .A2(n7358), .ZN(n7301) );
  NAND2_X1 U8977 ( .A1(n7335), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7300) );
  INV_X1 U8978 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U8979 ( .A1(n7303), .A2(n7302), .ZN(n7304) );
  NAND2_X1 U8980 ( .A1(n7319), .A2(n7304), .ZN(n7928) );
  OR2_X1 U8981 ( .A1(n7928), .A2(n7305), .ZN(n7311) );
  INV_X1 U8982 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7308) );
  NAND2_X1 U8983 ( .A1(n7322), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7307) );
  NAND2_X1 U8984 ( .A1(n6657), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7306) );
  OAI211_X1 U8985 ( .C1(n7308), .C2(n7325), .A(n7307), .B(n7306), .ZN(n7309)
         );
  INV_X1 U8986 ( .A(n7309), .ZN(n7310) );
  INV_X1 U8987 ( .A(n7625), .ZN(n8193) );
  NAND2_X1 U8988 ( .A1(n8175), .A2(n8193), .ZN(n7481) );
  INV_X1 U8989 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7630) );
  INV_X1 U8990 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7923) );
  MUX2_X1 U8991 ( .A(n7630), .B(n7923), .S(n7333), .Z(n7332) );
  XNOR2_X1 U8992 ( .A(n7332), .B(SI_28_), .ZN(n7329) );
  NAND2_X1 U8993 ( .A1(n7631), .A2(n7358), .ZN(n7317) );
  NAND2_X1 U8994 ( .A1(n7335), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7316) );
  NAND2_X1 U8995 ( .A1(n7319), .A2(n7318), .ZN(n7320) );
  INV_X1 U8996 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7326) );
  NAND2_X1 U8997 ( .A1(n6657), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U8998 ( .A1(n7322), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7323) );
  OAI211_X1 U8999 ( .C1(n7326), .C2(n7325), .A(n7324), .B(n7323), .ZN(n7327)
         );
  AOI21_X1 U9000 ( .B1(n8158), .B2(n7328), .A(n7327), .ZN(n8145) );
  NAND2_X1 U9001 ( .A1(n8424), .A2(n8145), .ZN(n7486) );
  INV_X1 U9002 ( .A(SI_28_), .ZN(n7331) );
  INV_X1 U9003 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8540) );
  INV_X1 U9004 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8682) );
  MUX2_X1 U9005 ( .A(n8540), .B(n8682), .S(n7333), .Z(n7340) );
  XNOR2_X1 U9006 ( .A(n7340), .B(SI_29_), .ZN(n7334) );
  NAND2_X1 U9007 ( .A1(n8681), .A2(n7358), .ZN(n7337) );
  NAND2_X1 U9008 ( .A1(n7335), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7336) );
  NAND2_X1 U9009 ( .A1(n8421), .A2(n7623), .ZN(n7368) );
  INV_X1 U9010 ( .A(SI_29_), .ZN(n7339) );
  AND2_X1 U9011 ( .A1(n7340), .A2(n7339), .ZN(n7343) );
  INV_X1 U9012 ( .A(n7340), .ZN(n7341) );
  NAND2_X1 U9013 ( .A1(n7341), .A2(SI_29_), .ZN(n7342) );
  MUX2_X1 U9014 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7355), .Z(n7351) );
  NAND2_X1 U9015 ( .A1(n8744), .A2(n7358), .ZN(n7346) );
  INV_X1 U9016 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7921) );
  OR2_X1 U9017 ( .A1(n7359), .A2(n7921), .ZN(n7345) );
  OAI211_X1 U9018 ( .C1(n7348), .C2(n8416), .A(n8116), .B(n7367), .ZN(n7347)
         );
  INV_X1 U9019 ( .A(n7347), .ZN(n7364) );
  INV_X1 U9020 ( .A(n7348), .ZN(n7361) );
  INV_X1 U9021 ( .A(SI_30_), .ZN(n7349) );
  NAND2_X1 U9022 ( .A1(n7352), .A2(n7351), .ZN(n7353) );
  MUX2_X1 U9023 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7355), .Z(n7356) );
  XNOR2_X1 U9024 ( .A(n7356), .B(SI_31_), .ZN(n7357) );
  OR2_X1 U9025 ( .A1(n7359), .A2(n5137), .ZN(n7360) );
  NAND2_X1 U9026 ( .A1(n8416), .A2(n8143), .ZN(n7490) );
  NAND2_X1 U9027 ( .A1(n7362), .A2(n8116), .ZN(n7498) );
  AND2_X1 U9028 ( .A1(n8228), .A2(n7369), .ZN(n7468) );
  NAND2_X1 U9029 ( .A1(n7371), .A2(n7370), .ZN(n7377) );
  OAI21_X1 U9030 ( .B1(n7539), .B2(n7377), .A(n7372), .ZN(n7374) );
  INV_X1 U9031 ( .A(n7376), .ZN(n7373) );
  AOI21_X1 U9032 ( .B1(n7374), .B2(n7378), .A(n7373), .ZN(n7381) );
  NAND3_X1 U9033 ( .A1(n7377), .A2(n7376), .A3(n7375), .ZN(n7379) );
  AND2_X1 U9034 ( .A1(n7379), .A2(n7378), .ZN(n7380) );
  MUX2_X1 U9035 ( .A(n7381), .B(n7380), .S(n4262), .Z(n7386) );
  INV_X1 U9036 ( .A(n7396), .ZN(n7384) );
  NAND2_X1 U9037 ( .A1(n7382), .A2(n7387), .ZN(n7383) );
  MUX2_X1 U9038 ( .A(n7384), .B(n7383), .S(n4262), .Z(n7398) );
  NOR3_X1 U9039 ( .A1(n7386), .A2(n7385), .A3(n7398), .ZN(n7394) );
  INV_X1 U9040 ( .A(n7387), .ZN(n7390) );
  INV_X1 U9041 ( .A(n7398), .ZN(n7388) );
  OAI21_X1 U9042 ( .B1(n7390), .B2(n7389), .A(n7388), .ZN(n7392) );
  AOI21_X1 U9043 ( .B1(n7392), .B2(n7391), .A(n4262), .ZN(n7393) );
  OAI21_X1 U9044 ( .B1(n7394), .B2(n7393), .A(n7399), .ZN(n7404) );
  AOI22_X1 U9045 ( .A1(n7398), .A2(n7397), .B1(n7396), .B2(n7395), .ZN(n7400)
         );
  OAI21_X1 U9046 ( .B1(n7400), .B2(n4676), .A(n4262), .ZN(n7403) );
  NOR3_X1 U9047 ( .A1(n8067), .A2(n7401), .A3(n7477), .ZN(n7402) );
  AOI211_X1 U9048 ( .C1(n7404), .C2(n7403), .A(n7402), .B(n7512), .ZN(n7413)
         );
  MUX2_X1 U9049 ( .A(n7406), .B(n7405), .S(n4262), .Z(n7407) );
  NAND2_X1 U9050 ( .A1(n7407), .A2(n7514), .ZN(n7412) );
  NAND2_X1 U9051 ( .A1(n7408), .A2(n4262), .ZN(n7410) );
  NAND2_X1 U9052 ( .A1(n9735), .A2(n7477), .ZN(n7409) );
  MUX2_X1 U9053 ( .A(n7410), .B(n7409), .S(n8065), .Z(n7411) );
  OAI211_X1 U9054 ( .C1(n7413), .C2(n7412), .A(n7415), .B(n7411), .ZN(n7420)
         );
  INV_X1 U9055 ( .A(n7418), .ZN(n7414) );
  AOI21_X1 U9056 ( .B1(n7420), .B2(n7415), .A(n7414), .ZN(n7417) );
  INV_X1 U9057 ( .A(n7421), .ZN(n7416) );
  OAI211_X1 U9058 ( .C1(n7417), .C2(n7416), .A(n7427), .B(n7419), .ZN(n7424)
         );
  NAND3_X1 U9059 ( .A1(n7420), .A2(n7419), .A3(n7418), .ZN(n7422) );
  NAND3_X1 U9060 ( .A1(n7422), .A2(n7425), .A3(n7421), .ZN(n7423) );
  MUX2_X1 U9061 ( .A(n7424), .B(n7423), .S(n4262), .Z(n7429) );
  NAND3_X1 U9062 ( .A1(n7429), .A2(n7430), .A3(n7425), .ZN(n7426) );
  NAND3_X1 U9063 ( .A1(n7429), .A2(n7428), .A3(n7427), .ZN(n7431) );
  MUX2_X1 U9064 ( .A(n7433), .B(n7432), .S(n4262), .Z(n7434) );
  NAND2_X1 U9065 ( .A1(n7439), .A2(n8354), .ZN(n8373) );
  INV_X1 U9066 ( .A(n8373), .ZN(n8382) );
  NAND2_X1 U9067 ( .A1(n8495), .A2(n7436), .ZN(n7437) );
  MUX2_X1 U9068 ( .A(n7437), .B(n8380), .S(n4262), .Z(n7438) );
  MUX2_X1 U9069 ( .A(n7439), .B(n8354), .S(n4262), .Z(n7440) );
  NAND3_X1 U9070 ( .A1(n7441), .A2(n8356), .A3(n7440), .ZN(n7451) );
  INV_X1 U9071 ( .A(n7442), .ZN(n7444) );
  INV_X1 U9072 ( .A(n8334), .ZN(n7443) );
  MUX2_X1 U9073 ( .A(n7444), .B(n7443), .S(n4262), .Z(n7445) );
  NOR2_X1 U9074 ( .A1(n7445), .A2(n8335), .ZN(n7450) );
  NAND2_X1 U9075 ( .A1(n7452), .A2(n7446), .ZN(n7447) );
  MUX2_X1 U9076 ( .A(n7448), .B(n7447), .S(n4262), .Z(n7449) );
  AOI21_X1 U9077 ( .B1(n7451), .B2(n7450), .A(n7449), .ZN(n7456) );
  INV_X1 U9078 ( .A(n7452), .ZN(n7453) );
  OAI211_X1 U9079 ( .C1(n7456), .C2(n7453), .A(n7459), .B(n7457), .ZN(n7455)
         );
  INV_X1 U9080 ( .A(n7456), .ZN(n7458) );
  AOI21_X1 U9081 ( .B1(n7458), .B2(n7457), .A(n8294), .ZN(n7463) );
  NAND2_X1 U9082 ( .A1(n7460), .A2(n7459), .ZN(n7462) );
  MUX2_X1 U9083 ( .A(n8244), .B(n7465), .S(n4262), .Z(n7466) );
  OAI21_X1 U9084 ( .B1(n7468), .B2(n7477), .A(n7467), .ZN(n7471) );
  AOI21_X1 U9085 ( .B1(n7470), .B2(n8229), .A(n4262), .ZN(n7469) );
  AOI21_X1 U9086 ( .B1(n7471), .B2(n7470), .A(n7469), .ZN(n7475) );
  OAI21_X1 U9087 ( .B1(n4262), .B2(n7472), .A(n8207), .ZN(n7474) );
  NAND3_X1 U9088 ( .A1(n8216), .A2(n4262), .A3(n8192), .ZN(n7473) );
  OAI211_X1 U9089 ( .C1(n7475), .C2(n7474), .A(n7480), .B(n7473), .ZN(n7479)
         );
  OAI21_X1 U9090 ( .B1(n8216), .B2(n8192), .A(n7478), .ZN(n7476) );
  AOI22_X1 U9091 ( .A1(n7479), .A2(n7478), .B1(n7477), .B2(n7476), .ZN(n7485)
         );
  INV_X1 U9092 ( .A(n8176), .ZN(n7527) );
  OAI21_X1 U9093 ( .B1(n4262), .B2(n7480), .A(n7527), .ZN(n7484) );
  NAND2_X1 U9094 ( .A1(n8428), .A2(n7625), .ZN(n7482) );
  MUX2_X1 U9095 ( .A(n7482), .B(n7481), .S(n4262), .Z(n7483) );
  OAI211_X1 U9096 ( .C1(n7485), .C2(n7484), .A(n7529), .B(n7483), .ZN(n7489)
         );
  MUX2_X1 U9097 ( .A(n7487), .B(n7486), .S(n4262), .Z(n7488) );
  NAND3_X1 U9098 ( .A1(n7489), .A2(n8140), .A3(n7488), .ZN(n7491) );
  NAND2_X1 U9099 ( .A1(n7491), .A2(n7490), .ZN(n7493) );
  INV_X1 U9100 ( .A(n7533), .ZN(n7492) );
  OAI22_X1 U9101 ( .A1(n7493), .A2(n7531), .B1(n7492), .B2(n7477), .ZN(n7494)
         );
  INV_X1 U9102 ( .A(n7531), .ZN(n7495) );
  AOI21_X1 U9103 ( .B1(n7498), .B2(n7495), .A(n4262), .ZN(n7496) );
  INV_X1 U9104 ( .A(n7497), .ZN(n7499) );
  INV_X1 U9105 ( .A(n7498), .ZN(n7532) );
  MUX2_X1 U9106 ( .A(n7499), .B(n7532), .S(n4262), .Z(n7500) );
  INV_X1 U9107 ( .A(n7537), .ZN(n7542) );
  OAI21_X1 U9108 ( .B1(n7535), .B2(n7536), .A(n9865), .ZN(n7541) );
  INV_X1 U9109 ( .A(n8228), .ZN(n8219) );
  INV_X1 U9110 ( .A(n7503), .ZN(n8325) );
  NOR2_X1 U9111 ( .A1(n7505), .A2(n7504), .ZN(n7510) );
  NAND4_X1 U9112 ( .A1(n7510), .A2(n7509), .A3(n7508), .A4(n7507), .ZN(n7513)
         );
  NOR3_X1 U9113 ( .A1(n7513), .A2(n7512), .A3(n7511), .ZN(n7517) );
  NAND4_X1 U9114 ( .A1(n7517), .A2(n7516), .A3(n7515), .A4(n7514), .ZN(n7518)
         );
  NOR2_X1 U9115 ( .A1(n7518), .A2(n8126), .ZN(n7519) );
  NAND4_X1 U9116 ( .A1(n7521), .A2(n7520), .A3(n9773), .A4(n7519), .ZN(n7522)
         );
  NOR3_X1 U9117 ( .A1(n8373), .A2(n8400), .A3(n7522), .ZN(n7523) );
  NAND4_X1 U9118 ( .A1(n8325), .A2(n4836), .A3(n8356), .A4(n7523), .ZN(n7524)
         );
  NOR3_X1 U9119 ( .A1(n8295), .A2(n8305), .A3(n7524), .ZN(n7525) );
  NAND4_X1 U9120 ( .A1(n8246), .A2(n8263), .A3(n8281), .A4(n7525), .ZN(n7526)
         );
  NOR4_X1 U9121 ( .A1(n8185), .A2(n8204), .A3(n8219), .A4(n7526), .ZN(n7528)
         );
  NAND4_X1 U9122 ( .A1(n8140), .A2(n7529), .A3(n7528), .A4(n7527), .ZN(n7530)
         );
  NOR4_X1 U9123 ( .A1(n7533), .A2(n7532), .A3(n7531), .A4(n7530), .ZN(n7534)
         );
  XNOR2_X1 U9124 ( .A(n7534), .B(n8198), .ZN(n7540) );
  AOI21_X1 U9125 ( .B1(n7537), .B2(n7536), .A(n7535), .ZN(n7538) );
  INV_X1 U9126 ( .A(n7543), .ZN(n8114) );
  NAND4_X1 U9127 ( .A1(n7545), .A2(n8114), .A3(n7544), .A4(n9778), .ZN(n7546)
         );
  OAI211_X1 U9128 ( .C1(n7547), .C2(n7549), .A(n7546), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7548) );
  INV_X1 U9129 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8745) );
  INV_X1 U9130 ( .A(n8744), .ZN(n7919) );
  OAI222_X1 U9131 ( .A1(n9478), .A2(n8745), .B1(n7551), .B2(n7919), .C1(
        P1_U3084), .C2(n7550), .ZN(P1_U3323) );
  OR2_X1 U9132 ( .A1(n7553), .A2(n7552), .ZN(n8038) );
  AOI22_X1 U9133 ( .A1(n9748), .A2(n7554), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8038), .ZN(n7559) );
  OAI21_X1 U9134 ( .B1(n7555), .B2(n5765), .A(n9823), .ZN(n7556) );
  NAND3_X1 U9135 ( .A1(n9730), .A2(n7557), .A3(n7556), .ZN(n7558) );
  OAI211_X1 U9136 ( .C1(n8046), .C2(n7560), .A(n7559), .B(n7558), .ZN(P2_U3234) );
  INV_X1 U9137 ( .A(n8158), .ZN(n7628) );
  XNOR2_X1 U9138 ( .A(n8216), .B(n7607), .ZN(n7601) );
  INV_X1 U9139 ( .A(n7601), .ZN(n7967) );
  INV_X1 U9140 ( .A(n8008), .ZN(n7600) );
  NOR2_X1 U9141 ( .A1(n8210), .A2(n5765), .ZN(n8007) );
  INV_X1 U9142 ( .A(n8007), .ZN(n7599) );
  XNOR2_X1 U9143 ( .A(n8483), .B(n7612), .ZN(n7561) );
  OR2_X1 U9144 ( .A1(n8061), .A2(n5765), .ZN(n7562) );
  NAND2_X1 U9145 ( .A1(n7561), .A2(n7562), .ZN(n7567) );
  INV_X1 U9146 ( .A(n7561), .ZN(n7564) );
  INV_X1 U9147 ( .A(n7562), .ZN(n7563) );
  NAND2_X1 U9148 ( .A1(n7564), .A2(n7563), .ZN(n7565) );
  NAND2_X1 U9149 ( .A1(n7567), .A2(n7565), .ZN(n7982) );
  XNOR2_X1 U9150 ( .A(n8480), .B(n7607), .ZN(n7568) );
  NOR2_X1 U9151 ( .A1(n8358), .A2(n5765), .ZN(n7569) );
  XNOR2_X1 U9152 ( .A(n7568), .B(n7569), .ZN(n7998) );
  INV_X1 U9153 ( .A(n7568), .ZN(n7571) );
  INV_X1 U9154 ( .A(n7569), .ZN(n7570) );
  XNOR2_X1 U9155 ( .A(n8473), .B(n7607), .ZN(n7574) );
  NAND2_X1 U9156 ( .A1(n8338), .A2(n7602), .ZN(n7572) );
  XNOR2_X1 U9157 ( .A(n7574), .B(n7572), .ZN(n8043) );
  INV_X1 U9158 ( .A(n7572), .ZN(n7573) );
  NAND2_X1 U9159 ( .A1(n7574), .A2(n7573), .ZN(n7575) );
  XNOR2_X1 U9160 ( .A(n8470), .B(n7612), .ZN(n7576) );
  OR2_X1 U9161 ( .A1(n8135), .A2(n5765), .ZN(n7577) );
  NAND2_X1 U9162 ( .A1(n7576), .A2(n7577), .ZN(n8016) );
  INV_X1 U9163 ( .A(n7576), .ZN(n7579) );
  INV_X1 U9164 ( .A(n7577), .ZN(n7578) );
  NAND2_X1 U9165 ( .A1(n7579), .A2(n7578), .ZN(n7580) );
  NAND2_X1 U9166 ( .A1(n8016), .A2(n7580), .ZN(n7940) );
  XNOR2_X1 U9167 ( .A(n8463), .B(n7607), .ZN(n7586) );
  NOR2_X1 U9168 ( .A1(n8308), .A2(n5765), .ZN(n7585) );
  AND2_X1 U9169 ( .A1(n7586), .A2(n7585), .ZN(n7587) );
  OR2_X1 U9170 ( .A1(n7940), .A2(n7587), .ZN(n7954) );
  XNOR2_X1 U9171 ( .A(n8279), .B(n7607), .ZN(n7584) );
  INV_X1 U9172 ( .A(n7584), .ZN(n7581) );
  NOR2_X1 U9173 ( .A1(n8267), .A2(n5765), .ZN(n7583) );
  XNOR2_X1 U9174 ( .A(n7584), .B(n7583), .ZN(n7958) );
  XNOR2_X1 U9175 ( .A(n8453), .B(n7612), .ZN(n7592) );
  XNOR2_X1 U9176 ( .A(n7590), .B(n7592), .ZN(n8028) );
  OR2_X1 U9177 ( .A1(n8060), .A2(n5765), .ZN(n8027) );
  NAND2_X1 U9178 ( .A1(n8028), .A2(n8027), .ZN(n8026) );
  OR2_X1 U9179 ( .A1(n4326), .A2(n7591), .ZN(n7593) );
  NAND2_X1 U9180 ( .A1(n7593), .A2(n7592), .ZN(n7594) );
  NAND2_X1 U9181 ( .A1(n8026), .A2(n7594), .ZN(n7598) );
  XNOR2_X1 U9182 ( .A(n8448), .B(n7607), .ZN(n7597) );
  INV_X1 U9183 ( .A(n8210), .ZN(n8248) );
  NOR2_X1 U9184 ( .A1(n8268), .A2(n5765), .ZN(n8006) );
  NAND2_X1 U9185 ( .A1(n8192), .A2(n7602), .ZN(n7966) );
  XNOR2_X1 U9186 ( .A(n8188), .B(n7612), .ZN(n7604) );
  AND2_X1 U9187 ( .A1(n8179), .A2(n7602), .ZN(n7603) );
  NAND2_X1 U9188 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  OAI21_X1 U9189 ( .B1(n7604), .B2(n7603), .A(n7605), .ZN(n8052) );
  INV_X1 U9190 ( .A(n7605), .ZN(n7606) );
  XNOR2_X1 U9191 ( .A(n8428), .B(n7607), .ZN(n7609) );
  NOR2_X1 U9192 ( .A1(n7625), .A2(n5765), .ZN(n7608) );
  NAND2_X1 U9193 ( .A1(n7609), .A2(n7608), .ZN(n7610) );
  OAI21_X1 U9194 ( .B1(n7609), .B2(n7608), .A(n7610), .ZN(n7926) );
  NOR2_X1 U9195 ( .A1(n7927), .A2(n7926), .ZN(n7925) );
  INV_X1 U9196 ( .A(n7610), .ZN(n7611) );
  NOR2_X1 U9197 ( .A1(n7925), .A2(n7611), .ZN(n7622) );
  OR2_X1 U9198 ( .A1(n8145), .A2(n5765), .ZN(n7613) );
  XNOR2_X1 U9199 ( .A(n7613), .B(n7612), .ZN(n7616) );
  NOR3_X1 U9200 ( .A1(n8160), .A2(n7616), .A3(n9876), .ZN(n7614) );
  AOI21_X1 U9201 ( .B1(n7616), .B2(n8160), .A(n7614), .ZN(n7621) );
  NAND3_X1 U9202 ( .A1(n8424), .A2(n9863), .A3(n7616), .ZN(n7615) );
  OAI21_X1 U9203 ( .B1(n8424), .B2(n7616), .A(n7615), .ZN(n7620) );
  INV_X1 U9204 ( .A(n7617), .ZN(n7618) );
  NAND4_X1 U9205 ( .A1(n8424), .A2(P2_STATE_REG_SCAN_IN), .A3(n7618), .A4(
        n9876), .ZN(n7619) );
  OR2_X1 U9206 ( .A1(n7623), .A2(n8404), .ZN(n7624) );
  OAI21_X1 U9207 ( .B1(n7625), .B2(n8402), .A(n7624), .ZN(n8163) );
  AOI22_X1 U9208 ( .A1(n8163), .A2(n9741), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7626) );
  OAI211_X1 U9209 ( .C1(n7628), .C2(n9752), .A(n7627), .B(n7626), .ZN(P2_U3222) );
  INV_X1 U9210 ( .A(n7631), .ZN(n7922) );
  OAI222_X1 U9211 ( .A1(n8539), .A2(n7630), .B1(P2_U3152), .B2(n7629), .C1(
        n8543), .C2(n7922), .ZN(P2_U3330) );
  NAND2_X1 U9212 ( .A1(n7631), .A2(n8760), .ZN(n7633) );
  OR2_X1 U9213 ( .A1(n8758), .A2(n7923), .ZN(n7632) );
  NAND2_X1 U9214 ( .A1(n9393), .A2(n5357), .ZN(n7649) );
  INV_X1 U9215 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7700) );
  INV_X1 U9216 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7737) );
  INV_X1 U9217 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8574) );
  INV_X1 U9218 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8635) );
  INV_X1 U9219 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7840) );
  INV_X1 U9220 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7640) );
  INV_X1 U9221 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7639) );
  OAI21_X1 U9222 ( .B1(n7882), .B2(n7640), .A(n7639), .ZN(n7642) );
  NAND2_X1 U9223 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7641) );
  NAND2_X1 U9224 ( .A1(n9145), .A2(n7897), .ZN(n7647) );
  INV_X1 U9225 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U9226 ( .A1(n7898), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9227 ( .A1(n8748), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7643) );
  OAI211_X1 U9228 ( .C1(n8753), .C2(n10011), .A(n7644), .B(n7643), .ZN(n7645)
         );
  INV_X1 U9229 ( .A(n7645), .ZN(n7646) );
  NAND2_X1 U9230 ( .A1(n7647), .A2(n7646), .ZN(n9123) );
  NAND2_X1 U9231 ( .A1(n9123), .A2(n4264), .ZN(n7648) );
  NAND2_X1 U9232 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  XNOR2_X1 U9233 ( .A(n7650), .B(n5361), .ZN(n7652) );
  AOI22_X1 U9234 ( .A1(n9393), .A2(n7891), .B1(n5377), .B2(n9123), .ZN(n7651)
         );
  XNOR2_X1 U9235 ( .A(n7652), .B(n7651), .ZN(n7912) );
  NOR2_X1 U9236 ( .A1(n7912), .A2(n8664), .ZN(n7910) );
  NAND2_X1 U9237 ( .A1(n7653), .A2(n8760), .ZN(n7656) );
  OR2_X1 U9238 ( .A1(n8758), .A2(n7654), .ZN(n7655) );
  INV_X1 U9239 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7657) );
  NAND2_X1 U9240 ( .A1(n7799), .A2(n7657), .ZN(n7658) );
  NAND2_X1 U9241 ( .A1(n7820), .A2(n7658), .ZN(n9223) );
  OR2_X1 U9242 ( .A1(n9223), .A2(n7863), .ZN(n7664) );
  INV_X1 U9243 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9244 ( .A1(n7898), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9245 ( .A1(n5393), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7659) );
  OAI211_X1 U9246 ( .C1(n7824), .C2(n7661), .A(n7660), .B(n7659), .ZN(n7662)
         );
  INV_X1 U9247 ( .A(n7662), .ZN(n7663) );
  NAND2_X1 U9248 ( .A1(n7664), .A2(n7663), .ZN(n9234) );
  INV_X1 U9249 ( .A(n9234), .ZN(n9090) );
  INV_X1 U9250 ( .A(n5377), .ZN(n7806) );
  OAI22_X1 U9251 ( .A1(n9217), .A2(n5700), .B1(n9090), .B2(n7806), .ZN(n8558)
         );
  INV_X1 U9252 ( .A(n7676), .ZN(n7666) );
  NAND2_X1 U9253 ( .A1(n7666), .A2(n4290), .ZN(n7674) );
  NAND2_X1 U9254 ( .A1(n9506), .A2(n7889), .ZN(n7668) );
  NAND2_X1 U9255 ( .A1(n9342), .A2(n7891), .ZN(n7667) );
  NAND2_X1 U9256 ( .A1(n7668), .A2(n7667), .ZN(n7669) );
  XNOR2_X1 U9257 ( .A(n7669), .B(n5361), .ZN(n7677) );
  INV_X1 U9258 ( .A(n7670), .ZN(n7672) );
  NAND2_X1 U9259 ( .A1(n7672), .A2(n7671), .ZN(n7675) );
  AND2_X1 U9260 ( .A1(n7677), .A2(n7675), .ZN(n7673) );
  NAND2_X1 U9261 ( .A1(n7676), .A2(n7675), .ZN(n7680) );
  INV_X1 U9262 ( .A(n7677), .ZN(n7678) );
  AND2_X1 U9263 ( .A1(n7678), .A2(n4290), .ZN(n7679) );
  NAND2_X1 U9264 ( .A1(n7680), .A2(n7679), .ZN(n8672) );
  NAND2_X1 U9265 ( .A1(n9506), .A2(n7891), .ZN(n7682) );
  NAND2_X1 U9266 ( .A1(n5377), .A2(n9342), .ZN(n7681) );
  NAND2_X1 U9267 ( .A1(n7682), .A2(n7681), .ZN(n8673) );
  NAND2_X1 U9268 ( .A1(n7683), .A2(n8760), .ZN(n7685) );
  AOI22_X1 U9269 ( .A1(n7734), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7733), .B2(
        n9599), .ZN(n7684) );
  NAND2_X1 U9270 ( .A1(n9360), .A2(n7889), .ZN(n7687) );
  NAND2_X1 U9271 ( .A1(n9328), .A2(n4264), .ZN(n7686) );
  NAND2_X1 U9272 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  XNOR2_X1 U9273 ( .A(n7688), .B(n7872), .ZN(n7690) );
  AND2_X1 U9274 ( .A1(n5377), .A2(n9328), .ZN(n7689) );
  AOI21_X1 U9275 ( .B1(n9360), .B2(n7891), .A(n7689), .ZN(n7691) );
  NAND2_X1 U9276 ( .A1(n7690), .A2(n7691), .ZN(n7695) );
  INV_X1 U9277 ( .A(n7690), .ZN(n7693) );
  INV_X1 U9278 ( .A(n7691), .ZN(n7692) );
  NAND2_X1 U9279 ( .A1(n7693), .A2(n7692), .ZN(n7694) );
  AND2_X1 U9280 ( .A1(n7695), .A2(n7694), .ZN(n8592) );
  NAND2_X1 U9281 ( .A1(n7696), .A2(n8760), .ZN(n7698) );
  AOI22_X1 U9282 ( .A1(n7734), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7733), .B2(
        n9610), .ZN(n7697) );
  NAND2_X1 U9283 ( .A1(n9448), .A2(n7889), .ZN(n7708) );
  NAND2_X1 U9284 ( .A1(n8748), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7706) );
  INV_X1 U9285 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7699) );
  OR2_X1 U9286 ( .A1(n7783), .A2(n7699), .ZN(n7705) );
  INV_X1 U9287 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9055) );
  OR2_X1 U9288 ( .A1(n8753), .A2(n9055), .ZN(n7704) );
  NAND2_X1 U9289 ( .A1(n7701), .A2(n7700), .ZN(n7702) );
  NAND2_X1 U9290 ( .A1(n7719), .A2(n7702), .ZN(n9319) );
  OR2_X1 U9291 ( .A1(n7863), .A2(n9319), .ZN(n7703) );
  NAND4_X1 U9292 ( .A1(n7706), .A2(n7705), .A3(n7704), .A4(n7703), .ZN(n9302)
         );
  NAND2_X1 U9293 ( .A1(n9302), .A2(n7891), .ZN(n7707) );
  NAND2_X1 U9294 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  XNOR2_X1 U9295 ( .A(n7709), .B(n5361), .ZN(n7711) );
  AND2_X1 U9296 ( .A1(n5377), .A2(n9302), .ZN(n7710) );
  AOI21_X1 U9297 ( .B1(n9448), .B2(n7891), .A(n7710), .ZN(n7712) );
  XNOR2_X1 U9298 ( .A(n7711), .B(n7712), .ZN(n8605) );
  INV_X1 U9299 ( .A(n7711), .ZN(n7713) );
  NAND2_X1 U9300 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  NAND2_X1 U9301 ( .A1(n7715), .A2(n8760), .ZN(n7717) );
  AOI22_X1 U9302 ( .A1(n7734), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7733), .B2(
        n9627), .ZN(n7716) );
  NAND2_X1 U9303 ( .A1(n9311), .A2(n7889), .ZN(n7726) );
  NAND2_X1 U9304 ( .A1(n8748), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7724) );
  INV_X1 U9305 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U9306 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  NAND2_X1 U9307 ( .A1(n7738), .A2(n7720), .ZN(n9309) );
  OR2_X1 U9308 ( .A1(n9309), .A2(n7863), .ZN(n7723) );
  INV_X1 U9309 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9057) );
  OR2_X1 U9310 ( .A1(n8753), .A2(n9057), .ZN(n7722) );
  INV_X1 U9311 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9044) );
  OR2_X1 U9312 ( .A1(n7783), .A2(n9044), .ZN(n7721) );
  NAND4_X1 U9313 ( .A1(n7724), .A2(n7723), .A3(n7722), .A4(n7721), .ZN(n9330)
         );
  NAND2_X1 U9314 ( .A1(n9330), .A2(n7891), .ZN(n7725) );
  NAND2_X1 U9315 ( .A1(n7726), .A2(n7725), .ZN(n7727) );
  XNOR2_X1 U9316 ( .A(n7727), .B(n7872), .ZN(n7730) );
  NAND2_X1 U9317 ( .A1(n9311), .A2(n4264), .ZN(n7729) );
  NAND2_X1 U9318 ( .A1(n5377), .A2(n9330), .ZN(n7728) );
  NAND2_X1 U9319 ( .A1(n7729), .A2(n7728), .ZN(n8643) );
  NAND2_X1 U9320 ( .A1(n7732), .A2(n8760), .ZN(n7736) );
  AOI22_X1 U9321 ( .A1(n7734), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5586), .B2(
        n7733), .ZN(n7735) );
  NAND2_X1 U9322 ( .A1(n9436), .A2(n7889), .ZN(n7746) );
  NAND2_X1 U9323 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  NAND2_X1 U9324 ( .A1(n7759), .A2(n7739), .ZN(n9286) );
  INV_X1 U9325 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9059) );
  OR2_X1 U9326 ( .A1(n8753), .A2(n9059), .ZN(n7742) );
  INV_X1 U9327 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n7740) );
  OR2_X1 U9328 ( .A1(n7824), .A2(n7740), .ZN(n7741) );
  AND2_X1 U9329 ( .A1(n7742), .A2(n7741), .ZN(n7744) );
  NAND2_X1 U9330 ( .A1(n7898), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7743) );
  OAI211_X1 U9331 ( .C1(n9286), .C2(n7863), .A(n7744), .B(n7743), .ZN(n9303)
         );
  NAND2_X1 U9332 ( .A1(n9303), .A2(n4264), .ZN(n7745) );
  NAND2_X1 U9333 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  XNOR2_X1 U9334 ( .A(n7747), .B(n7872), .ZN(n7749) );
  AND2_X1 U9335 ( .A1(n9303), .A2(n5377), .ZN(n7748) );
  AOI21_X1 U9336 ( .B1(n9436), .B2(n4264), .A(n7748), .ZN(n7750) );
  NAND2_X1 U9337 ( .A1(n7749), .A2(n7750), .ZN(n8622) );
  INV_X1 U9338 ( .A(n7749), .ZN(n7752) );
  INV_X1 U9339 ( .A(n7750), .ZN(n7751) );
  NAND2_X1 U9340 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  NAND2_X1 U9341 ( .A1(n7754), .A2(n8760), .ZN(n7757) );
  OR2_X1 U9342 ( .A1(n8758), .A2(n7755), .ZN(n7756) );
  NAND2_X1 U9343 ( .A1(n9430), .A2(n7889), .ZN(n7765) );
  INV_X1 U9344 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n7763) );
  INV_X1 U9345 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U9346 ( .A1(n7759), .A2(n7758), .ZN(n7760) );
  NAND2_X1 U9347 ( .A1(n7779), .A2(n7760), .ZN(n9265) );
  OR2_X1 U9348 ( .A1(n9265), .A2(n7863), .ZN(n7762) );
  AOI22_X1 U9349 ( .A1(n5393), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n8748), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n7761) );
  OAI211_X1 U9350 ( .C1(n7783), .C2(n7763), .A(n7762), .B(n7761), .ZN(n9250)
         );
  NAND2_X1 U9351 ( .A1(n9250), .A2(n7891), .ZN(n7764) );
  NAND2_X1 U9352 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  XNOR2_X1 U9353 ( .A(n7766), .B(n7872), .ZN(n7768) );
  AND2_X1 U9354 ( .A1(n9250), .A2(n5377), .ZN(n7767) );
  AOI21_X1 U9355 ( .B1(n9430), .B2(n4264), .A(n7767), .ZN(n7769) );
  NAND2_X1 U9356 ( .A1(n7768), .A2(n7769), .ZN(n7773) );
  INV_X1 U9357 ( .A(n7768), .ZN(n7771) );
  INV_X1 U9358 ( .A(n7769), .ZN(n7770) );
  NAND2_X1 U9359 ( .A1(n7771), .A2(n7770), .ZN(n7772) );
  NAND2_X1 U9360 ( .A1(n7773), .A2(n7772), .ZN(n8621) );
  INV_X1 U9361 ( .A(n7773), .ZN(n7774) );
  NAND2_X1 U9362 ( .A1(n7775), .A2(n8760), .ZN(n7778) );
  OR2_X1 U9363 ( .A1(n8758), .A2(n7776), .ZN(n7777) );
  NAND2_X1 U9364 ( .A1(n7779), .A2(n8574), .ZN(n7780) );
  NAND2_X1 U9365 ( .A1(n7797), .A2(n7780), .ZN(n9258) );
  OR2_X1 U9366 ( .A1(n9258), .A2(n7863), .ZN(n7786) );
  INV_X1 U9367 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U9368 ( .A1(n5393), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U9369 ( .A1(n8748), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7781) );
  OAI211_X1 U9370 ( .C1(n9259), .C2(n7783), .A(n7782), .B(n7781), .ZN(n7784)
         );
  INV_X1 U9371 ( .A(n7784), .ZN(n7785) );
  NAND2_X1 U9372 ( .A1(n7786), .A2(n7785), .ZN(n9271) );
  AOI22_X1 U9373 ( .A1(n9426), .A2(n7891), .B1(n5377), .B2(n9271), .ZN(n7791)
         );
  NAND2_X1 U9374 ( .A1(n9426), .A2(n7889), .ZN(n7788) );
  NAND2_X1 U9375 ( .A1(n9271), .A2(n7891), .ZN(n7787) );
  NAND2_X1 U9376 ( .A1(n7788), .A2(n7787), .ZN(n7789) );
  XNOR2_X1 U9377 ( .A(n7789), .B(n5361), .ZN(n7790) );
  XOR2_X1 U9378 ( .A(n7791), .B(n7790), .Z(n8572) );
  INV_X1 U9379 ( .A(n7790), .ZN(n7792) );
  NAND2_X1 U9380 ( .A1(n7793), .A2(n8760), .ZN(n7796) );
  OR2_X1 U9381 ( .A1(n8758), .A2(n7794), .ZN(n7795) );
  NAND2_X1 U9382 ( .A1(n7797), .A2(n8635), .ZN(n7798) );
  NAND2_X1 U9383 ( .A1(n7799), .A2(n7798), .ZN(n8638) );
  INV_X1 U9384 ( .A(n8638), .ZN(n9236) );
  NAND2_X1 U9385 ( .A1(n9236), .A2(n7897), .ZN(n7805) );
  INV_X1 U9386 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U9387 ( .A1(n7898), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U9388 ( .A1(n8748), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7800) );
  OAI211_X1 U9389 ( .C1(n8753), .C2(n7802), .A(n7801), .B(n7800), .ZN(n7803)
         );
  INV_X1 U9390 ( .A(n7803), .ZN(n7804) );
  OAI22_X1 U9391 ( .A1(n9231), .A2(n5700), .B1(n9088), .B2(n7806), .ZN(n7810)
         );
  NAND2_X1 U9392 ( .A1(n7811), .A2(n7810), .ZN(n8632) );
  NAND2_X1 U9393 ( .A1(n9415), .A2(n7889), .ZN(n7808) );
  NAND2_X1 U9394 ( .A1(n9234), .A2(n7891), .ZN(n7807) );
  NAND2_X1 U9395 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  XNOR2_X1 U9396 ( .A(n7809), .B(n7872), .ZN(n7813) );
  OR2_X1 U9397 ( .A1(n7811), .A2(n7810), .ZN(n8631) );
  AOI22_X1 U9398 ( .A1(n9420), .A2(n5357), .B1(n4264), .B2(n9251), .ZN(n7812)
         );
  XOR2_X1 U9399 ( .A(n5361), .B(n7812), .Z(n8634) );
  NAND2_X1 U9400 ( .A1(n8631), .A2(n8634), .ZN(n7814) );
  AOI21_X2 U9401 ( .B1(n7814), .B2(n8632), .A(n7813), .ZN(n8556) );
  NAND2_X1 U9402 ( .A1(n7815), .A2(n8760), .ZN(n7818) );
  OR2_X1 U9403 ( .A1(n8758), .A2(n7816), .ZN(n7817) );
  NAND2_X1 U9404 ( .A1(n9411), .A2(n7889), .ZN(n7829) );
  INV_X1 U9405 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U9406 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  NAND2_X1 U9407 ( .A1(n7841), .A2(n7821), .ZN(n8615) );
  OR2_X1 U9408 ( .A1(n8615), .A2(n7863), .ZN(n7827) );
  INV_X1 U9409 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U9410 ( .A1(n5393), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U9411 ( .A1(n7898), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7822) );
  OAI211_X1 U9412 ( .C1(n7824), .C2(n9979), .A(n7823), .B(n7822), .ZN(n7825)
         );
  INV_X1 U9413 ( .A(n7825), .ZN(n7826) );
  NAND2_X1 U9414 ( .A1(n7827), .A2(n7826), .ZN(n9221) );
  NAND2_X1 U9415 ( .A1(n9221), .A2(n7891), .ZN(n7828) );
  NAND2_X1 U9416 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  XNOR2_X1 U9417 ( .A(n7830), .B(n5361), .ZN(n7834) );
  NAND2_X1 U9418 ( .A1(n9411), .A2(n4264), .ZN(n7832) );
  NAND2_X1 U9419 ( .A1(n9221), .A2(n5377), .ZN(n7831) );
  NAND2_X1 U9420 ( .A1(n7832), .A2(n7831), .ZN(n7833) );
  AOI21_X1 U9421 ( .B1(n7834), .B2(n7833), .A(n7835), .ZN(n8612) );
  INV_X1 U9422 ( .A(n7835), .ZN(n7836) );
  OR2_X1 U9423 ( .A1(n8758), .A2(n7838), .ZN(n7839) );
  NAND2_X1 U9424 ( .A1(n9094), .A2(n7889), .ZN(n7850) );
  NAND2_X1 U9425 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  NAND2_X1 U9426 ( .A1(n9192), .A2(n7897), .ZN(n7848) );
  INV_X1 U9427 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U9428 ( .A1(n7898), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U9429 ( .A1(n8748), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7843) );
  OAI211_X1 U9430 ( .C1(n8753), .C2(n7845), .A(n7844), .B(n7843), .ZN(n7846)
         );
  INV_X1 U9431 ( .A(n7846), .ZN(n7847) );
  NAND2_X1 U9432 ( .A1(n7848), .A2(n7847), .ZN(n9207) );
  NAND2_X1 U9433 ( .A1(n9207), .A2(n7891), .ZN(n7849) );
  NAND2_X1 U9434 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  AOI22_X1 U9435 ( .A1(n9094), .A2(n7891), .B1(n5377), .B2(n9207), .ZN(n7852)
         );
  XNOR2_X1 U9436 ( .A(n7854), .B(n7852), .ZN(n8583) );
  INV_X1 U9437 ( .A(n7852), .ZN(n7853) );
  INV_X1 U9438 ( .A(n8654), .ZN(n7877) );
  OR2_X1 U9439 ( .A1(n8758), .A2(n7857), .ZN(n7858) );
  NAND2_X1 U9440 ( .A1(n9402), .A2(n5357), .ZN(n7871) );
  INV_X1 U9441 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U9442 ( .A1(n7861), .A2(n7860), .ZN(n7862) );
  NAND2_X1 U9443 ( .A1(n7882), .A2(n7862), .ZN(n9177) );
  INV_X1 U9444 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U9445 ( .A1(n7898), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U9446 ( .A1(n8748), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7864) );
  OAI211_X1 U9447 ( .C1(n8753), .C2(n7866), .A(n7865), .B(n7864), .ZN(n7867)
         );
  INV_X1 U9448 ( .A(n7867), .ZN(n7868) );
  NAND2_X1 U9449 ( .A1(n9186), .A2(n4264), .ZN(n7870) );
  NAND2_X1 U9450 ( .A1(n7871), .A2(n7870), .ZN(n7873) );
  XNOR2_X1 U9451 ( .A(n7873), .B(n7872), .ZN(n7876) );
  AND2_X1 U9452 ( .A1(n9186), .A2(n5377), .ZN(n7874) );
  AOI21_X1 U9453 ( .B1(n9402), .B2(n7891), .A(n7874), .ZN(n7875) );
  NOR2_X1 U9454 ( .A1(n7876), .A2(n7875), .ZN(n8655) );
  NAND2_X1 U9455 ( .A1(n7876), .A2(n7875), .ZN(n8656) );
  OR2_X1 U9456 ( .A1(n8758), .A2(n7879), .ZN(n7880) );
  XNOR2_X1 U9457 ( .A(n7882), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U9458 ( .A1(n9159), .A2(n7897), .ZN(n7888) );
  INV_X1 U9459 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U9460 ( .A1(n7898), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U9461 ( .A1(n8748), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7883) );
  OAI211_X1 U9462 ( .C1(n8753), .C2(n7885), .A(n7884), .B(n7883), .ZN(n7886)
         );
  INV_X1 U9463 ( .A(n7886), .ZN(n7887) );
  NAND2_X1 U9464 ( .A1(n7888), .A2(n7887), .ZN(n9097) );
  AOI22_X1 U9465 ( .A1(n9397), .A2(n7889), .B1(n7891), .B2(n9097), .ZN(n7890)
         );
  XNOR2_X1 U9466 ( .A(n7890), .B(n5361), .ZN(n8545) );
  NAND2_X1 U9467 ( .A1(n9397), .A2(n4264), .ZN(n7893) );
  NAND2_X1 U9468 ( .A1(n9097), .A2(n5377), .ZN(n7892) );
  NAND2_X1 U9469 ( .A1(n7893), .A2(n7892), .ZN(n8546) );
  INV_X1 U9470 ( .A(n8546), .ZN(n7894) );
  AOI21_X1 U9471 ( .B1(n8549), .B2(n8545), .A(n7894), .ZN(n7895) );
  INV_X1 U9472 ( .A(n7895), .ZN(n7916) );
  INV_X1 U9473 ( .A(n9145), .ZN(n7906) );
  INV_X1 U9474 ( .A(n7896), .ZN(n9127) );
  NAND2_X1 U9475 ( .A1(n9127), .A2(n7897), .ZN(n7904) );
  INV_X1 U9476 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U9477 ( .A1(n7898), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U9478 ( .A1(n8748), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7899) );
  OAI211_X1 U9479 ( .C1(n8753), .C2(n7901), .A(n7900), .B(n7899), .ZN(n7902)
         );
  INV_X1 U9480 ( .A(n7902), .ZN(n7903) );
  NAND2_X1 U9481 ( .A1(n7904), .A2(n7903), .ZN(n8987) );
  AOI22_X1 U9482 ( .A1(n8987), .A2(n8659), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7905) );
  OAI21_X1 U9483 ( .B1(n8671), .B2(n7906), .A(n7905), .ZN(n7907) );
  AOI21_X1 U9484 ( .B1(n8668), .B2(n9097), .A(n7907), .ZN(n7908) );
  OAI21_X1 U9485 ( .B1(n9148), .B2(n8653), .A(n7908), .ZN(n7909) );
  AOI21_X1 U9486 ( .B1(n7911), .B2(n7910), .A(n7909), .ZN(n7915) );
  INV_X1 U9487 ( .A(n7911), .ZN(n7914) );
  AND2_X1 U9488 ( .A1(n7912), .A2(n8647), .ZN(n7913) );
  OAI222_X1 U9489 ( .A1(n8533), .A2(n7921), .B1(n7920), .B2(n7919), .C1(n7918), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U9490 ( .A1(n9478), .A2(n7923), .B1(n4258), .B2(n9011), .C1(n7922), 
        .C2(n7551), .ZN(P1_U3325) );
  INV_X1 U9491 ( .A(n8681), .ZN(n8542) );
  OAI222_X1 U9492 ( .A1(n9478), .A2(n8682), .B1(n7551), .B2(n8542), .C1(n7924), 
        .C2(n4258), .ZN(P1_U3324) );
  AOI211_X1 U9493 ( .C1(n7927), .C2(n7926), .A(n9744), .B(n7925), .ZN(n7932)
         );
  INV_X1 U9494 ( .A(n8145), .ZN(n8178) );
  AOI22_X1 U9495 ( .A1(n8178), .A2(n9721), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n7930) );
  INV_X1 U9496 ( .A(n7928), .ZN(n8173) );
  AOI22_X1 U9497 ( .A1(n9724), .A2(n8179), .B1(n8173), .B2(n8054), .ZN(n7929)
         );
  OAI211_X1 U9498 ( .C1(n8175), .C2(n9734), .A(n7930), .B(n7929), .ZN(n7931)
         );
  OR2_X1 U9499 ( .A1(n7932), .A2(n7931), .ZN(P2_U3216) );
  XNOR2_X1 U9500 ( .A(n7933), .B(n8006), .ZN(n7938) );
  OAI22_X1 U9501 ( .A1(n8046), .A2(n8210), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7934), .ZN(n7936) );
  OAI22_X1 U9502 ( .A1(n8021), .A2(n8060), .B1(n9752), .B2(n8240), .ZN(n7935)
         );
  AOI211_X1 U9503 ( .C1(n8448), .C2(n9748), .A(n7936), .B(n7935), .ZN(n7937)
         );
  OAI21_X1 U9504 ( .B1(n7938), .B2(n9744), .A(n7937), .ZN(P2_U3218) );
  OR2_X1 U9505 ( .A1(n7955), .A2(n7940), .ZN(n8017) );
  INV_X1 U9506 ( .A(n8017), .ZN(n7939) );
  AOI21_X1 U9507 ( .B1(n7955), .B2(n7940), .A(n7939), .ZN(n7945) );
  AOI22_X1 U9508 ( .A1(n9724), .A2(n8338), .B1(n8311), .B2(n8054), .ZN(n7942)
         );
  OAI211_X1 U9509 ( .C1(n8046), .C2(n8308), .A(n7942), .B(n7941), .ZN(n7943)
         );
  AOI21_X1 U9510 ( .B1(n8470), .B2(n9748), .A(n7943), .ZN(n7944) );
  OAI21_X1 U9511 ( .B1(n7945), .B2(n9744), .A(n7944), .ZN(P2_U3221) );
  AOI22_X1 U9512 ( .A1(n9724), .A2(n8072), .B1(n9721), .B2(n9723), .ZN(n7953)
         );
  AOI22_X1 U9513 ( .A1(n9748), .A2(n7946), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8038), .ZN(n7952) );
  OAI21_X1 U9514 ( .B1(n7949), .B2(n7948), .A(n7947), .ZN(n7950) );
  NAND2_X1 U9515 ( .A1(n7950), .A2(n9730), .ZN(n7951) );
  NAND3_X1 U9516 ( .A1(n7953), .A2(n7952), .A3(n7951), .ZN(P2_U3224) );
  OR2_X1 U9517 ( .A1(n7955), .A2(n7954), .ZN(n7957) );
  AND2_X1 U9518 ( .A1(n7957), .A2(n7956), .ZN(n7959) );
  XNOR2_X1 U9519 ( .A(n7959), .B(n7958), .ZN(n7965) );
  OAI22_X1 U9520 ( .A1(n8046), .A2(n8060), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7960), .ZN(n7963) );
  INV_X1 U9521 ( .A(n8277), .ZN(n7961) );
  OAI22_X1 U9522 ( .A1(n8021), .A2(n8308), .B1(n7961), .B2(n9752), .ZN(n7962)
         );
  AOI211_X1 U9523 ( .C1(n8458), .C2(n9748), .A(n7963), .B(n7962), .ZN(n7964)
         );
  OAI21_X1 U9524 ( .B1(n7965), .B2(n9744), .A(n7964), .ZN(P2_U3225) );
  XNOR2_X1 U9525 ( .A(n7967), .B(n7966), .ZN(n7968) );
  XNOR2_X1 U9526 ( .A(n7969), .B(n7968), .ZN(n7974) );
  OAI22_X1 U9527 ( .A1(n8021), .A2(n8210), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10013), .ZN(n7972) );
  INV_X1 U9528 ( .A(n8213), .ZN(n7970) );
  OAI22_X1 U9529 ( .A1(n8046), .A2(n8211), .B1(n9752), .B2(n7970), .ZN(n7971)
         );
  AOI211_X1 U9530 ( .C1(n8440), .C2(n9748), .A(n7972), .B(n7971), .ZN(n7973)
         );
  OAI21_X1 U9531 ( .B1(n7974), .B2(n9744), .A(n7973), .ZN(P2_U3227) );
  OR2_X1 U9532 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  NAND2_X1 U9533 ( .A1(n7978), .A2(n7977), .ZN(n7981) );
  INV_X1 U9534 ( .A(n7979), .ZN(n7980) );
  AOI21_X1 U9535 ( .B1(n7982), .B2(n7981), .A(n7980), .ZN(n7986) );
  INV_X1 U9536 ( .A(n8405), .ZN(n8062) );
  AOI22_X1 U9537 ( .A1(n9724), .A2(n8062), .B1(n8366), .B2(n8054), .ZN(n7983)
         );
  NAND2_X1 U9538 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8076) );
  OAI211_X1 U9539 ( .C1(n8046), .C2(n8358), .A(n7983), .B(n8076), .ZN(n7984)
         );
  AOI21_X1 U9540 ( .B1(n8483), .B2(n9748), .A(n7984), .ZN(n7985) );
  OAI21_X1 U9541 ( .B1(n7986), .B2(n9744), .A(n7985), .ZN(P2_U3228) );
  OAI211_X1 U9542 ( .C1(n7989), .C2(n7988), .A(n7987), .B(n9730), .ZN(n7997)
         );
  AOI22_X1 U9543 ( .A1(n9724), .A2(n9720), .B1(n7990), .B2(n8054), .ZN(n7996)
         );
  OAI22_X1 U9544 ( .A1(n8046), .A2(n7992), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7991), .ZN(n7993) );
  AOI21_X1 U9545 ( .B1(n9748), .B2(n7994), .A(n7993), .ZN(n7995) );
  NAND3_X1 U9546 ( .A1(n7997), .A2(n7996), .A3(n7995), .ZN(P2_U3229) );
  XNOR2_X1 U9547 ( .A(n7999), .B(n7998), .ZN(n8004) );
  OAI22_X1 U9548 ( .A1(n8046), .A2(n8307), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9989), .ZN(n8002) );
  INV_X1 U9549 ( .A(n8345), .ZN(n8000) );
  OAI22_X1 U9550 ( .A1(n8021), .A2(n8061), .B1(n8000), .B2(n9752), .ZN(n8001)
         );
  AOI211_X1 U9551 ( .C1(n8480), .C2(n9748), .A(n8002), .B(n8001), .ZN(n8003)
         );
  OAI21_X1 U9552 ( .B1(n8004), .B2(n9744), .A(n8003), .ZN(P2_U3230) );
  AOI21_X1 U9553 ( .B1(n8006), .B2(n7933), .A(n8005), .ZN(n8010) );
  XNOR2_X1 U9554 ( .A(n8008), .B(n8007), .ZN(n8009) );
  XNOR2_X1 U9555 ( .A(n8010), .B(n8009), .ZN(n8015) );
  OAI22_X1 U9556 ( .A1(n8046), .A2(n8232), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8011), .ZN(n8013) );
  OAI22_X1 U9557 ( .A1(n8021), .A2(n8268), .B1(n8223), .B2(n9752), .ZN(n8012)
         );
  AOI211_X1 U9558 ( .C1(n8443), .C2(n9748), .A(n8013), .B(n8012), .ZN(n8014)
         );
  OAI21_X1 U9559 ( .B1(n8015), .B2(n9744), .A(n8014), .ZN(P2_U3231) );
  NAND2_X1 U9560 ( .A1(n8017), .A2(n8016), .ZN(n8019) );
  XNOR2_X1 U9561 ( .A(n8019), .B(n8018), .ZN(n8025) );
  OAI22_X1 U9562 ( .A1(n8046), .A2(n8267), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10010), .ZN(n8023) );
  INV_X1 U9563 ( .A(n8291), .ZN(n8020) );
  OAI22_X1 U9564 ( .A1(n8021), .A2(n8135), .B1(n8020), .B2(n9752), .ZN(n8022)
         );
  AOI211_X1 U9565 ( .C1(n8463), .C2(n9748), .A(n8023), .B(n8022), .ZN(n8024)
         );
  OAI21_X1 U9566 ( .B1(n8025), .B2(n9744), .A(n8024), .ZN(P2_U3235) );
  OAI21_X1 U9567 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8032) );
  INV_X1 U9568 ( .A(n8453), .ZN(n8261) );
  INV_X1 U9569 ( .A(n8268), .ZN(n8059) );
  AOI22_X1 U9570 ( .A1(n9721), .A2(n8059), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8030) );
  INV_X1 U9571 ( .A(n8267), .ZN(n8297) );
  AOI22_X1 U9572 ( .A1(n9724), .A2(n8297), .B1(n8259), .B2(n8054), .ZN(n8029)
         );
  OAI211_X1 U9573 ( .C1(n8261), .C2(n9734), .A(n8030), .B(n8029), .ZN(n8031)
         );
  AOI21_X1 U9574 ( .B1(n8032), .B2(n9730), .A(n8031), .ZN(n8033) );
  INV_X1 U9575 ( .A(n8033), .ZN(P2_U3237) );
  AND2_X1 U9576 ( .A1(n7947), .A2(n8034), .ZN(n8037) );
  OAI211_X1 U9577 ( .C1(n8037), .C2(n8036), .A(n8035), .B(n9730), .ZN(n8042)
         );
  AOI22_X1 U9578 ( .A1(n9721), .A2(n8069), .B1(n9724), .B2(n8070), .ZN(n8041)
         );
  AOI22_X1 U9579 ( .A1(n9748), .A2(n8039), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8038), .ZN(n8040) );
  NAND3_X1 U9580 ( .A1(n8042), .A2(n8041), .A3(n8040), .ZN(P2_U3239) );
  XNOR2_X1 U9581 ( .A(n8044), .B(n8043), .ZN(n8049) );
  INV_X1 U9582 ( .A(n8358), .ZN(n8326) );
  AOI22_X1 U9583 ( .A1(n9724), .A2(n8326), .B1(n8321), .B2(n8054), .ZN(n8045)
         );
  NAND2_X1 U9584 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8105) );
  OAI211_X1 U9585 ( .C1(n8046), .C2(n8135), .A(n8045), .B(n8105), .ZN(n8047)
         );
  AOI21_X1 U9586 ( .B1(n8473), .B2(n9748), .A(n8047), .ZN(n8048) );
  OAI21_X1 U9587 ( .B1(n8049), .B2(n9744), .A(n8048), .ZN(P2_U3240) );
  AOI211_X1 U9588 ( .C1(n8052), .C2(n8051), .A(n9744), .B(n8050), .ZN(n8058)
         );
  AOI22_X1 U9589 ( .A1(n8193), .A2(n9721), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8056) );
  INV_X1 U9590 ( .A(n8053), .ZN(n8197) );
  AOI22_X1 U9591 ( .A1(n9724), .A2(n8192), .B1(n8197), .B2(n8054), .ZN(n8055)
         );
  OAI211_X1 U9592 ( .C1(n8188), .C2(n9734), .A(n8056), .B(n8055), .ZN(n8057)
         );
  OR2_X1 U9593 ( .A1(n8058), .A2(n8057), .ZN(P2_U3242) );
  MUX2_X1 U9594 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8178), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9595 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8193), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9596 ( .A(n8179), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8071), .Z(
        P2_U3578) );
  MUX2_X1 U9597 ( .A(n8192), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8071), .Z(
        P2_U3577) );
  MUX2_X1 U9598 ( .A(n8248), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8071), .Z(
        P2_U3576) );
  MUX2_X1 U9599 ( .A(n8059), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8071), .Z(
        P2_U3575) );
  INV_X1 U9600 ( .A(n8060), .ZN(n8283) );
  MUX2_X1 U9601 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8283), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9602 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8297), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U9603 ( .A(n8308), .ZN(n8282) );
  MUX2_X1 U9604 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8282), .S(P2_U3966), .Z(
        P2_U3572) );
  INV_X1 U9605 ( .A(n8135), .ZN(n8327) );
  MUX2_X1 U9606 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8327), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9607 ( .A(n8338), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8071), .Z(
        P2_U3570) );
  MUX2_X1 U9608 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8326), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U9609 ( .A(n8061), .ZN(n8385) );
  MUX2_X1 U9610 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8385), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9611 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8062), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9612 ( .A(n8384), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8071), .Z(
        P2_U3566) );
  MUX2_X1 U9613 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8123), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9614 ( .A(n9776), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8071), .Z(
        P2_U3564) );
  MUX2_X1 U9615 ( .A(n8063), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8071), .Z(
        P2_U3563) );
  MUX2_X1 U9616 ( .A(n9777), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8071), .Z(
        P2_U3562) );
  MUX2_X1 U9617 ( .A(n8064), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8071), .Z(
        P2_U3561) );
  MUX2_X1 U9618 ( .A(n8065), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8071), .Z(
        P2_U3560) );
  MUX2_X1 U9619 ( .A(n8066), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8071), .Z(
        P2_U3559) );
  MUX2_X1 U9620 ( .A(n8067), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8071), .Z(
        P2_U3558) );
  MUX2_X1 U9621 ( .A(n8068), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8071), .Z(
        P2_U3557) );
  MUX2_X1 U9622 ( .A(n9720), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8071), .Z(
        P2_U3556) );
  MUX2_X1 U9623 ( .A(n8069), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8071), .Z(
        P2_U3555) );
  MUX2_X1 U9624 ( .A(n9723), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8071), .Z(
        P2_U3554) );
  MUX2_X1 U9625 ( .A(n8070), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8071), .Z(
        P2_U3553) );
  MUX2_X1 U9626 ( .A(n8072), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8071), .Z(
        P2_U3552) );
  AOI21_X1 U9627 ( .B1(n8075), .B2(n8074), .A(n8073), .ZN(n8084) );
  INV_X1 U9628 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9952) );
  OAI21_X1 U9629 ( .B1(n8106), .B2(n9952), .A(n8076), .ZN(n8081) );
  AOI211_X1 U9630 ( .C1(n8079), .C2(n8078), .A(n8091), .B(n8077), .ZN(n8080)
         );
  AOI211_X1 U9631 ( .C1(n8109), .C2(n8082), .A(n8081), .B(n8080), .ZN(n8083)
         );
  OAI21_X1 U9632 ( .B1(n8084), .B2(n9759), .A(n8083), .ZN(P2_U3261) );
  XNOR2_X1 U9633 ( .A(n8086), .B(n8085), .ZN(n8096) );
  NOR2_X1 U9634 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9989), .ZN(n8087) );
  AOI21_X1 U9635 ( .B1(n9754), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8087), .ZN(
        n8088) );
  OAI21_X1 U9636 ( .B1(n9757), .B2(n8089), .A(n8088), .ZN(n8095) );
  AOI211_X1 U9637 ( .C1(n8093), .C2(n8092), .A(n8091), .B(n8090), .ZN(n8094)
         );
  AOI211_X1 U9638 ( .C1(n8096), .C2(n9753), .A(n8095), .B(n8094), .ZN(n8097)
         );
  INV_X1 U9639 ( .A(n8097), .ZN(P2_U3262) );
  AOI21_X1 U9640 ( .B1(n8100), .B2(n8099), .A(n8098), .ZN(n8112) );
  OAI21_X1 U9641 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8104) );
  NAND2_X1 U9642 ( .A1(n8104), .A2(n4352), .ZN(n8111) );
  OAI21_X1 U9643 ( .B1(n8106), .B2(n10084), .A(n8105), .ZN(n8107) );
  AOI21_X1 U9644 ( .B1(n8109), .B2(n8108), .A(n8107), .ZN(n8110) );
  OAI211_X1 U9645 ( .C1(n8112), .C2(n9759), .A(n8111), .B(n8110), .ZN(P2_U3263) );
  INV_X1 U9646 ( .A(n8495), .ZN(n8399) );
  NAND2_X1 U9647 ( .A1(n8392), .A2(n8399), .ZN(n8393) );
  INV_X1 U9648 ( .A(n8480), .ZN(n8348) );
  INV_X1 U9649 ( .A(n8473), .ZN(n8323) );
  NOR2_X1 U9650 ( .A1(n8416), .A2(n8147), .ZN(n8113) );
  XOR2_X1 U9651 ( .A(n7362), .B(n8113), .Z(n8414) );
  NAND2_X1 U9652 ( .A1(n8114), .A2(P2_B_REG_SCAN_IN), .ZN(n8115) );
  NAND2_X1 U9653 ( .A1(n9775), .A2(n8115), .ZN(n8144) );
  NOR2_X1 U9654 ( .A1(n8116), .A2(n8144), .ZN(n8415) );
  INV_X1 U9655 ( .A(n8415), .ZN(n8117) );
  NOR2_X1 U9656 ( .A1(n8117), .A2(n9813), .ZN(n8120) );
  AOI21_X1 U9657 ( .B1(n9813), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8120), .ZN(
        n8119) );
  NAND2_X1 U9658 ( .A1(n7362), .A2(n9803), .ZN(n8118) );
  OAI211_X1 U9659 ( .C1(n8414), .C2(n8369), .A(n8119), .B(n8118), .ZN(P2_U3265) );
  XNOR2_X1 U9660 ( .A(n8416), .B(n8147), .ZN(n8418) );
  AOI21_X1 U9661 ( .B1(n9813), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8120), .ZN(
        n8122) );
  NAND2_X1 U9662 ( .A1(n8416), .A2(n9803), .ZN(n8121) );
  OAI211_X1 U9663 ( .C1(n8418), .C2(n8369), .A(n8122), .B(n8121), .ZN(P2_U3266) );
  INV_X1 U9664 ( .A(n8463), .ZN(n8293) );
  INV_X1 U9665 ( .A(n8470), .ZN(n8136) );
  NAND2_X1 U9666 ( .A1(n9493), .A2(n8123), .ZN(n8129) );
  INV_X1 U9667 ( .A(n8129), .ZN(n8124) );
  INV_X1 U9668 ( .A(n8490), .ZN(n8379) );
  NAND2_X1 U9669 ( .A1(n8379), .A2(n8405), .ZN(n8133) );
  NAND2_X1 U9670 ( .A1(n8372), .A2(n8133), .ZN(n8351) );
  NAND2_X1 U9671 ( .A1(n8473), .A2(n8338), .ZN(n8134) );
  AOI22_X1 U9672 ( .A1(n8317), .A2(n8134), .B1(n8323), .B2(n8307), .ZN(n8303)
         );
  NAND2_X1 U9673 ( .A1(n8303), .A2(n8305), .ZN(n8302) );
  NAND2_X1 U9674 ( .A1(n8279), .A2(n8267), .ZN(n8137) );
  INV_X1 U9675 ( .A(n8448), .ZN(n8243) );
  NAND2_X1 U9676 ( .A1(n8203), .A2(n8138), .ZN(n8186) );
  NAND2_X1 U9677 ( .A1(n8169), .A2(n8176), .ZN(n8168) );
  NAND2_X1 U9678 ( .A1(n8175), .A2(n7625), .ZN(n8139) );
  INV_X1 U9679 ( .A(n8421), .ZN(n8150) );
  NOR2_X1 U9680 ( .A1(n8419), .A2(n8369), .ZN(n8152) );
  AOI22_X1 U9681 ( .A1(n8148), .A2(n9802), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9813), .ZN(n8149) );
  OAI21_X1 U9682 ( .B1(n8150), .B2(n8398), .A(n8149), .ZN(n8151) );
  AOI211_X1 U9683 ( .C1(n8420), .C2(n9783), .A(n8152), .B(n8151), .ZN(n8153)
         );
  OAI21_X1 U9684 ( .B1(n8422), .B2(n8412), .A(n8153), .ZN(P2_U3267) );
  OAI21_X1 U9685 ( .B1(n8155), .B2(n8161), .A(n8154), .ZN(n8156) );
  INV_X1 U9686 ( .A(n8156), .ZN(n8427) );
  INV_X1 U9687 ( .A(n8171), .ZN(n8157) );
  AOI211_X1 U9688 ( .C1(n8424), .C2(n8157), .A(n9865), .B(n4537), .ZN(n8423)
         );
  AOI22_X1 U9689 ( .A1(n8158), .A2(n9802), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9813), .ZN(n8159) );
  OAI21_X1 U9690 ( .B1(n8160), .B2(n8398), .A(n8159), .ZN(n8166) );
  XNOR2_X1 U9691 ( .A(n8162), .B(n8161), .ZN(n8164) );
  NOR2_X1 U9692 ( .A1(n8426), .A2(n9813), .ZN(n8165) );
  AOI211_X1 U9693 ( .C1(n8423), .C2(n8344), .A(n8166), .B(n8165), .ZN(n8167)
         );
  OAI21_X1 U9694 ( .B1(n8427), .B2(n8412), .A(n8167), .ZN(P2_U3268) );
  OAI21_X1 U9695 ( .B1(n8169), .B2(n8176), .A(n8168), .ZN(n8170) );
  INV_X1 U9696 ( .A(n8170), .ZN(n8432) );
  INV_X1 U9697 ( .A(n8195), .ZN(n8172) );
  AOI21_X1 U9698 ( .B1(n8428), .B2(n8172), .A(n8171), .ZN(n8429) );
  AOI22_X1 U9699 ( .A1(n8173), .A2(n9802), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9813), .ZN(n8174) );
  OAI21_X1 U9700 ( .B1(n8175), .B2(n8398), .A(n8174), .ZN(n8182) );
  XOR2_X1 U9701 ( .A(n8177), .B(n8176), .Z(n8180) );
  AOI222_X1 U9702 ( .A1(n9771), .A2(n8180), .B1(n8179), .B2(n9778), .C1(n8178), 
        .C2(n9775), .ZN(n8431) );
  NOR2_X1 U9703 ( .A1(n8431), .A2(n9813), .ZN(n8181) );
  AOI211_X1 U9704 ( .C1(n8429), .C2(n9809), .A(n8182), .B(n8181), .ZN(n8183)
         );
  OAI21_X1 U9705 ( .B1(n8432), .B2(n8412), .A(n8183), .ZN(P2_U3269) );
  OAI21_X1 U9706 ( .B1(n8186), .B2(n8185), .A(n8184), .ZN(n8187) );
  INV_X1 U9707 ( .A(n8187), .ZN(n8437) );
  NOR2_X1 U9708 ( .A1(n8188), .A2(n8398), .ZN(n8201) );
  OAI21_X1 U9709 ( .B1(n8191), .B2(n8190), .A(n8189), .ZN(n8194) );
  AOI222_X1 U9710 ( .A1(n9771), .A2(n8194), .B1(n8193), .B2(n9775), .C1(n8192), 
        .C2(n9778), .ZN(n8436) );
  INV_X1 U9711 ( .A(n8212), .ZN(n8196) );
  AOI211_X1 U9712 ( .C1(n8434), .C2(n8196), .A(n9865), .B(n8195), .ZN(n8433)
         );
  AOI22_X1 U9713 ( .A1(n8433), .A2(n8198), .B1(n9802), .B2(n8197), .ZN(n8199)
         );
  AOI21_X1 U9714 ( .B1(n8436), .B2(n8199), .A(n9813), .ZN(n8200) );
  AOI211_X1 U9715 ( .C1(n9813), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8201), .B(
        n8200), .ZN(n8202) );
  OAI21_X1 U9716 ( .B1(n8437), .B2(n8412), .A(n8202), .ZN(P2_U3270) );
  OAI21_X1 U9717 ( .B1(n8205), .B2(n8204), .A(n8203), .ZN(n8206) );
  INV_X1 U9718 ( .A(n8206), .ZN(n8442) );
  XNOR2_X1 U9719 ( .A(n8208), .B(n8207), .ZN(n8209) );
  OAI222_X1 U9720 ( .A1(n8404), .A2(n8211), .B1(n8402), .B2(n8210), .C1(n8209), 
        .C2(n9795), .ZN(n8438) );
  AOI211_X1 U9721 ( .C1(n8440), .C2(n8221), .A(n9865), .B(n8212), .ZN(n8439)
         );
  NAND2_X1 U9722 ( .A1(n8439), .A2(n8344), .ZN(n8215) );
  AOI22_X1 U9723 ( .A1(n9813), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8213), .B2(
        n9802), .ZN(n8214) );
  OAI211_X1 U9724 ( .C1(n8216), .C2(n8398), .A(n8215), .B(n8214), .ZN(n8217)
         );
  AOI21_X1 U9725 ( .B1(n8438), .B2(n9783), .A(n8217), .ZN(n8218) );
  OAI21_X1 U9726 ( .B1(n8442), .B2(n8412), .A(n8218), .ZN(P2_U3271) );
  XNOR2_X1 U9727 ( .A(n8220), .B(n8219), .ZN(n8447) );
  INV_X1 U9728 ( .A(n8221), .ZN(n8222) );
  AOI21_X1 U9729 ( .B1(n8443), .B2(n8239), .A(n8222), .ZN(n8444) );
  INV_X1 U9730 ( .A(n8443), .ZN(n8226) );
  INV_X1 U9731 ( .A(n8223), .ZN(n8224) );
  AOI22_X1 U9732 ( .A1(n9813), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8224), .B2(
        n9802), .ZN(n8225) );
  OAI21_X1 U9733 ( .B1(n8226), .B2(n8398), .A(n8225), .ZN(n8236) );
  INV_X1 U9734 ( .A(n8227), .ZN(n8231) );
  AOI21_X1 U9735 ( .B1(n8245), .B2(n8229), .A(n8228), .ZN(n8230) );
  NOR3_X1 U9736 ( .A1(n8231), .A2(n8230), .A3(n9795), .ZN(n8234) );
  OAI22_X1 U9737 ( .A1(n8232), .A2(n8404), .B1(n8268), .B2(n8402), .ZN(n8233)
         );
  NOR2_X1 U9738 ( .A1(n8234), .A2(n8233), .ZN(n8446) );
  NOR2_X1 U9739 ( .A1(n8446), .A2(n9813), .ZN(n8235) );
  AOI211_X1 U9740 ( .C1(n8444), .C2(n9809), .A(n8236), .B(n8235), .ZN(n8237)
         );
  OAI21_X1 U9741 ( .B1(n8447), .B2(n8412), .A(n8237), .ZN(P2_U3272) );
  XNOR2_X1 U9742 ( .A(n8238), .B(n8246), .ZN(n8452) );
  AOI21_X1 U9743 ( .B1(n8448), .B2(n8257), .A(n4557), .ZN(n8449) );
  INV_X1 U9744 ( .A(n8240), .ZN(n8241) );
  AOI22_X1 U9745 ( .A1(n9813), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8241), .B2(
        n9802), .ZN(n8242) );
  OAI21_X1 U9746 ( .B1(n8243), .B2(n8398), .A(n8242), .ZN(n8251) );
  AND2_X1 U9747 ( .A1(n8262), .A2(n8244), .ZN(n8247) );
  OAI21_X1 U9748 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8249) );
  AOI222_X1 U9749 ( .A1(n9771), .A2(n8249), .B1(n8283), .B2(n9778), .C1(n8248), 
        .C2(n9775), .ZN(n8451) );
  NOR2_X1 U9750 ( .A1(n8451), .A2(n9813), .ZN(n8250) );
  AOI211_X1 U9751 ( .C1(n8449), .C2(n9809), .A(n8251), .B(n8250), .ZN(n8252)
         );
  OAI21_X1 U9752 ( .B1(n8452), .B2(n8412), .A(n8252), .ZN(P2_U3273) );
  OAI21_X1 U9753 ( .B1(n8255), .B2(n8254), .A(n8253), .ZN(n8256) );
  INV_X1 U9754 ( .A(n8256), .ZN(n8457) );
  INV_X1 U9755 ( .A(n8275), .ZN(n8258) );
  AOI21_X1 U9756 ( .B1(n8453), .B2(n8258), .A(n4558), .ZN(n8454) );
  AOI22_X1 U9757 ( .A1(n9813), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8259), .B2(
        n9802), .ZN(n8260) );
  OAI21_X1 U9758 ( .B1(n8261), .B2(n8398), .A(n8260), .ZN(n8272) );
  INV_X1 U9759 ( .A(n8262), .ZN(n8266) );
  AOI21_X1 U9760 ( .B1(n8280), .B2(n8264), .A(n8263), .ZN(n8265) );
  NOR3_X1 U9761 ( .A1(n8266), .A2(n8265), .A3(n9795), .ZN(n8270) );
  OAI22_X1 U9762 ( .A1(n8268), .A2(n8404), .B1(n8267), .B2(n8402), .ZN(n8269)
         );
  NOR2_X1 U9763 ( .A1(n8270), .A2(n8269), .ZN(n8456) );
  NOR2_X1 U9764 ( .A1(n8456), .A2(n9813), .ZN(n8271) );
  AOI211_X1 U9765 ( .C1(n8454), .C2(n9809), .A(n8272), .B(n8271), .ZN(n8273)
         );
  OAI21_X1 U9766 ( .B1(n8457), .B2(n8412), .A(n8273), .ZN(P2_U3274) );
  XOR2_X1 U9767 ( .A(n8281), .B(n8274), .Z(n8462) );
  INV_X1 U9768 ( .A(n8290), .ZN(n8276) );
  AOI21_X1 U9769 ( .B1(n8458), .B2(n8276), .A(n8275), .ZN(n8459) );
  AOI22_X1 U9770 ( .A1(n9813), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8277), .B2(
        n9802), .ZN(n8278) );
  OAI21_X1 U9771 ( .B1(n8279), .B2(n8398), .A(n8278), .ZN(n8286) );
  OAI21_X1 U9772 ( .B1(n4282), .B2(n8281), .A(n8280), .ZN(n8284) );
  AOI222_X1 U9773 ( .A1(n9771), .A2(n8284), .B1(n8283), .B2(n9775), .C1(n8282), 
        .C2(n9778), .ZN(n8461) );
  NOR2_X1 U9774 ( .A1(n8461), .A2(n9813), .ZN(n8285) );
  AOI211_X1 U9775 ( .C1(n8459), .C2(n9809), .A(n8286), .B(n8285), .ZN(n8287)
         );
  OAI21_X1 U9776 ( .B1(n8412), .B2(n8462), .A(n8287), .ZN(P2_U3275) );
  OAI21_X1 U9777 ( .B1(n8289), .B2(n8295), .A(n8288), .ZN(n8467) );
  AOI21_X1 U9778 ( .B1(n8463), .B2(n8309), .A(n8290), .ZN(n8464) );
  AOI22_X1 U9779 ( .A1(n9813), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8291), .B2(
        n9802), .ZN(n8292) );
  OAI21_X1 U9780 ( .B1(n8293), .B2(n8398), .A(n8292), .ZN(n8300) );
  NOR2_X1 U9781 ( .A1(n4284), .A2(n8294), .ZN(n8296) );
  XNOR2_X1 U9782 ( .A(n8296), .B(n8295), .ZN(n8298) );
  AOI222_X1 U9783 ( .A1(n9771), .A2(n8298), .B1(n8297), .B2(n9775), .C1(n8327), 
        .C2(n9778), .ZN(n8466) );
  NOR2_X1 U9784 ( .A1(n8466), .A2(n9813), .ZN(n8299) );
  AOI211_X1 U9785 ( .C1(n8464), .C2(n9809), .A(n8300), .B(n8299), .ZN(n8301)
         );
  OAI21_X1 U9786 ( .B1(n8412), .B2(n8467), .A(n8301), .ZN(P2_U3276) );
  OAI21_X1 U9787 ( .B1(n8303), .B2(n8305), .A(n8302), .ZN(n8472) );
  AOI22_X1 U9788 ( .A1(n8470), .A2(n9803), .B1(n9813), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8316) );
  AOI21_X1 U9789 ( .B1(n8305), .B2(n8304), .A(n4284), .ZN(n8306) );
  OAI222_X1 U9790 ( .A1(n8404), .A2(n8308), .B1(n8402), .B2(n8307), .C1(n9795), 
        .C2(n8306), .ZN(n8468) );
  INV_X1 U9791 ( .A(n8309), .ZN(n8310) );
  AOI211_X1 U9792 ( .C1(n8470), .C2(n8318), .A(n9865), .B(n8310), .ZN(n8469)
         );
  INV_X1 U9793 ( .A(n8469), .ZN(n8313) );
  INV_X1 U9794 ( .A(n8311), .ZN(n8312) );
  OAI22_X1 U9795 ( .A1(n8313), .A2(n4643), .B1(n9788), .B2(n8312), .ZN(n8314)
         );
  OAI21_X1 U9796 ( .B1(n8468), .B2(n8314), .A(n9783), .ZN(n8315) );
  OAI211_X1 U9797 ( .C1(n8472), .C2(n8412), .A(n8316), .B(n8315), .ZN(P2_U3277) );
  XNOR2_X1 U9798 ( .A(n8317), .B(n8325), .ZN(n8477) );
  INV_X1 U9799 ( .A(n8342), .ZN(n8320) );
  INV_X1 U9800 ( .A(n8318), .ZN(n8319) );
  AOI21_X1 U9801 ( .B1(n8473), .B2(n8320), .A(n8319), .ZN(n8474) );
  AOI22_X1 U9802 ( .A1(n9813), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8321), .B2(
        n9802), .ZN(n8322) );
  OAI21_X1 U9803 ( .B1(n8323), .B2(n8398), .A(n8322), .ZN(n8330) );
  XNOR2_X1 U9804 ( .A(n8324), .B(n8325), .ZN(n8328) );
  AOI222_X1 U9805 ( .A1(n9771), .A2(n8328), .B1(n8327), .B2(n9775), .C1(n8326), 
        .C2(n9778), .ZN(n8476) );
  NOR2_X1 U9806 ( .A1(n8476), .A2(n9813), .ZN(n8329) );
  AOI211_X1 U9807 ( .C1(n8474), .C2(n9809), .A(n8330), .B(n8329), .ZN(n8331)
         );
  OAI21_X1 U9808 ( .B1(n8477), .B2(n8412), .A(n8331), .ZN(P2_U3278) );
  OAI21_X1 U9809 ( .B1(n4330), .B2(n8335), .A(n8332), .ZN(n8333) );
  INV_X1 U9810 ( .A(n8333), .ZN(n8482) );
  NAND3_X1 U9811 ( .A1(n8336), .A2(n8335), .A3(n8334), .ZN(n8337) );
  NAND2_X1 U9812 ( .A1(n8337), .A2(n9771), .ZN(n8340) );
  AOI22_X1 U9813 ( .A1(n8385), .A2(n9778), .B1(n9775), .B2(n8338), .ZN(n8339)
         );
  OAI21_X1 U9814 ( .B1(n8341), .B2(n8340), .A(n8339), .ZN(n8478) );
  INV_X1 U9815 ( .A(n8364), .ZN(n8343) );
  AOI211_X1 U9816 ( .C1(n8480), .C2(n8343), .A(n9865), .B(n8342), .ZN(n8479)
         );
  NAND2_X1 U9817 ( .A1(n8479), .A2(n8344), .ZN(n8347) );
  AOI22_X1 U9818 ( .A1(n9813), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8345), .B2(
        n9802), .ZN(n8346) );
  OAI211_X1 U9819 ( .C1(n8348), .C2(n8398), .A(n8347), .B(n8346), .ZN(n8349)
         );
  AOI21_X1 U9820 ( .B1(n8478), .B2(n9783), .A(n8349), .ZN(n8350) );
  OAI21_X1 U9821 ( .B1(n8482), .B2(n8412), .A(n8350), .ZN(P2_U3279) );
  AND2_X1 U9822 ( .A1(n8351), .A2(n8356), .ZN(n8352) );
  OR2_X1 U9823 ( .A1(n8353), .A2(n8352), .ZN(n8363) );
  OR2_X1 U9824 ( .A1(n8363), .A2(n9790), .ZN(n8362) );
  AND2_X1 U9825 ( .A1(n8355), .A2(n8354), .ZN(n8357) );
  XNOR2_X1 U9826 ( .A(n8357), .B(n4834), .ZN(n8360) );
  OAI22_X1 U9827 ( .A1(n8405), .A2(n8402), .B1(n8358), .B2(n8404), .ZN(n8359)
         );
  AOI21_X1 U9828 ( .B1(n8360), .B2(n9771), .A(n8359), .ZN(n8361) );
  INV_X1 U9829 ( .A(n8363), .ZN(n8487) );
  AND2_X1 U9830 ( .A1(n4337), .A2(n8483), .ZN(n8365) );
  OR2_X1 U9831 ( .A1(n8365), .A2(n8364), .ZN(n8485) );
  AOI22_X1 U9832 ( .A1(n9813), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8366), .B2(
        n9802), .ZN(n8368) );
  NAND2_X1 U9833 ( .A1(n8483), .A2(n9803), .ZN(n8367) );
  OAI211_X1 U9834 ( .C1(n8485), .C2(n8369), .A(n8368), .B(n8367), .ZN(n8370)
         );
  AOI21_X1 U9835 ( .B1(n8487), .B2(n9810), .A(n8370), .ZN(n8371) );
  OAI21_X1 U9836 ( .B1(n8488), .B2(n9813), .A(n8371), .ZN(P2_U3280) );
  OAI21_X1 U9837 ( .B1(n8374), .B2(n8373), .A(n8372), .ZN(n8375) );
  INV_X1 U9838 ( .A(n8375), .ZN(n8494) );
  INV_X1 U9839 ( .A(n4337), .ZN(n8376) );
  AOI21_X1 U9840 ( .B1(n8490), .B2(n8393), .A(n8376), .ZN(n8491) );
  AOI22_X1 U9841 ( .A1(n9813), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8377), .B2(
        n9802), .ZN(n8378) );
  OAI21_X1 U9842 ( .B1(n8379), .B2(n8398), .A(n8378), .ZN(n8389) );
  NAND2_X1 U9843 ( .A1(n8407), .A2(n8380), .ZN(n8383) );
  NAND2_X1 U9844 ( .A1(n8383), .A2(n8382), .ZN(n8381) );
  OAI211_X1 U9845 ( .C1(n8383), .C2(n8382), .A(n8381), .B(n9771), .ZN(n8387)
         );
  AOI22_X1 U9846 ( .A1(n8385), .A2(n9775), .B1(n9778), .B2(n8384), .ZN(n8386)
         );
  AND2_X1 U9847 ( .A1(n8387), .A2(n8386), .ZN(n8493) );
  NOR2_X1 U9848 ( .A1(n8493), .A2(n9813), .ZN(n8388) );
  AOI211_X1 U9849 ( .C1(n8491), .C2(n9809), .A(n8389), .B(n8388), .ZN(n8390)
         );
  OAI21_X1 U9850 ( .B1(n8494), .B2(n8412), .A(n8390), .ZN(P2_U3281) );
  XNOR2_X1 U9851 ( .A(n8391), .B(n8400), .ZN(n8499) );
  INV_X1 U9852 ( .A(n8392), .ZN(n8395) );
  INV_X1 U9853 ( .A(n8393), .ZN(n8394) );
  AOI21_X1 U9854 ( .B1(n8495), .B2(n8395), .A(n8394), .ZN(n8496) );
  AOI22_X1 U9855 ( .A1(n9813), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8396), .B2(
        n9802), .ZN(n8397) );
  OAI21_X1 U9856 ( .B1(n8399), .B2(n8398), .A(n8397), .ZN(n8410) );
  AOI21_X1 U9857 ( .B1(n8401), .B2(n8400), .A(n9795), .ZN(n8408) );
  OAI22_X1 U9858 ( .A1(n8405), .A2(n8404), .B1(n8403), .B2(n8402), .ZN(n8406)
         );
  AOI21_X1 U9859 ( .B1(n8408), .B2(n8407), .A(n8406), .ZN(n8498) );
  NOR2_X1 U9860 ( .A1(n8498), .A2(n9813), .ZN(n8409) );
  AOI211_X1 U9861 ( .C1(n8496), .C2(n9809), .A(n8410), .B(n8409), .ZN(n8411)
         );
  OAI21_X1 U9862 ( .B1(n8499), .B2(n8412), .A(n8411), .ZN(P2_U3282) );
  AOI21_X1 U9863 ( .B1(n7362), .B2(n9876), .A(n8415), .ZN(n8413) );
  OAI21_X1 U9864 ( .B1(n8414), .B2(n9865), .A(n8413), .ZN(n8512) );
  MUX2_X1 U9865 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8512), .S(n9889), .Z(
        P2_U3551) );
  AOI21_X1 U9866 ( .B1(n8416), .B2(n9876), .A(n8415), .ZN(n8417) );
  OAI21_X1 U9867 ( .B1(n8418), .B2(n9865), .A(n8417), .ZN(n8513) );
  MUX2_X1 U9868 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8513), .S(n9889), .Z(
        P2_U3550) );
  AOI21_X1 U9869 ( .B1(n8424), .B2(n9876), .A(n8423), .ZN(n8425) );
  OAI211_X1 U9870 ( .C1(n8427), .C2(n9829), .A(n8426), .B(n8425), .ZN(n8514)
         );
  MUX2_X1 U9871 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8514), .S(n9889), .Z(
        P2_U3548) );
  AOI22_X1 U9872 ( .A1(n8429), .A2(n9878), .B1(n8428), .B2(n9876), .ZN(n8430)
         );
  OAI211_X1 U9873 ( .C1(n8432), .C2(n9829), .A(n8431), .B(n8430), .ZN(n8515)
         );
  MUX2_X1 U9874 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8515), .S(n9889), .Z(
        P2_U3547) );
  AOI21_X1 U9875 ( .B1(n8434), .B2(n9876), .A(n8433), .ZN(n8435) );
  OAI211_X1 U9876 ( .C1(n8437), .C2(n9829), .A(n8436), .B(n8435), .ZN(n8516)
         );
  MUX2_X1 U9877 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8516), .S(n9889), .Z(
        P2_U3546) );
  AOI211_X1 U9878 ( .C1(n8440), .C2(n9876), .A(n8439), .B(n8438), .ZN(n8441)
         );
  OAI21_X1 U9879 ( .B1(n8442), .B2(n9829), .A(n8441), .ZN(n8517) );
  MUX2_X1 U9880 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8517), .S(n9889), .Z(
        P2_U3545) );
  AOI22_X1 U9881 ( .A1(n8444), .A2(n9878), .B1(n8443), .B2(n9876), .ZN(n8445)
         );
  OAI211_X1 U9882 ( .C1(n8447), .C2(n9829), .A(n8446), .B(n8445), .ZN(n8518)
         );
  MUX2_X1 U9883 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8518), .S(n9889), .Z(
        P2_U3544) );
  AOI22_X1 U9884 ( .A1(n8449), .A2(n9878), .B1(n8448), .B2(n9876), .ZN(n8450)
         );
  OAI211_X1 U9885 ( .C1(n8452), .C2(n9829), .A(n8451), .B(n8450), .ZN(n8519)
         );
  MUX2_X1 U9886 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8519), .S(n9889), .Z(
        P2_U3543) );
  AOI22_X1 U9887 ( .A1(n8454), .A2(n9878), .B1(n8453), .B2(n9876), .ZN(n8455)
         );
  OAI211_X1 U9888 ( .C1(n8457), .C2(n9829), .A(n8456), .B(n8455), .ZN(n8520)
         );
  MUX2_X1 U9889 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8520), .S(n9889), .Z(
        P2_U3542) );
  AOI22_X1 U9890 ( .A1(n8459), .A2(n9878), .B1(n8458), .B2(n9876), .ZN(n8460)
         );
  OAI211_X1 U9891 ( .C1(n8462), .C2(n9829), .A(n8461), .B(n8460), .ZN(n8521)
         );
  MUX2_X1 U9892 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8521), .S(n9889), .Z(
        P2_U3541) );
  AOI22_X1 U9893 ( .A1(n8464), .A2(n9878), .B1(n8463), .B2(n9876), .ZN(n8465)
         );
  OAI211_X1 U9894 ( .C1(n8467), .C2(n9829), .A(n8466), .B(n8465), .ZN(n8522)
         );
  MUX2_X1 U9895 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8522), .S(n9889), .Z(
        P2_U3540) );
  AOI211_X1 U9896 ( .C1(n8470), .C2(n9876), .A(n8469), .B(n8468), .ZN(n8471)
         );
  OAI21_X1 U9897 ( .B1(n9829), .B2(n8472), .A(n8471), .ZN(n8523) );
  MUX2_X1 U9898 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8523), .S(n9889), .Z(
        P2_U3539) );
  AOI22_X1 U9899 ( .A1(n8474), .A2(n9878), .B1(n8473), .B2(n9876), .ZN(n8475)
         );
  OAI211_X1 U9900 ( .C1(n8477), .C2(n9829), .A(n8476), .B(n8475), .ZN(n8524)
         );
  MUX2_X1 U9901 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8524), .S(n9889), .Z(
        P2_U3538) );
  AOI211_X1 U9902 ( .C1(n8480), .C2(n9876), .A(n8479), .B(n8478), .ZN(n8481)
         );
  OAI21_X1 U9903 ( .B1(n8482), .B2(n9829), .A(n8481), .ZN(n8525) );
  MUX2_X1 U9904 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8525), .S(n9889), .Z(
        P2_U3537) );
  INV_X1 U9905 ( .A(n8511), .ZN(n9860) );
  INV_X1 U9906 ( .A(n8483), .ZN(n8484) );
  OAI22_X1 U9907 ( .A1(n8485), .A2(n9865), .B1(n8484), .B2(n9863), .ZN(n8486)
         );
  AOI21_X1 U9908 ( .B1(n8487), .B2(n9860), .A(n8486), .ZN(n8489) );
  NAND2_X1 U9909 ( .A1(n8489), .A2(n8488), .ZN(n8526) );
  MUX2_X1 U9910 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8526), .S(n9889), .Z(
        P2_U3536) );
  AOI22_X1 U9911 ( .A1(n8491), .A2(n9878), .B1(n8490), .B2(n9876), .ZN(n8492)
         );
  OAI211_X1 U9912 ( .C1(n8494), .C2(n9829), .A(n8493), .B(n8492), .ZN(n8527)
         );
  MUX2_X1 U9913 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8527), .S(n9889), .Z(
        P2_U3535) );
  AOI22_X1 U9914 ( .A1(n8496), .A2(n9878), .B1(n8495), .B2(n9876), .ZN(n8497)
         );
  OAI211_X1 U9915 ( .C1(n8499), .C2(n9829), .A(n8498), .B(n8497), .ZN(n8528)
         );
  MUX2_X1 U9916 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8528), .S(n9889), .Z(
        P2_U3534) );
  AOI21_X1 U9917 ( .B1(n8501), .B2(n9876), .A(n8500), .ZN(n8502) );
  OAI211_X1 U9918 ( .C1(n8504), .C2(n9829), .A(n8503), .B(n8502), .ZN(n8529)
         );
  MUX2_X1 U9919 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8529), .S(n9889), .Z(
        P2_U3532) );
  INV_X1 U9920 ( .A(n8505), .ZN(n8509) );
  AOI22_X1 U9921 ( .A1(n8507), .A2(n9878), .B1(n8506), .B2(n9876), .ZN(n8508)
         );
  OAI211_X1 U9922 ( .C1(n8511), .C2(n8510), .A(n8509), .B(n8508), .ZN(n8530)
         );
  MUX2_X1 U9923 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8530), .S(n9889), .Z(
        P2_U3530) );
  MUX2_X1 U9924 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8512), .S(n10073), .Z(
        P2_U3519) );
  MUX2_X1 U9925 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8513), .S(n10073), .Z(
        P2_U3518) );
  MUX2_X1 U9926 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8514), .S(n10073), .Z(
        P2_U3516) );
  MUX2_X1 U9927 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8515), .S(n10073), .Z(
        P2_U3515) );
  MUX2_X1 U9928 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8516), .S(n10073), .Z(
        P2_U3514) );
  MUX2_X1 U9929 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8517), .S(n10073), .Z(
        P2_U3513) );
  MUX2_X1 U9930 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8518), .S(n10073), .Z(
        P2_U3512) );
  MUX2_X1 U9931 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8519), .S(n10073), .Z(
        P2_U3511) );
  MUX2_X1 U9932 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8520), .S(n10073), .Z(
        P2_U3510) );
  MUX2_X1 U9933 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8521), .S(n10073), .Z(
        P2_U3509) );
  MUX2_X1 U9934 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8522), .S(n10073), .Z(
        P2_U3508) );
  MUX2_X1 U9935 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8523), .S(n10073), .Z(
        P2_U3507) );
  MUX2_X1 U9936 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8524), .S(n10073), .Z(
        P2_U3505) );
  MUX2_X1 U9937 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8525), .S(n10073), .Z(
        P2_U3502) );
  MUX2_X1 U9938 ( .A(n8526), .B(P2_REG0_REG_16__SCAN_IN), .S(n10071), .Z(
        P2_U3499) );
  MUX2_X1 U9939 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8527), .S(n10073), .Z(
        P2_U3496) );
  MUX2_X1 U9940 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8528), .S(n10073), .Z(
        P2_U3493) );
  MUX2_X1 U9941 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8529), .S(n10073), .Z(
        P2_U3487) );
  MUX2_X1 U9942 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n8530), .S(n10073), .Z(
        P2_U3481) );
  INV_X1 U9943 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8532) );
  NAND3_X1 U9944 ( .A1(n8532), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8534) );
  OAI22_X1 U9945 ( .A1(n8535), .A2(n8534), .B1(n5137), .B2(n8533), .ZN(n8536)
         );
  AOI21_X1 U9946 ( .B1(n8531), .B2(n8537), .A(n8536), .ZN(n8538) );
  INV_X1 U9947 ( .A(n8538), .ZN(P2_U3327) );
  OAI222_X1 U9948 ( .A1(n8543), .A2(n8542), .B1(P2_U3152), .B2(n8541), .C1(
        n8540), .C2(n8539), .ZN(P2_U3329) );
  MUX2_X1 U9949 ( .A(n8544), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U9950 ( .A(n8545), .ZN(n8547) );
  XNOR2_X1 U9951 ( .A(n8547), .B(n8546), .ZN(n8548) );
  XNOR2_X1 U9952 ( .A(n8549), .B(n8548), .ZN(n8554) );
  AOI22_X1 U9953 ( .A1(n9186), .A2(n8668), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        n4258), .ZN(n8551) );
  NAND2_X1 U9954 ( .A1(n9159), .A2(n8618), .ZN(n8550) );
  OAI211_X1 U9955 ( .C1(n9157), .C2(n8666), .A(n8551), .B(n8550), .ZN(n8552)
         );
  AOI21_X1 U9956 ( .B1(n9397), .B2(n8679), .A(n8552), .ZN(n8553) );
  OAI21_X1 U9957 ( .B1(n8554), .B2(n8664), .A(n8553), .ZN(P1_U3212) );
  INV_X1 U9958 ( .A(n8555), .ZN(n8557) );
  NOR2_X1 U9959 ( .A1(n8557), .A2(n8556), .ZN(n8559) );
  XNOR2_X1 U9960 ( .A(n8559), .B(n8558), .ZN(n8564) );
  AOI22_X1 U9961 ( .A1(n9251), .A2(n8668), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        n4258), .ZN(n8561) );
  NAND2_X1 U9962 ( .A1(n9221), .A2(n8659), .ZN(n8560) );
  OAI211_X1 U9963 ( .C1(n8671), .C2(n9223), .A(n8561), .B(n8560), .ZN(n8562)
         );
  AOI21_X1 U9964 ( .B1(n9415), .B2(n8679), .A(n8562), .ZN(n8563) );
  OAI21_X1 U9965 ( .B1(n8564), .B2(n8664), .A(n8563), .ZN(P1_U3214) );
  INV_X1 U9966 ( .A(n9436), .ZN(n9291) );
  INV_X1 U9967 ( .A(n8623), .ZN(n8567) );
  NOR3_X1 U9968 ( .A1(n8642), .A2(n8646), .A3(n8565), .ZN(n8566) );
  OAI21_X1 U9969 ( .B1(n8567), .B2(n8566), .A(n8647), .ZN(n8571) );
  INV_X1 U9970 ( .A(n9250), .ZN(n9283) );
  NAND2_X1 U9971 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9067) );
  OAI21_X1 U9972 ( .B1(n8666), .B2(n9283), .A(n9067), .ZN(n8569) );
  NOR2_X1 U9973 ( .A1(n8671), .A2(n9286), .ZN(n8568) );
  AOI211_X1 U9974 ( .C1(n8668), .C2(n9330), .A(n8569), .B(n8568), .ZN(n8570)
         );
  OAI211_X1 U9975 ( .C1(n9291), .C2(n8653), .A(n8571), .B(n8570), .ZN(P1_U3217) );
  AOI21_X1 U9976 ( .B1(n8573), .B2(n8572), .A(n4306), .ZN(n8579) );
  OAI22_X1 U9977 ( .A1(n9088), .A2(n8666), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8574), .ZN(n8575) );
  AOI21_X1 U9978 ( .B1(n8668), .B2(n9250), .A(n8575), .ZN(n8576) );
  OAI21_X1 U9979 ( .B1(n8671), .B2(n9258), .A(n8576), .ZN(n8577) );
  AOI21_X1 U9980 ( .B1(n9426), .B2(n8679), .A(n8577), .ZN(n8578) );
  OAI21_X1 U9981 ( .B1(n8579), .B2(n8664), .A(n8578), .ZN(P1_U3221) );
  INV_X1 U9982 ( .A(n8580), .ZN(n8589) );
  NAND2_X1 U9983 ( .A1(n9094), .A2(n9456), .ZN(n9407) );
  OAI21_X1 U9984 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8584) );
  NAND2_X1 U9985 ( .A1(n8584), .A2(n8647), .ZN(n8588) );
  AOI22_X1 U9986 ( .A1(n9221), .A2(n8668), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8585) );
  OAI21_X1 U9987 ( .B1(n9095), .B2(n8666), .A(n8585), .ZN(n8586) );
  AOI21_X1 U9988 ( .B1(n9192), .B2(n8618), .A(n8586), .ZN(n8587) );
  OAI211_X1 U9989 ( .C1(n8589), .C2(n9407), .A(n8588), .B(n8587), .ZN(P1_U3223) );
  INV_X1 U9990 ( .A(n8590), .ZN(n8594) );
  AOI21_X1 U9991 ( .B1(n8591), .B2(n8675), .A(n8592), .ZN(n8593) );
  OAI21_X1 U9992 ( .B1(n8594), .B2(n8593), .A(n8647), .ZN(n8602) );
  INV_X1 U9993 ( .A(n9353), .ZN(n8600) );
  INV_X1 U9994 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8595) );
  NOR2_X1 U9995 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8595), .ZN(n9598) );
  AOI21_X1 U9996 ( .B1(n8659), .B2(n9302), .A(n9598), .ZN(n8596) );
  OAI21_X1 U9997 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8599) );
  AOI21_X1 U9998 ( .B1(n8600), .B2(n8618), .A(n8599), .ZN(n8601) );
  OAI211_X1 U9999 ( .C1(n4613), .C2(n8653), .A(n8602), .B(n8601), .ZN(P1_U3224) );
  INV_X1 U10000 ( .A(n9448), .ZN(n9322) );
  OAI21_X1 U10001 ( .B1(n8605), .B2(n8604), .A(n8603), .ZN(n8606) );
  NAND2_X1 U10002 ( .A1(n8606), .A2(n8647), .ZN(n8610) );
  INV_X1 U10003 ( .A(n9330), .ZN(n9281) );
  NAND2_X1 U10004 ( .A1(n4258), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9611) );
  OAI21_X1 U10005 ( .B1(n8666), .B2(n9281), .A(n9611), .ZN(n8608) );
  NOR2_X1 U10006 ( .A1(n8671), .A2(n9319), .ZN(n8607) );
  AOI211_X1 U10007 ( .C1(n8668), .C2(n9328), .A(n8608), .B(n8607), .ZN(n8609)
         );
  OAI211_X1 U10008 ( .C1(n9322), .C2(n8653), .A(n8610), .B(n8609), .ZN(
        P1_U3226) );
  INV_X1 U10009 ( .A(n9411), .ZN(n9203) );
  OAI21_X1 U10010 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8614) );
  NAND2_X1 U10011 ( .A1(n8614), .A2(n8647), .ZN(n8620) );
  INV_X1 U10012 ( .A(n8615), .ZN(n9201) );
  AOI22_X1 U10013 ( .A1(n9234), .A2(n8668), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        n4258), .ZN(n8616) );
  OAI21_X1 U10014 ( .B1(n9173), .B2(n8666), .A(n8616), .ZN(n8617) );
  AOI21_X1 U10015 ( .B1(n9201), .B2(n8618), .A(n8617), .ZN(n8619) );
  OAI211_X1 U10016 ( .C1(n9203), .C2(n8653), .A(n8620), .B(n8619), .ZN(
        P1_U3227) );
  AND3_X1 U10017 ( .A1(n8623), .A2(n8622), .A3(n8621), .ZN(n8624) );
  OAI21_X1 U10018 ( .B1(n8625), .B2(n8624), .A(n8647), .ZN(n8630) );
  AOI22_X1 U10019 ( .A1(n9271), .A2(n8659), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8627) );
  NAND2_X1 U10020 ( .A1(n8668), .A2(n9303), .ZN(n8626) );
  OAI211_X1 U10021 ( .C1(n8671), .C2(n9265), .A(n8627), .B(n8626), .ZN(n8628)
         );
  AOI21_X1 U10022 ( .B1(n9430), .B2(n8679), .A(n8628), .ZN(n8629) );
  NAND2_X1 U10023 ( .A1(n8630), .A2(n8629), .ZN(P1_U3231) );
  NAND2_X1 U10024 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  XOR2_X1 U10025 ( .A(n8634), .B(n8633), .Z(n8641) );
  OAI22_X1 U10026 ( .A1(n9090), .A2(n8666), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8635), .ZN(n8636) );
  AOI21_X1 U10027 ( .B1(n8668), .B2(n9271), .A(n8636), .ZN(n8637) );
  OAI21_X1 U10028 ( .B1(n8671), .B2(n8638), .A(n8637), .ZN(n8639) );
  AOI21_X1 U10029 ( .B1(n9420), .B2(n8679), .A(n8639), .ZN(n8640) );
  OAI21_X1 U10030 ( .B1(n8641), .B2(n8664), .A(n8640), .ZN(P1_U3233) );
  INV_X1 U10031 ( .A(n9311), .ZN(n9442) );
  OAI21_X1 U10032 ( .B1(n8644), .B2(n8646), .A(n8643), .ZN(n8645) );
  OAI21_X1 U10033 ( .B1(n4858), .B2(n8646), .A(n8645), .ZN(n8648) );
  NAND2_X1 U10034 ( .A1(n8648), .A2(n8647), .ZN(n8652) );
  INV_X1 U10035 ( .A(n9303), .ZN(n9085) );
  NAND2_X1 U10036 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9629) );
  OAI21_X1 U10037 ( .B1(n8666), .B2(n9085), .A(n9629), .ZN(n8650) );
  NOR2_X1 U10038 ( .A1(n8671), .A2(n9309), .ZN(n8649) );
  AOI211_X1 U10039 ( .C1(n8668), .C2(n9302), .A(n8650), .B(n8649), .ZN(n8651)
         );
  OAI211_X1 U10040 ( .C1(n9442), .C2(n8653), .A(n8652), .B(n8651), .ZN(
        P1_U3236) );
  INV_X1 U10041 ( .A(n8655), .ZN(n8657) );
  NAND2_X1 U10042 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  XNOR2_X1 U10043 ( .A(n8654), .B(n8658), .ZN(n8665) );
  NAND2_X1 U10044 ( .A1(n9097), .A2(n8659), .ZN(n8661) );
  AOI22_X1 U10045 ( .A1(n9207), .A2(n8668), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8660) );
  OAI211_X1 U10046 ( .C1(n8671), .C2(n9177), .A(n8661), .B(n8660), .ZN(n8662)
         );
  AOI21_X1 U10047 ( .B1(n9402), .B2(n8679), .A(n8662), .ZN(n8663) );
  OAI21_X1 U10048 ( .B1(n8665), .B2(n8664), .A(n8663), .ZN(P1_U3238) );
  AND2_X1 U10049 ( .A1(n4258), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9587) );
  INV_X1 U10050 ( .A(n9328), .ZN(n8708) );
  NOR2_X1 U10051 ( .A1(n8666), .A2(n8708), .ZN(n8667) );
  AOI211_X1 U10052 ( .C1(n8668), .C2(n8988), .A(n9587), .B(n8667), .ZN(n8669)
         );
  OAI21_X1 U10053 ( .B1(n8671), .B2(n8670), .A(n8669), .ZN(n8678) );
  INV_X1 U10054 ( .A(n8591), .ZN(n8676) );
  AOI21_X1 U10055 ( .B1(n8675), .B2(n8672), .A(n8673), .ZN(n8674) );
  AOI211_X1 U10056 ( .C1(n8676), .C2(n8675), .A(n8664), .B(n8674), .ZN(n8677)
         );
  AOI211_X1 U10057 ( .C1(n8679), .C2(n9506), .A(n8678), .B(n8677), .ZN(n8680)
         );
  INV_X1 U10058 ( .A(n8680), .ZN(P1_U3239) );
  NAND2_X1 U10059 ( .A1(n8681), .A2(n8760), .ZN(n8684) );
  OR2_X1 U10060 ( .A1(n8758), .A2(n8682), .ZN(n8683) );
  INV_X1 U10061 ( .A(n8987), .ZN(n9141) );
  NAND2_X1 U10062 ( .A1(n9389), .A2(n9141), .ZN(n8930) );
  INV_X1 U10063 ( .A(n8930), .ZN(n8755) );
  NAND2_X1 U10064 ( .A1(n9393), .A2(n9157), .ZN(n9117) );
  NAND2_X1 U10065 ( .A1(n9138), .A2(n9114), .ZN(n8685) );
  NAND3_X1 U10066 ( .A1(n9117), .A2(n8879), .A3(n8685), .ZN(n8921) );
  INV_X1 U10067 ( .A(n8921), .ZN(n8743) );
  NOR2_X1 U10068 ( .A1(n9231), .A2(n9251), .ZN(n9109) );
  INV_X1 U10069 ( .A(n9271), .ZN(n8686) );
  OR2_X1 U10070 ( .A1(n9426), .A2(n8686), .ZN(n8935) );
  AND2_X1 U10071 ( .A1(n9430), .A2(n9283), .ZN(n9107) );
  NAND2_X1 U10072 ( .A1(n8935), .A2(n9107), .ZN(n8687) );
  NAND2_X1 U10073 ( .A1(n9426), .A2(n8686), .ZN(n9108) );
  NAND2_X1 U10074 ( .A1(n8687), .A2(n9108), .ZN(n8688) );
  OR2_X1 U10075 ( .A1(n9109), .A2(n8688), .ZN(n8731) );
  NAND2_X1 U10076 ( .A1(n9311), .A2(n9281), .ZN(n9103) );
  INV_X1 U10077 ( .A(n9302), .ZN(n9346) );
  NAND2_X1 U10078 ( .A1(n9448), .A2(n9346), .ZN(n9102) );
  NAND2_X1 U10079 ( .A1(n9103), .A2(n9102), .ZN(n8841) );
  NAND2_X1 U10080 ( .A1(n9360), .A2(n8708), .ZN(n8938) );
  AND2_X1 U10081 ( .A1(n8938), .A2(n9337), .ZN(n9100) );
  NAND2_X1 U10082 ( .A1(n8690), .A2(n8689), .ZN(n8808) );
  NAND2_X1 U10083 ( .A1(n8808), .A2(n8691), .ZN(n8822) );
  INV_X1 U10084 ( .A(n8822), .ZN(n8696) );
  NAND2_X1 U10085 ( .A1(n8798), .A2(n8692), .ZN(n8819) );
  NAND2_X1 U10086 ( .A1(n8794), .A2(n8793), .ZN(n8693) );
  NAND2_X1 U10087 ( .A1(n8693), .A2(n8701), .ZN(n8805) );
  NAND3_X1 U10088 ( .A1(n8805), .A2(n8800), .A3(n8785), .ZN(n8694) );
  NOR2_X1 U10089 ( .A1(n8819), .A2(n8694), .ZN(n8695) );
  NAND3_X1 U10090 ( .A1(n9100), .A2(n8696), .A3(n8695), .ZN(n8711) );
  NAND2_X1 U10091 ( .A1(n8818), .A2(n8697), .ZN(n8698) );
  NAND2_X1 U10092 ( .A1(n8698), .A2(n8798), .ZN(n8699) );
  NAND2_X1 U10093 ( .A1(n8807), .A2(n8699), .ZN(n8816) );
  NAND2_X1 U10094 ( .A1(n4623), .A2(n8701), .ZN(n8796) );
  INV_X1 U10095 ( .A(n8702), .ZN(n8703) );
  OR2_X1 U10096 ( .A1(n8796), .A2(n8703), .ZN(n8801) );
  NAND2_X1 U10097 ( .A1(n8801), .A2(n8805), .ZN(n8704) );
  NOR2_X1 U10098 ( .A1(n8819), .A2(n8704), .ZN(n8705) );
  NOR2_X1 U10099 ( .A1(n8816), .A2(n8705), .ZN(n8706) );
  OAI21_X1 U10100 ( .B1(n8822), .B2(n8706), .A(n8814), .ZN(n8707) );
  NAND2_X1 U10101 ( .A1(n9100), .A2(n8707), .ZN(n8709) );
  OR2_X1 U10102 ( .A1(n9360), .A2(n8708), .ZN(n8939) );
  NAND2_X1 U10103 ( .A1(n8939), .A2(n9336), .ZN(n8833) );
  NAND2_X1 U10104 ( .A1(n8833), .A2(n8938), .ZN(n9101) );
  AND2_X1 U10105 ( .A1(n8709), .A2(n9101), .ZN(n8710) );
  OR2_X1 U10106 ( .A1(n8841), .A2(n8710), .ZN(n8714) );
  OAI21_X1 U10107 ( .B1(n8841), .B2(n8711), .A(n8714), .ZN(n8712) );
  NAND2_X1 U10108 ( .A1(n9436), .A2(n9085), .ZN(n9105) );
  NAND2_X1 U10109 ( .A1(n8712), .A2(n9105), .ZN(n8713) );
  NOR2_X1 U10110 ( .A1(n8731), .A2(n8713), .ZN(n8912) );
  INV_X1 U10111 ( .A(n8912), .ZN(n8736) );
  NAND2_X1 U10112 ( .A1(n8714), .A2(n8789), .ZN(n8913) );
  INV_X1 U10113 ( .A(n8715), .ZN(n8717) );
  NAND2_X1 U10114 ( .A1(n9002), .A2(n4598), .ZN(n8716) );
  NAND3_X1 U10115 ( .A1(n8717), .A2(n8968), .A3(n8716), .ZN(n8719) );
  NAND2_X1 U10116 ( .A1(n8719), .A2(n8718), .ZN(n8721) );
  OAI21_X1 U10117 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(n8723) );
  NAND2_X1 U10118 ( .A1(n8723), .A2(n8904), .ZN(n8729) );
  AND2_X1 U10119 ( .A1(n8774), .A2(n8724), .ZN(n8725) );
  NAND2_X1 U10120 ( .A1(n8728), .A2(n8725), .ZN(n8947) );
  INV_X1 U10121 ( .A(n8947), .ZN(n8910) );
  NAND2_X1 U10122 ( .A1(n8726), .A2(n8905), .ZN(n8727) );
  AOI22_X1 U10123 ( .A1(n8729), .A2(n8910), .B1(n8728), .B2(n8727), .ZN(n8730)
         );
  NOR2_X1 U10124 ( .A1(n8913), .A2(n8730), .ZN(n8735) );
  NAND2_X1 U10125 ( .A1(n9231), .A2(n9251), .ZN(n9110) );
  NAND2_X1 U10126 ( .A1(n8731), .A2(n9110), .ZN(n8855) );
  NAND2_X1 U10127 ( .A1(n9110), .A2(n8935), .ZN(n8858) );
  NAND2_X1 U10128 ( .A1(n9105), .A2(n9103), .ZN(n8846) );
  OR2_X1 U10129 ( .A1(n9311), .A2(n9281), .ZN(n8937) );
  OR2_X1 U10130 ( .A1(n9448), .A2(n9346), .ZN(n8836) );
  AND2_X1 U10131 ( .A1(n8937), .A2(n8836), .ZN(n8840) );
  NOR2_X1 U10132 ( .A1(n8846), .A2(n8840), .ZN(n8733) );
  NOR2_X1 U10133 ( .A1(n9430), .A2(n9283), .ZN(n9106) );
  OR2_X1 U10134 ( .A1(n9436), .A2(n9085), .ZN(n8936) );
  INV_X1 U10135 ( .A(n8936), .ZN(n8732) );
  OR2_X1 U10136 ( .A1(n9106), .A2(n8732), .ZN(n8848) );
  OR3_X1 U10137 ( .A1(n8858), .A2(n8733), .A3(n8848), .ZN(n8734) );
  NAND2_X1 U10138 ( .A1(n8855), .A2(n8734), .ZN(n8915) );
  OAI21_X1 U10139 ( .B1(n8736), .B2(n8735), .A(n8915), .ZN(n8737) );
  NAND2_X1 U10140 ( .A1(n9415), .A2(n9090), .ZN(n8863) );
  INV_X1 U10141 ( .A(n9221), .ZN(n9092) );
  OR2_X1 U10142 ( .A1(n9411), .A2(n9092), .ZN(n8933) );
  OR2_X1 U10143 ( .A1(n9415), .A2(n9090), .ZN(n9111) );
  AND2_X1 U10144 ( .A1(n8933), .A2(n9111), .ZN(n8916) );
  INV_X1 U10145 ( .A(n8916), .ZN(n8764) );
  AOI21_X1 U10146 ( .B1(n8737), .B2(n8863), .A(n8764), .ZN(n8741) );
  NAND2_X1 U10147 ( .A1(n9411), .A2(n9092), .ZN(n9184) );
  INV_X1 U10148 ( .A(n9113), .ZN(n8740) );
  OR2_X1 U10149 ( .A1(n9402), .A2(n9095), .ZN(n8738) );
  NAND2_X1 U10150 ( .A1(n9138), .A2(n9115), .ZN(n8918) );
  INV_X1 U10151 ( .A(n8918), .ZN(n8739) );
  OAI21_X1 U10152 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n8742) );
  NAND2_X1 U10153 ( .A1(n8931), .A2(n8881), .ZN(n8924) );
  AOI21_X1 U10154 ( .B1(n8743), .B2(n8742), .A(n8924), .ZN(n8754) );
  NAND2_X1 U10155 ( .A1(n8744), .A2(n8760), .ZN(n8747) );
  OR2_X1 U10156 ( .A1(n8758), .A2(n8745), .ZN(n8746) );
  INV_X1 U10157 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U10158 ( .A1(n8748), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8751) );
  INV_X1 U10159 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8749) );
  OR2_X1 U10160 ( .A1(n7783), .A2(n8749), .ZN(n8750) );
  OAI211_X1 U10161 ( .C1(n8753), .C2(n8752), .A(n8751), .B(n8750), .ZN(n9121)
         );
  INV_X1 U10162 ( .A(n9121), .ZN(n8756) );
  NOR2_X1 U10163 ( .A1(n9077), .A2(n8756), .ZN(n8965) );
  INV_X1 U10164 ( .A(n8965), .ZN(n8885) );
  OAI21_X1 U10165 ( .B1(n8755), .B2(n8754), .A(n8885), .ZN(n8757) );
  NAND2_X1 U10166 ( .A1(n9077), .A2(n8756), .ZN(n8963) );
  NAND2_X1 U10167 ( .A1(n8757), .A2(n8963), .ZN(n8762) );
  NOR2_X1 U10168 ( .A1(n8758), .A2(n10022), .ZN(n8759) );
  INV_X1 U10169 ( .A(n9379), .ZN(n8886) );
  INV_X1 U10170 ( .A(n9073), .ZN(n8892) );
  AND2_X1 U10171 ( .A1(n8886), .A2(n8892), .ZN(n8966) );
  INV_X1 U10172 ( .A(n8966), .ZN(n8761) );
  NAND2_X1 U10173 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  AND2_X1 U10174 ( .A1(n9379), .A2(n9073), .ZN(n8967) );
  INV_X1 U10175 ( .A(n8967), .ZN(n8897) );
  AND2_X1 U10176 ( .A1(n8763), .A2(n8897), .ZN(n8976) );
  NOR2_X1 U10177 ( .A1(n8976), .A2(n9256), .ZN(n8975) );
  NAND2_X1 U10178 ( .A1(n8764), .A2(n9184), .ZN(n8765) );
  NAND2_X1 U10179 ( .A1(n9166), .A2(n8765), .ZN(n8769) );
  INV_X1 U10180 ( .A(n8863), .ZN(n8766) );
  NAND2_X1 U10181 ( .A1(n8933), .A2(n8766), .ZN(n8767) );
  AND2_X1 U10182 ( .A1(n9113), .A2(n8767), .ZN(n8920) );
  INV_X1 U10183 ( .A(n8920), .ZN(n8768) );
  INV_X1 U10184 ( .A(n8884), .ZN(n8891) );
  MUX2_X1 U10185 ( .A(n8769), .B(n8768), .S(n8891), .Z(n8770) );
  INV_X1 U10186 ( .A(n8770), .ZN(n8867) );
  NAND2_X1 U10187 ( .A1(n8771), .A2(n8774), .ZN(n8772) );
  NAND2_X1 U10188 ( .A1(n8783), .A2(n8774), .ZN(n8903) );
  INV_X1 U10189 ( .A(n8903), .ZN(n8775) );
  NAND2_X1 U10190 ( .A1(n8782), .A2(n8775), .ZN(n8776) );
  NAND2_X1 U10191 ( .A1(n8776), .A2(n8781), .ZN(n8777) );
  NAND2_X1 U10192 ( .A1(n8777), .A2(n8891), .ZN(n8779) );
  NAND2_X1 U10193 ( .A1(n8779), .A2(n8778), .ZN(n8788) );
  NAND3_X1 U10194 ( .A1(n8788), .A2(n8908), .A3(n8789), .ZN(n8780) );
  NAND2_X1 U10195 ( .A1(n8780), .A2(n8785), .ZN(n8792) );
  NAND3_X1 U10196 ( .A1(n8782), .A2(n8905), .A3(n8781), .ZN(n8784) );
  NAND2_X1 U10197 ( .A1(n8784), .A2(n8783), .ZN(n8787) );
  NAND2_X1 U10198 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  NOR2_X1 U10199 ( .A1(n8804), .A2(n8801), .ZN(n8831) );
  AND2_X1 U10200 ( .A1(n8793), .A2(n8800), .ZN(n8795) );
  OAI211_X1 U10201 ( .C1(n8796), .C2(n8795), .A(n8884), .B(n8794), .ZN(n8797)
         );
  NOR2_X1 U10202 ( .A1(n8797), .A2(n8950), .ZN(n8799) );
  NAND2_X1 U10203 ( .A1(n8822), .A2(n8814), .ZN(n8815) );
  NAND4_X1 U10204 ( .A1(n8955), .A2(n8799), .A3(n8798), .A4(n8815), .ZN(n8830)
         );
  INV_X1 U10205 ( .A(n8800), .ZN(n8803) );
  INV_X1 U10206 ( .A(n8801), .ZN(n8802) );
  OAI21_X1 U10207 ( .B1(n8804), .B2(n8803), .A(n8802), .ZN(n8806) );
  NAND2_X1 U10208 ( .A1(n8806), .A2(n8805), .ZN(n8813) );
  NAND2_X1 U10209 ( .A1(n8814), .A2(n8807), .ZN(n8809) );
  NAND2_X1 U10210 ( .A1(n8809), .A2(n8808), .ZN(n8820) );
  NAND4_X1 U10211 ( .A1(n8820), .A2(n8891), .A3(n8810), .A4(n8818), .ZN(n8811)
         );
  NOR2_X1 U10212 ( .A1(n8823), .A2(n8811), .ZN(n8812) );
  NAND2_X1 U10213 ( .A1(n8813), .A2(n8812), .ZN(n8829) );
  INV_X1 U10214 ( .A(n9100), .ZN(n8827) );
  INV_X1 U10215 ( .A(n8814), .ZN(n8817) );
  OAI211_X1 U10216 ( .C1(n8817), .C2(n8816), .A(n8815), .B(n8884), .ZN(n8825)
         );
  AND2_X1 U10217 ( .A1(n8819), .A2(n8818), .ZN(n8821) );
  OAI211_X1 U10218 ( .C1(n8822), .C2(n8821), .A(n8820), .B(n8891), .ZN(n8824)
         );
  AOI21_X1 U10219 ( .B1(n8825), .B2(n8824), .A(n8823), .ZN(n8826) );
  AOI21_X1 U10220 ( .B1(n8827), .B2(n8891), .A(n8826), .ZN(n8828) );
  OAI211_X1 U10221 ( .C1(n8831), .C2(n8830), .A(n8829), .B(n8828), .ZN(n8832)
         );
  NAND2_X1 U10222 ( .A1(n8832), .A2(n8939), .ZN(n8835) );
  NAND2_X1 U10223 ( .A1(n8833), .A2(n8884), .ZN(n8834) );
  NAND2_X1 U10224 ( .A1(n8835), .A2(n8834), .ZN(n8839) );
  NAND2_X1 U10225 ( .A1(n8836), .A2(n9102), .ZN(n9324) );
  NOR2_X1 U10226 ( .A1(n8938), .A2(n8891), .ZN(n8837) );
  NOR2_X1 U10227 ( .A1(n9324), .A2(n8837), .ZN(n8838) );
  NAND2_X1 U10228 ( .A1(n8839), .A2(n8838), .ZN(n8845) );
  INV_X1 U10229 ( .A(n8840), .ZN(n8842) );
  MUX2_X1 U10230 ( .A(n8842), .B(n8841), .S(n8891), .Z(n8843) );
  INV_X1 U10231 ( .A(n8843), .ZN(n8844) );
  NAND2_X1 U10232 ( .A1(n8845), .A2(n8844), .ZN(n8851) );
  INV_X1 U10233 ( .A(n8846), .ZN(n8847) );
  NAND2_X1 U10234 ( .A1(n8851), .A2(n8847), .ZN(n8850) );
  INV_X1 U10235 ( .A(n8848), .ZN(n8849) );
  NAND2_X1 U10236 ( .A1(n8850), .A2(n8849), .ZN(n8854) );
  NAND3_X1 U10237 ( .A1(n8851), .A2(n8937), .A3(n8936), .ZN(n8852) );
  INV_X1 U10238 ( .A(n9107), .ZN(n9245) );
  NAND3_X1 U10239 ( .A1(n8852), .A2(n9245), .A3(n9105), .ZN(n8853) );
  OAI21_X1 U10240 ( .B1(n8857), .B2(n8858), .A(n8855), .ZN(n8862) );
  INV_X1 U10241 ( .A(n9106), .ZN(n8856) );
  NAND2_X1 U10242 ( .A1(n8857), .A2(n8856), .ZN(n8859) );
  AOI21_X1 U10243 ( .B1(n8859), .B2(n9108), .A(n8858), .ZN(n8860) );
  OAI21_X1 U10244 ( .B1(n8860), .B2(n9109), .A(n8933), .ZN(n8861) );
  MUX2_X1 U10245 ( .A(n8862), .B(n8861), .S(n8891), .Z(n8865) );
  NAND2_X1 U10246 ( .A1(n9220), .A2(n9184), .ZN(n8864) );
  OR2_X1 U10247 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  NAND2_X1 U10248 ( .A1(n8867), .A2(n8866), .ZN(n8877) );
  NAND2_X1 U10249 ( .A1(n8877), .A2(n9166), .ZN(n8868) );
  AOI21_X1 U10250 ( .B1(n8868), .B2(n9181), .A(n9186), .ZN(n8871) );
  NAND2_X1 U10251 ( .A1(n8877), .A2(n8932), .ZN(n8869) );
  AOI21_X1 U10252 ( .B1(n8869), .B2(n9095), .A(n9402), .ZN(n8870) );
  NAND2_X1 U10253 ( .A1(n9402), .A2(n9166), .ZN(n8872) );
  NAND2_X1 U10254 ( .A1(n8879), .A2(n8872), .ZN(n8875) );
  NAND2_X1 U10255 ( .A1(n8932), .A2(n9186), .ZN(n8873) );
  NAND2_X1 U10256 ( .A1(n9138), .A2(n8873), .ZN(n8874) );
  MUX2_X1 U10257 ( .A(n8875), .B(n8874), .S(n8884), .Z(n8876) );
  OAI21_X1 U10258 ( .B1(n8877), .B2(n9116), .A(n8876), .ZN(n8878) );
  MUX2_X1 U10259 ( .A(n8879), .B(n9138), .S(n8891), .Z(n8880) );
  MUX2_X1 U10260 ( .A(n9117), .B(n8881), .S(n8891), .Z(n8882) );
  NOR3_X1 U10261 ( .A1(n8898), .A2(n8987), .A3(n9389), .ZN(n8883) );
  AOI21_X1 U10262 ( .B1(n8987), .B2(n8884), .A(n8883), .ZN(n8902) );
  NAND2_X1 U10263 ( .A1(n8885), .A2(n9073), .ZN(n8887) );
  NAND2_X1 U10264 ( .A1(n8887), .A2(n8886), .ZN(n8928) );
  INV_X1 U10265 ( .A(n8928), .ZN(n8890) );
  INV_X1 U10266 ( .A(n8888), .ZN(n8889) );
  AND2_X1 U10267 ( .A1(n9389), .A2(n8891), .ZN(n8896) );
  NAND2_X1 U10268 ( .A1(n9077), .A2(n8892), .ZN(n8893) );
  AND2_X1 U10269 ( .A1(n8963), .A2(n8893), .ZN(n8923) );
  INV_X1 U10270 ( .A(n8923), .ZN(n8895) );
  NAND3_X1 U10271 ( .A1(n8923), .A2(n8898), .A3(n8987), .ZN(n8894) );
  OAI211_X1 U10272 ( .C1(n8896), .C2(n8895), .A(n8894), .B(n8928), .ZN(n8901)
         );
  NAND2_X1 U10273 ( .A1(n8897), .A2(n8968), .ZN(n8926) );
  INV_X1 U10274 ( .A(n8926), .ZN(n8900) );
  NAND4_X1 U10275 ( .A1(n8928), .A2(n8983), .A3(n9389), .A4(n8898), .ZN(n8899)
         );
  NAND3_X1 U10276 ( .A1(n8902), .A2(n8983), .A3(n8928), .ZN(n8973) );
  AOI21_X1 U10277 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8907) );
  NOR2_X1 U10278 ( .A1(n8907), .A2(n8906), .ZN(n8943) );
  INV_X1 U10279 ( .A(n8943), .ZN(n8909) );
  AOI22_X1 U10280 ( .A1(n8911), .A2(n8910), .B1(n8909), .B2(n8908), .ZN(n8914)
         );
  OAI21_X1 U10281 ( .B1(n8914), .B2(n8913), .A(n8912), .ZN(n8917) );
  NAND3_X1 U10282 ( .A1(n8917), .A2(n8916), .A3(n8915), .ZN(n8919) );
  AOI21_X1 U10283 ( .B1(n8920), .B2(n8919), .A(n8918), .ZN(n8922) );
  NOR2_X1 U10284 ( .A1(n8922), .A2(n8921), .ZN(n8925) );
  OAI211_X1 U10285 ( .C1(n8925), .C2(n8924), .A(n8923), .B(n8930), .ZN(n8927)
         );
  AOI21_X1 U10286 ( .B1(n8928), .B2(n8927), .A(n8926), .ZN(n8929) );
  NOR2_X1 U10287 ( .A1(n8929), .A2(n5586), .ZN(n8971) );
  XNOR2_X1 U10288 ( .A(n9402), .B(n9095), .ZN(n9168) );
  INV_X1 U10289 ( .A(n9110), .ZN(n8934) );
  NOR2_X1 U10290 ( .A1(n9109), .A2(n8934), .ZN(n9232) );
  INV_X1 U10291 ( .A(n9243), .ZN(n9246) );
  OR2_X1 U10292 ( .A1(n9106), .A2(n9107), .ZN(n9269) );
  NAND2_X1 U10293 ( .A1(n8936), .A2(n9105), .ZN(n9278) );
  NAND2_X1 U10294 ( .A1(n8937), .A2(n9103), .ZN(n9294) );
  INV_X1 U10295 ( .A(n9294), .ZN(n9298) );
  NAND2_X1 U10296 ( .A1(n8939), .A2(n8938), .ZN(n9351) );
  NAND4_X1 U10297 ( .A1(n8943), .A2(n8942), .A3(n8941), .A4(n8940), .ZN(n8946)
         );
  OR4_X1 U10298 ( .A1(n8947), .A2(n8946), .A3(n8945), .A4(n8944), .ZN(n8951)
         );
  NOR4_X1 U10299 ( .A1(n8951), .A2(n8950), .A3(n8949), .A4(n8948), .ZN(n8952)
         );
  NAND4_X1 U10300 ( .A1(n8955), .A2(n8954), .A3(n8953), .A4(n8952), .ZN(n8957)
         );
  NOR4_X1 U10301 ( .A1(n9324), .A2(n9351), .A3(n8957), .A4(n8956), .ZN(n8958)
         );
  NAND2_X1 U10302 ( .A1(n9298), .A2(n8958), .ZN(n8959) );
  NOR4_X1 U10303 ( .A1(n9246), .A2(n9269), .A3(n9278), .A4(n8959), .ZN(n8960)
         );
  NAND4_X1 U10304 ( .A1(n9206), .A2(n9220), .A3(n9232), .A4(n8960), .ZN(n8961)
         );
  NOR4_X1 U10305 ( .A1(n9116), .A2(n9168), .A3(n9188), .A4(n8961), .ZN(n8962)
         );
  NAND4_X1 U10306 ( .A1(n8963), .A2(n9137), .A3(n9118), .A4(n8962), .ZN(n8964)
         );
  NOR4_X1 U10307 ( .A1(n8967), .A2(n8966), .A3(n8965), .A4(n8964), .ZN(n8969)
         );
  NOR2_X1 U10308 ( .A1(n8969), .A2(n8968), .ZN(n8970) );
  MUX2_X1 U10309 ( .A(n8971), .B(n5586), .S(n8970), .Z(n8972) );
  INV_X1 U10310 ( .A(n8976), .ZN(n8979) );
  OAI21_X1 U10311 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n8985) );
  NAND2_X1 U10312 ( .A1(n8980), .A2(n9013), .ZN(n8981) );
  OAI211_X1 U10313 ( .C1(n8983), .C2(n8982), .A(n8981), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8984) );
  OAI21_X1 U10314 ( .B1(n8986), .B2(n8985), .A(n8984), .ZN(P1_U3240) );
  MUX2_X1 U10315 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9121), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10316 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8987), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10317 ( .A(n9123), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9001), .Z(
        P1_U3583) );
  MUX2_X1 U10318 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9097), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10319 ( .A(n9186), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9001), .Z(
        P1_U3581) );
  MUX2_X1 U10320 ( .A(n9207), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9001), .Z(
        P1_U3580) );
  MUX2_X1 U10321 ( .A(n9221), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9001), .Z(
        P1_U3579) );
  MUX2_X1 U10322 ( .A(n9234), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9001), .Z(
        P1_U3578) );
  MUX2_X1 U10323 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9251), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10324 ( .A(n9271), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9001), .Z(
        P1_U3576) );
  MUX2_X1 U10325 ( .A(n9250), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9001), .Z(
        P1_U3575) );
  MUX2_X1 U10326 ( .A(n9303), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9001), .Z(
        P1_U3574) );
  MUX2_X1 U10327 ( .A(n9330), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9001), .Z(
        P1_U3573) );
  MUX2_X1 U10328 ( .A(n9302), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9001), .Z(
        P1_U3572) );
  MUX2_X1 U10329 ( .A(n9328), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9001), .Z(
        P1_U3571) );
  MUX2_X1 U10330 ( .A(n9342), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9001), .Z(
        P1_U3570) );
  MUX2_X1 U10331 ( .A(n8988), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9001), .Z(
        P1_U3569) );
  MUX2_X1 U10332 ( .A(n8989), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9001), .Z(
        P1_U3568) );
  MUX2_X1 U10333 ( .A(n8990), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9001), .Z(
        P1_U3567) );
  MUX2_X1 U10334 ( .A(n8991), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9001), .Z(
        P1_U3566) );
  MUX2_X1 U10335 ( .A(n8992), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9001), .Z(
        P1_U3565) );
  MUX2_X1 U10336 ( .A(n8993), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9001), .Z(
        P1_U3564) );
  MUX2_X1 U10337 ( .A(n8994), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9001), .Z(
        P1_U3563) );
  MUX2_X1 U10338 ( .A(n8995), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9001), .Z(
        P1_U3562) );
  MUX2_X1 U10339 ( .A(n8996), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9001), .Z(
        P1_U3561) );
  MUX2_X1 U10340 ( .A(n8997), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9001), .Z(
        P1_U3560) );
  MUX2_X1 U10341 ( .A(n8998), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9001), .Z(
        P1_U3559) );
  MUX2_X1 U10342 ( .A(n8999), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9001), .Z(
        P1_U3558) );
  MUX2_X1 U10343 ( .A(n9000), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9001), .Z(
        P1_U3557) );
  MUX2_X1 U10344 ( .A(n9002), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9001), .Z(
        P1_U3556) );
  INV_X1 U10345 ( .A(n9003), .ZN(n9004) );
  NOR2_X1 U10346 ( .A1(n9005), .A2(n9004), .ZN(n9008) );
  AOI211_X1 U10347 ( .C1(n9008), .C2(n9007), .A(n9006), .B(n9638), .ZN(n9009)
         );
  AOI21_X1 U10348 ( .B1(n9628), .B2(n9010), .A(n9009), .ZN(n9024) );
  AOI22_X1 U10349 ( .A1(n9544), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n4258), .ZN(n9023) );
  AOI21_X1 U10350 ( .B1(n9013), .B2(n9012), .A(n9011), .ZN(n9543) );
  MUX2_X1 U10351 ( .A(n9015), .B(n9014), .S(n9071), .Z(n9017) );
  NAND2_X1 U10352 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  OAI211_X1 U10353 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9543), .A(n9018), .B(
        P1_U4006), .ZN(n9563) );
  OAI211_X1 U10354 ( .C1(n9021), .C2(n9020), .A(n9553), .B(n9019), .ZN(n9022)
         );
  NAND4_X1 U10355 ( .A1(n9024), .A2(n9023), .A3(n9563), .A4(n9022), .ZN(
        P1_U3243) );
  OAI21_X1 U10356 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n9029) );
  AOI22_X1 U10357 ( .A1(n9553), .A2(n9029), .B1(n9628), .B2(n9028), .ZN(n9036)
         );
  AOI21_X1 U10358 ( .B1(n9544), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9030), .ZN(
        n9035) );
  OAI211_X1 U10359 ( .C1(n9033), .C2(n9032), .A(n9616), .B(n9031), .ZN(n9034)
         );
  NAND3_X1 U10360 ( .A1(n9036), .A2(n9035), .A3(n9034), .ZN(P1_U3249) );
  NAND2_X1 U10361 ( .A1(n9037), .A2(n9049), .ZN(n9039) );
  NAND2_X1 U10362 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9599), .ZN(n9041) );
  OAI21_X1 U10363 ( .B1(n9599), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9041), .ZN(
        n9595) );
  NOR2_X1 U10364 ( .A1(n9596), .A2(n9595), .ZN(n9594) );
  AOI21_X1 U10365 ( .B1(n9599), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9594), .ZN(
        n9605) );
  OR2_X1 U10366 ( .A1(n9610), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U10367 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9610), .ZN(n9042) );
  NAND2_X1 U10368 ( .A1(n9043), .A2(n9042), .ZN(n9606) );
  NOR2_X1 U10369 ( .A1(n9605), .A2(n9606), .ZN(n9607) );
  OR2_X1 U10370 ( .A1(n9627), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U10371 ( .A1(n9627), .A2(n9044), .ZN(n9045) );
  AND2_X1 U10372 ( .A1(n9046), .A2(n9045), .ZN(n9623) );
  XNOR2_X1 U10373 ( .A(n9627), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9636) );
  INV_X1 U10374 ( .A(n9610), .ZN(n9056) );
  XOR2_X1 U10375 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9610), .Z(n9618) );
  INV_X1 U10376 ( .A(n9599), .ZN(n9054) );
  MUX2_X1 U10377 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9047), .S(n9599), .Z(n9601) );
  AOI21_X1 U10378 ( .B1(n9518), .B2(n9049), .A(n9048), .ZN(n9050) );
  XNOR2_X1 U10379 ( .A(n9050), .B(n9588), .ZN(n9589) );
  INV_X1 U10380 ( .A(n9050), .ZN(n9051) );
  OAI22_X1 U10381 ( .A1(n9589), .A2(n9053), .B1(n9052), .B2(n9051), .ZN(n9602)
         );
  NAND2_X1 U10382 ( .A1(n9601), .A2(n9602), .ZN(n9600) );
  OAI21_X1 U10383 ( .B1(n9054), .B2(n9047), .A(n9600), .ZN(n9617) );
  NAND2_X1 U10384 ( .A1(n9618), .A2(n9617), .ZN(n9615) );
  OAI21_X1 U10385 ( .B1(n9056), .B2(n9055), .A(n9615), .ZN(n9635) );
  NOR2_X1 U10386 ( .A1(n9636), .A2(n9635), .ZN(n9634) );
  AOI21_X1 U10387 ( .B1(n9058), .B2(n9057), .A(n9634), .ZN(n9060) );
  XOR2_X1 U10388 ( .A(n9060), .B(n9059), .Z(n9062) );
  OAI22_X1 U10389 ( .A1(n9061), .A2(n9632), .B1(n9062), .B2(n9638), .ZN(n9066)
         );
  NAND2_X1 U10390 ( .A1(n9061), .A2(n9541), .ZN(n9064) );
  AOI21_X1 U10391 ( .B1(n9062), .B2(n9616), .A(n9628), .ZN(n9063) );
  NAND2_X1 U10392 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  MUX2_X1 U10393 ( .A(n9066), .B(n9065), .S(n5586), .Z(n9069) );
  OAI21_X1 U10394 ( .B1(n9641), .B2(n5042), .A(n9067), .ZN(n9068) );
  INV_X1 U10395 ( .A(n9426), .ZN(n9260) );
  NAND2_X1 U10396 ( .A1(n9384), .A2(n9126), .ZN(n9381) );
  NAND2_X1 U10397 ( .A1(n9378), .A2(n9372), .ZN(n9075) );
  INV_X1 U10398 ( .A(P1_B_REG_SCAN_IN), .ZN(n9070) );
  NOR2_X1 U10399 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  NOR2_X1 U10400 ( .A1(n9345), .A2(n9072), .ZN(n9122) );
  NAND2_X1 U10401 ( .A1(n9122), .A2(n9073), .ZN(n9382) );
  NOR2_X1 U10402 ( .A1(n9364), .A2(n9382), .ZN(n9078) );
  AOI21_X1 U10403 ( .B1(n9364), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9078), .ZN(
        n9074) );
  OAI211_X1 U10404 ( .C1(n9379), .C2(n9369), .A(n9075), .B(n9074), .ZN(
        P1_U3261) );
  INV_X1 U10405 ( .A(n9126), .ZN(n9076) );
  NAND2_X1 U10406 ( .A1(n9077), .A2(n9076), .ZN(n9380) );
  NAND3_X1 U10407 ( .A1(n9381), .A2(n9372), .A3(n9380), .ZN(n9080) );
  AOI21_X1 U10408 ( .B1(n9364), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9078), .ZN(
        n9079) );
  OAI211_X1 U10409 ( .C1(n9384), .C2(n9369), .A(n9080), .B(n9079), .ZN(
        P1_U3262) );
  NAND2_X1 U10410 ( .A1(n9506), .A2(n9342), .ZN(n9082) );
  NAND2_X1 U10411 ( .A1(n9083), .A2(n9082), .ZN(n9350) );
  AND2_X1 U10412 ( .A1(n9360), .A2(n9328), .ZN(n9084) );
  INV_X1 U10413 ( .A(n9430), .ZN(n9268) );
  AOI21_X1 U10414 ( .B1(n9426), .B2(n9271), .A(n9241), .ZN(n9227) );
  NOR2_X1 U10415 ( .A1(n9420), .A2(n9251), .ZN(n9089) );
  NAND2_X1 U10416 ( .A1(n9217), .A2(n9090), .ZN(n9091) );
  NAND2_X1 U10417 ( .A1(n9203), .A2(n9092), .ZN(n9093) );
  INV_X1 U10418 ( .A(n9094), .ZN(n9194) );
  NAND2_X1 U10419 ( .A1(n9181), .A2(n9095), .ZN(n9096) );
  NOR2_X1 U10420 ( .A1(n9397), .A2(n9097), .ZN(n9098) );
  AOI21_X1 U10421 ( .B1(n9151), .B2(n9116), .A(n9098), .ZN(n9135) );
  NAND2_X1 U10422 ( .A1(n9135), .A2(n9134), .ZN(n9133) );
  OAI21_X1 U10423 ( .B1(n9148), .B2(n9157), .A(n9133), .ZN(n9099) );
  XNOR2_X1 U10424 ( .A(n9099), .B(n9118), .ZN(n9386) );
  INV_X1 U10425 ( .A(n9386), .ZN(n9132) );
  INV_X1 U10426 ( .A(n9103), .ZN(n9104) );
  INV_X1 U10427 ( .A(n9111), .ZN(n9112) );
  NAND2_X1 U10428 ( .A1(n9136), .A2(n9117), .ZN(n9120) );
  INV_X1 U10429 ( .A(n9118), .ZN(n9119) );
  XNOR2_X1 U10430 ( .A(n9120), .B(n9119), .ZN(n9125) );
  AOI22_X1 U10431 ( .A1(n9123), .A2(n9343), .B1(n9122), .B2(n9121), .ZN(n9124)
         );
  OAI21_X1 U10432 ( .B1(n9125), .B2(n9280), .A(n9124), .ZN(n9387) );
  AOI211_X1 U10433 ( .C1(n9389), .C2(n9142), .A(n9696), .B(n9126), .ZN(n9388)
         );
  NAND2_X1 U10434 ( .A1(n9388), .A2(n9211), .ZN(n9129) );
  AOI22_X1 U10435 ( .A1(n9127), .A2(n9287), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9364), .ZN(n9128) );
  OAI211_X1 U10436 ( .C1(n4605), .C2(n9369), .A(n9129), .B(n9128), .ZN(n9130)
         );
  AOI21_X1 U10437 ( .B1(n9387), .B2(n6776), .A(n9130), .ZN(n9131) );
  OAI21_X1 U10438 ( .B1(n9132), .B2(n9335), .A(n9131), .ZN(P1_U3355) );
  INV_X1 U10439 ( .A(n9136), .ZN(n9140) );
  AOI21_X1 U10440 ( .B1(n9152), .B2(n9138), .A(n9137), .ZN(n9139) );
  INV_X1 U10441 ( .A(n9158), .ZN(n9144) );
  INV_X1 U10442 ( .A(n9142), .ZN(n9143) );
  AOI211_X1 U10443 ( .C1(n9393), .C2(n9144), .A(n9696), .B(n9143), .ZN(n9392)
         );
  NAND2_X1 U10444 ( .A1(n9392), .A2(n9211), .ZN(n9147) );
  AOI22_X1 U10445 ( .A1(n9145), .A2(n9287), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9364), .ZN(n9146) );
  OAI211_X1 U10446 ( .C1(n9148), .C2(n9369), .A(n9147), .B(n9146), .ZN(n9149)
         );
  AOI21_X1 U10447 ( .B1(n9391), .B2(n6776), .A(n9149), .ZN(n9150) );
  OAI21_X1 U10448 ( .B1(n9394), .B2(n9335), .A(n9150), .ZN(P1_U3263) );
  XNOR2_X1 U10449 ( .A(n9151), .B(n9153), .ZN(n9399) );
  OAI211_X1 U10450 ( .C1(n9154), .C2(n9153), .A(n9152), .B(n9348), .ZN(n9156)
         );
  NAND2_X1 U10451 ( .A1(n9186), .A2(n9343), .ZN(n9155) );
  OAI211_X1 U10452 ( .C1(n9157), .C2(n9345), .A(n9156), .B(n9155), .ZN(n9395)
         );
  INV_X1 U10453 ( .A(n9397), .ZN(n9162) );
  NAND2_X1 U10454 ( .A1(n9396), .A2(n9211), .ZN(n9161) );
  AOI22_X1 U10455 ( .A1(n9159), .A2(n9287), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9364), .ZN(n9160) );
  OAI211_X1 U10456 ( .C1(n9162), .C2(n9369), .A(n9161), .B(n9160), .ZN(n9163)
         );
  AOI21_X1 U10457 ( .B1(n9395), .B2(n6776), .A(n9163), .ZN(n9164) );
  OAI21_X1 U10458 ( .B1(n9399), .B2(n9335), .A(n9164), .ZN(P1_U3264) );
  XNOR2_X1 U10459 ( .A(n9165), .B(n9168), .ZN(n9404) );
  NAND2_X1 U10460 ( .A1(n9167), .A2(n9166), .ZN(n9170) );
  INV_X1 U10461 ( .A(n9168), .ZN(n9169) );
  XNOR2_X1 U10462 ( .A(n9170), .B(n9169), .ZN(n9171) );
  OAI222_X1 U10463 ( .A1(n9282), .A2(n9173), .B1(n9345), .B2(n9172), .C1(n9171), .C2(n9280), .ZN(n9400) );
  INV_X1 U10464 ( .A(n9174), .ZN(n9191) );
  INV_X1 U10465 ( .A(n9175), .ZN(n9176) );
  AOI211_X1 U10466 ( .C1(n9402), .C2(n9191), .A(n9696), .B(n9176), .ZN(n9401)
         );
  NAND2_X1 U10467 ( .A1(n9401), .A2(n9211), .ZN(n9180) );
  INV_X1 U10468 ( .A(n9177), .ZN(n9178) );
  AOI22_X1 U10469 ( .A1(n9178), .A2(n9287), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9364), .ZN(n9179) );
  OAI211_X1 U10470 ( .C1(n9181), .C2(n9369), .A(n9180), .B(n9179), .ZN(n9182)
         );
  AOI21_X1 U10471 ( .B1(n9400), .B2(n6776), .A(n9182), .ZN(n9183) );
  OAI21_X1 U10472 ( .B1(n9404), .B2(n9335), .A(n9183), .ZN(P1_U3265) );
  NAND2_X1 U10473 ( .A1(n9204), .A2(n9184), .ZN(n9185) );
  XOR2_X1 U10474 ( .A(n9188), .B(n9185), .Z(n9187) );
  AOI222_X1 U10475 ( .A1(n9348), .A2(n9187), .B1(n9221), .B2(n9343), .C1(n9186), .C2(n9329), .ZN(n9408) );
  XNOR2_X1 U10476 ( .A(n9189), .B(n9188), .ZN(n9405) );
  NAND2_X1 U10477 ( .A1(n9405), .A2(n9352), .ZN(n9198) );
  INV_X1 U10478 ( .A(n9190), .ZN(n9200) );
  OAI211_X1 U10479 ( .C1(n9194), .C2(n9200), .A(n9191), .B(n9673), .ZN(n9406)
         );
  INV_X1 U10480 ( .A(n9406), .ZN(n9196) );
  AOI22_X1 U10481 ( .A1(n9192), .A2(n9287), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9364), .ZN(n9193) );
  OAI21_X1 U10482 ( .B1(n9194), .B2(n9369), .A(n9193), .ZN(n9195) );
  AOI21_X1 U10483 ( .B1(n9196), .B2(n9211), .A(n9195), .ZN(n9197) );
  OAI211_X1 U10484 ( .C1(n9364), .C2(n9408), .A(n9198), .B(n9197), .ZN(
        P1_U3266) );
  XNOR2_X1 U10485 ( .A(n9199), .B(n9206), .ZN(n9414) );
  AOI211_X1 U10486 ( .C1(n9411), .C2(n4603), .A(n9696), .B(n9200), .ZN(n9410)
         );
  AOI22_X1 U10487 ( .A1(n9201), .A2(n9287), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9364), .ZN(n9202) );
  OAI21_X1 U10488 ( .B1(n9203), .B2(n9369), .A(n9202), .ZN(n9210) );
  OAI21_X1 U10489 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9208) );
  AOI222_X1 U10490 ( .A1(n9348), .A2(n9208), .B1(n9207), .B2(n9329), .C1(n9234), .C2(n9343), .ZN(n9413) );
  NOR2_X1 U10491 ( .A1(n9413), .A2(n9364), .ZN(n9209) );
  AOI211_X1 U10492 ( .C1(n9410), .C2(n9211), .A(n9210), .B(n9209), .ZN(n9212)
         );
  OAI21_X1 U10493 ( .B1(n9414), .B2(n9335), .A(n9212), .ZN(P1_U3267) );
  XOR2_X1 U10494 ( .A(n9220), .B(n9213), .Z(n9419) );
  AND2_X1 U10495 ( .A1(n9228), .A2(n9415), .ZN(n9214) );
  NOR2_X1 U10496 ( .A1(n9215), .A2(n9214), .ZN(n9416) );
  INV_X1 U10497 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9216) );
  OAI22_X1 U10498 ( .A1(n9217), .A2(n9369), .B1(n9216), .B2(n6776), .ZN(n9218)
         );
  AOI21_X1 U10499 ( .B1(n9416), .B2(n9372), .A(n9218), .ZN(n9226) );
  XOR2_X1 U10500 ( .A(n9220), .B(n9219), .Z(n9222) );
  AOI222_X1 U10501 ( .A1(n9348), .A2(n9222), .B1(n9221), .B2(n9329), .C1(n9251), .C2(n9343), .ZN(n9418) );
  OAI21_X1 U10502 ( .B1(n9223), .B2(n9367), .A(n9418), .ZN(n9224) );
  NAND2_X1 U10503 ( .A1(n9224), .A2(n6776), .ZN(n9225) );
  OAI211_X1 U10504 ( .C1(n9419), .C2(n9335), .A(n9226), .B(n9225), .ZN(
        P1_U3268) );
  XNOR2_X1 U10505 ( .A(n9227), .B(n9232), .ZN(n9424) );
  INV_X1 U10506 ( .A(n9228), .ZN(n9229) );
  AOI21_X1 U10507 ( .B1(n9420), .B2(n9253), .A(n9229), .ZN(n9421) );
  INV_X1 U10508 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9230) );
  OAI22_X1 U10509 ( .A1(n9231), .A2(n9369), .B1(n9230), .B2(n6776), .ZN(n9239)
         );
  XNOR2_X1 U10510 ( .A(n9233), .B(n9232), .ZN(n9235) );
  AOI222_X1 U10511 ( .A1(n9348), .A2(n9235), .B1(n9234), .B2(n9329), .C1(n9271), .C2(n9343), .ZN(n9423) );
  NAND2_X1 U10512 ( .A1(n9236), .A2(n9287), .ZN(n9237) );
  AOI21_X1 U10513 ( .B1(n9423), .B2(n9237), .A(n9364), .ZN(n9238) );
  AOI211_X1 U10514 ( .C1(n9421), .C2(n9372), .A(n9239), .B(n9238), .ZN(n9240)
         );
  OAI21_X1 U10515 ( .B1(n9424), .B2(n9335), .A(n9240), .ZN(P1_U3269) );
  AOI21_X1 U10516 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9244) );
  INV_X1 U10517 ( .A(n9244), .ZN(n9429) );
  NAND2_X1 U10518 ( .A1(n9246), .A2(n9245), .ZN(n9248) );
  OAI21_X1 U10519 ( .B1(n9249), .B2(n9248), .A(n9247), .ZN(n9252) );
  AOI222_X1 U10520 ( .A1(n9348), .A2(n9252), .B1(n9251), .B2(n9329), .C1(n9250), .C2(n9343), .ZN(n9428) );
  INV_X1 U10521 ( .A(n9264), .ZN(n9255) );
  INV_X1 U10522 ( .A(n9253), .ZN(n9254) );
  AOI211_X1 U10523 ( .C1(n9426), .C2(n9255), .A(n9696), .B(n9254), .ZN(n9425)
         );
  NAND2_X1 U10524 ( .A1(n9425), .A2(n9256), .ZN(n9257) );
  OAI211_X1 U10525 ( .C1(n9367), .C2(n9258), .A(n9428), .B(n9257), .ZN(n9262)
         );
  OAI22_X1 U10526 ( .A1(n9260), .A2(n9369), .B1(n6776), .B2(n9259), .ZN(n9261)
         );
  AOI21_X1 U10527 ( .B1(n9262), .B2(n6776), .A(n9261), .ZN(n9263) );
  OAI21_X1 U10528 ( .B1(n9429), .B2(n9335), .A(n9263), .ZN(P1_U3270) );
  XOR2_X1 U10529 ( .A(n9269), .B(n4329), .Z(n9434) );
  AOI21_X1 U10530 ( .B1(n9430), .B2(n9284), .A(n9264), .ZN(n9431) );
  INV_X1 U10531 ( .A(n9265), .ZN(n9266) );
  AOI22_X1 U10532 ( .A1(n9364), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9266), .B2(
        n9287), .ZN(n9267) );
  OAI21_X1 U10533 ( .B1(n9268), .B2(n9369), .A(n9267), .ZN(n9274) );
  XNOR2_X1 U10534 ( .A(n9270), .B(n9269), .ZN(n9272) );
  AOI222_X1 U10535 ( .A1(n9348), .A2(n9272), .B1(n9271), .B2(n9329), .C1(n9303), .C2(n9343), .ZN(n9433) );
  NOR2_X1 U10536 ( .A1(n9433), .A2(n9364), .ZN(n9273) );
  AOI211_X1 U10537 ( .C1(n9431), .C2(n9372), .A(n9274), .B(n9273), .ZN(n9275)
         );
  OAI21_X1 U10538 ( .B1(n9434), .B2(n9335), .A(n9275), .ZN(P1_U3271) );
  XOR2_X1 U10539 ( .A(n9276), .B(n9278), .Z(n9440) );
  AOI21_X1 U10540 ( .B1(n4340), .B2(n9278), .A(n9277), .ZN(n9279) );
  OAI222_X1 U10541 ( .A1(n9345), .A2(n9283), .B1(n9282), .B2(n9281), .C1(n9280), .C2(n9279), .ZN(n9435) );
  INV_X1 U10542 ( .A(n9284), .ZN(n9285) );
  AOI21_X1 U10543 ( .B1(n9436), .B2(n9307), .A(n9285), .ZN(n9437) );
  NAND2_X1 U10544 ( .A1(n9437), .A2(n9372), .ZN(n9290) );
  INV_X1 U10545 ( .A(n9286), .ZN(n9288) );
  AOI22_X1 U10546 ( .A1(n9364), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9288), .B2(
        n9287), .ZN(n9289) );
  OAI211_X1 U10547 ( .C1(n9291), .C2(n9369), .A(n9290), .B(n9289), .ZN(n9292)
         );
  AOI21_X1 U10548 ( .B1(n9435), .B2(n6776), .A(n9292), .ZN(n9293) );
  OAI21_X1 U10549 ( .B1(n9440), .B2(n9335), .A(n9293), .ZN(P1_U3272) );
  NOR2_X1 U10550 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  OR2_X1 U10551 ( .A1(n9297), .A2(n9296), .ZN(n9441) );
  NOR2_X1 U10552 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  OAI21_X1 U10553 ( .B1(n9301), .B2(n9300), .A(n9348), .ZN(n9305) );
  AOI22_X1 U10554 ( .A1(n9329), .A2(n9303), .B1(n9343), .B2(n9302), .ZN(n9304)
         );
  NAND2_X1 U10555 ( .A1(n9305), .A2(n9304), .ZN(n9445) );
  OR2_X1 U10556 ( .A1(n9318), .A2(n9442), .ZN(n9306) );
  NAND2_X1 U10557 ( .A1(n9307), .A2(n9306), .ZN(n9443) );
  NAND2_X1 U10558 ( .A1(n9364), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9308) );
  OAI21_X1 U10559 ( .B1(n9367), .B2(n9309), .A(n9308), .ZN(n9310) );
  AOI21_X1 U10560 ( .B1(n9311), .B2(n9361), .A(n9310), .ZN(n9312) );
  OAI21_X1 U10561 ( .B1(n9443), .B2(n9313), .A(n9312), .ZN(n9314) );
  AOI21_X1 U10562 ( .B1(n9445), .B2(n6776), .A(n9314), .ZN(n9316) );
  OAI21_X1 U10563 ( .B1(n9441), .B2(n9335), .A(n9316), .ZN(P1_U3273) );
  XOR2_X1 U10564 ( .A(n9324), .B(n9317), .Z(n9452) );
  AOI21_X1 U10565 ( .B1(n9448), .B2(n9356), .A(n9318), .ZN(n9449) );
  NOR2_X1 U10566 ( .A1(n9319), .A2(n9367), .ZN(n9320) );
  AOI21_X1 U10567 ( .B1(n9364), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9320), .ZN(
        n9321) );
  OAI21_X1 U10568 ( .B1(n9322), .B2(n9369), .A(n9321), .ZN(n9333) );
  INV_X1 U10569 ( .A(n9323), .ZN(n9327) );
  INV_X1 U10570 ( .A(n9324), .ZN(n9326) );
  OAI21_X1 U10571 ( .B1(n9327), .B2(n9326), .A(n9325), .ZN(n9331) );
  AOI222_X1 U10572 ( .A1(n9348), .A2(n9331), .B1(n9330), .B2(n9329), .C1(n9328), .C2(n9343), .ZN(n9451) );
  NOR2_X1 U10573 ( .A1(n9451), .A2(n9364), .ZN(n9332) );
  AOI211_X1 U10574 ( .C1(n9449), .C2(n9372), .A(n9333), .B(n9332), .ZN(n9334)
         );
  OAI21_X1 U10575 ( .B1(n9335), .B2(n9452), .A(n9334), .ZN(P1_U3274) );
  INV_X1 U10576 ( .A(n9336), .ZN(n9338) );
  OAI21_X1 U10577 ( .B1(n9339), .B2(n9338), .A(n9337), .ZN(n9341) );
  INV_X1 U10578 ( .A(n9351), .ZN(n9340) );
  XNOR2_X1 U10579 ( .A(n9341), .B(n9340), .ZN(n9349) );
  NAND2_X1 U10580 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  OAI21_X1 U10581 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(n9347) );
  AOI21_X1 U10582 ( .B1(n9349), .B2(n9348), .A(n9347), .ZN(n9503) );
  XOR2_X1 U10583 ( .A(n9351), .B(n9350), .Z(n9505) );
  NAND2_X1 U10584 ( .A1(n9505), .A2(n9352), .ZN(n9363) );
  OAI22_X1 U10585 ( .A1(n6776), .A2(n9354), .B1(n9353), .B2(n9367), .ZN(n9359)
         );
  OAI211_X1 U10586 ( .C1(n4614), .C2(n4613), .A(n9673), .B(n9356), .ZN(n9502)
         );
  NOR2_X1 U10587 ( .A1(n9502), .A2(n9357), .ZN(n9358) );
  AOI211_X1 U10588 ( .C1(n9361), .C2(n9360), .A(n9359), .B(n9358), .ZN(n9362)
         );
  OAI211_X1 U10589 ( .C1(n9364), .C2(n9503), .A(n9363), .B(n9362), .ZN(
        P1_U3275) );
  MUX2_X1 U10590 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9365), .S(n6776), .Z(n9366)
         );
  INV_X1 U10591 ( .A(n9366), .ZN(n9377) );
  OAI22_X1 U10592 ( .A1(n9369), .A2(n9368), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9367), .ZN(n9370) );
  AOI21_X1 U10593 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(n9376) );
  NAND2_X1 U10594 ( .A1(n9374), .A2(n9373), .ZN(n9375) );
  NAND3_X1 U10595 ( .A1(n9377), .A2(n9376), .A3(n9375), .ZN(P1_U3288) );
  MUX2_X1 U10596 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9459), .S(n9716), .Z(
        P1_U3554) );
  NAND3_X1 U10597 ( .A1(n9381), .A2(n9673), .A3(n9380), .ZN(n9383) );
  OAI211_X1 U10598 ( .C1(n9384), .C2(n9694), .A(n9383), .B(n9382), .ZN(n9460)
         );
  MUX2_X1 U10599 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9460), .S(n9716), .Z(
        P1_U3553) );
  NAND2_X1 U10600 ( .A1(n9385), .A2(n9653), .ZN(n9700) );
  NAND2_X1 U10601 ( .A1(n9386), .A2(n9700), .ZN(n9390) );
  MUX2_X1 U10602 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9461), .S(n9716), .Z(
        P1_U3552) );
  MUX2_X1 U10603 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9462), .S(n9716), .Z(
        P1_U3551) );
  AOI211_X1 U10604 ( .C1(n9456), .C2(n9397), .A(n9396), .B(n9395), .ZN(n9398)
         );
  OAI21_X1 U10605 ( .B1(n9399), .B2(n9678), .A(n9398), .ZN(n9463) );
  MUX2_X1 U10606 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9463), .S(n9716), .Z(
        P1_U3550) );
  OAI21_X1 U10607 ( .B1(n9404), .B2(n9678), .A(n9403), .ZN(n9464) );
  MUX2_X1 U10608 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9464), .S(n9716), .Z(
        P1_U3549) );
  NAND2_X1 U10609 ( .A1(n9405), .A2(n9700), .ZN(n9409) );
  NAND4_X1 U10610 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(n9465)
         );
  MUX2_X1 U10611 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9465), .S(n9716), .Z(
        P1_U3548) );
  AOI21_X1 U10612 ( .B1(n9456), .B2(n9411), .A(n9410), .ZN(n9412) );
  OAI211_X1 U10613 ( .C1(n9414), .C2(n9678), .A(n9413), .B(n9412), .ZN(n9466)
         );
  MUX2_X1 U10614 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9466), .S(n9716), .Z(
        P1_U3547) );
  AOI22_X1 U10615 ( .A1(n9416), .A2(n9673), .B1(n9456), .B2(n9415), .ZN(n9417)
         );
  OAI211_X1 U10616 ( .C1(n9419), .C2(n9678), .A(n9418), .B(n9417), .ZN(n9467)
         );
  MUX2_X1 U10617 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9467), .S(n9716), .Z(
        P1_U3546) );
  AOI22_X1 U10618 ( .A1(n9421), .A2(n9673), .B1(n9456), .B2(n9420), .ZN(n9422)
         );
  OAI211_X1 U10619 ( .C1(n9424), .C2(n9678), .A(n9423), .B(n9422), .ZN(n9468)
         );
  MUX2_X1 U10620 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9468), .S(n9716), .Z(
        P1_U3545) );
  AOI21_X1 U10621 ( .B1(n9456), .B2(n9426), .A(n9425), .ZN(n9427) );
  OAI211_X1 U10622 ( .C1(n9429), .C2(n9678), .A(n9428), .B(n9427), .ZN(n9469)
         );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9469), .S(n9716), .Z(
        P1_U3544) );
  AOI22_X1 U10624 ( .A1(n9431), .A2(n9673), .B1(n9456), .B2(n9430), .ZN(n9432)
         );
  OAI211_X1 U10625 ( .C1(n9434), .C2(n9678), .A(n9433), .B(n9432), .ZN(n9470)
         );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9470), .S(n9716), .Z(
        P1_U3543) );
  INV_X1 U10627 ( .A(n9435), .ZN(n9439) );
  AOI22_X1 U10628 ( .A1(n9437), .A2(n9673), .B1(n9456), .B2(n9436), .ZN(n9438)
         );
  OAI211_X1 U10629 ( .C1(n9440), .C2(n9678), .A(n9439), .B(n9438), .ZN(n9471)
         );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9471), .S(n9716), .Z(
        P1_U3542) );
  OAI22_X1 U10631 ( .A1(n9443), .A2(n9696), .B1(n9442), .B2(n9694), .ZN(n9444)
         );
  NOR2_X1 U10632 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  NAND2_X1 U10633 ( .A1(n9447), .A2(n9446), .ZN(n9472) );
  MUX2_X1 U10634 ( .A(n9472), .B(P1_REG1_REG_18__SCAN_IN), .S(n9713), .Z(
        P1_U3541) );
  AOI22_X1 U10635 ( .A1(n9449), .A2(n9673), .B1(n9456), .B2(n9448), .ZN(n9450)
         );
  OAI211_X1 U10636 ( .C1(n9452), .C2(n9678), .A(n9451), .B(n9450), .ZN(n9473)
         );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9473), .S(n9716), .Z(
        P1_U3540) );
  AOI211_X1 U10638 ( .C1(n9456), .C2(n9455), .A(n9454), .B(n9453), .ZN(n9457)
         );
  OAI21_X1 U10639 ( .B1(n9678), .B2(n9458), .A(n9457), .ZN(n9474) );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9474), .S(n9716), .Z(
        P1_U3535) );
  MUX2_X1 U10641 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9460), .S(n9704), .Z(
        P1_U3521) );
  MUX2_X1 U10642 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9461), .S(n9704), .Z(
        P1_U3520) );
  MUX2_X1 U10643 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9462), .S(n9704), .Z(
        P1_U3519) );
  MUX2_X1 U10644 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9463), .S(n9704), .Z(
        P1_U3518) );
  MUX2_X1 U10645 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9464), .S(n9704), .Z(
        P1_U3517) );
  MUX2_X1 U10646 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9465), .S(n9704), .Z(
        P1_U3516) );
  MUX2_X1 U10647 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9466), .S(n9704), .Z(
        P1_U3515) );
  MUX2_X1 U10648 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9467), .S(n9704), .Z(
        P1_U3514) );
  MUX2_X1 U10649 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9468), .S(n9704), .Z(
        P1_U3513) );
  MUX2_X1 U10650 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9469), .S(n9704), .Z(
        P1_U3512) );
  MUX2_X1 U10651 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9470), .S(n9704), .Z(
        P1_U3511) );
  MUX2_X1 U10652 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9471), .S(n9704), .Z(
        P1_U3510) );
  MUX2_X1 U10653 ( .A(n9472), .B(P1_REG0_REG_18__SCAN_IN), .S(n9702), .Z(
        P1_U3508) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9473), .S(n9704), .Z(
        P1_U3505) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9474), .S(n9704), .Z(
        P1_U3490) );
  MUX2_X1 U10656 ( .A(P1_D_REG_1__SCAN_IN), .B(n9475), .S(n9648), .Z(P1_U3441)
         );
  NAND3_X1 U10657 ( .A1(n9477), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9479) );
  OAI22_X1 U10658 ( .A1(n9476), .A2(n9479), .B1(n10022), .B2(n9478), .ZN(n9480) );
  AOI21_X1 U10659 ( .B1(n8531), .B2(n9481), .A(n9480), .ZN(n9482) );
  INV_X1 U10660 ( .A(n9482), .ZN(P1_U3322) );
  MUX2_X1 U10661 ( .A(n9483), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10662 ( .A(n9653), .ZN(n9658) );
  OAI21_X1 U10663 ( .B1(n9485), .B2(n9694), .A(n9484), .ZN(n9486) );
  AOI21_X1 U10664 ( .B1(n9487), .B2(n9658), .A(n9486), .ZN(n9488) );
  AND2_X1 U10665 ( .A1(n9489), .A2(n9488), .ZN(n9492) );
  INV_X1 U10666 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9490) );
  AOI22_X1 U10667 ( .A1(n9704), .A2(n9492), .B1(n9490), .B2(n9702), .ZN(
        P1_U3484) );
  AOI22_X1 U10668 ( .A1(n9716), .A2(n9492), .B1(n9491), .B2(n9713), .ZN(
        P1_U3533) );
  INV_X1 U10669 ( .A(n9493), .ZN(n9494) );
  OAI22_X1 U10670 ( .A1(n9495), .A2(n9865), .B1(n9494), .B2(n9863), .ZN(n9497)
         );
  AOI211_X1 U10671 ( .C1(n9860), .C2(n9498), .A(n9497), .B(n9496), .ZN(n9501)
         );
  AOI22_X1 U10672 ( .A1(n9889), .A2(n9501), .B1(n9499), .B2(n9887), .ZN(
        P2_U3533) );
  INV_X1 U10673 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9500) );
  AOI22_X1 U10674 ( .A1(n10073), .A2(n9501), .B1(n9500), .B2(n10071), .ZN(
        P2_U3490) );
  OAI211_X1 U10675 ( .C1(n4613), .C2(n9694), .A(n9503), .B(n9502), .ZN(n9504)
         );
  AOI21_X1 U10676 ( .B1(n9505), .B2(n9700), .A(n9504), .ZN(n9533) );
  AOI22_X1 U10677 ( .A1(n9716), .A2(n9533), .B1(n9047), .B2(n9713), .ZN(
        P1_U3539) );
  INV_X1 U10678 ( .A(n9506), .ZN(n9507) );
  OAI22_X1 U10679 ( .A1(n9508), .A2(n9696), .B1(n9507), .B2(n9694), .ZN(n9509)
         );
  AOI21_X1 U10680 ( .B1(n9510), .B2(n9658), .A(n9509), .ZN(n9511) );
  AND2_X1 U10681 ( .A1(n9512), .A2(n9511), .ZN(n9534) );
  AOI22_X1 U10682 ( .A1(n9716), .A2(n9534), .B1(n9053), .B2(n9713), .ZN(
        P1_U3538) );
  OAI21_X1 U10683 ( .B1(n9514), .B2(n9694), .A(n9513), .ZN(n9515) );
  AOI211_X1 U10684 ( .C1(n9517), .C2(n9700), .A(n9516), .B(n9515), .ZN(n9536)
         );
  AOI22_X1 U10685 ( .A1(n9716), .A2(n9536), .B1(n9518), .B2(n9713), .ZN(
        P1_U3537) );
  OAI22_X1 U10686 ( .A1(n9520), .A2(n9696), .B1(n9519), .B2(n9694), .ZN(n9521)
         );
  AOI21_X1 U10687 ( .B1(n9522), .B2(n9658), .A(n9521), .ZN(n9523) );
  AND2_X1 U10688 ( .A1(n9524), .A2(n9523), .ZN(n9538) );
  AOI22_X1 U10689 ( .A1(n9716), .A2(n9538), .B1(n9525), .B2(n9713), .ZN(
        P1_U3536) );
  OAI22_X1 U10690 ( .A1(n9527), .A2(n9696), .B1(n9526), .B2(n9694), .ZN(n9529)
         );
  AOI211_X1 U10691 ( .C1(n9700), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9540)
         );
  AOI22_X1 U10692 ( .A1(n9716), .A2(n9540), .B1(n9531), .B2(n9713), .ZN(
        P1_U3534) );
  INV_X1 U10693 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9532) );
  AOI22_X1 U10694 ( .A1(n9704), .A2(n9533), .B1(n9532), .B2(n9702), .ZN(
        P1_U3502) );
  INV_X1 U10695 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U10696 ( .A1(n9704), .A2(n9534), .B1(n9994), .B2(n9702), .ZN(
        P1_U3499) );
  INV_X1 U10697 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9535) );
  AOI22_X1 U10698 ( .A1(n9704), .A2(n9536), .B1(n9535), .B2(n9702), .ZN(
        P1_U3496) );
  INV_X1 U10699 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9537) );
  AOI22_X1 U10700 ( .A1(n9704), .A2(n9538), .B1(n9537), .B2(n9702), .ZN(
        P1_U3493) );
  INV_X1 U10701 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9539) );
  AOI22_X1 U10702 ( .A1(n9704), .A2(n9540), .B1(n9539), .B2(n9702), .ZN(
        P1_U3487) );
  XNOR2_X1 U10703 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10704 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10705 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9542), .A(n9541), .ZN(
        n9548) );
  XNOR2_X1 U10706 ( .A(n9543), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9547) );
  AOI22_X1 U10707 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9544), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n9546) );
  NAND3_X1 U10708 ( .A1(n9616), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5141), .ZN(
        n9545) );
  OAI211_X1 U10709 ( .C1(n9548), .C2(n9547), .A(n9546), .B(n9545), .ZN(
        P1_U3241) );
  INV_X1 U10710 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9565) );
  XNOR2_X1 U10711 ( .A(n9550), .B(n9549), .ZN(n9552) );
  AOI22_X1 U10712 ( .A1(n9553), .A2(n9552), .B1(n9628), .B2(n9551), .ZN(n9562)
         );
  INV_X1 U10713 ( .A(n9554), .ZN(n9558) );
  MUX2_X1 U10714 ( .A(n5521), .B(P1_REG1_REG_4__SCAN_IN), .S(n9555), .Z(n9557)
         );
  OAI21_X1 U10715 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9560) );
  AOI21_X1 U10716 ( .B1(n9616), .B2(n9560), .A(n9559), .ZN(n9561) );
  AND2_X1 U10717 ( .A1(n9562), .A2(n9561), .ZN(n9564) );
  OAI211_X1 U10718 ( .C1(n9565), .C2(n9641), .A(n9564), .B(n9563), .ZN(
        P1_U3245) );
  INV_X1 U10719 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U10720 ( .A1(n9567), .A2(n9566), .ZN(n9570) );
  INV_X1 U10721 ( .A(n9568), .ZN(n9569) );
  NAND2_X1 U10722 ( .A1(n9570), .A2(n9569), .ZN(n9575) );
  NAND2_X1 U10723 ( .A1(n9628), .A2(n9571), .ZN(n9574) );
  INV_X1 U10724 ( .A(n9572), .ZN(n9573) );
  OAI211_X1 U10725 ( .C1(n9632), .C2(n9575), .A(n9574), .B(n9573), .ZN(n9576)
         );
  INV_X1 U10726 ( .A(n9576), .ZN(n9582) );
  AOI21_X1 U10727 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9580) );
  OR2_X1 U10728 ( .A1(n9580), .A2(n9638), .ZN(n9581) );
  OAI211_X1 U10729 ( .C1(n9583), .C2(n9641), .A(n9582), .B(n9581), .ZN(
        P1_U3254) );
  INV_X1 U10730 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9593) );
  AOI211_X1 U10731 ( .C1(n7055), .C2(n9585), .A(n9632), .B(n9584), .ZN(n9586)
         );
  AOI211_X1 U10732 ( .C1(n9628), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9592)
         );
  XNOR2_X1 U10733 ( .A(n9589), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U10734 ( .A1(n9590), .A2(n9616), .ZN(n9591) );
  OAI211_X1 U10735 ( .C1(n9593), .C2(n9641), .A(n9592), .B(n9591), .ZN(
        P1_U3256) );
  INV_X1 U10736 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9958) );
  AOI211_X1 U10737 ( .C1(n9596), .C2(n9595), .A(n9594), .B(n9632), .ZN(n9597)
         );
  AOI211_X1 U10738 ( .C1(n9628), .C2(n9599), .A(n9598), .B(n9597), .ZN(n9604)
         );
  OAI211_X1 U10739 ( .C1(n9602), .C2(n9601), .A(n9616), .B(n9600), .ZN(n9603)
         );
  OAI211_X1 U10740 ( .C1(n9958), .C2(n9641), .A(n9604), .B(n9603), .ZN(
        P1_U3257) );
  INV_X1 U10741 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U10742 ( .A1(n9606), .A2(n9605), .ZN(n9609) );
  INV_X1 U10743 ( .A(n9607), .ZN(n9608) );
  NAND2_X1 U10744 ( .A1(n9609), .A2(n9608), .ZN(n9613) );
  NAND2_X1 U10745 ( .A1(n9628), .A2(n9610), .ZN(n9612) );
  OAI211_X1 U10746 ( .C1(n9632), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9614)
         );
  INV_X1 U10747 ( .A(n9614), .ZN(n9620) );
  OAI211_X1 U10748 ( .C1(n9618), .C2(n9617), .A(n9616), .B(n9615), .ZN(n9619)
         );
  OAI211_X1 U10749 ( .C1(n9621), .C2(n9641), .A(n9620), .B(n9619), .ZN(
        P1_U3258) );
  INV_X1 U10750 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U10751 ( .A1(n9623), .A2(n9622), .ZN(n9626) );
  INV_X1 U10752 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U10753 ( .A1(n9626), .A2(n9625), .ZN(n9631) );
  NAND2_X1 U10754 ( .A1(n9628), .A2(n9627), .ZN(n9630) );
  OAI211_X1 U10755 ( .C1(n9632), .C2(n9631), .A(n9630), .B(n9629), .ZN(n9633)
         );
  INV_X1 U10756 ( .A(n9633), .ZN(n9640) );
  AOI21_X1 U10757 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9637) );
  OR2_X1 U10758 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  OAI211_X1 U10759 ( .C1(n9642), .C2(n9641), .A(n9640), .B(n9639), .ZN(
        P1_U3259) );
  NAND2_X1 U10760 ( .A1(n9643), .A2(n9648), .ZN(n9645) );
  AND2_X1 U10761 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9645), .ZN(P1_U3292) );
  AND2_X1 U10762 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9645), .ZN(P1_U3293) );
  AND2_X1 U10763 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9645), .ZN(P1_U3294) );
  INV_X1 U10764 ( .A(n9645), .ZN(n9644) );
  INV_X1 U10765 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U10766 ( .A1(n9644), .A2(n10008), .ZN(P1_U3295) );
  AND2_X1 U10767 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9645), .ZN(P1_U3296) );
  AND2_X1 U10768 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9645), .ZN(P1_U3297) );
  AND2_X1 U10769 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9645), .ZN(P1_U3298) );
  AND2_X1 U10770 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9645), .ZN(P1_U3299) );
  AND2_X1 U10771 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9645), .ZN(P1_U3300) );
  AND2_X1 U10772 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9645), .ZN(P1_U3301) );
  INV_X1 U10773 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U10774 ( .A1(n9644), .A2(n10028), .ZN(P1_U3302) );
  AND2_X1 U10775 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9645), .ZN(P1_U3303) );
  AND2_X1 U10776 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9645), .ZN(P1_U3304) );
  AND2_X1 U10777 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9645), .ZN(P1_U3305) );
  AND2_X1 U10778 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9645), .ZN(P1_U3306) );
  INV_X1 U10779 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9956) );
  NOR2_X1 U10780 ( .A1(n9644), .A2(n9956), .ZN(P1_U3307) );
  AND2_X1 U10781 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9645), .ZN(P1_U3308) );
  AND2_X1 U10782 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9645), .ZN(P1_U3309) );
  AND2_X1 U10783 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9645), .ZN(P1_U3310) );
  INV_X1 U10784 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U10785 ( .A1(n9644), .A2(n9955), .ZN(P1_U3311) );
  AND2_X1 U10786 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9645), .ZN(P1_U3312) );
  INV_X1 U10787 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U10788 ( .A1(n9644), .A2(n10032), .ZN(P1_U3313) );
  AND2_X1 U10789 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9645), .ZN(P1_U3314) );
  AND2_X1 U10790 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9645), .ZN(P1_U3315) );
  AND2_X1 U10791 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9645), .ZN(P1_U3316) );
  AND2_X1 U10792 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9645), .ZN(P1_U3317) );
  AND2_X1 U10793 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9645), .ZN(P1_U3318) );
  AND2_X1 U10794 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9645), .ZN(P1_U3319) );
  AND2_X1 U10795 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9645), .ZN(P1_U3320) );
  AND2_X1 U10796 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9645), .ZN(P1_U3321) );
  INV_X1 U10797 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U10798 ( .A1(n9646), .A2(n9648), .ZN(n9647) );
  OAI21_X1 U10799 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(P1_U3440) );
  INV_X1 U10800 ( .A(n9650), .ZN(n9652) );
  OAI211_X1 U10801 ( .C1(n9654), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9655)
         );
  NOR2_X1 U10802 ( .A1(n9656), .A2(n9655), .ZN(n9705) );
  INV_X1 U10803 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9657) );
  AOI22_X1 U10804 ( .A1(n9704), .A2(n9705), .B1(n9657), .B2(n9702), .ZN(
        P1_U3457) );
  NAND2_X1 U10805 ( .A1(n9659), .A2(n9658), .ZN(n9661) );
  OAI211_X1 U10806 ( .C1(n9662), .C2(n9694), .A(n9661), .B(n9660), .ZN(n9663)
         );
  NOR2_X1 U10807 ( .A1(n9664), .A2(n9663), .ZN(n9707) );
  INV_X1 U10808 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9665) );
  AOI22_X1 U10809 ( .A1(n9704), .A2(n9707), .B1(n9665), .B2(n9702), .ZN(
        P1_U3460) );
  OAI211_X1 U10810 ( .C1(n9668), .C2(n9694), .A(n9667), .B(n9666), .ZN(n9670)
         );
  AOI211_X1 U10811 ( .C1(n9700), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9708)
         );
  AOI22_X1 U10812 ( .A1(n9704), .A2(n9708), .B1(n5544), .B2(n9702), .ZN(
        P1_U3469) );
  AOI21_X1 U10813 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9675) );
  OAI211_X1 U10814 ( .C1(n9678), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9679)
         );
  INV_X1 U10815 ( .A(n9679), .ZN(n9710) );
  INV_X1 U10816 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9680) );
  AOI22_X1 U10817 ( .A1(n9704), .A2(n9710), .B1(n9680), .B2(n9702), .ZN(
        P1_U3472) );
  OAI21_X1 U10818 ( .B1(n9682), .B2(n9694), .A(n9681), .ZN(n9684) );
  AOI211_X1 U10819 ( .C1(n9700), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9711)
         );
  INV_X1 U10820 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9686) );
  AOI22_X1 U10821 ( .A1(n9704), .A2(n9711), .B1(n9686), .B2(n9702), .ZN(
        P1_U3475) );
  INV_X1 U10822 ( .A(n9687), .ZN(n9688) );
  OAI21_X1 U10823 ( .B1(n9689), .B2(n9696), .A(n9688), .ZN(n9690) );
  AOI211_X1 U10824 ( .C1(n9692), .C2(n9700), .A(n9691), .B(n9690), .ZN(n9712)
         );
  INV_X1 U10825 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9693) );
  AOI22_X1 U10826 ( .A1(n9704), .A2(n9712), .B1(n9693), .B2(n9702), .ZN(
        P1_U3478) );
  OAI22_X1 U10827 ( .A1(n9697), .A2(n9696), .B1(n9695), .B2(n9694), .ZN(n9699)
         );
  AOI211_X1 U10828 ( .C1(n9701), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9715)
         );
  INV_X1 U10829 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9703) );
  AOI22_X1 U10830 ( .A1(n9704), .A2(n9715), .B1(n9703), .B2(n9702), .ZN(
        P1_U3481) );
  AOI22_X1 U10831 ( .A1(n9716), .A2(n9705), .B1(n5264), .B2(n9713), .ZN(
        P1_U3524) );
  INV_X1 U10832 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9706) );
  AOI22_X1 U10833 ( .A1(n9716), .A2(n9707), .B1(n9706), .B2(n9713), .ZN(
        P1_U3525) );
  AOI22_X1 U10834 ( .A1(n9716), .A2(n9708), .B1(n5545), .B2(n9713), .ZN(
        P1_U3528) );
  AOI22_X1 U10835 ( .A1(n9716), .A2(n9710), .B1(n9709), .B2(n9713), .ZN(
        P1_U3529) );
  AOI22_X1 U10836 ( .A1(n9716), .A2(n9711), .B1(n5859), .B2(n9713), .ZN(
        P1_U3530) );
  AOI22_X1 U10837 ( .A1(n9716), .A2(n9712), .B1(n5960), .B2(n9713), .ZN(
        P1_U3531) );
  AOI22_X1 U10838 ( .A1(n9716), .A2(n9715), .B1(n9714), .B2(n9713), .ZN(
        P1_U3532) );
  OAI211_X1 U10839 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n9730), .ZN(n9727)
         );
  AOI22_X1 U10840 ( .A1(n9721), .A2(n9720), .B1(P2_U3152), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n9726) );
  AOI22_X1 U10841 ( .A1(n9724), .A2(n9723), .B1(n9748), .B2(n9722), .ZN(n9725)
         );
  AND3_X1 U10842 ( .A1(n9727), .A2(n9726), .A3(n9725), .ZN(n9728) );
  OAI21_X1 U10843 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n9752), .A(n9728), .ZN(
        P2_U3220) );
  AOI22_X1 U10844 ( .A1(n9741), .A2(n9729), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n9738) );
  OAI211_X1 U10845 ( .C1(n6400), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9733)
         );
  OAI21_X1 U10846 ( .B1(n9735), .B2(n9734), .A(n9733), .ZN(n9736) );
  INV_X1 U10847 ( .A(n9736), .ZN(n9737) );
  OAI211_X1 U10848 ( .C1(n9752), .C2(n9739), .A(n9738), .B(n9737), .ZN(
        P2_U3223) );
  AOI22_X1 U10849 ( .A1(n9741), .A2(n9740), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n9750) );
  NAND2_X1 U10850 ( .A1(n9743), .A2(n9742), .ZN(n9745) );
  AOI21_X1 U10851 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9747) );
  AOI21_X1 U10852 ( .B1(n9748), .B2(n9877), .A(n9747), .ZN(n9749) );
  OAI211_X1 U10853 ( .C1(n9752), .C2(n9751), .A(n9750), .B(n9749), .ZN(
        P2_U3241) );
  AOI22_X1 U10854 ( .A1(n4352), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9753), .ZN(n9763) );
  AOI22_X1 U10855 ( .A1(n9754), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9762) );
  NAND2_X1 U10856 ( .A1(n4352), .A2(n9755), .ZN(n9758) );
  OAI211_X1 U10857 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9759), .A(n9758), .B(
        n9757), .ZN(n9760) );
  NAND2_X1 U10858 ( .A1(n9760), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9761) );
  OAI211_X1 U10859 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9763), .A(n9762), .B(
        n9761), .ZN(P2_U3245) );
  INV_X1 U10860 ( .A(n9764), .ZN(n9767) );
  INV_X1 U10861 ( .A(n9765), .ZN(n9864) );
  OAI21_X1 U10862 ( .B1(n9767), .B2(n9864), .A(n9766), .ZN(n9866) );
  INV_X1 U10863 ( .A(n9866), .ZN(n9768) );
  AOI22_X1 U10864 ( .A1(n9768), .A2(n9809), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n9813), .ZN(n9786) );
  XNOR2_X1 U10865 ( .A(n9769), .B(n9773), .ZN(n9869) );
  NAND2_X1 U10866 ( .A1(n9869), .A2(n9770), .ZN(n9781) );
  OAI211_X1 U10867 ( .C1(n9774), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9780)
         );
  AOI22_X1 U10868 ( .A1(n9778), .A2(n9777), .B1(n9776), .B2(n9775), .ZN(n9779)
         );
  AND2_X1 U10869 ( .A1(n9780), .A2(n9779), .ZN(n9862) );
  OAI211_X1 U10870 ( .C1(n9864), .C2(n9782), .A(n9781), .B(n9862), .ZN(n9784)
         );
  NAND2_X1 U10871 ( .A1(n9784), .A2(n9783), .ZN(n9785) );
  OAI211_X1 U10872 ( .C1(n9788), .C2(n9787), .A(n9786), .B(n9785), .ZN(
        P2_U3285) );
  OAI21_X1 U10873 ( .B1(n4342), .B2(n9797), .A(n9789), .ZN(n9859) );
  INV_X1 U10874 ( .A(n9790), .ZN(n9800) );
  NAND2_X1 U10875 ( .A1(n9792), .A2(n9791), .ZN(n9796) );
  INV_X1 U10876 ( .A(n9793), .ZN(n9794) );
  AOI211_X1 U10877 ( .C1(n9797), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9798)
         );
  AOI211_X1 U10878 ( .C1(n9859), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9856)
         );
  AOI222_X1 U10879 ( .A1(n9804), .A2(n9803), .B1(P2_REG2_REG_9__SCAN_IN), .B2(
        n9813), .C1(n9802), .C2(n9801), .ZN(n9812) );
  INV_X1 U10880 ( .A(n9805), .ZN(n9806) );
  OAI21_X1 U10881 ( .B1(n9854), .B2(n9807), .A(n9806), .ZN(n9855) );
  INV_X1 U10882 ( .A(n9855), .ZN(n9808) );
  AOI22_X1 U10883 ( .A1(n9859), .A2(n9810), .B1(n9809), .B2(n9808), .ZN(n9811)
         );
  OAI211_X1 U10884 ( .C1(n9813), .C2(n9856), .A(n9812), .B(n9811), .ZN(
        P2_U3287) );
  NOR2_X1 U10885 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  AND2_X1 U10886 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9819), .ZN(P2_U3297) );
  AND2_X1 U10887 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9819), .ZN(P2_U3298) );
  INV_X1 U10888 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U10889 ( .A1(n9816), .A2(n10052), .ZN(P2_U3299) );
  INV_X1 U10890 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U10891 ( .A1(n9816), .A2(n10029), .ZN(P2_U3300) );
  AND2_X1 U10892 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9819), .ZN(P2_U3301) );
  AND2_X1 U10893 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9819), .ZN(P2_U3302) );
  AND2_X1 U10894 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9819), .ZN(P2_U3303) );
  AND2_X1 U10895 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9819), .ZN(P2_U3304) );
  AND2_X1 U10896 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9819), .ZN(P2_U3305) );
  AND2_X1 U10897 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9819), .ZN(P2_U3306) );
  AND2_X1 U10898 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9819), .ZN(P2_U3307) );
  AND2_X1 U10899 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9819), .ZN(P2_U3308) );
  AND2_X1 U10900 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9819), .ZN(P2_U3309) );
  AND2_X1 U10901 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9819), .ZN(P2_U3310) );
  AND2_X1 U10902 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9819), .ZN(P2_U3311) );
  AND2_X1 U10903 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9819), .ZN(P2_U3312) );
  AND2_X1 U10904 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9819), .ZN(P2_U3313) );
  INV_X1 U10905 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U10906 ( .A1(n9816), .A2(n10051), .ZN(P2_U3314) );
  AND2_X1 U10907 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9819), .ZN(P2_U3315) );
  AND2_X1 U10908 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9819), .ZN(P2_U3316) );
  INV_X1 U10909 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U10910 ( .A1(n9816), .A2(n9990), .ZN(P2_U3317) );
  AND2_X1 U10911 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9819), .ZN(P2_U3318) );
  AND2_X1 U10912 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9819), .ZN(P2_U3319) );
  AND2_X1 U10913 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9819), .ZN(P2_U3320) );
  AND2_X1 U10914 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9819), .ZN(P2_U3321) );
  AND2_X1 U10915 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9819), .ZN(P2_U3322) );
  AND2_X1 U10916 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9819), .ZN(P2_U3323) );
  AND2_X1 U10917 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9819), .ZN(P2_U3324) );
  AND2_X1 U10918 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9819), .ZN(P2_U3325) );
  INV_X1 U10919 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U10920 ( .A1(n9816), .A2(n10026), .ZN(P2_U3326) );
  AOI22_X1 U10921 ( .A1(n9818), .A2(n9821), .B1(n9817), .B2(n9819), .ZN(
        P2_U3437) );
  AOI22_X1 U10922 ( .A1(n9822), .A2(n9821), .B1(n9820), .B2(n9819), .ZN(
        P2_U3438) );
  OAI22_X1 U10923 ( .A1(n9825), .A2(n9829), .B1(n9824), .B2(n9823), .ZN(n9826)
         );
  NOR2_X1 U10924 ( .A1(n9827), .A2(n9826), .ZN(n9871) );
  INV_X1 U10925 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10926 ( .A1(n10073), .A2(n9871), .B1(n9828), .B2(n10071), .ZN(
        P2_U3451) );
  INV_X1 U10927 ( .A(n9829), .ZN(n9883) );
  OAI21_X1 U10928 ( .B1(n9831), .B2(n9863), .A(n9830), .ZN(n9833) );
  AOI211_X1 U10929 ( .C1(n9883), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9872)
         );
  INV_X1 U10930 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9835) );
  AOI22_X1 U10931 ( .A1(n10073), .A2(n9872), .B1(n9835), .B2(n10071), .ZN(
        P2_U3454) );
  OAI22_X1 U10932 ( .A1(n9837), .A2(n9865), .B1(n9836), .B2(n9863), .ZN(n9839)
         );
  AOI211_X1 U10933 ( .C1(n9860), .C2(n9840), .A(n9839), .B(n9838), .ZN(n9873)
         );
  INV_X1 U10934 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U10935 ( .A1(n10073), .A2(n9873), .B1(n9841), .B2(n10071), .ZN(
        P2_U3460) );
  OAI211_X1 U10936 ( .C1(n9844), .C2(n9863), .A(n9843), .B(n9842), .ZN(n9845)
         );
  AOI21_X1 U10937 ( .B1(n9883), .B2(n9846), .A(n9845), .ZN(n9875) );
  INV_X1 U10938 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U10939 ( .A1(n10073), .A2(n9875), .B1(n9847), .B2(n10071), .ZN(
        P2_U3466) );
  OAI22_X1 U10940 ( .A1(n9849), .A2(n9865), .B1(n9848), .B2(n9863), .ZN(n9850)
         );
  AOI211_X1 U10941 ( .C1(n9852), .C2(n9883), .A(n9851), .B(n9850), .ZN(n9885)
         );
  INV_X1 U10942 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U10943 ( .A1(n10073), .A2(n9885), .B1(n9853), .B2(n10071), .ZN(
        P2_U3472) );
  OAI22_X1 U10944 ( .A1(n9855), .A2(n9865), .B1(n9854), .B2(n9863), .ZN(n9858)
         );
  INV_X1 U10945 ( .A(n9856), .ZN(n9857) );
  AOI211_X1 U10946 ( .C1(n9860), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9886)
         );
  INV_X1 U10947 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U10948 ( .A1(n10073), .A2(n9886), .B1(n9861), .B2(n10071), .ZN(
        P2_U3478) );
  INV_X1 U10949 ( .A(n9862), .ZN(n9868) );
  OAI22_X1 U10950 ( .A1(n9866), .A2(n9865), .B1(n9864), .B2(n9863), .ZN(n9867)
         );
  AOI211_X1 U10951 ( .C1(n9869), .C2(n9883), .A(n9868), .B(n9867), .ZN(n9888)
         );
  INV_X1 U10952 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U10953 ( .A1(n10073), .A2(n9888), .B1(n10038), .B2(n10071), .ZN(
        P2_U3484) );
  AOI22_X1 U10954 ( .A1(n9889), .A2(n9871), .B1(n9870), .B2(n9887), .ZN(
        P2_U3520) );
  AOI22_X1 U10955 ( .A1(n9889), .A2(n9872), .B1(n6081), .B2(n9887), .ZN(
        P2_U3521) );
  AOI22_X1 U10956 ( .A1(n9889), .A2(n9873), .B1(n10016), .B2(n9887), .ZN(
        P2_U3523) );
  AOI22_X1 U10957 ( .A1(n9889), .A2(n9875), .B1(n9874), .B2(n9887), .ZN(
        P2_U3525) );
  AOI22_X1 U10958 ( .A1(n9879), .A2(n9878), .B1(n9877), .B2(n9876), .ZN(n9880)
         );
  NAND2_X1 U10959 ( .A1(n9881), .A2(n9880), .ZN(n9882) );
  AOI21_X1 U10960 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n10070) );
  AOI22_X1 U10961 ( .A1(n9889), .A2(n10070), .B1(n6080), .B2(n9887), .ZN(
        P2_U3526) );
  AOI22_X1 U10962 ( .A1(n9889), .A2(n9885), .B1(n6078), .B2(n9887), .ZN(
        P2_U3527) );
  AOI22_X1 U10963 ( .A1(n9889), .A2(n9886), .B1(n6077), .B2(n9887), .ZN(
        P2_U3529) );
  AOI22_X1 U10964 ( .A1(n9889), .A2(n9888), .B1(n6075), .B2(n9887), .ZN(
        P2_U3531) );
  INV_X1 U10965 ( .A(n9890), .ZN(n9891) );
  NAND2_X1 U10966 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  XNOR2_X1 U10967 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9893), .ZN(ADD_1071_U5) );
  INV_X1 U10968 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9964) );
  INV_X1 U10969 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9894) );
  AOI22_X1 U10970 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9964), .B2(n9894), .ZN(ADD_1071_U46) );
  OAI21_X1 U10971 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(ADD_1071_U56) );
  OAI21_X1 U10972 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(ADD_1071_U57) );
  OAI21_X1 U10973 ( .B1(n9903), .B2(n9902), .A(n9901), .ZN(ADD_1071_U58) );
  OAI21_X1 U10974 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(ADD_1071_U59) );
  OAI21_X1 U10975 ( .B1(n9909), .B2(n9908), .A(n9907), .ZN(ADD_1071_U60) );
  OAI21_X1 U10976 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(ADD_1071_U61) );
  AOI21_X1 U10977 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(ADD_1071_U62) );
  AOI21_X1 U10978 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(ADD_1071_U63) );
  NAND2_X1 U10979 ( .A1(keyinput13), .A2(keyinput56), .ZN(n9922) );
  NOR3_X1 U10980 ( .A1(keyinput25), .A2(keyinput51), .A3(keyinput23), .ZN(
        n9920) );
  NOR3_X1 U10981 ( .A1(keyinput45), .A2(keyinput57), .A3(keyinput50), .ZN(
        n9919) );
  NAND4_X1 U10982 ( .A1(keyinput2), .A2(n9920), .A3(keyinput35), .A4(n9919), 
        .ZN(n9921) );
  NOR4_X1 U10983 ( .A1(keyinput58), .A2(keyinput38), .A3(n9922), .A4(n9921), 
        .ZN(n9924) );
  INV_X1 U10984 ( .A(keyinput20), .ZN(n9923) );
  NAND4_X1 U10985 ( .A1(keyinput21), .A2(keyinput33), .A3(n9924), .A4(n9923), 
        .ZN(n9949) );
  NOR3_X1 U10986 ( .A1(keyinput54), .A2(keyinput30), .A3(keyinput36), .ZN(
        n9947) );
  NOR2_X1 U10987 ( .A1(keyinput52), .A2(keyinput3), .ZN(n9925) );
  NAND3_X1 U10988 ( .A1(keyinput47), .A2(keyinput53), .A3(n9925), .ZN(n9929)
         );
  NOR2_X1 U10989 ( .A1(keyinput34), .A2(keyinput48), .ZN(n9926) );
  NAND3_X1 U10990 ( .A1(keyinput39), .A2(keyinput17), .A3(n9926), .ZN(n9928)
         );
  NAND3_X1 U10991 ( .A1(keyinput37), .A2(keyinput32), .A3(keyinput62), .ZN(
        n9927) );
  NOR4_X1 U10992 ( .A1(keyinput41), .A2(n9929), .A3(n9928), .A4(n9927), .ZN(
        n9946) );
  NOR2_X1 U10993 ( .A1(keyinput49), .A2(keyinput19), .ZN(n9935) );
  NAND2_X1 U10994 ( .A1(keyinput31), .A2(keyinput14), .ZN(n9933) );
  NOR3_X1 U10995 ( .A1(keyinput27), .A2(keyinput4), .A3(keyinput5), .ZN(n9931)
         );
  NOR3_X1 U10996 ( .A1(keyinput10), .A2(keyinput44), .A3(keyinput12), .ZN(
        n9930) );
  NAND4_X1 U10997 ( .A1(keyinput26), .A2(n9931), .A3(keyinput18), .A4(n9930), 
        .ZN(n9932) );
  NOR4_X1 U10998 ( .A1(keyinput29), .A2(keyinput15), .A3(n9933), .A4(n9932), 
        .ZN(n9934) );
  NAND4_X1 U10999 ( .A1(keyinput9), .A2(keyinput46), .A3(n9935), .A4(n9934), 
        .ZN(n9944) );
  NOR2_X1 U11000 ( .A1(keyinput16), .A2(keyinput43), .ZN(n9936) );
  NAND3_X1 U11001 ( .A1(keyinput28), .A2(keyinput63), .A3(n9936), .ZN(n9943)
         );
  INV_X1 U11002 ( .A(keyinput40), .ZN(n9937) );
  NAND4_X1 U11003 ( .A1(keyinput0), .A2(keyinput42), .A3(keyinput11), .A4(
        n9937), .ZN(n9942) );
  NOR2_X1 U11004 ( .A1(keyinput6), .A2(keyinput24), .ZN(n9940) );
  INV_X1 U11005 ( .A(keyinput7), .ZN(n9938) );
  NOR4_X1 U11006 ( .A1(keyinput61), .A2(keyinput22), .A3(keyinput1), .A4(n9938), .ZN(n9939) );
  NAND4_X1 U11007 ( .A1(keyinput59), .A2(keyinput55), .A3(n9940), .A4(n9939), 
        .ZN(n9941) );
  NOR4_X1 U11008 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9945)
         );
  NAND4_X1 U11009 ( .A1(keyinput8), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(
        n9948) );
  OAI21_X1 U11010 ( .B1(n9949), .B2(n9948), .A(keyinput60), .ZN(n10069) );
  AOI22_X1 U11011 ( .A1(keyinput21), .A2(P1_U3084), .B1(keyinput60), .B2(n6612), .ZN(n9950) );
  OAI21_X1 U11012 ( .B1(n4258), .B2(keyinput21), .A(n9950), .ZN(n9962) );
  AOI22_X1 U11013 ( .A1(n9953), .A2(keyinput20), .B1(keyinput13), .B2(n9952), 
        .ZN(n9951) );
  OAI221_X1 U11014 ( .B1(n9953), .B2(keyinput20), .C1(n9952), .C2(keyinput13), 
        .A(n9951), .ZN(n9961) );
  AOI22_X1 U11015 ( .A1(n9956), .A2(keyinput58), .B1(keyinput56), .B2(n9955), 
        .ZN(n9954) );
  OAI221_X1 U11016 ( .B1(n9956), .B2(keyinput58), .C1(n9955), .C2(keyinput56), 
        .A(n9954), .ZN(n9960) );
  AOI22_X1 U11017 ( .A1(n9047), .A2(keyinput38), .B1(keyinput2), .B2(n9958), 
        .ZN(n9957) );
  OAI221_X1 U11018 ( .B1(n9047), .B2(keyinput38), .C1(n9958), .C2(keyinput2), 
        .A(n9957), .ZN(n9959) );
  NOR4_X1 U11019 ( .A1(n9962), .A2(n9961), .A3(n9960), .A4(n9959), .ZN(n10006)
         );
  AOI22_X1 U11020 ( .A1(n9965), .A2(keyinput50), .B1(keyinput34), .B2(n9964), 
        .ZN(n9963) );
  OAI221_X1 U11021 ( .B1(n9965), .B2(keyinput50), .C1(n9964), .C2(keyinput34), 
        .A(n9963), .ZN(n9974) );
  XNOR2_X1 U11022 ( .A(keyinput35), .B(n9966), .ZN(n9973) );
  XNOR2_X1 U11023 ( .A(keyinput57), .B(n5681), .ZN(n9972) );
  XNOR2_X1 U11024 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput25), .ZN(n9970)
         );
  XNOR2_X1 U11025 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput51), .ZN(n9969) );
  XNOR2_X1 U11026 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput45), .ZN(n9968) );
  XNOR2_X1 U11027 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput23), .ZN(n9967) );
  NAND4_X1 U11028 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n9967), .ZN(n9971)
         );
  NOR4_X1 U11029 ( .A1(n9974), .A2(n9973), .A3(n9972), .A4(n9971), .ZN(n10005)
         );
  AOI22_X1 U11030 ( .A1(n9976), .A2(keyinput3), .B1(keyinput47), .B2(n5680), 
        .ZN(n9975) );
  OAI221_X1 U11031 ( .B1(n9976), .B2(keyinput3), .C1(n5680), .C2(keyinput47), 
        .A(n9975), .ZN(n9987) );
  AOI22_X1 U11032 ( .A1(n9979), .A2(keyinput48), .B1(n9978), .B2(keyinput39), 
        .ZN(n9977) );
  OAI221_X1 U11033 ( .B1(n9979), .B2(keyinput48), .C1(n9978), .C2(keyinput39), 
        .A(n9977), .ZN(n9986) );
  XOR2_X1 U11034 ( .A(n9980), .B(keyinput17), .Z(n9984) );
  XOR2_X1 U11035 ( .A(n7055), .B(keyinput41), .Z(n9983) );
  XNOR2_X1 U11036 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput52), .ZN(n9982) );
  XNOR2_X1 U11037 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput53), .ZN(n9981) );
  NAND4_X1 U11038 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(n9985)
         );
  NOR3_X1 U11039 ( .A1(n9987), .A2(n9986), .A3(n9985), .ZN(n10004) );
  AOI22_X1 U11040 ( .A1(n9990), .A2(keyinput37), .B1(keyinput32), .B2(n9989), 
        .ZN(n9988) );
  OAI221_X1 U11041 ( .B1(n9990), .B2(keyinput37), .C1(n9989), .C2(keyinput32), 
        .A(n9988), .ZN(n10002) );
  INV_X1 U11042 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11043 ( .A1(n9993), .A2(keyinput62), .B1(n9992), .B2(keyinput8), 
        .ZN(n9991) );
  OAI221_X1 U11044 ( .B1(n9993), .B2(keyinput62), .C1(n9992), .C2(keyinput8), 
        .A(n9991), .ZN(n10001) );
  XOR2_X1 U11045 ( .A(n9994), .B(keyinput54), .Z(n9999) );
  INV_X1 U11046 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9995) );
  XOR2_X1 U11047 ( .A(n9995), .B(keyinput9), .Z(n9998) );
  XNOR2_X1 U11048 ( .A(SI_2_), .B(keyinput30), .ZN(n9997) );
  XNOR2_X1 U11049 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput36), .ZN(n9996) );
  NAND4_X1 U11050 ( .A1(n9999), .A2(n9998), .A3(n9997), .A4(n9996), .ZN(n10000) );
  NOR3_X1 U11051 ( .A1(n10002), .A2(n10001), .A3(n10000), .ZN(n10003) );
  NAND4_X1 U11052 ( .A1(n10006), .A2(n10005), .A3(n10004), .A4(n10003), .ZN(
        n10068) );
  AOI22_X1 U11053 ( .A1(n9259), .A2(keyinput12), .B1(n10008), .B2(keyinput29), 
        .ZN(n10007) );
  OAI221_X1 U11054 ( .B1(n9259), .B2(keyinput12), .C1(n10008), .C2(keyinput29), 
        .A(n10007), .ZN(n10020) );
  AOI22_X1 U11055 ( .A1(n10011), .A2(keyinput44), .B1(keyinput18), .B2(n10010), 
        .ZN(n10009) );
  OAI221_X1 U11056 ( .B1(n10011), .B2(keyinput44), .C1(n10010), .C2(keyinput18), .A(n10009), .ZN(n10019) );
  INV_X1 U11057 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10014) );
  AOI22_X1 U11058 ( .A1(n10014), .A2(keyinput14), .B1(keyinput16), .B2(n10013), 
        .ZN(n10012) );
  OAI221_X1 U11059 ( .B1(n10014), .B2(keyinput14), .C1(n10013), .C2(keyinput16), .A(n10012), .ZN(n10018) );
  AOI22_X1 U11060 ( .A1(n10016), .A2(keyinput31), .B1(n4507), .B2(keyinput15), 
        .ZN(n10015) );
  OAI221_X1 U11061 ( .B1(n10016), .B2(keyinput31), .C1(n4507), .C2(keyinput15), 
        .A(n10015), .ZN(n10017) );
  NOR4_X1 U11062 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10066) );
  INV_X1 U11063 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10023) );
  AOI22_X1 U11064 ( .A1(n10023), .A2(keyinput46), .B1(keyinput27), .B2(n10022), 
        .ZN(n10021) );
  OAI221_X1 U11065 ( .B1(n10023), .B2(keyinput46), .C1(n10022), .C2(keyinput27), .A(n10021), .ZN(n10036) );
  AOI22_X1 U11066 ( .A1(n10026), .A2(keyinput49), .B1(keyinput19), .B2(n10025), 
        .ZN(n10024) );
  OAI221_X1 U11067 ( .B1(n10026), .B2(keyinput49), .C1(n10025), .C2(keyinput19), .A(n10024), .ZN(n10035) );
  AOI22_X1 U11068 ( .A1(n10029), .A2(keyinput5), .B1(n10028), .B2(keyinput10), 
        .ZN(n10027) );
  OAI221_X1 U11069 ( .B1(n10029), .B2(keyinput5), .C1(n10028), .C2(keyinput10), 
        .A(n10027), .ZN(n10034) );
  AOI22_X1 U11070 ( .A1(n10032), .A2(keyinput4), .B1(keyinput26), .B2(n10031), 
        .ZN(n10030) );
  OAI221_X1 U11071 ( .B1(n10032), .B2(keyinput4), .C1(n10031), .C2(keyinput26), 
        .A(n10030), .ZN(n10033) );
  NOR4_X1 U11072 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(
        n10065) );
  AOI22_X1 U11073 ( .A1(n7318), .A2(keyinput55), .B1(keyinput61), .B2(n10038), 
        .ZN(n10037) );
  OAI221_X1 U11074 ( .B1(n7318), .B2(keyinput55), .C1(n10038), .C2(keyinput61), 
        .A(n10037), .ZN(n10049) );
  INV_X1 U11075 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11076 ( .A1(n10041), .A2(keyinput24), .B1(keyinput59), .B2(n10040), 
        .ZN(n10039) );
  OAI221_X1 U11077 ( .B1(n10041), .B2(keyinput24), .C1(n10040), .C2(keyinput59), .A(n10039), .ZN(n10048) );
  INV_X1 U11078 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10042) );
  XOR2_X1 U11079 ( .A(n10042), .B(keyinput1), .Z(n10046) );
  XNOR2_X1 U11080 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput33), .ZN(n10045) );
  XNOR2_X1 U11081 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput22), .ZN(n10044)
         );
  XNOR2_X1 U11082 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput7), .ZN(n10043) );
  NAND4_X1 U11083 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10047) );
  NOR3_X1 U11084 ( .A1(n10049), .A2(n10048), .A3(n10047), .ZN(n10064) );
  AOI22_X1 U11085 ( .A1(n10052), .A2(keyinput28), .B1(keyinput43), .B2(n10051), 
        .ZN(n10050) );
  OAI221_X1 U11086 ( .B1(n10052), .B2(keyinput28), .C1(n10051), .C2(keyinput43), .A(n10050), .ZN(n10062) );
  AOI22_X1 U11087 ( .A1(n9477), .A2(keyinput63), .B1(n4914), .B2(keyinput42), 
        .ZN(n10053) );
  OAI221_X1 U11088 ( .B1(n9477), .B2(keyinput63), .C1(n4914), .C2(keyinput42), 
        .A(n10053), .ZN(n10061) );
  AOI22_X1 U11089 ( .A1(n10056), .A2(keyinput40), .B1(n10055), .B2(keyinput6), 
        .ZN(n10054) );
  OAI221_X1 U11090 ( .B1(n10056), .B2(keyinput40), .C1(n10055), .C2(keyinput6), 
        .A(n10054), .ZN(n10060) );
  XNOR2_X1 U11091 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput0), .ZN(n10058) );
  XNOR2_X1 U11092 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput11), .ZN(n10057)
         );
  NAND2_X1 U11093 ( .A1(n10058), .A2(n10057), .ZN(n10059) );
  NOR4_X1 U11094 ( .A1(n10062), .A2(n10061), .A3(n10060), .A4(n10059), .ZN(
        n10063) );
  NAND4_X1 U11095 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10067) );
  AOI211_X1 U11096 ( .C1(P1_REG3_REG_13__SCAN_IN), .C2(n10069), .A(n10068), 
        .B(n10067), .ZN(n10075) );
  INV_X1 U11097 ( .A(n10070), .ZN(n10072) );
  AOI22_X1 U11098 ( .A1(n10073), .A2(n10072), .B1(P2_REG0_REG_6__SCAN_IN), 
        .B2(n10071), .ZN(n10074) );
  XNOR2_X1 U11099 ( .A(n10075), .B(n10074), .ZN(P2_U3469) );
  XOR2_X1 U11100 ( .A(n10076), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11101 ( .A(n10077), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  NOR2_X1 U11102 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  XOR2_X1 U11103 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10080), .Z(ADD_1071_U51) );
  XOR2_X1 U11104 ( .A(n10081), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11105 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10085) );
  XNOR2_X1 U11106 ( .A(n10085), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11107 ( .A(n10087), .B(n10086), .Z(ADD_1071_U54) );
  AOI21_X1 U11108 ( .B1(n10090), .B2(n10089), .A(n10088), .ZN(ADD_1071_U47) );
  XOR2_X1 U11109 ( .A(n10092), .B(n10091), .Z(ADD_1071_U53) );
  XNOR2_X1 U11110 ( .A(n10094), .B(n10093), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4778 ( .A(n5533), .Z(n8758) );
  CLKBUF_X1 U4788 ( .A(n5348), .Z(n4259) );
  INV_X2 U6188 ( .A(n9364), .ZN(n6776) );
endmodule

