

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9597, n9598, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670;

  INV_X1 U11028 ( .A(n19641), .ZN(n19713) );
  NOR2_X1 U11029 ( .A1(n13809), .A2(n13816), .ZN(n13808) );
  INV_X1 U11030 ( .A(n18294), .ZN(n17806) );
  NAND2_X1 U11031 ( .A1(n12769), .A2(n12768), .ZN(n13406) );
  BUF_X2 U11032 ( .A(n15259), .Z(n16619) );
  INV_X1 U11034 ( .A(n9585), .ZN(n15236) );
  CLKBUF_X1 U11035 ( .A(n14956), .Z(n9588) );
  CLKBUF_X2 U11036 ( .A(n15067), .Z(n16804) );
  CLKBUF_X1 U11037 ( .A(n15067), .Z(n16786) );
  CLKBUF_X1 U11038 ( .A(n15274), .Z(n15251) );
  INV_X1 U11039 ( .A(n15188), .ZN(n16797) );
  CLKBUF_X1 U11040 ( .A(n15259), .Z(n16801) );
  BUF_X1 U11041 ( .A(n14956), .Z(n9587) );
  CLKBUF_X2 U11042 ( .A(n11570), .Z(n9593) );
  AND2_X1 U11043 ( .A1(n10754), .A2(n15934), .ZN(n10455) );
  CLKBUF_X2 U11044 ( .A(n10253), .Z(n10752) );
  INV_X1 U11045 ( .A(n11907), .ZN(n10095) );
  CLKBUF_X2 U11046 ( .A(n11688), .Z(n11760) );
  AND2_X1 U11047 ( .A1(n11025), .A2(n11022), .ZN(n11537) );
  BUF_X2 U11048 ( .A(n11634), .Z(n11820) );
  BUF_X1 U11049 ( .A(n11040), .Z(n11775) );
  AND2_X1 U11050 ( .A1(n11023), .A2(n12483), .ZN(n11634) );
  AND2_X1 U11051 ( .A1(n11022), .A2(n14111), .ZN(n11040) );
  CLKBUF_X2 U11052 ( .A(n10278), .Z(n10294) );
  INV_X4 U11053 ( .A(n17712), .ZN(n9597) );
  AND2_X2 U11054 ( .A1(n14111), .A2(n12484), .ZN(n11707) );
  OAI21_X1 U11055 ( .B1(n9894), .B2(n12426), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11150) );
  NOR2_X1 U11056 ( .A1(n11296), .A2(n20401), .ZN(n11898) );
  CLKBUF_X2 U11057 ( .A(n10390), .Z(n9608) );
  INV_X1 U11059 ( .A(n10524), .ZN(n10957) );
  INV_X1 U11061 ( .A(n9645), .ZN(n14160) );
  NAND2_X1 U11062 ( .A1(n10207), .A2(n15934), .ZN(n10208) );
  NOR3_X2 U11063 ( .A1(n17321), .A2(n17323), .A3(n17308), .ZN(n17281) );
  CLKBUF_X2 U11064 ( .A(n14956), .Z(n9586) );
  NAND2_X1 U11065 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18425), .ZN(
        n14943) );
  NAND2_X1 U11066 ( .A1(n11907), .A2(n12469), .ZN(n13702) );
  AND4_X1 U11068 ( .A1(n11124), .A2(n11123), .A3(n11122), .A4(n11121), .ZN(
        n11140) );
  INV_X1 U11069 ( .A(n12416), .ZN(n19875) );
  AOI21_X1 U11070 ( .B1(n10999), .B2(n14185), .A(n14164), .ZN(n14635) );
  INV_X1 U11072 ( .A(n12889), .ZN(n19871) );
  NAND2_X1 U11073 ( .A1(n12697), .A2(n12696), .ZN(n13098) );
  INV_X1 U11075 ( .A(n12719), .ZN(n12734) );
  CLKBUF_X3 U11076 ( .A(n10160), .Z(n19592) );
  NAND2_X1 U11077 ( .A1(n17689), .A2(n17594), .ZN(n17631) );
  INV_X1 U11078 ( .A(n17488), .ZN(n17457) );
  INV_X1 U11079 ( .A(n18861), .ZN(n18859) );
  INV_X1 U11080 ( .A(n19667), .ZN(n15480) );
  OR3_X1 U11081 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18425), .A3(
        n18299), .ZN(n9584) );
  AND2_X2 U11082 ( .A1(n10246), .A2(n10245), .ZN(n10160) );
  OR2_X1 U11083 ( .A1(n14946), .A2(n18285), .ZN(n9585) );
  AND2_X2 U11084 ( .A1(n9772), .A2(n12767), .ZN(n12768) );
  AND2_X2 U11085 ( .A1(n9770), .A2(n12746), .ZN(n12769) );
  NOR2_X2 U11086 ( .A1(n17443), .A2(n15290), .ZN(n17428) );
  NAND2_X2 U11087 ( .A1(n10260), .A2(n10259), .ZN(n12779) );
  NOR3_X2 U11088 ( .A1(n17263), .A2(n17557), .A3(n17254), .ZN(n17207) );
  NOR2_X4 U11089 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14922) );
  AOI211_X2 U11090 ( .C1(n15148), .C2(n15147), .A(n15161), .B(n15160), .ZN(
        n15206) );
  INV_X4 U11091 ( .A(n9647), .ZN(n16779) );
  INV_X1 U11092 ( .A(n18884), .ZN(n12777) );
  NOR2_X2 U11093 ( .A1(n12615), .A2(n12855), .ZN(n12845) );
  NOR3_X2 U11094 ( .A1(n16820), .A2(n20629), .A3(n16826), .ZN(n16795) );
  INV_X4 U11095 ( .A(n9646), .ZN(n16800) );
  NAND2_X4 U11096 ( .A1(n10209), .A2(n10208), .ZN(n18913) );
  XNOR2_X2 U11097 ( .A(n11274), .B(n11273), .ZN(n19931) );
  NAND2_X2 U11098 ( .A1(n11219), .A2(n11218), .ZN(n11274) );
  NAND2_X2 U11099 ( .A1(n9731), .A2(n9757), .ZN(n16612) );
  OR2_X1 U11100 ( .A1(n12558), .A2(n9669), .ZN(n13028) );
  NAND2_X1 U11101 ( .A1(n12673), .A2(n10094), .ZN(n12558) );
  AND2_X1 U11102 ( .A1(n14809), .A2(n9698), .ZN(n14797) );
  NOR2_X2 U11103 ( .A1(n16732), .A2(n16757), .ZN(n16746) );
  CLKBUF_X1 U11105 ( .A(n12631), .Z(n20230) );
  BUF_X1 U11106 ( .A(n16496), .Z(n9609) );
  CLKBUF_X1 U11107 ( .A(n11169), .Z(n11290) );
  NAND2_X1 U11108 ( .A1(n9895), .A2(n11150), .ZN(n11169) );
  NAND2_X1 U11109 ( .A1(n9933), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10329) );
  OR2_X1 U11110 ( .A1(n12421), .A2(n11921), .ZN(n12383) );
  OR2_X1 U11111 ( .A1(n11870), .A2(n11918), .ZN(n12439) );
  NAND2_X1 U11112 ( .A1(n11914), .A2(n11918), .ZN(n13472) );
  BUF_X2 U11113 ( .A(n10294), .Z(n18899) );
  CLKBUF_X2 U11114 ( .A(n11141), .Z(n19883) );
  INV_X2 U11116 ( .A(n16901), .ZN(n17864) );
  INV_X2 U11117 ( .A(n16857), .ZN(n17857) );
  NAND2_X2 U11118 ( .A1(n10160), .A2(n12779), .ZN(n12939) );
  NAND2_X1 U11119 ( .A1(n10182), .A2(n15934), .ZN(n10183) );
  AND4_X1 U11120 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11049) );
  CLKBUF_X2 U11121 ( .A(n11537), .Z(n11659) );
  CLKBUF_X2 U11122 ( .A(n14991), .Z(n16802) );
  CLKBUF_X2 U11123 ( .A(n11298), .Z(n11633) );
  CLKBUF_X2 U11125 ( .A(n10239), .Z(n10226) );
  BUF_X4 U11127 ( .A(n15095), .Z(n9589) );
  INV_X4 U11128 ( .A(n9648), .ZN(n9590) );
  BUF_X4 U11129 ( .A(n15275), .Z(n9591) );
  BUF_X4 U11130 ( .A(n15186), .Z(n9592) );
  AND2_X2 U11131 ( .A1(n14902), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10390) );
  NOR2_X4 U11132 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12483) );
  INV_X2 U11133 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11260) );
  OR2_X1 U11134 ( .A1(n9800), .A2(n9795), .ZN(n9794) );
  AND2_X1 U11135 ( .A1(n9784), .A2(n9783), .ZN(n15750) );
  NAND2_X1 U11136 ( .A1(n9800), .A2(n9798), .ZN(n14442) );
  NAND2_X1 U11137 ( .A1(n14497), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14705) );
  OR2_X1 U11138 ( .A1(n13779), .A2(n9954), .ZN(n9950) );
  INV_X1 U11139 ( .A(n14490), .ZN(n14497) );
  OAI22_X1 U11140 ( .A1(n9953), .A2(n9692), .B1(n9957), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U11141 ( .A1(n10703), .A2(n10701), .ZN(n14263) );
  OR2_X1 U11142 ( .A1(n15771), .A2(n14784), .ZN(n15760) );
  INV_X1 U11143 ( .A(n10703), .ZN(n9910) );
  AND2_X1 U11144 ( .A1(n9884), .A2(n9883), .ZN(n13809) );
  OR2_X1 U11145 ( .A1(n10699), .A2(n10700), .ZN(n10703) );
  AND2_X1 U11146 ( .A1(n9881), .A2(n10117), .ZN(n13816) );
  NAND2_X1 U11147 ( .A1(n13882), .A2(n13881), .ZN(n13880) );
  NAND2_X1 U11148 ( .A1(n9767), .A2(n13423), .ZN(n15801) );
  NAND2_X1 U11149 ( .A1(n10115), .A2(n15515), .ZN(n13882) );
  NAND2_X1 U11150 ( .A1(n13417), .A2(n13416), .ZN(n14588) );
  NAND3_X1 U11151 ( .A1(n9824), .A2(n9825), .A3(n9821), .ZN(n10115) );
  OR2_X1 U11152 ( .A1(n10652), .A2(n10651), .ZN(n10152) );
  NAND2_X1 U11153 ( .A1(n13400), .A2(n9938), .ZN(n14639) );
  NAND2_X1 U11154 ( .A1(n14876), .A2(n14874), .ZN(n14878) );
  NOR3_X2 U11155 ( .A1(n14299), .A2(n9942), .A3(n9939), .ZN(n14268) );
  OR2_X2 U11156 ( .A1(n14308), .A2(n14297), .ZN(n14299) );
  NAND2_X1 U11157 ( .A1(n9776), .A2(n12941), .ZN(n13242) );
  NAND2_X1 U11158 ( .A1(n9835), .A2(n18664), .ZN(n13251) );
  XNOR2_X1 U11159 ( .A(n13419), .B(n13418), .ZN(n13411) );
  NAND2_X1 U11160 ( .A1(n9668), .A2(n9745), .ZN(n9926) );
  AOI21_X1 U11161 ( .B1(n9840), .B2(n9842), .A(n9838), .ZN(n9837) );
  NAND2_X1 U11162 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16625), .ZN(n16605) );
  XNOR2_X1 U11163 ( .A(n13408), .B(n13254), .ZN(n13409) );
  NOR2_X1 U11164 ( .A1(n17144), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17143) );
  AND2_X1 U11165 ( .A1(n13278), .A2(n13277), .ZN(n13418) );
  NAND2_X1 U11166 ( .A1(n10387), .A2(n10386), .ZN(n12673) );
  AND4_X1 U11167 ( .A1(n12748), .A2(n12761), .A3(n12747), .A4(n12764), .ZN(
        n9618) );
  AND3_X1 U11168 ( .A1(n13229), .A2(n13231), .A3(n13230), .ZN(n9769) );
  NAND2_X2 U11169 ( .A1(n13137), .A2(n13136), .ZN(n9615) );
  AND4_X1 U11170 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        n12743) );
  NOR2_X1 U11171 ( .A1(n16901), .A2(n16895), .ZN(n16891) );
  AND4_X1 U11172 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12742) );
  AND2_X1 U11173 ( .A1(n10385), .A2(n10384), .ZN(n10386) );
  OAI21_X1 U11174 ( .B1(n13224), .B2(n12759), .A(n9773), .ZN(n12760) );
  NOR2_X1 U11175 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17176), .ZN(
        n17175) );
  OR2_X1 U11176 ( .A1(n12753), .A2(n12709), .ZN(n12710) );
  NAND2_X1 U11177 ( .A1(n11255), .A2(n11254), .ZN(n11256) );
  AND2_X1 U11178 ( .A1(n17205), .A2(n9743), .ZN(n17263) );
  INV_X1 U11179 ( .A(n17477), .ZN(n17492) );
  OR2_X1 U11180 ( .A1(n12736), .A2(n12723), .ZN(n13224) );
  NAND2_X1 U11181 ( .A1(n11311), .A2(n11310), .ZN(n19992) );
  CLKBUF_X2 U11182 ( .A(n12713), .Z(n12728) );
  AND2_X1 U11183 ( .A1(n11250), .A2(n11249), .ZN(n12504) );
  CLKBUF_X1 U11184 ( .A(n16276), .Z(n16531) );
  NAND2_X1 U11185 ( .A1(n12411), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12679) );
  AND2_X1 U11186 ( .A1(n15907), .A2(n9700), .ZN(n14834) );
  NAND2_X2 U11187 ( .A1(n19728), .A2(n12469), .ZN(n13696) );
  NAND2_X1 U11188 ( .A1(n18690), .A2(n12706), .ZN(n12733) );
  CLKBUF_X1 U11189 ( .A(n12871), .Z(n20111) );
  OAI21_X1 U11190 ( .B1(n19931), .B2(n12689), .A(n12410), .ZN(n12411) );
  AND2_X1 U11191 ( .A1(n16901), .A2(n16856), .ZN(n16996) );
  NAND2_X1 U11192 ( .A1(n10947), .A2(n10946), .ZN(n14860) );
  NOR2_X1 U11193 ( .A1(n15414), .A2(n17060), .ZN(n16940) );
  NAND2_X2 U11194 ( .A1(n10357), .A2(n10356), .ZN(n13035) );
  INV_X1 U11195 ( .A(n10349), .ZN(n10357) );
  AND2_X1 U11196 ( .A1(n12048), .A2(n10338), .ZN(n12050) );
  NAND2_X1 U11197 ( .A1(n19960), .A2(n11243), .ZN(n11246) );
  CLKBUF_X1 U11198 ( .A(n11276), .Z(n19961) );
  AND2_X1 U11199 ( .A1(n10353), .A2(n9932), .ZN(n10349) );
  OR2_X1 U11200 ( .A1(n10337), .A2(n10336), .ZN(n12048) );
  NOR2_X1 U11201 ( .A1(n17410), .A2(n17737), .ZN(n17409) );
  AOI221_X2 U11202 ( .B1(n17834), .B2(n15167), .C1(n17063), .C2(n15167), .A(
        n15163), .ZN(n15412) );
  NOR2_X2 U11203 ( .A1(n18866), .A2(n19162), .ZN(n18867) );
  NOR2_X2 U11204 ( .A1(n18878), .A2(n19162), .ZN(n18879) );
  NOR2_X2 U11205 ( .A1(n18882), .A2(n19162), .ZN(n18883) );
  AOI21_X1 U11206 ( .B1(n11290), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11170), .ZN(n11179) );
  CLKBUF_X2 U11207 ( .A(n18286), .Z(n9600) );
  OAI211_X1 U11208 ( .C1(n13398), .C2(n14614), .A(n10332), .B(n10331), .ZN(
        n10337) );
  OR2_X1 U11209 ( .A1(n10322), .A2(n10333), .ZN(n9932) );
  INV_X1 U11210 ( .A(n10329), .ZN(n10308) );
  CLKBUF_X3 U11211 ( .A(n10329), .Z(n13398) );
  NOR2_X1 U11212 ( .A1(n12780), .A2(n10813), .ZN(n15943) );
  CLKBUF_X1 U11213 ( .A(n10323), .Z(n12803) );
  NAND2_X1 U11214 ( .A1(n17644), .A2(n15295), .ZN(n17359) );
  AOI21_X1 U11215 ( .B1(n14912), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10315), 
        .ZN(n10316) );
  NAND2_X1 U11216 ( .A1(n15149), .A2(n18280), .ZN(n15200) );
  AND2_X1 U11217 ( .A1(n12280), .A2(n12279), .ZN(n12282) );
  OAI22_X1 U11218 ( .A1(n17465), .A2(n10016), .B1(n10019), .B2(n15288), .ZN(
        n17445) );
  OAI22_X1 U11219 ( .A1(n10836), .A2(n18868), .B1(n10282), .B2(n12805), .ZN(
        n10291) );
  OR2_X1 U11220 ( .A1(n12022), .A2(n12254), .ZN(n10301) );
  NAND2_X1 U11221 ( .A1(n12374), .A2(n12383), .ZN(n12426) );
  AND2_X1 U11222 ( .A1(n10814), .A2(n10273), .ZN(n9904) );
  NAND2_X1 U11223 ( .A1(n10038), .A2(n11143), .ZN(n11849) );
  OR2_X1 U11224 ( .A1(n12470), .A2(n11149), .ZN(n12456) );
  AND2_X1 U11225 ( .A1(n11120), .A2(n19871), .ZN(n10100) );
  NAND2_X1 U11226 ( .A1(n10274), .A2(n10297), .ZN(n12787) );
  AND2_X1 U11227 ( .A1(n10282), .A2(n10261), .ZN(n14916) );
  NOR2_X1 U11228 ( .A1(n10295), .A2(n10294), .ZN(n10296) );
  NOR2_X1 U11229 ( .A1(n15177), .A2(n15148), .ZN(n18279) );
  INV_X2 U11230 ( .A(n16087), .ZN(n16105) );
  NAND2_X1 U11231 ( .A1(n10283), .A2(n11000), .ZN(n12806) );
  NOR2_X1 U11232 ( .A1(n10263), .A2(n10160), .ZN(n10840) );
  AND3_X1 U11233 ( .A1(n18892), .A2(n10278), .A3(n18903), .ZN(n10283) );
  INV_X1 U11234 ( .A(n12429), .ZN(n11141) );
  NAND2_X2 U11235 ( .A1(n9651), .A2(n9617), .ZN(n9919) );
  NAND3_X1 U11236 ( .A1(n17281), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17266) );
  NOR2_X2 U11237 ( .A1(n19851), .A2(n19849), .ZN(n19850) );
  AND4_X1 U11238 ( .A1(n11039), .A2(n11038), .A3(n11037), .A4(n11036), .ZN(
        n11051) );
  AND4_X1 U11239 ( .A1(n11035), .A2(n11034), .A3(n11033), .A4(n11032), .ZN(
        n11052) );
  NAND2_X1 U11240 ( .A1(n10177), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10184) );
  INV_X1 U11241 ( .A(n18888), .ZN(n9594) );
  AND4_X1 U11242 ( .A1(n11115), .A2(n11114), .A3(n11113), .A4(n11112), .ZN(
        n11116) );
  AND4_X1 U11243 ( .A1(n11107), .A2(n11106), .A3(n11105), .A4(n11104), .ZN(
        n11118) );
  AND4_X1 U11244 ( .A1(n11103), .A2(n11102), .A3(n11101), .A4(n11100), .ZN(
        n11119) );
  AND4_X1 U11245 ( .A1(n11136), .A2(n11135), .A3(n11134), .A4(n11133), .ZN(
        n11137) );
  AND4_X1 U11246 ( .A1(n11132), .A2(n11131), .A3(n11130), .A4(n11129), .ZN(
        n11138) );
  AND4_X1 U11247 ( .A1(n11128), .A2(n11127), .A3(n11126), .A4(n11125), .ZN(
        n11139) );
  AND4_X1 U11248 ( .A1(n11044), .A2(n11043), .A3(n11042), .A4(n11041), .ZN(
        n11050) );
  AND4_X1 U11249 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10238) );
  AND4_X1 U11250 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  CLKBUF_X1 U11251 ( .A(n11228), .Z(n11706) );
  AOI21_X1 U11253 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18091), .A(
        n14977), .ZN(n14984) );
  INV_X2 U11254 ( .A(n18355), .ZN(n9595) );
  NAND2_X2 U11255 ( .A1(n18482), .A2(n18349), .ZN(n18395) );
  INV_X2 U11256 ( .A(n15601), .ZN(n12502) );
  INV_X2 U11257 ( .A(n19730), .ZN(n19759) );
  CLKBUF_X2 U11258 ( .A(n11297), .Z(n11639) );
  INV_X2 U11259 ( .A(n15188), .ZN(n16785) );
  NAND2_X2 U11260 ( .A1(n19606), .A2(n19485), .ZN(n19534) );
  BUF_X4 U11262 ( .A(n11040), .Z(n11818) );
  NAND2_X2 U11263 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19606), .ZN(n19531) );
  INV_X2 U11264 ( .A(n16138), .ZN(U215) );
  BUF_X2 U11265 ( .A(n11634), .Z(n11660) );
  NOR2_X1 U11266 ( .A1(n10373), .A2(n19554), .ZN(n19448) );
  NAND3_X1 U11267 ( .A1(n16442), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17421) );
  NOR3_X2 U11268 ( .A1(n18166), .A2(n18091), .A3(n17949), .ZN(n17927) );
  AND2_X1 U11269 ( .A1(n11023), .A2(n11022), .ZN(n11297) );
  AND2_X1 U11270 ( .A1(n11022), .A2(n14110), .ZN(n11688) );
  BUF_X4 U11271 ( .A(n11827), .Z(n9598) );
  BUF_X4 U11272 ( .A(n10390), .Z(n9607) );
  BUF_X2 U11274 ( .A(n10390), .Z(n9606) );
  OR2_X1 U11275 ( .A1(n18277), .A2(n14946), .ZN(n15188) );
  OR2_X1 U11276 ( .A1(n18299), .A2(n14943), .ZN(n9648) );
  NOR2_X1 U11277 ( .A1(n14946), .A2(n18299), .ZN(n15259) );
  AND2_X1 U11278 ( .A1(n15156), .A2(n15155), .ZN(n14977) );
  OR2_X1 U11279 ( .A1(n14943), .A2(n18285), .ZN(n9647) );
  INV_X2 U11280 ( .A(n16141), .ZN(n16143) );
  AND2_X1 U11281 ( .A1(n12495), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11024) );
  AND2_X1 U11282 ( .A1(n14914), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9604) );
  NAND2_X1 U11283 ( .A1(n18443), .A2(n18436), .ZN(n18277) );
  NAND2_X1 U11284 ( .A1(n18425), .A2(n18450), .ZN(n14946) );
  NAND2_X1 U11285 ( .A1(n18443), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18285) );
  NAND2_X1 U11286 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18436), .ZN(
        n18283) );
  AND2_X1 U11287 ( .A1(n14112), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11023) );
  AND2_X2 U11288 ( .A1(n14914), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9605) );
  AND2_X1 U11289 ( .A1(n10037), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11022) );
  INV_X1 U11290 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12495) );
  INV_X2 U11291 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18450) );
  NAND2_X2 U11292 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18299) );
  NAND2_X1 U11293 ( .A1(n10267), .A2(n10287), .ZN(n10268) );
  AND2_X1 U11294 ( .A1(n11023), .A2(n11024), .ZN(n11570) );
  XNOR2_X2 U11295 ( .A(n14460), .B(n14459), .ZN(n14658) );
  INV_X1 U11296 ( .A(n12713), .ZN(n9935) );
  NAND2_X1 U11297 ( .A1(n12742), .A2(n12743), .ZN(n9770) );
  NAND2_X1 U11298 ( .A1(n9654), .A2(n9618), .ZN(n9772) );
  AND4_X1 U11299 ( .A1(n12762), .A2(n12749), .A3(n12763), .A4(n12750), .ZN(
        n9654) );
  NOR2_X2 U11300 ( .A1(n13555), .A2(n13665), .ZN(n15435) );
  NAND2_X1 U11301 ( .A1(n9620), .A2(n9816), .ZN(n14495) );
  NAND2_X1 U11302 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  NAND2_X1 U11303 ( .A1(n10849), .A2(n10263), .ZN(n10976) );
  AND2_X1 U11304 ( .A1(n14496), .A2(n9774), .ZN(n14448) );
  AND2_X4 U11305 ( .A1(n15741), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14496) );
  OAI21_X2 U11306 ( .B1(n13162), .B2(n10112), .A(n10109), .ZN(n13910) );
  NAND2_X2 U11307 ( .A1(n10801), .A2(n12939), .ZN(n10832) );
  NOR4_X2 U11308 ( .A1(n16932), .A2(n17015), .A3(n17017), .A4(n16855), .ZN(
        n16896) );
  NOR2_X2 U11309 ( .A1(n17226), .A2(n17266), .ZN(n17241) );
  NOR2_X2 U11310 ( .A1(n10150), .A2(n12722), .ZN(n19010) );
  NOR2_X1 U11311 ( .A1(n12736), .A2(n12735), .ZN(n12737) );
  NAND2_X1 U11312 ( .A1(n15825), .A2(n13404), .ZN(n14896) );
  NAND2_X1 U11313 ( .A1(n10266), .A2(n10265), .ZN(n10281) );
  AND3_X1 U11314 ( .A1(n10266), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10160), 
        .ZN(n10697) );
  INV_X2 U11315 ( .A(n18903), .ZN(n10266) );
  OAI21_X2 U11316 ( .B1(n14457), .B2(n14456), .A(n14671), .ZN(n14460) );
  NAND2_X2 U11317 ( .A1(n14468), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14671) );
  XNOR2_X2 U11318 ( .A(n14455), .B(n14456), .ZN(n14468) );
  NAND2_X2 U11319 ( .A1(n14454), .A2(n14453), .ZN(n14455) );
  NAND2_X1 U11320 ( .A1(n9594), .A2(n18884), .ZN(n12815) );
  AND3_X1 U11321 ( .A1(n18892), .A2(n18884), .A3(n18888), .ZN(n10297) );
  BUF_X4 U11322 ( .A(n10239), .Z(n10641) );
  NOR2_X1 U11323 ( .A1(n18472), .A2(n16152), .ZN(n17477) );
  NAND2_X1 U11324 ( .A1(n14916), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U11325 ( .A1(n14916), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U11326 ( .A1(n14916), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12125) );
  AND3_X2 U11327 ( .A1(n10274), .A2(n12779), .A3(n10297), .ZN(n10314) );
  NOR2_X4 U11328 ( .A1(n19692), .A2(n11937), .ZN(n15642) );
  OR2_X2 U11329 ( .A1(n19690), .A2(n19689), .ZN(n19692) );
  NOR2_X2 U11330 ( .A1(n10269), .A2(n10268), .ZN(n12021) );
  AOI21_X2 U11331 ( .B1(n14690), .B2(n14705), .A(n9616), .ZN(n14693) );
  OR2_X1 U11332 ( .A1(n12713), .A2(n18830), .ZN(n12720) );
  NOR2_X2 U11333 ( .A1(n17421), .A2(n17422), .ZN(n17391) );
  AND2_X1 U11334 ( .A1(n14914), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10392) );
  INV_X2 U11335 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10776) );
  NOR3_X4 U11336 ( .A1(n16550), .A2(n16549), .A3(n16605), .ZN(n16600) );
  INV_X4 U11337 ( .A(n16612), .ZN(n16778) );
  XOR2_X1 U11338 ( .A(n16174), .B(n15998), .Z(n16496) );
  NAND2_X1 U11339 ( .A1(n16901), .A2(n16856), .ZN(n9610) );
  NAND3_X2 U11340 ( .A1(n14955), .A2(n14954), .A3(n14953), .ZN(n16901) );
  NAND2_X1 U11341 ( .A1(n9820), .A2(n9828), .ZN(n13198) );
  OR2_X1 U11342 ( .A1(n9991), .A2(n9990), .ZN(n9820) );
  NOR2_X1 U11343 ( .A1(n9662), .A2(n9823), .ZN(n9822) );
  INV_X1 U11344 ( .A(n14454), .ZN(n9847) );
  NOR2_X1 U11345 ( .A1(n14452), .A2(n9799), .ZN(n9798) );
  NOR2_X1 U11346 ( .A1(n14458), .A2(n9844), .ZN(n9799) );
  NOR2_X1 U11347 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9844) );
  INV_X1 U11348 ( .A(n13420), .ZN(n13386) );
  INV_X1 U11349 ( .A(n11257), .ZN(n9831) );
  INV_X1 U11350 ( .A(n11256), .ZN(n9832) );
  OR2_X1 U11351 ( .A1(n13274), .A2(n13273), .ZN(n13278) );
  INV_X1 U11352 ( .A(n10904), .ZN(n9791) );
  AOI22_X1 U11353 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n17818), .B2(n18436), .ZN(
        n14983) );
  NOR2_X1 U11354 ( .A1(n10049), .A2(n9903), .ZN(n9902) );
  INV_X1 U11355 ( .A(n13582), .ZN(n9903) );
  NAND2_X1 U11356 ( .A1(n13557), .A2(n10050), .ZN(n10049) );
  NOR2_X1 U11357 ( .A1(n10051), .A2(n13664), .ZN(n10050) );
  INV_X1 U11358 ( .A(n11836), .ZN(n11809) );
  NOR2_X1 U11359 ( .A1(n12456), .A2(n20401), .ZN(n11836) );
  CLKBUF_X1 U11360 ( .A(n11313), .Z(n12878) );
  INV_X1 U11361 ( .A(n11313), .ZN(n11812) );
  NAND2_X1 U11362 ( .A1(n9878), .A2(n13999), .ZN(n9877) );
  NAND2_X1 U11363 ( .A1(n13910), .A2(n9624), .ZN(n9824) );
  NOR2_X1 U11364 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10116) );
  OR2_X1 U11365 ( .A1(n11206), .A2(n11205), .ZN(n13139) );
  INV_X1 U11366 ( .A(n13139), .ZN(n11240) );
  NAND2_X1 U11367 ( .A1(n10087), .A2(n14284), .ZN(n10086) );
  OR2_X1 U11368 ( .A1(n10598), .A2(n10623), .ZN(n10085) );
  NOR2_X1 U11369 ( .A1(n14433), .A2(n9797), .ZN(n9796) );
  INV_X1 U11370 ( .A(n14441), .ZN(n9797) );
  AND2_X1 U11371 ( .A1(n14458), .A2(n14659), .ZN(n9801) );
  NAND2_X1 U11372 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  NAND2_X1 U11373 ( .A1(n14456), .A2(n14674), .ZN(n9846) );
  OR2_X1 U11374 ( .A1(n13380), .A2(n14690), .ZN(n13381) );
  NAND2_X1 U11375 ( .A1(n13289), .A2(n10140), .ZN(n10139) );
  NOR2_X1 U11376 ( .A1(n15805), .A2(n14591), .ZN(n10140) );
  AND2_X1 U11377 ( .A1(n10298), .A2(n19571), .ZN(n10849) );
  NAND2_X1 U11378 ( .A1(n18830), .A2(n10370), .ZN(n10377) );
  NOR2_X1 U11379 ( .A1(n10389), .A2(n10378), .ZN(n10381) );
  NOR2_X1 U11380 ( .A1(n14945), .A2(n18285), .ZN(n15274) );
  NOR2_X1 U11381 ( .A1(n18283), .A2(n14944), .ZN(n15275) );
  NOR2_X1 U11382 ( .A1(n14946), .A2(n18283), .ZN(n14956) );
  AND3_X1 U11383 ( .A1(n16857), .A2(n17853), .A3(n18279), .ZN(n15153) );
  NOR2_X1 U11384 ( .A1(n12454), .A2(n12442), .ZN(n13450) );
  AND2_X1 U11385 ( .A1(n13450), .A2(n13456), .ZN(n12381) );
  AND4_X1 U11386 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n11117) );
  NOR2_X1 U11387 ( .A1(n13456), .A2(n19610), .ZN(n12466) );
  NOR3_X2 U11388 ( .A1(n13530), .A2(n13498), .A3(n10053), .ZN(n11842) );
  OR2_X1 U11389 ( .A1(n9615), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9834) );
  INV_X1 U11390 ( .A(n13200), .ZN(n9833) );
  OR2_X1 U11391 ( .A1(n9615), .A2(n14089), .ZN(n13901) );
  NAND2_X1 U11392 ( .A1(n13162), .A2(n13161), .ZN(n10113) );
  AND2_X1 U11393 ( .A1(n13368), .A2(n9649), .ZN(n13391) );
  AND2_X1 U11394 ( .A1(n10462), .A2(n12864), .ZN(n10089) );
  AND2_X1 U11395 ( .A1(n12986), .A2(n12985), .ZN(n10462) );
  NAND2_X1 U11396 ( .A1(n10416), .A2(n9908), .ZN(n9907) );
  INV_X1 U11397 ( .A(n12851), .ZN(n9908) );
  XNOR2_X1 U11398 ( .A(n10597), .B(n10622), .ZN(n14292) );
  AND2_X1 U11399 ( .A1(n9916), .A2(n9699), .ZN(n9915) );
  INV_X1 U11400 ( .A(n10092), .ZN(n10090) );
  INV_X1 U11401 ( .A(n12670), .ZN(n10062) );
  AND2_X1 U11402 ( .A1(n14137), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14135) );
  AND2_X1 U11403 ( .A1(n15967), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n10370) );
  NOR2_X1 U11404 ( .A1(n14484), .A2(n10145), .ZN(n10144) );
  INV_X1 U11405 ( .A(n10147), .ZN(n10145) );
  INV_X1 U11406 ( .A(n15767), .ZN(n10132) );
  NAND2_X1 U11407 ( .A1(n9786), .A2(n9785), .ZN(n14506) );
  AND2_X1 U11408 ( .A1(n14564), .A2(n14574), .ZN(n9785) );
  OAI21_X1 U11409 ( .B1(n10126), .B2(n10131), .A(n9787), .ZN(n9786) );
  NAND2_X1 U11410 ( .A1(n14878), .A2(n14875), .ZN(n13415) );
  AND2_X1 U11411 ( .A1(n12799), .A2(n12798), .ZN(n12834) );
  NAND2_X1 U11412 ( .A1(n12348), .A2(n12349), .ZN(n12350) );
  INV_X1 U11413 ( .A(n15536), .ZN(n19810) );
  NOR2_X2 U11414 ( .A1(n15373), .A2(n19610), .ZN(n19795) );
  OR2_X1 U11415 ( .A1(n14639), .A2(n18656), .ZN(n9987) );
  INV_X1 U11416 ( .A(n17804), .ZN(n17793) );
  NAND2_X1 U11417 ( .A1(n10281), .A2(n12778), .ZN(n10816) );
  AND2_X1 U11418 ( .A1(n11375), .A2(n11374), .ZN(n11382) );
  INV_X1 U11419 ( .A(n9690), .ZN(n9968) );
  AND2_X1 U11420 ( .A1(n9979), .A2(n9978), .ZN(n9977) );
  NAND2_X1 U11421 ( .A1(n10281), .A2(n18888), .ZN(n10287) );
  INV_X1 U11422 ( .A(n17163), .ZN(n10032) );
  INV_X1 U11423 ( .A(n10029), .ZN(n10023) );
  NOR2_X1 U11424 ( .A1(n15291), .A2(n16977), .ZN(n15294) );
  NOR2_X1 U11425 ( .A1(n16984), .A2(n15271), .ZN(n15270) );
  NAND2_X1 U11426 ( .A1(n15306), .A2(n9919), .ZN(n15271) );
  NAND2_X1 U11427 ( .A1(n17487), .A2(n9919), .ZN(n15305) );
  NOR2_X1 U11428 ( .A1(n18299), .A2(n14944), .ZN(n15256) );
  NAND2_X1 U11429 ( .A1(n11654), .A2(n10052), .ZN(n10051) );
  INV_X1 U11430 ( .A(n13669), .ZN(n10052) );
  INV_X1 U11431 ( .A(n13619), .ZN(n10044) );
  NAND2_X1 U11432 ( .A1(n10047), .A2(n11504), .ZN(n10046) );
  INV_X1 U11433 ( .A(n13762), .ZN(n10047) );
  OR2_X1 U11434 ( .A1(n13180), .A2(n13632), .ZN(n11457) );
  OR2_X1 U11435 ( .A1(n13180), .A2(n13179), .ZN(n13633) );
  INV_X1 U11436 ( .A(n13063), .ZN(n10043) );
  AND2_X1 U11437 ( .A1(n10043), .A2(n13089), .ZN(n10042) );
  XNOR2_X1 U11438 ( .A(n13137), .B(n11386), .ZN(n13123) );
  INV_X1 U11439 ( .A(n13006), .ZN(n11397) );
  AND2_X1 U11440 ( .A1(n11258), .A2(n13133), .ZN(n10118) );
  INV_X1 U11441 ( .A(n13999), .ZN(n9879) );
  NAND2_X1 U11442 ( .A1(n10114), .A2(n9615), .ZN(n9825) );
  NAND2_X1 U11443 ( .A1(n9827), .A2(n9826), .ZN(n9821) );
  OR2_X1 U11444 ( .A1(n10114), .A2(n9615), .ZN(n9826) );
  NAND2_X1 U11445 ( .A1(n9868), .A2(n13681), .ZN(n9867) );
  INV_X1 U11446 ( .A(n11973), .ZN(n9868) );
  NAND2_X1 U11447 ( .A1(n13164), .A2(n9658), .ZN(n10112) );
  INV_X1 U11448 ( .A(n10112), .ZN(n10111) );
  AND2_X1 U11449 ( .A1(n13122), .A2(n15556), .ZN(n9872) );
  INV_X1 U11450 ( .A(n13115), .ZN(n9873) );
  NAND2_X1 U11451 ( .A1(n10104), .A2(n13105), .ZN(n10103) );
  NAND2_X1 U11452 ( .A1(n19803), .A2(n12688), .ZN(n13096) );
  INV_X1 U11453 ( .A(n20489), .ZN(n13140) );
  OR2_X1 U11454 ( .A1(n13469), .A2(n13471), .ZN(n12012) );
  INV_X1 U11455 ( .A(n11843), .ZN(n10038) );
  AND2_X1 U11456 ( .A1(n11242), .A2(n11241), .ZN(n11251) );
  NAND2_X1 U11457 ( .A1(n11225), .A2(n11224), .ZN(n11253) );
  NOR2_X1 U11458 ( .A1(n11256), .A2(n11257), .ZN(n9964) );
  NOR2_X1 U11459 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n19854), .ZN(n19858) );
  OAI22_X1 U11460 ( .A1(n10790), .A2(n10778), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15934), .ZN(n10806) );
  AND2_X1 U11461 ( .A1(n9640), .A2(n20558), .ZN(n9973) );
  NAND2_X1 U11462 ( .A1(n13368), .A2(n13337), .ZN(n13327) );
  NAND2_X1 U11463 ( .A1(n13303), .A2(n9969), .ZN(n13314) );
  NOR2_X1 U11464 ( .A1(n13280), .A2(n13279), .ZN(n13287) );
  NAND2_X1 U11465 ( .A1(n14274), .A2(n10152), .ZN(n10670) );
  AND2_X1 U11466 ( .A1(n9685), .A2(n14335), .ZN(n9916) );
  INV_X1 U11467 ( .A(n13020), .ZN(n10059) );
  NOR2_X1 U11468 ( .A1(n10932), .A2(n10931), .ZN(n13238) );
  INV_X1 U11469 ( .A(n10697), .ZN(n10389) );
  NAND2_X1 U11470 ( .A1(n10252), .A2(n15934), .ZN(n10260) );
  INV_X1 U11471 ( .A(n12988), .ZN(n9936) );
  AND2_X1 U11472 ( .A1(n10011), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10009) );
  NOR2_X1 U11473 ( .A1(n15822), .A2(n10008), .ZN(n10011) );
  NOR2_X1 U11474 ( .A1(n15666), .A2(n13420), .ZN(n13379) );
  NAND2_X1 U11475 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  INV_X1 U11476 ( .A(n14281), .ZN(n9940) );
  NOR2_X1 U11477 ( .A1(n14293), .A2(n9943), .ZN(n9941) );
  OR3_X1 U11478 ( .A1(n13378), .A2(n13420), .A3(n14697), .ZN(n14475) );
  INV_X1 U11479 ( .A(n14732), .ZN(n9843) );
  AOI21_X1 U11480 ( .B1(n18547), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14539) );
  AND2_X1 U11481 ( .A1(n9632), .A2(n15846), .ZN(n10058) );
  NOR2_X1 U11482 ( .A1(n10131), .A2(n10129), .ZN(n10128) );
  INV_X1 U11483 ( .A(n14574), .ZN(n10129) );
  AND2_X1 U11484 ( .A1(n13405), .A2(n12767), .ZN(n9771) );
  NAND4_X1 U11485 ( .A1(n9790), .A2(n10903), .A3(n10905), .A4(n10906), .ZN(
        n12232) );
  NOR2_X1 U11486 ( .A1(n10902), .A2(n10901), .ZN(n10914) );
  NAND2_X1 U11487 ( .A1(n10348), .A2(n10318), .ZN(n10327) );
  INV_X1 U11488 ( .A(n12803), .ZN(n14917) );
  NOR2_X1 U11489 ( .A1(n18450), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n15155) );
  NOR2_X1 U11491 ( .A1(n14943), .A2(n18283), .ZN(n15095) );
  NAND2_X1 U11492 ( .A1(n15250), .A2(n15244), .ZN(n9734) );
  INV_X1 U11493 ( .A(n15247), .ZN(n9735) );
  INV_X1 U11494 ( .A(n15246), .ZN(n9739) );
  NAND2_X1 U11495 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n9738) );
  XNOR2_X1 U11496 ( .A(n9919), .B(n15306), .ZN(n15285) );
  NOR2_X1 U11497 ( .A1(n17409), .A2(n15298), .ZN(n15337) );
  INV_X1 U11498 ( .A(n10021), .ZN(n15296) );
  AND2_X1 U11499 ( .A1(n15328), .A2(n15326), .ZN(n9746) );
  NOR2_X1 U11500 ( .A1(n15328), .A2(n17737), .ZN(n9752) );
  NOR2_X1 U11501 ( .A1(n15320), .A2(n17431), .ZN(n15322) );
  XNOR2_X1 U11502 ( .A(n15294), .B(n9927), .ZN(n15292) );
  NAND2_X1 U11503 ( .A1(n15270), .A2(n15300), .ZN(n15291) );
  NOR2_X1 U11504 ( .A1(n17453), .A2(n15314), .ZN(n15316) );
  XNOR2_X1 U11505 ( .A(n15306), .B(n15305), .ZN(n15307) );
  AOI21_X1 U11506 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n15181) );
  NAND2_X1 U11507 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n9766) );
  NAND2_X1 U11508 ( .A1(n15154), .A2(n9600), .ZN(n15167) );
  AND2_X1 U11509 ( .A1(n11610), .A2(n11609), .ZN(n13582) );
  AND2_X1 U11510 ( .A1(n13678), .A2(n13677), .ZN(n13680) );
  AND2_X1 U11511 ( .A1(n15384), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U11512 ( .A1(n19871), .A2(n12443), .ZN(n20489) );
  OR2_X1 U11513 ( .A1(n13530), .A2(n10053), .ZN(n13508) );
  AOI21_X1 U11514 ( .B1(n11749), .B2(n11748), .A(n11747), .ZN(n13531) );
  AND2_X1 U11515 ( .A1(n13824), .A2(n12878), .ZN(n11747) );
  OR2_X1 U11516 ( .A1(n15427), .A2(n11812), .ZN(n11684) );
  XNOR2_X1 U11517 ( .A(n9615), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13881) );
  INV_X1 U11518 ( .A(n13546), .ZN(n9863) );
  NAND2_X1 U11519 ( .A1(n13881), .A2(n9994), .ZN(n9993) );
  INV_X1 U11520 ( .A(n13936), .ZN(n9994) );
  AND2_X1 U11521 ( .A1(n9992), .A2(n9615), .ZN(n9991) );
  OR2_X1 U11522 ( .A1(n15515), .A2(n9993), .ZN(n9992) );
  NAND2_X1 U11523 ( .A1(n9718), .A2(n9963), .ZN(n9962) );
  NOR2_X1 U11524 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9963) );
  OR2_X1 U11525 ( .A1(n12450), .A2(n12448), .ZN(n13933) );
  INV_X1 U11526 ( .A(n13912), .ZN(n9983) );
  OR2_X1 U11527 ( .A1(n12450), .A2(n12449), .ZN(n19812) );
  NAND2_X1 U11528 ( .A1(n14128), .A2(n20401), .ZN(n12407) );
  NAND2_X1 U11529 ( .A1(n13132), .A2(n15544), .ZN(n13162) );
  AND2_X1 U11530 ( .A1(n19932), .A2(n19931), .ZN(n20162) );
  OR2_X1 U11531 ( .A1(n19932), .A2(n19931), .ZN(n20141) );
  OR2_X1 U11532 ( .A1(n19932), .A2(n19853), .ZN(n20225) );
  AND2_X1 U11533 ( .A1(n11906), .A2(n11905), .ZN(n13456) );
  NAND2_X1 U11534 ( .A1(n13212), .A2(n13213), .ZN(n13376) );
  NAND2_X1 U11535 ( .A1(n13373), .A2(n13374), .ZN(n13382) );
  INV_X1 U11536 ( .A(n13376), .ZN(n13373) );
  AND2_X1 U11537 ( .A1(n12790), .A2(n12798), .ZN(n12928) );
  AND2_X1 U11538 ( .A1(n9716), .A2(n14202), .ZN(n10069) );
  INV_X1 U11539 ( .A(n10999), .ZN(n10070) );
  NOR2_X1 U11540 ( .A1(n10078), .A2(n10082), .ZN(n10077) );
  INV_X1 U11541 ( .A(n14251), .ZN(n10078) );
  INV_X1 U11542 ( .A(n10080), .ZN(n10079) );
  OAI22_X1 U11543 ( .A1(n14251), .A2(n10081), .B1(n10744), .B2(n10082), .ZN(
        n10080) );
  NAND2_X1 U11544 ( .A1(n10744), .A2(n10082), .ZN(n10081) );
  NOR2_X1 U11545 ( .A1(n14300), .A2(n9611), .ZN(n10598) );
  NAND2_X1 U11546 ( .A1(n9914), .A2(n9913), .ZN(n10597) );
  NOR2_X1 U11547 ( .A1(n10918), .A2(n10064), .ZN(n10063) );
  INV_X1 U11548 ( .A(n12658), .ZN(n10064) );
  NAND2_X1 U11549 ( .A1(n14310), .A2(n14309), .ZN(n14308) );
  NOR2_X1 U11550 ( .A1(n18625), .A2(n12958), .ZN(n12961) );
  NAND2_X1 U11551 ( .A1(n14268), .A2(n14209), .ZN(n14211) );
  XNOR2_X1 U11552 ( .A(n13379), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10142) );
  NAND2_X1 U11553 ( .A1(n10149), .A2(n14709), .ZN(n10147) );
  NAND2_X1 U11554 ( .A1(n14493), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10148) );
  AOI21_X1 U11555 ( .B1(n9841), .B2(n9613), .A(n9708), .ZN(n9840) );
  NOR2_X1 U11556 ( .A1(n14514), .A2(n9805), .ZN(n10124) );
  NAND2_X1 U11557 ( .A1(n10125), .A2(n10133), .ZN(n9805) );
  INV_X1 U11558 ( .A(n14516), .ZN(n10133) );
  AND2_X1 U11559 ( .A1(n9655), .A2(n10128), .ZN(n10125) );
  NAND2_X1 U11560 ( .A1(n10127), .A2(n10128), .ZN(n14579) );
  INV_X1 U11561 ( .A(n14827), .ZN(n9848) );
  INV_X1 U11562 ( .A(n14824), .ZN(n9849) );
  OR2_X1 U11563 ( .A1(n18603), .A2(n13305), .ZN(n14825) );
  NOR2_X1 U11564 ( .A1(n14844), .A2(n10138), .ZN(n10137) );
  INV_X1 U11565 ( .A(n10157), .ZN(n10138) );
  NAND3_X1 U11566 ( .A1(n9888), .A2(n13414), .A3(n9886), .ZN(n14599) );
  AND3_X1 U11567 ( .A1(n10864), .A2(n10863), .A3(n10862), .ZN(n12670) );
  NAND2_X1 U11568 ( .A1(n10060), .A2(n10063), .ZN(n12668) );
  OAI21_X1 U11569 ( .B1(n13035), .B2(n12233), .A(n10359), .ZN(n10360) );
  AOI21_X1 U11570 ( .B1(n12719), .B2(n10370), .A(n10352), .ZN(n12348) );
  INV_X1 U11571 ( .A(n12345), .ZN(n10379) );
  INV_X1 U11572 ( .A(n19550), .ZN(n19355) );
  AND2_X1 U11573 ( .A1(n19160), .A2(n19127), .ZN(n19098) );
  NAND2_X1 U11574 ( .A1(n19555), .A2(n19565), .ZN(n19235) );
  OR2_X1 U11575 ( .A1(n19555), .A2(n19563), .ZN(n19352) );
  OR2_X1 U11576 ( .A1(n19160), .A2(n19127), .ZN(n19353) );
  NAND2_X1 U11577 ( .A1(n10202), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10209) );
  INV_X1 U11578 ( .A(n19405), .ZN(n19162) );
  INV_X1 U11579 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n20564) );
  OAI221_X1 U11580 ( .B1(n15412), .B2(n15411), .C1(n15412), .C2(n15410), .A(
        n18470), .ZN(n15414) );
  NOR2_X1 U11581 ( .A1(n17466), .A2(n17467), .ZN(n17465) );
  INV_X1 U11582 ( .A(n17834), .ZN(n18472) );
  NAND2_X1 U11583 ( .A1(n9744), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16037) );
  INV_X1 U11584 ( .A(n9926), .ZN(n9744) );
  AND2_X1 U11585 ( .A1(n9926), .A2(n9925), .ZN(n17131) );
  NAND2_X1 U11586 ( .A1(n17272), .A2(n17359), .ZN(n17205) );
  NOR2_X1 U11587 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17388), .ZN(
        n17261) );
  NAND2_X1 U11588 ( .A1(n17273), .A2(n17607), .ZN(n17272) );
  NAND2_X1 U11589 ( .A1(n9759), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9758) );
  INV_X1 U11590 ( .A(n9760), .ZN(n9759) );
  OR3_X1 U11591 ( .A1(n17691), .A2(n17329), .A3(n9760), .ZN(n17305) );
  INV_X1 U11592 ( .A(n17359), .ZN(n17388) );
  NAND2_X1 U11593 ( .A1(n9756), .A2(n9754), .ZN(n17403) );
  AND2_X1 U11594 ( .A1(n9612), .A2(n15326), .ZN(n9754) );
  XNOR2_X1 U11595 ( .A(n15292), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17415) );
  NOR2_X1 U11596 ( .A1(n17415), .A2(n10026), .ZN(n10025) );
  INV_X1 U11597 ( .A(n10028), .ZN(n10026) );
  NAND2_X1 U11598 ( .A1(n17429), .A2(n10030), .ZN(n10028) );
  AND2_X1 U11599 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15289), .ZN(
        n15290) );
  NOR2_X1 U11600 ( .A1(n17445), .A2(n17444), .ZN(n17443) );
  INV_X1 U11601 ( .A(n17465), .ZN(n10018) );
  XNOR2_X1 U11602 ( .A(n13474), .B(n13473), .ZN(n13929) );
  INV_X1 U11603 ( .A(n13764), .ZN(n13774) );
  XNOR2_X1 U11604 ( .A(n13206), .B(n13205), .ZN(n13700) );
  AND2_X1 U11605 ( .A1(n13917), .A2(n12501), .ZN(n15536) );
  NAND2_X1 U11606 ( .A1(n9956), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9954) );
  INV_X1 U11607 ( .A(n13929), .ZN(n9855) );
  OR2_X1 U11608 ( .A1(n12407), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15601) );
  INV_X1 U11609 ( .A(n19834), .ZN(n19825) );
  NOR2_X1 U11610 ( .A1(n14174), .A2(n14437), .ZN(n14173) );
  NAND2_X1 U11611 ( .A1(n18653), .A2(n9996), .ZN(n9995) );
  INV_X1 U11612 ( .A(n14444), .ZN(n9996) );
  INV_X1 U11613 ( .A(n18669), .ZN(n18653) );
  OAI21_X2 U11614 ( .B1(n14263), .B2(n9911), .A(n9909), .ZN(n14252) );
  NAND2_X1 U11615 ( .A1(n9912), .A2(n9717), .ZN(n9911) );
  NAND2_X1 U11616 ( .A1(n9910), .A2(n9717), .ZN(n9909) );
  INV_X1 U11617 ( .A(n14262), .ZN(n9912) );
  INV_X1 U11618 ( .A(n9907), .ZN(n9905) );
  AND2_X1 U11619 ( .A1(n10089), .A2(n10159), .ZN(n10088) );
  XNOR2_X1 U11620 ( .A(n12923), .B(n20511), .ZN(n13402) );
  NAND2_X1 U11621 ( .A1(n14135), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12923) );
  INV_X1 U11622 ( .A(n15833), .ZN(n18810) );
  INV_X1 U11623 ( .A(n15824), .ZN(n18817) );
  AND2_X1 U11624 ( .A1(n15833), .A2(n19562), .ZN(n18819) );
  INV_X1 U11625 ( .A(n15816), .ZN(n18814) );
  XNOR2_X1 U11626 ( .A(n9775), .B(n14622), .ZN(n14628) );
  NAND2_X1 U11627 ( .A1(n14496), .A2(n9644), .ZN(n9775) );
  NAND2_X1 U11628 ( .A1(n9794), .A2(n9792), .ZN(n13394) );
  OR2_X1 U11629 ( .A1(n14181), .A2(n12131), .ZN(n9938) );
  XNOR2_X1 U11630 ( .A(n14435), .B(n14434), .ZN(n14643) );
  NAND2_X1 U11631 ( .A1(n14442), .A2(n14441), .ZN(n14432) );
  OR2_X1 U11632 ( .A1(n14791), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9891) );
  NAND2_X1 U11633 ( .A1(n9893), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9892) );
  NAND2_X1 U11634 ( .A1(n18854), .A2(n14790), .ZN(n9893) );
  AND2_X1 U11635 ( .A1(n12834), .A2(n12821), .ZN(n18836) );
  INV_X1 U11636 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19578) );
  INV_X1 U11637 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19570) );
  INV_X1 U11638 ( .A(n19563), .ZN(n19565) );
  INV_X1 U11639 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19554) );
  NAND2_X1 U11640 ( .A1(n18921), .A2(n19571), .ZN(n19550) );
  NOR2_X2 U11641 ( .A1(n18419), .A2(n16529), .ZN(n16533) );
  AOI211_X1 U11642 ( .C1(n16619), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n14952), .B(n14951), .ZN(n14953) );
  INV_X1 U11643 ( .A(n16940), .ZN(n16995) );
  NOR2_X1 U11644 ( .A1(n18269), .A2(n15414), .ZN(n16993) );
  INV_X1 U11645 ( .A(n15414), .ZN(n16856) );
  NOR2_X2 U11646 ( .A1(n17491), .A2(n17646), .ZN(n17342) );
  NAND2_X1 U11647 ( .A1(n9930), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9929) );
  NAND2_X1 U11648 ( .A1(n15400), .A2(n16022), .ZN(n9930) );
  NAND2_X1 U11649 ( .A1(n10036), .A2(n15976), .ZN(n16005) );
  OR2_X1 U11650 ( .A1(n15398), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10036) );
  INV_X1 U11651 ( .A(n16037), .ZN(n17132) );
  NAND3_X1 U11652 ( .A1(n15197), .A2(n15196), .A3(n15195), .ZN(n17644) );
  INV_X1 U11653 ( .A(n17644), .ZN(n17646) );
  INV_X1 U11654 ( .A(n17727), .ZN(n17681) );
  OAI21_X2 U11655 ( .B1(n15185), .B2(n15184), .A(n18470), .ZN(n17804) );
  NOR2_X1 U11656 ( .A1(n17804), .A2(n18261), .ZN(n17811) );
  INV_X1 U11657 ( .A(n9825), .ZN(n9823) );
  NOR2_X1 U11658 ( .A1(n9959), .A2(n11154), .ZN(n9958) );
  OAI21_X1 U11659 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18436), .A(
        n14978), .ZN(n14979) );
  NAND2_X1 U11660 ( .A1(n10095), .A2(n11142), .ZN(n11148) );
  AOI21_X1 U11661 ( .B1(n10117), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10114) );
  OR2_X1 U11662 ( .A1(n11333), .A2(n11332), .ZN(n13108) );
  INV_X1 U11663 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10037) );
  INV_X1 U11664 ( .A(n9901), .ZN(n12377) );
  OAI21_X1 U11665 ( .B1(n12470), .B2(n12429), .A(n11155), .ZN(n9901) );
  NAND2_X1 U11666 ( .A1(n11095), .A2(n19875), .ZN(n11097) );
  OR2_X1 U11667 ( .A1(n11309), .A2(n11308), .ZN(n13107) );
  NAND2_X1 U11668 ( .A1(n10098), .A2(n11152), .ZN(n10097) );
  NAND2_X1 U11669 ( .A1(n11169), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10098) );
  OR3_X1 U11670 ( .A1(n11894), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n19848), .ZN(n11896) );
  NOR2_X1 U11671 ( .A1(n9970), .A2(n13311), .ZN(n9969) );
  NAND2_X1 U11672 ( .A1(n13255), .A2(n13254), .ZN(n13419) );
  INV_X1 U11673 ( .A(n13408), .ZN(n13255) );
  INV_X1 U11674 ( .A(n12815), .ZN(n10819) );
  OAI21_X1 U11675 ( .B1(n9603), .B2(n10310), .A(n10309), .ZN(n10311) );
  INV_X1 U11676 ( .A(n12806), .ZN(n10282) );
  INV_X1 U11677 ( .A(n10160), .ZN(n10298) );
  AOI22_X1 U11678 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U11679 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10206) );
  AND2_X1 U11680 ( .A1(n10797), .A2(n10775), .ZN(n10794) );
  OR2_X1 U11681 ( .A1(n10796), .A2(n10795), .ZN(n10797) );
  NAND2_X1 U11682 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18450), .ZN(
        n14945) );
  NAND2_X1 U11683 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14944) );
  NOR2_X1 U11684 ( .A1(n16981), .A2(n15315), .ZN(n15302) );
  AOI21_X1 U11685 ( .B1(n15138), .B2(n17853), .A(n15177), .ZN(n15135) );
  NOR2_X1 U11686 ( .A1(n15199), .A2(n16151), .ZN(n15159) );
  AND4_X1 U11687 ( .A1(n11160), .A2(n11159), .A3(n11158), .A4(n12438), .ZN(
        n11164) );
  XNOR2_X1 U11688 ( .A(n9981), .B(n11363), .ZN(n13106) );
  AND2_X1 U11689 ( .A1(n19992), .A2(n11343), .ZN(n9830) );
  NAND2_X1 U11690 ( .A1(n13509), .A2(n10054), .ZN(n10053) );
  INV_X1 U11691 ( .A(n13519), .ZN(n10054) );
  AND2_X1 U11692 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11376), .ZN(
        n11387) );
  NOR2_X1 U11693 ( .A1(n11357), .A2(n19670), .ZN(n11376) );
  NAND2_X1 U11694 ( .A1(n12681), .A2(n12680), .ZN(n12687) );
  NAND2_X1 U11695 ( .A1(n10039), .A2(n11443), .ZN(n11286) );
  NAND2_X1 U11696 ( .A1(n10040), .A2(n11288), .ZN(n10039) );
  AND2_X1 U11697 ( .A1(n11258), .A2(n11514), .ZN(n10040) );
  INV_X1 U11698 ( .A(n13510), .ZN(n9859) );
  INV_X1 U11699 ( .A(n13533), .ZN(n9862) );
  NAND2_X1 U11700 ( .A1(n9961), .A2(n13189), .ZN(n13890) );
  INV_X1 U11701 ( .A(n13902), .ZN(n9961) );
  OR2_X1 U11702 ( .A1(n9615), .A2(n13197), .ZN(n13911) );
  OR2_X1 U11703 ( .A1(n9615), .A2(n13196), .ZN(n13913) );
  NAND2_X1 U11704 ( .A1(n19883), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13134) );
  AND2_X1 U11705 ( .A1(n19992), .A2(n9701), .ZN(n9829) );
  INV_X1 U11706 ( .A(n11382), .ZN(n11383) );
  OAI211_X1 U11707 ( .C1(n12006), .C2(P1_EBX_REG_1__SCAN_IN), .A(n11913), .B(
        n9852), .ZN(n9851) );
  NAND2_X1 U11708 ( .A1(n12013), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n9852) );
  INV_X1 U11709 ( .A(n13702), .ZN(n11259) );
  OR2_X1 U11710 ( .A1(n11238), .A2(n11237), .ZN(n12506) );
  INV_X1 U11711 ( .A(n13134), .ZN(n11248) );
  OR2_X1 U11712 ( .A1(n11253), .A2(n11252), .ZN(n11254) );
  OR2_X1 U11713 ( .A1(n12441), .A2(n11850), .ZN(n12454) );
  INV_X1 U11714 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20163) );
  AOI21_X1 U11715 ( .B1(n20494), .B2(n15664), .A(n15388), .ZN(n19854) );
  AND2_X1 U11716 ( .A1(n11296), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11879) );
  NAND2_X1 U11717 ( .A1(n10271), .A2(n10298), .ZN(n10801) );
  INV_X1 U11718 ( .A(n13359), .ZN(n9975) );
  AND2_X1 U11719 ( .A1(n13211), .A2(n13328), .ZN(n9971) );
  NAND2_X1 U11720 ( .A1(n13326), .A2(n10265), .ZN(n9814) );
  AND2_X1 U11721 ( .A1(n13327), .A2(n13328), .ZN(n13326) );
  NAND2_X1 U11722 ( .A1(n13303), .A2(n9614), .ZN(n13336) );
  NAND2_X1 U11723 ( .A1(n13303), .A2(n9661), .ZN(n13337) );
  AND2_X1 U11724 ( .A1(n9977), .A2(n12026), .ZN(n9976) );
  NAND2_X1 U11725 ( .A1(n9660), .A2(n13368), .ZN(n13303) );
  AND2_X1 U11726 ( .A1(n13287), .A2(n9977), .ZN(n13300) );
  AND2_X1 U11727 ( .A1(n13285), .A2(n9980), .ZN(n9979) );
  INV_X1 U11728 ( .A(n12972), .ZN(n9980) );
  NAND2_X1 U11729 ( .A1(n9811), .A2(n9810), .ZN(n13280) );
  AND3_X1 U11730 ( .A1(n9807), .A2(n13245), .A3(n9806), .ZN(n9810) );
  INV_X1 U11731 ( .A(n13240), .ZN(n9806) );
  INV_X1 U11732 ( .A(n12773), .ZN(n9811) );
  NAND2_X1 U11733 ( .A1(n9967), .A2(n9966), .ZN(n12774) );
  NAND2_X1 U11734 ( .A1(n18899), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n9966) );
  OR2_X1 U11735 ( .A1(n12772), .A2(n18899), .ZN(n9967) );
  NAND2_X1 U11736 ( .A1(n12244), .A2(n12245), .ZN(n12773) );
  INV_X1 U11737 ( .A(n10762), .ZN(n10082) );
  NOR2_X1 U11738 ( .A1(n14269), .A2(n10671), .ZN(n10699) );
  NOR2_X1 U11739 ( .A1(n14389), .A2(n14378), .ZN(n10056) );
  NAND2_X1 U11740 ( .A1(n10517), .A2(n10093), .ZN(n10092) );
  INV_X1 U11741 ( .A(n14322), .ZN(n10093) );
  INV_X1 U11742 ( .A(n14343), .ZN(n9917) );
  NOR2_X1 U11743 ( .A1(n10944), .A2(n10943), .ZN(n13276) );
  OR2_X1 U11744 ( .A1(n10788), .A2(n10787), .ZN(n12765) );
  NAND2_X1 U11745 ( .A1(n12806), .A2(n9594), .ZN(n10279) );
  AND2_X1 U11746 ( .A1(n10298), .A2(n18884), .ZN(n12788) );
  NOR2_X1 U11747 ( .A1(n14487), .A2(n10014), .ZN(n10013) );
  AND2_X1 U11748 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  INV_X1 U11749 ( .A(n14318), .ZN(n9947) );
  NOR2_X1 U11750 ( .A1(n14543), .A2(n10003), .ZN(n10002) );
  INV_X1 U11751 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10003) );
  NOR2_X1 U11752 ( .A1(n18591), .A2(n10007), .ZN(n10006) );
  INV_X1 U11753 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10007) );
  INV_X1 U11754 ( .A(n12859), .ZN(n9937) );
  NOR2_X1 U11755 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  INV_X1 U11756 ( .A(n10144), .ZN(n10143) );
  AND2_X1 U11757 ( .A1(n9643), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10120) );
  NOR2_X1 U11758 ( .A1(n14620), .A2(n14709), .ZN(n10121) );
  INV_X1 U11759 ( .A(n14719), .ZN(n9838) );
  INV_X1 U11760 ( .A(n10130), .ZN(n9818) );
  NOR2_X1 U11761 ( .A1(n9839), .A2(n9679), .ZN(n9817) );
  INV_X1 U11762 ( .A(n9840), .ZN(n9839) );
  INV_X1 U11763 ( .A(n13398), .ZN(n12124) );
  INV_X1 U11764 ( .A(n14407), .ZN(n14741) );
  AND2_X1 U11765 ( .A1(n14228), .A2(n14415), .ZN(n10065) );
  AND2_X1 U11766 ( .A1(n14336), .A2(n14327), .ZN(n9948) );
  NOR2_X1 U11767 ( .A1(n14504), .A2(n9788), .ZN(n9787) );
  NAND2_X1 U11768 ( .A1(n14575), .A2(n15767), .ZN(n9788) );
  INV_X1 U11769 ( .A(n12025), .ZN(n12126) );
  NOR2_X1 U11770 ( .A1(n12978), .A2(n10068), .ZN(n10067) );
  INV_X1 U11771 ( .A(n15906), .ZN(n10068) );
  INV_X1 U11772 ( .A(n14590), .ZN(n13289) );
  OR2_X1 U11773 ( .A1(n13419), .A2(n13412), .ZN(n13424) );
  INV_X1 U11774 ( .A(n13411), .ZN(n9887) );
  AND2_X1 U11775 ( .A1(n13411), .A2(n14875), .ZN(n9889) );
  NAND2_X1 U11776 ( .A1(n13409), .A2(n13420), .ZN(n9835) );
  INV_X1 U11777 ( .A(n10976), .ZN(n10964) );
  OAI21_X1 U11778 ( .B1(n10286), .B2(n10285), .A(n10284), .ZN(n10288) );
  OR2_X2 U11779 ( .A1(n13035), .A2(n12706), .ZN(n12726) );
  NAND2_X1 U11780 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10227) );
  NAND2_X1 U11781 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10228) );
  NAND2_X1 U11782 ( .A1(n10225), .A2(n10224), .ZN(n10231) );
  AOI22_X1 U11783 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10217) );
  OR2_X1 U11784 ( .A1(n18277), .A2(n14944), .ZN(n9646) );
  NOR2_X1 U11785 ( .A1(n18283), .A2(n14945), .ZN(n15067) );
  NAND2_X1 U11786 ( .A1(n15256), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10015) );
  INV_X1 U11787 ( .A(n17143), .ZN(n9745) );
  NAND2_X1 U11788 ( .A1(n9741), .A2(n17359), .ZN(n15338) );
  AND2_X1 U11789 ( .A1(n9709), .A2(n17733), .ZN(n9742) );
  INV_X1 U11790 ( .A(n14944), .ZN(n9757) );
  INV_X1 U11791 ( .A(n18285), .ZN(n9731) );
  NAND2_X1 U11792 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n9760) );
  AND2_X1 U11793 ( .A1(n15294), .A2(n15299), .ZN(n15295) );
  AOI21_X1 U11794 ( .B1(n10025), .B2(n10023), .A(n15293), .ZN(n10022) );
  INV_X1 U11795 ( .A(n10025), .ZN(n10024) );
  AND2_X1 U11796 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15292), .ZN(
        n15293) );
  INV_X1 U11797 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20625) );
  INV_X1 U11798 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19670) );
  INV_X1 U11799 ( .A(n13465), .ZN(n13462) );
  OR2_X1 U11800 ( .A1(n20496), .A2(n12880), .ZN(n19646) );
  OR2_X1 U11801 ( .A1(n13663), .A2(n13559), .ZN(n13561) );
  NOR3_X1 U11802 ( .A1(n15472), .A2(n9676), .A3(n11973), .ZN(n13682) );
  AND3_X1 U11803 ( .A1(n11410), .A2(n11409), .A3(n11408), .ZN(n13063) );
  AOI21_X1 U11804 ( .B1(n12515), .B2(n11985), .A(n9851), .ZN(n12612) );
  AND2_X1 U11805 ( .A1(n11594), .A2(n11593), .ZN(n13677) );
  INV_X1 U11806 ( .A(n11443), .ZN(n13202) );
  NOR2_X1 U11807 ( .A1(n11789), .A2(n13796), .ZN(n11790) );
  OR2_X1 U11808 ( .A1(n11752), .A2(n13520), .ZN(n11789) );
  NAND2_X1 U11809 ( .A1(n13680), .A2(n9686), .ZN(n13530) );
  NAND2_X1 U11810 ( .A1(n11725), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11726) );
  OR2_X1 U11811 ( .A1(n11726), .A2(n13832), .ZN(n11750) );
  AND2_X1 U11812 ( .A1(n13680), .A2(n9633), .ZN(n13543) );
  AND2_X1 U11813 ( .A1(n13845), .A2(n11313), .ZN(n11703) );
  INV_X1 U11814 ( .A(n10050), .ZN(n10048) );
  INV_X1 U11815 ( .A(n11650), .ZN(n11649) );
  NOR2_X1 U11816 ( .A1(n11587), .A2(n13600), .ZN(n11588) );
  OR2_X1 U11817 ( .A1(n11555), .A2(n11554), .ZN(n11587) );
  NAND2_X1 U11818 ( .A1(n11536), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11555) );
  INV_X1 U11819 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11554) );
  NOR2_X1 U11820 ( .A1(n11522), .A2(n15466), .ZN(n11536) );
  NOR2_X1 U11821 ( .A1(n9693), .A2(n9898), .ZN(n9897) );
  INV_X1 U11822 ( .A(n11487), .ZN(n9898) );
  OR2_X1 U11823 ( .A1(n11505), .A2(n15476), .ZN(n11522) );
  NOR2_X1 U11824 ( .A1(n13638), .A2(n10046), .ZN(n13618) );
  INV_X1 U11825 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15476) );
  INV_X1 U11826 ( .A(n13638), .ZN(n10045) );
  NOR2_X1 U11827 ( .A1(n11471), .A2(n11472), .ZN(n11489) );
  INV_X1 U11828 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11472) );
  AND2_X1 U11829 ( .A1(n11440), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11441) );
  AND2_X1 U11830 ( .A1(n10042), .A2(n13150), .ZN(n10041) );
  NAND2_X1 U11831 ( .A1(n11411), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11435) );
  NOR2_X1 U11832 ( .A1(n13011), .A2(n9900), .ZN(n9899) );
  INV_X1 U11833 ( .A(n12844), .ZN(n9900) );
  NAND2_X1 U11834 ( .A1(n11397), .A2(n11396), .ZN(n13062) );
  NAND2_X1 U11835 ( .A1(n12845), .A2(n12844), .ZN(n13012) );
  NOR2_X1 U11836 ( .A1(n11315), .A2(n11314), .ZN(n11338) );
  INV_X1 U11837 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U11838 ( .A1(n11323), .A2(n11322), .ZN(n12616) );
  OR2_X1 U11839 ( .A1(n20107), .A2(n11438), .ZN(n11323) );
  NAND2_X1 U11840 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11315) );
  NAND2_X1 U11841 ( .A1(n11288), .A2(n10118), .ZN(n12686) );
  XNOR2_X1 U11842 ( .A(n11286), .B(n11284), .ZN(n12564) );
  OR2_X1 U11843 ( .A1(n13454), .A2(n13456), .ZN(n15373) );
  AND2_X1 U11844 ( .A1(n12498), .A2(n12499), .ZN(n12563) );
  NAND2_X1 U11845 ( .A1(n9881), .A2(n9880), .ZN(n9874) );
  NOR2_X1 U11846 ( .A1(n9615), .A2(n13966), .ZN(n9880) );
  NOR3_X1 U11847 ( .A1(n13561), .A2(n9856), .A3(n9858), .ZN(n13512) );
  NAND2_X1 U11848 ( .A1(n13523), .A2(n9857), .ZN(n9856) );
  OR2_X1 U11849 ( .A1(n9862), .A2(n9859), .ZN(n9858) );
  INV_X1 U11850 ( .A(n13547), .ZN(n9857) );
  NOR2_X1 U11851 ( .A1(n9861), .A2(n9860), .ZN(n13521) );
  NAND2_X1 U11852 ( .A1(n13848), .A2(n13999), .ZN(n9884) );
  INV_X1 U11853 ( .A(n13848), .ZN(n13827) );
  NOR2_X1 U11854 ( .A1(n13828), .A2(n14029), .ZN(n13839) );
  NOR2_X1 U11855 ( .A1(n13673), .A2(n13572), .ZN(n13661) );
  OR2_X1 U11856 ( .A1(n13671), .A2(n13670), .ZN(n13673) );
  NAND2_X1 U11857 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  INV_X1 U11858 ( .A(n9867), .ZN(n9866) );
  NOR2_X1 U11859 ( .A1(n9676), .A2(n13583), .ZN(n9865) );
  NOR2_X1 U11860 ( .A1(n13891), .A2(n13888), .ZN(n15515) );
  NOR2_X1 U11861 ( .A1(n15472), .A2(n11973), .ZN(n13621) );
  OR2_X1 U11862 ( .A1(n13692), .A2(n13693), .ZN(n15472) );
  NOR2_X1 U11863 ( .A1(n15488), .A2(n15487), .ZN(n15490) );
  NAND2_X1 U11864 ( .A1(n15490), .A2(n13645), .ZN(n13692) );
  AND2_X1 U11865 ( .A1(n13187), .A2(n13901), .ZN(n9819) );
  NAND2_X1 U11866 ( .A1(n9850), .A2(n9715), .ZN(n15488) );
  NAND2_X1 U11867 ( .A1(n10113), .A2(n10111), .ZN(n14093) );
  AOI21_X1 U11868 ( .B1(n10111), .B2(n10110), .A(n9667), .ZN(n10109) );
  INV_X1 U11869 ( .A(n13161), .ZN(n10110) );
  AOI21_X1 U11870 ( .B1(n13122), .B2(n9873), .A(n9665), .ZN(n9870) );
  AND2_X1 U11871 ( .A1(n12612), .A2(n12611), .ZN(n12619) );
  XNOR2_X1 U11872 ( .A(n9851), .B(n12433), .ZN(n12515) );
  INV_X1 U11873 ( .A(n13933), .ZN(n13170) );
  AND2_X1 U11874 ( .A1(n12424), .A2(n12423), .ZN(n12450) );
  NAND2_X1 U11875 ( .A1(n11223), .A2(n11222), .ZN(n11273) );
  NAND2_X1 U11876 ( .A1(n11295), .A2(n11294), .ZN(n19993) );
  NAND2_X1 U11877 ( .A1(n9964), .A2(n19992), .ZN(n11344) );
  INV_X1 U11878 ( .A(n9964), .ZN(n11288) );
  BUF_X1 U11879 ( .A(n11303), .Z(n11736) );
  NOR2_X1 U11880 ( .A1(n12389), .A2(n12388), .ZN(n15360) );
  INV_X1 U11881 ( .A(n20081), .ZN(n20076) );
  INV_X1 U11882 ( .A(n20111), .ZN(n20294) );
  INV_X1 U11883 ( .A(n20141), .ZN(n20257) );
  INV_X1 U11884 ( .A(n20162), .ZN(n20289) );
  OR2_X1 U11885 ( .A1(n20105), .A2(n12839), .ZN(n20290) );
  INV_X1 U11886 ( .A(n20290), .ZN(n20258) );
  INV_X1 U11887 ( .A(n20201), .ZN(n20075) );
  AOI21_X1 U11888 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20259), .A(n19999), 
        .ZN(n20344) );
  OR3_X1 U11889 ( .A1(n20232), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n19854), 
        .ZN(n19896) );
  NAND2_X1 U11890 ( .A1(n9789), .A2(n12156), .ZN(n12243) );
  NAND2_X1 U11891 ( .A1(n12232), .A2(n12200), .ZN(n9789) );
  NAND2_X1 U11892 ( .A1(n10808), .A2(n10807), .ZN(n12160) );
  OR2_X1 U11893 ( .A1(n10806), .A2(n10805), .ZN(n10808) );
  NAND2_X1 U11894 ( .A1(n10297), .A2(n10296), .ZN(n15941) );
  NOR2_X1 U11895 ( .A1(n14444), .A2(n14464), .ZN(n9998) );
  NAND2_X1 U11896 ( .A1(n14200), .A2(n14183), .ZN(n14185) );
  OR2_X1 U11897 ( .A1(n14219), .A2(n18653), .ZN(n10000) );
  NAND2_X1 U11898 ( .A1(n13391), .A2(n13372), .ZN(n15666) );
  NAND2_X1 U11899 ( .A1(n9803), .A2(n10263), .ZN(n13368) );
  INV_X1 U11900 ( .A(n12973), .ZN(n9803) );
  NAND2_X1 U11901 ( .A1(n13318), .A2(n13355), .ZN(n13360) );
  NAND2_X1 U11902 ( .A1(n13357), .A2(n13368), .ZN(n13318) );
  NAND2_X1 U11903 ( .A1(n13327), .A2(n9971), .ZN(n13323) );
  NOR2_X1 U11904 ( .A1(n9813), .A2(n9812), .ZN(n18547) );
  NAND2_X1 U11905 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  INV_X1 U11906 ( .A(n13321), .ZN(n9812) );
  OR2_X1 U11907 ( .A1(n13326), .A2(n13320), .ZN(n9815) );
  NOR2_X1 U11908 ( .A1(n14145), .A2(n14149), .ZN(n14152) );
  NAND2_X1 U11909 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14150), .ZN(
        n14149) );
  NAND2_X1 U11910 ( .A1(n13303), .A2(n12951), .ZN(n13312) );
  AND2_X1 U11911 ( .A1(n18899), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12972) );
  NAND2_X1 U11912 ( .A1(n13287), .A2(n9979), .ZN(n13294) );
  NAND2_X1 U11913 ( .A1(n9811), .A2(n9808), .ZN(n13248) );
  NOR2_X1 U11914 ( .A1(n12774), .A2(n9809), .ZN(n9808) );
  INV_X1 U11915 ( .A(n13245), .ZN(n9809) );
  AND2_X1 U11916 ( .A1(n9634), .A2(n12559), .ZN(n10094) );
  NAND2_X1 U11917 ( .A1(n10326), .A2(n10325), .ZN(n10353) );
  OR2_X1 U11918 ( .A1(n9602), .A2(n12203), .ZN(n10320) );
  NAND2_X1 U11919 ( .A1(n10056), .A2(n10055), .ZN(n14373) );
  INV_X1 U11920 ( .A(n14371), .ZN(n10055) );
  INV_X1 U11921 ( .A(n10056), .ZN(n14380) );
  XNOR2_X1 U11922 ( .A(n10652), .B(n10648), .ZN(n14276) );
  OR2_X1 U11923 ( .A1(n10556), .A2(n10555), .ZN(n14307) );
  AND2_X1 U11924 ( .A1(n14777), .A2(n14415), .ZN(n14417) );
  OR2_X1 U11925 ( .A1(n10505), .A2(n10504), .ZN(n14335) );
  NAND2_X1 U11926 ( .A1(n14809), .A2(n10058), .ZN(n15845) );
  NAND2_X1 U11927 ( .A1(n14809), .A2(n14810), .ZN(n14811) );
  NAND2_X1 U11928 ( .A1(n15907), .A2(n9681), .ZN(n15881) );
  INV_X1 U11929 ( .A(n18913), .ZN(n11000) );
  INV_X1 U11930 ( .A(n11011), .ZN(n18861) );
  OAI21_X1 U11931 ( .B1(n11010), .B2(n11009), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n11011) );
  AND2_X1 U11932 ( .A1(n14139), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14137) );
  AND2_X1 U11933 ( .A1(n14143), .A2(n10012), .ZN(n14139) );
  AND2_X1 U11934 ( .A1(n9638), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10012) );
  NAND2_X1 U11935 ( .A1(n14143), .A2(n9638), .ZN(n14158) );
  NAND2_X1 U11936 ( .A1(n14143), .A2(n10013), .ZN(n14156) );
  NAND2_X1 U11937 ( .A1(n14143), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14142) );
  NOR2_X1 U11938 ( .A1(n14153), .A2(n20563), .ZN(n14143) );
  NAND2_X1 U11939 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n14154), .ZN(
        n14153) );
  AND2_X1 U11940 ( .A1(n14152), .A2(n10001), .ZN(n14154) );
  AND2_X1 U11941 ( .A1(n9639), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10001) );
  NAND2_X1 U11942 ( .A1(n14152), .A2(n9639), .ZN(n14144) );
  AND2_X1 U11943 ( .A1(n14345), .A2(n9944), .ZN(n14310) );
  AND2_X1 U11944 ( .A1(n9946), .A2(n9945), .ZN(n9944) );
  INV_X1 U11945 ( .A(n14226), .ZN(n9945) );
  NAND2_X1 U11946 ( .A1(n14345), .A2(n9946), .ZN(n14320) );
  NAND2_X1 U11947 ( .A1(n14152), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14151) );
  OR2_X1 U11948 ( .A1(n13085), .A2(n13084), .ZN(n14346) );
  AND2_X1 U11949 ( .A1(n12962), .A2(n10005), .ZN(n14150) );
  AND2_X1 U11950 ( .A1(n9629), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10005) );
  NAND2_X1 U11951 ( .A1(n12962), .A2(n9629), .ZN(n14146) );
  INV_X1 U11952 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18591) );
  NAND2_X1 U11953 ( .A1(n12962), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13016) );
  NAND2_X1 U11954 ( .A1(n12866), .A2(n9680), .ZN(n12989) );
  NOR2_X1 U11955 ( .A1(n18602), .A2(n12960), .ZN(n12962) );
  NAND2_X1 U11956 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n12961), .ZN(
        n12960) );
  NAND2_X1 U11957 ( .A1(n10010), .A2(n9689), .ZN(n12958) );
  AND2_X1 U11958 ( .A1(n10010), .A2(n10009), .ZN(n12959) );
  AND2_X1 U11959 ( .A1(n12534), .A2(n12533), .ZN(n12556) );
  AND2_X1 U11960 ( .A1(n12526), .A2(n12527), .ZN(n12534) );
  NAND2_X1 U11961 ( .A1(n10010), .A2(n10011), .ZN(n12956) );
  NOR2_X1 U11962 ( .A1(n12954), .A2(n15822), .ZN(n12957) );
  NOR2_X1 U11963 ( .A1(n13434), .A2(n12477), .ZN(n12526) );
  NAND2_X1 U11964 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12955), .ZN(
        n12954) );
  OAI21_X1 U11965 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13241), .ZN(n13244) );
  NOR2_X1 U11966 ( .A1(n12922), .A2(n15834), .ZN(n12955) );
  NAND2_X1 U11967 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12922) );
  AND2_X1 U11968 ( .A1(n10120), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9774) );
  INV_X1 U11969 ( .A(n9796), .ZN(n9795) );
  AOI21_X1 U11970 ( .B1(n9796), .B2(n9793), .A(n9694), .ZN(n9792) );
  INV_X1 U11971 ( .A(n9798), .ZN(n9793) );
  INV_X1 U11972 ( .A(n14440), .ZN(n9802) );
  NOR2_X1 U11973 ( .A1(n14196), .A2(n14182), .ZN(n14181) );
  OR2_X1 U11974 ( .A1(n14215), .A2(n13420), .ZN(n14456) );
  OR2_X1 U11975 ( .A1(n14211), .A2(n14194), .ZN(n14196) );
  NAND2_X1 U11976 ( .A1(n14496), .A2(n10120), .ZN(n14451) );
  NOR2_X1 U11977 ( .A1(n14299), .A2(n9939), .ZN(n14277) );
  NAND2_X1 U11978 ( .A1(n14496), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14490) );
  AND2_X1 U11979 ( .A1(n14721), .A2(n14619), .ZN(n14698) );
  NOR3_X1 U11980 ( .A1(n14299), .A2(n14281), .A3(n14293), .ZN(n14282) );
  NOR2_X1 U11981 ( .A1(n14744), .A2(n14396), .ZN(n14398) );
  NAND2_X1 U11982 ( .A1(n14398), .A2(n14387), .ZN(n14389) );
  AND2_X1 U11983 ( .A1(n14777), .A2(n10065), .ZN(n14406) );
  AND2_X1 U11984 ( .A1(n9642), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10123) );
  AND2_X1 U11985 ( .A1(n14551), .A2(n9642), .ZN(n14542) );
  AND2_X1 U11986 ( .A1(n10848), .A2(n10847), .ZN(n14776) );
  NAND2_X1 U11987 ( .A1(n14345), .A2(n9948), .ZN(n14329) );
  AND2_X1 U11988 ( .A1(n14345), .A2(n14336), .ZN(n14338) );
  NAND2_X1 U11989 ( .A1(n14551), .A2(n14617), .ZN(n14771) );
  NAND2_X1 U11990 ( .A1(n14551), .A2(n9641), .ZN(n14769) );
  INV_X1 U11991 ( .A(n14798), .ZN(n10057) );
  AND2_X1 U11992 ( .A1(n13349), .A2(n13348), .ZN(n15756) );
  NAND2_X1 U11993 ( .A1(n10139), .A2(n10136), .ZN(n14824) );
  AND2_X1 U11994 ( .A1(n15784), .A2(n10137), .ZN(n10136) );
  NAND2_X1 U11995 ( .A1(n12866), .A2(n12865), .ZN(n12867) );
  AND2_X1 U11996 ( .A1(n12848), .A2(n12847), .ZN(n12866) );
  NAND2_X1 U11997 ( .A1(n12556), .A2(n12555), .ZN(n12624) );
  AND2_X1 U11998 ( .A1(n12037), .A2(n12036), .ZN(n12625) );
  NOR2_X1 U11999 ( .A1(n12625), .A2(n12624), .ZN(n12847) );
  AND2_X1 U12000 ( .A1(n15907), .A2(n10067), .ZN(n14851) );
  NAND2_X1 U12001 ( .A1(n15907), .A2(n15906), .ZN(n15905) );
  XNOR2_X1 U12002 ( .A(n13424), .B(n13420), .ZN(n14586) );
  XNOR2_X1 U12003 ( .A(n13251), .B(n9934), .ZN(n13250) );
  INV_X1 U12004 ( .A(n13409), .ZN(n13410) );
  NAND2_X1 U12005 ( .A1(n13409), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14875) );
  AOI21_X1 U12006 ( .B1(n12047), .B2(n12050), .A(n12049), .ZN(n13433) );
  INV_X1 U12007 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13033) );
  NAND2_X1 U12008 ( .A1(n12343), .A2(n10383), .ZN(n12395) );
  NOR2_X1 U12009 ( .A1(n12160), .A2(n12254), .ZN(n10813) );
  CLKBUF_X1 U12010 ( .A(n10814), .Z(n10815) );
  BUF_X1 U12011 ( .A(n13216), .Z(n19102) );
  NAND2_X1 U12012 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19405), .ZN(n18898) );
  OR2_X1 U12013 ( .A1(n19160), .A2(n19573), .ZN(n19297) );
  NOR2_X2 U12014 ( .A1(n18859), .A2(n18860), .ZN(n18917) );
  INV_X1 U12015 ( .A(n19352), .ZN(n19544) );
  INV_X1 U12016 ( .A(n15162), .ZN(n15149) );
  AOI21_X1 U12017 ( .B1(n15181), .B2(n15158), .A(n15157), .ZN(n18259) );
  NOR2_X1 U12018 ( .A1(n18276), .A2(n16169), .ZN(n18260) );
  NOR2_X1 U12019 ( .A1(n17146), .A2(n16236), .ZN(n16235) );
  NOR2_X1 U12020 ( .A1(n17185), .A2(n16270), .ZN(n16269) );
  NOR2_X1 U12021 ( .A1(n9739), .A2(n9737), .ZN(n9736) );
  INV_X1 U12022 ( .A(n15248), .ZN(n9740) );
  NOR2_X1 U12023 ( .A1(n9735), .A2(n9734), .ZN(n9733) );
  AND2_X1 U12024 ( .A1(n9923), .A2(n9921), .ZN(n9920) );
  AOI21_X1 U12025 ( .B1(n16734), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n9922), .ZN(n9921) );
  NAND2_X1 U12026 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9923) );
  OAI21_X1 U12027 ( .B1(n9648), .B2(n20625), .A(n10015), .ZN(n9922) );
  NOR2_X1 U12028 ( .A1(n17062), .A2(n17000), .ZN(n17028) );
  NOR2_X1 U12029 ( .A1(n17484), .A2(n15984), .ZN(n16010) );
  INV_X1 U12030 ( .A(n15333), .ZN(n17497) );
  NOR2_X1 U12031 ( .A1(n17156), .A2(n17157), .ZN(n17145) );
  NOR2_X1 U12032 ( .A1(n17533), .A2(n17177), .ZN(n17154) );
  OR2_X1 U12033 ( .A1(n17200), .A2(n16188), .ZN(n17155) );
  NAND4_X1 U12034 ( .A1(n17241), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17199) );
  INV_X1 U12035 ( .A(n17441), .ZN(n16442) );
  NAND2_X1 U12036 ( .A1(n17131), .A2(n17118), .ZN(n15394) );
  NAND2_X1 U12037 ( .A1(n17132), .A2(n17388), .ZN(n15395) );
  NAND2_X1 U12038 ( .A1(n17154), .A2(n17496), .ZN(n15333) );
  NAND2_X1 U12039 ( .A1(n9650), .A2(n15340), .ZN(n17533) );
  INV_X1 U12040 ( .A(n17219), .ZN(n9743) );
  NAND2_X1 U12041 ( .A1(n18301), .A2(n17806), .ZN(n17649) );
  AND2_X1 U12042 ( .A1(n15337), .A2(n17733), .ZN(n17387) );
  NOR2_X1 U12043 ( .A1(n15329), .A2(n17389), .ZN(n17691) );
  NAND2_X1 U12044 ( .A1(n17403), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15327) );
  NAND2_X1 U12045 ( .A1(n17646), .A2(n17784), .ZN(n17688) );
  AND4_X1 U12046 ( .A1(n9753), .A2(n9751), .A3(n9750), .A4(n9748), .ZN(n17390)
         );
  INV_X1 U12047 ( .A(n9749), .ZN(n9748) );
  NAND2_X1 U12048 ( .A1(n17418), .A2(n9755), .ZN(n9750) );
  NOR2_X1 U12049 ( .A1(n17390), .A2(n17733), .ZN(n17389) );
  XNOR2_X1 U12050 ( .A(n10021), .B(n9924), .ZN(n17410) );
  INV_X1 U12051 ( .A(n15297), .ZN(n9924) );
  NOR2_X1 U12052 ( .A1(n17439), .A2(n15318), .ZN(n17433) );
  XNOR2_X1 U12053 ( .A(n15316), .B(n15317), .ZN(n17440) );
  NOR2_X1 U12054 ( .A1(n17440), .A2(n17769), .ZN(n17439) );
  OR2_X1 U12055 ( .A1(n15288), .A2(n15286), .ZN(n10016) );
  INV_X1 U12056 ( .A(n15286), .ZN(n10017) );
  NOR2_X1 U12057 ( .A1(n17486), .A2(n17479), .ZN(n17478) );
  NAND2_X1 U12058 ( .A1(n14989), .A2(n14988), .ZN(n18265) );
  OR3_X1 U12059 ( .A1(n9765), .A2(n15281), .A3(n15280), .ZN(n17487) );
  AOI21_X1 U12060 ( .B1(n15153), .B2(n15152), .A(n16169), .ZN(n18286) );
  INV_X1 U12061 ( .A(n18266), .ZN(n18301) );
  NOR2_X1 U12062 ( .A1(n14976), .A2(n14975), .ZN(n17831) );
  NOR2_X2 U12063 ( .A1(n14966), .A2(n14965), .ZN(n17834) );
  INV_X1 U12064 ( .A(n15148), .ZN(n17843) );
  INV_X1 U12065 ( .A(n15142), .ZN(n17848) );
  BUF_X1 U12066 ( .A(n15986), .Z(n18205) );
  AOI21_X1 U12067 ( .B1(n18265), .B2(n15974), .A(n17619), .ZN(n18268) );
  NAND2_X1 U12068 ( .A1(n12466), .A2(n13463), .ZN(n12371) );
  INV_X1 U12069 ( .A(n12461), .ZN(n19610) );
  NAND2_X1 U12070 ( .A1(n12371), .A2(n12273), .ZN(n20496) );
  NAND2_X1 U12071 ( .A1(n12898), .A2(n12897), .ZN(n19695) );
  INV_X1 U12072 ( .A(n19693), .ZN(n19650) );
  NAND2_X1 U12073 ( .A1(n12898), .A2(n12896), .ZN(n19678) );
  INV_X1 U12074 ( .A(n19695), .ZN(n19708) );
  INV_X1 U12075 ( .A(n19678), .ZN(n19709) );
  AND2_X1 U12076 ( .A1(n19678), .A2(n19646), .ZN(n13640) );
  AND2_X1 U12077 ( .A1(n12898), .A2(n12891), .ZN(n19707) );
  NAND2_X2 U12078 ( .A1(n11911), .A2(n11910), .ZN(n19728) );
  INV_X1 U12079 ( .A(n13756), .ZN(n13750) );
  NAND2_X1 U12080 ( .A1(n12468), .A2(n12467), .ZN(n13764) );
  AOI21_X1 U12081 ( .B1(n12466), .B2(n12465), .A(n12464), .ZN(n12467) );
  OR2_X1 U12082 ( .A1(n13774), .A2(n12471), .ZN(n13766) );
  AOI21_X1 U12083 ( .B1(n15380), .B2(n12356), .A(n12355), .ZN(n19732) );
  INV_X2 U12084 ( .A(n12567), .ZN(n19786) );
  XNOR2_X1 U12085 ( .A(n11842), .B(n11841), .ZN(n13784) );
  INV_X1 U12086 ( .A(n13201), .ZN(n11841) );
  OAI21_X1 U12087 ( .B1(n10115), .B2(n9993), .A(n9991), .ZN(n13853) );
  NAND2_X1 U12088 ( .A1(n10113), .A2(n13164), .ZN(n13186) );
  NAND2_X1 U12089 ( .A1(n15555), .A2(n13115), .ZN(n15552) );
  NAND2_X1 U12090 ( .A1(n13098), .A2(n13097), .ZN(n19791) );
  OR2_X1 U12091 ( .A1(n12450), .A2(n12640), .ZN(n14058) );
  INV_X1 U12092 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20259) );
  INV_X1 U12093 ( .A(n12504), .ZN(n11267) );
  INV_X1 U12094 ( .A(n11266), .ZN(n11268) );
  INV_X1 U12095 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20226) );
  NAND2_X1 U12096 ( .A1(n11288), .A2(n11258), .ZN(n20105) );
  NAND2_X1 U12097 ( .A1(n11344), .A2(n11312), .ZN(n20107) );
  NAND2_X1 U12098 ( .A1(n11288), .A2(n12839), .ZN(n11312) );
  INV_X1 U12099 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19848) );
  NOR2_X1 U12100 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14128) );
  OAI211_X1 U12101 ( .C1(n20132), .C2(n20232), .A(n20167), .B(n20116), .ZN(
        n20134) );
  INV_X1 U12102 ( .A(n20193), .ZN(n20177) );
  OAI22_X1 U12103 ( .A1(n20236), .A2(n20235), .B1(n20287), .B2(n20234), .ZN(
        n20252) );
  NOR2_X2 U12104 ( .A1(n20290), .A2(n20225), .ZN(n20282) );
  NOR2_X2 U12105 ( .A1(n20290), .A2(n20289), .ZN(n20394) );
  NOR2_X1 U12106 ( .A1(n20232), .A2(n13456), .ZN(n15388) );
  INV_X1 U12107 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20400) );
  INV_X1 U12108 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20232) );
  INV_X1 U12109 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20401) );
  AND2_X1 U12110 ( .A1(n10000), .A2(n9999), .ZN(n14197) );
  AND2_X1 U12111 ( .A1(n13382), .A2(n13377), .ZN(n14206) );
  NAND2_X1 U12112 ( .A1(n9984), .A2(n18525), .ZN(n15350) );
  AND2_X1 U12113 ( .A1(n9986), .A2(n15749), .ZN(n9984) );
  NOR2_X1 U12114 ( .A1(n18527), .A2(n9985), .ZN(n15351) );
  AND2_X1 U12115 ( .A1(n19600), .A2(n12940), .ZN(n18639) );
  OR2_X1 U12116 ( .A1(n19600), .A2(n12932), .ZN(n18681) );
  NAND2_X1 U12117 ( .A1(n15964), .A2(n12928), .ZN(n18676) );
  INV_X1 U12118 ( .A(n18656), .ZN(n18689) );
  INV_X1 U12119 ( .A(n18663), .ZN(n18677) );
  INV_X1 U12120 ( .A(n19465), .ZN(n18678) );
  AND2_X1 U12121 ( .A1(n10075), .A2(n10079), .ZN(n10074) );
  INV_X1 U12122 ( .A(n10077), .ZN(n10075) );
  NAND2_X1 U12123 ( .A1(n10079), .A2(n10081), .ZN(n10076) );
  OR2_X1 U12124 ( .A1(n10461), .A2(n10460), .ZN(n12985) );
  OR2_X1 U12125 ( .A1(n10439), .A2(n10438), .ZN(n12864) );
  NOR2_X1 U12126 ( .A1(n10428), .A2(n10427), .ZN(n12851) );
  NAND2_X1 U12127 ( .A1(n12673), .A2(n9628), .ZN(n12532) );
  INV_X1 U12128 ( .A(n14344), .ZN(n14342) );
  XNOR2_X1 U12129 ( .A(n10071), .B(n9714), .ZN(n18696) );
  OAI211_X1 U12130 ( .C1(n14252), .C2(n10081), .A(n10079), .B(n10072), .ZN(
        n12024) );
  NOR2_X1 U12131 ( .A1(n14263), .A2(n14262), .ZN(n14261) );
  NOR2_X1 U12132 ( .A1(n14290), .A2(n10598), .ZN(n14285) );
  INV_X1 U12133 ( .A(n10597), .ZN(n14301) );
  INV_X1 U12134 ( .A(n18757), .ZN(n15723) );
  AND2_X1 U12135 ( .A1(n18755), .A2(n11013), .ZN(n18701) );
  NOR2_X1 U12136 ( .A1(n12663), .A2(n10061), .ZN(n14880) );
  NAND2_X1 U12137 ( .A1(n10063), .A2(n10062), .ZN(n10061) );
  NOR2_X1 U12138 ( .A1(n12663), .A2(n10918), .ZN(n12659) );
  NOR2_X1 U12139 ( .A1(n10360), .A2(n12286), .ZN(n19127) );
  INV_X1 U12140 ( .A(n18755), .ZN(n18756) );
  AND2_X1 U12141 ( .A1(n18755), .A2(n10877), .ZN(n18761) );
  AND2_X1 U12142 ( .A1(n18755), .A2(n11000), .ZN(n18757) );
  INV_X1 U12143 ( .A(n12935), .ZN(n12310) );
  NOR2_X1 U12144 ( .A1(n18817), .A2(n18545), .ZN(n9781) );
  INV_X1 U12145 ( .A(n15753), .ZN(n9780) );
  NAND2_X1 U12146 ( .A1(n15752), .A2(n18819), .ZN(n9782) );
  INV_X1 U12147 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18625) );
  INV_X1 U12148 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15822) );
  INV_X1 U12149 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15834) );
  INV_X1 U12150 ( .A(n18819), .ZN(n15828) );
  NAND2_X1 U12151 ( .A1(n12214), .A2(n12213), .ZN(n15833) );
  INV_X1 U12152 ( .A(n10142), .ZN(n14478) );
  AND2_X1 U12153 ( .A1(n10146), .A2(n10144), .ZN(n14476) );
  NAND2_X1 U12154 ( .A1(n10146), .A2(n10147), .ZN(n14485) );
  NAND2_X1 U12155 ( .A1(n9836), .A2(n9840), .ZN(n14720) );
  NAND2_X1 U12156 ( .A1(n10130), .A2(n9841), .ZN(n9836) );
  AOI21_X1 U12157 ( .B1(n10130), .B2(n10124), .A(n9613), .ZN(n14734) );
  NAND2_X1 U12158 ( .A1(n14768), .A2(n14767), .ZN(n9784) );
  INV_X1 U12159 ( .A(n14766), .ZN(n9783) );
  INV_X1 U12160 ( .A(n18853), .ZN(n15894) );
  AND2_X1 U12161 ( .A1(n10127), .A2(n9637), .ZN(n14577) );
  INV_X1 U12162 ( .A(n10126), .ZN(n14503) );
  AND2_X1 U12163 ( .A1(n10135), .A2(n10137), .ZN(n15782) );
  NAND2_X1 U12164 ( .A1(n10135), .A2(n10157), .ZN(n14845) );
  INV_X1 U12165 ( .A(n18832), .ZN(n18847) );
  AND2_X1 U12166 ( .A1(n12834), .A2(n19584), .ZN(n18846) );
  NAND2_X1 U12167 ( .A1(n14605), .A2(n14789), .ZN(n18854) );
  INV_X1 U12168 ( .A(n19127), .ZN(n19573) );
  INV_X1 U12169 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19560) );
  AND2_X1 U12170 ( .A1(n12351), .A2(n12350), .ZN(n19563) );
  NAND2_X1 U12171 ( .A1(n12343), .A2(n12346), .ZN(n19555) );
  OR2_X1 U12172 ( .A1(n18955), .A2(n19162), .ZN(n18974) );
  OAI21_X1 U12173 ( .B1(n19018), .B2(n19017), .A(n19016), .ZN(n19036) );
  AND2_X1 U12174 ( .A1(n19098), .A2(n19304), .ZN(n19094) );
  INV_X1 U12175 ( .A(n19183), .ZN(n19186) );
  NOR2_X1 U12176 ( .A1(n19297), .A2(n19161), .ZN(n19210) );
  OAI22_X1 U12177 ( .A1(n18896), .A2(n18909), .B1(n18895), .B2(n18907), .ZN(
        n19382) );
  OAI21_X1 U12178 ( .B1(n19364), .B2(n19363), .A(n19362), .ZN(n19393) );
  INV_X1 U12179 ( .A(n19367), .ZN(n19407) );
  INV_X1 U12180 ( .A(n19377), .ZN(n19423) );
  INV_X1 U12181 ( .A(n19456), .ZN(n19436) );
  INV_X1 U12182 ( .A(n19385), .ZN(n19435) );
  INV_X1 U12183 ( .A(n19390), .ZN(n19443) );
  NOR2_X1 U12184 ( .A1(n19353), .A2(n19352), .ZN(n19452) );
  NAND2_X1 U12185 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10837), .ZN(n19458) );
  NOR2_X1 U12186 ( .A1(n18260), .A2(n17062), .ZN(n18488) );
  NAND2_X1 U12187 ( .A1(n15177), .A2(n15150), .ZN(n16151) );
  NAND3_X1 U12188 ( .A1(n17853), .A2(n15149), .A3(n17001), .ZN(n17063) );
  NAND2_X1 U12189 ( .A1(n18470), .A2(n18259), .ZN(n17062) );
  NOR2_X1 U12190 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16344), .ZN(n16329) );
  NOR2_X1 U12191 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16413), .ZN(n16402) );
  NOR2_X1 U12192 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16437), .ZN(n16417) );
  INV_X1 U12193 ( .A(n16539), .ZN(n16525) );
  AND2_X1 U12194 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16610), .ZN(n16625) );
  NOR2_X1 U12195 ( .A1(n16777), .A2(n16774), .ZN(n16758) );
  NAND2_X1 U12196 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16758), .ZN(n16757) );
  INV_X1 U12197 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20519) );
  INV_X1 U12198 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20629) );
  AND2_X1 U12199 ( .A1(n16841), .A2(n16818), .ZN(n16827) );
  NAND2_X1 U12200 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16827), .ZN(n16826) );
  INV_X1 U12201 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16843) );
  INV_X1 U12202 ( .A(n16849), .ZN(n16841) );
  INV_X2 U12203 ( .A(n16850), .ZN(n16847) );
  NAND4_X1 U12204 ( .A1(n18470), .A2(n18472), .A3(n17001), .A4(n15410), .ZN(
        n16849) );
  INV_X1 U12205 ( .A(n16834), .ZN(n16850) );
  NOR2_X1 U12206 ( .A1(n17004), .A2(n16871), .ZN(n16864) );
  INV_X1 U12207 ( .A(n16876), .ZN(n16872) );
  NAND2_X1 U12208 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n16872), .ZN(n16871) );
  INV_X1 U12209 ( .A(n16890), .ZN(n16886) );
  INV_X1 U12210 ( .A(n16911), .ZN(n16907) );
  NOR2_X1 U12211 ( .A1(n17021), .A2(n16920), .ZN(n16915) );
  NAND2_X1 U12212 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n16921), .ZN(n16920) );
  NAND2_X1 U12213 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n16936), .ZN(n16932) );
  INV_X1 U12214 ( .A(n16879), .ZN(n16930) );
  INV_X1 U12215 ( .A(n16905), .ZN(n16931) );
  NOR2_X1 U12216 ( .A1(n15242), .A2(n15241), .ZN(n16984) );
  NOR2_X1 U12217 ( .A1(n18467), .A2(n17028), .ZN(n17047) );
  INV_X1 U12219 ( .A(n17110), .ZN(n17101) );
  NOR2_X1 U12220 ( .A1(n17125), .A2(n17126), .ZN(n16008) );
  INV_X1 U12221 ( .A(n17292), .ZN(n17212) );
  NOR2_X1 U12222 ( .A1(n17199), .A2(n17200), .ZN(n17195) );
  INV_X1 U12223 ( .A(n17117), .ZN(n17399) );
  NAND2_X1 U12224 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17441) );
  NOR2_X1 U12225 ( .A1(n17457), .A2(n17318), .ZN(n17485) );
  NAND2_X1 U12226 ( .A1(n17267), .A2(n17346), .ZN(n17480) );
  OAI21_X1 U12227 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18469), .A(n16152), 
        .ZN(n17488) );
  INV_X1 U12228 ( .A(n17481), .ZN(n17491) );
  INV_X1 U12229 ( .A(n17688), .ZN(n17725) );
  NOR2_X1 U12230 ( .A1(n17649), .A2(n18282), .ZN(n17722) );
  AOI21_X1 U12231 ( .B1(n15333), .B2(n18264), .A(n9762), .ZN(n17509) );
  NAND2_X1 U12232 ( .A1(n9764), .A2(n9763), .ZN(n9762) );
  NOR3_X1 U12233 ( .A1(n17519), .A2(n17500), .A3(n17499), .ZN(n9763) );
  OR2_X1 U12234 ( .A1(n17498), .A2(n17688), .ZN(n9764) );
  INV_X1 U12235 ( .A(n17205), .ZN(n17233) );
  NAND2_X1 U12236 ( .A1(n9747), .A2(n9755), .ZN(n17404) );
  NAND2_X1 U12237 ( .A1(n10027), .A2(n10028), .ZN(n17416) );
  AND2_X1 U12238 ( .A1(n10027), .A2(n10025), .ZN(n17414) );
  NAND2_X1 U12239 ( .A1(n17428), .A2(n10029), .ZN(n10027) );
  INV_X1 U12240 ( .A(n10020), .ZN(n17452) );
  AND2_X1 U12241 ( .A1(n10020), .A2(n10019), .ZN(n17450) );
  NAND2_X1 U12242 ( .A1(n10018), .A2(n10017), .ZN(n10020) );
  NOR2_X1 U12243 ( .A1(n17829), .A2(n15166), .ZN(n18451) );
  INV_X1 U12244 ( .A(n18315), .ZN(n18470) );
  NOR2_X1 U12245 ( .A1(n18475), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18326) );
  AND2_X1 U12246 ( .A1(n12146), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19852)
         );
  INV_X1 U12248 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20527) );
  AOI21_X1 U12249 ( .B1(n13700), .B2(n19794), .A(n13209), .ZN(n13210) );
  INV_X1 U12250 ( .A(n13953), .ZN(n9853) );
  NAND2_X1 U12251 ( .A1(n9855), .A2(n19825), .ZN(n9854) );
  OAI21_X1 U12252 ( .B1(n14173), .B2(n9988), .A(n9664), .ZN(P2_U2825) );
  INV_X1 U12253 ( .A(n9989), .ZN(n9988) );
  AOI21_X1 U12254 ( .B1(n14174), .B2(n14437), .A(n19465), .ZN(n9989) );
  OAI211_X1 U12255 ( .C1(n14631), .C2(n15817), .A(n10119), .B(n9653), .ZN(
        P2_U2983) );
  AOI21_X1 U12256 ( .B1(n14627), .B2(n18819), .A(n13431), .ZN(n10119) );
  OAI21_X1 U12257 ( .B1(n14643), .B2(n15817), .A(n9724), .ZN(P2_U2984) );
  AOI21_X1 U12258 ( .B1(n14641), .B2(n18814), .A(n9725), .ZN(n9724) );
  NAND2_X1 U12259 ( .A1(n9623), .A2(n9710), .ZN(n9725) );
  OAI21_X1 U12260 ( .B1(n15750), .B2(n15817), .A(n9777), .ZN(P2_U2996) );
  AOI21_X1 U12261 ( .B1(n15751), .B2(n18814), .A(n9778), .ZN(n9777) );
  NAND2_X1 U12262 ( .A1(n9782), .A2(n9779), .ZN(n9778) );
  NOR2_X1 U12263 ( .A1(n9781), .A2(n9780), .ZN(n9779) );
  OAI21_X1 U12264 ( .B1(n14804), .B2(n9892), .A(n9891), .ZN(n14795) );
  AOI211_X1 U12265 ( .C1(n9720), .C2(n16472), .A(n9597), .B(n16471), .ZN(
        n16478) );
  AOI21_X1 U12266 ( .B1(n16994), .B2(BUF2_REG_1__SCAN_IN), .A(n9918), .ZN(
        n16998) );
  OAI21_X1 U12267 ( .B1(n16005), .B2(n17402), .A(n10033), .ZN(P3_U2800) );
  AOI21_X1 U12268 ( .B1(n10035), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10034), .ZN(n10033) );
  OR2_X1 U12269 ( .A1(n16017), .A2(n16015), .ZN(n10035) );
  OAI21_X1 U12270 ( .B1(n16005), .B2(n17727), .A(n9659), .ZN(P3_U2832) );
  NAND2_X1 U12271 ( .A1(n9597), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n9928) );
  OR2_X1 U12272 ( .A1(n15399), .A2(n16004), .ZN(n9931) );
  AND2_X1 U12273 ( .A1(n16046), .A2(n16048), .ZN(n9732) );
  OR2_X1 U12274 ( .A1(n10622), .A2(n14302), .ZN(n9611) );
  OR2_X1 U12275 ( .A1(n15322), .A2(n15323), .ZN(n9612) );
  NAND2_X1 U12276 ( .A1(n9663), .A2(n9622), .ZN(n9613) );
  NAND2_X1 U12277 ( .A1(n10484), .A2(n9916), .ZN(n14325) );
  NAND2_X1 U12278 ( .A1(n10484), .A2(n10483), .ZN(n13083) );
  AND2_X1 U12279 ( .A1(n9619), .A2(n9968), .ZN(n9614) );
  NAND2_X1 U12280 ( .A1(n10045), .A2(n11504), .ZN(n13688) );
  NAND2_X1 U12281 ( .A1(n13289), .A2(n13288), .ZN(n14589) );
  AND2_X1 U12282 ( .A1(n14496), .A2(n10121), .ZN(n9616) );
  AND4_X1 U12283 ( .A1(n15255), .A2(n15254), .A3(n15253), .A4(n15252), .ZN(
        n9617) );
  AND2_X1 U12284 ( .A1(n9969), .A2(n9688), .ZN(n9619) );
  OR2_X1 U12285 ( .A1(n9837), .A2(n9679), .ZN(n9620) );
  AND4_X1 U12286 ( .A1(n13237), .A2(n13236), .A3(n13235), .A4(n13234), .ZN(
        n9621) );
  NOR2_X1 U12287 ( .A1(n14513), .A2(n14515), .ZN(n9622) );
  AOI21_X1 U12288 ( .B1(n13890), .B2(n13195), .A(n9691), .ZN(n13194) );
  INV_X1 U12289 ( .A(n13194), .ZN(n9827) );
  OR2_X1 U12290 ( .A1(n14639), .A2(n15828), .ZN(n9623) );
  OR2_X1 U12291 ( .A1(n9615), .A2(n10116), .ZN(n9624) );
  OR2_X1 U12292 ( .A1(n17346), .A2(n16196), .ZN(n9625) );
  AND2_X1 U12293 ( .A1(n9680), .A2(n9936), .ZN(n9626) );
  AND2_X1 U12294 ( .A1(n10063), .A2(n9657), .ZN(n9627) );
  INV_X1 U12295 ( .A(n9615), .ZN(n10117) );
  NAND2_X1 U12296 ( .A1(n9906), .A2(n10416), .ZN(n12623) );
  AND2_X1 U12297 ( .A1(n10484), .A2(n9685), .ZN(n14334) );
  AND2_X1 U12298 ( .A1(n12672), .A2(n9711), .ZN(n9628) );
  AND2_X1 U12299 ( .A1(n10006), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9629) );
  AND2_X1 U12300 ( .A1(n9971), .A2(n12090), .ZN(n9630) );
  INV_X1 U12301 ( .A(n10091), .ZN(n14321) );
  OR3_X1 U12302 ( .A1(n15472), .A2(n9867), .A3(n9676), .ZN(n9631) );
  AND2_X1 U12303 ( .A1(n10059), .A2(n14810), .ZN(n9632) );
  AND2_X1 U12304 ( .A1(n9902), .A2(n13545), .ZN(n9633) );
  AND2_X1 U12305 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9634)
         );
  AND2_X1 U12306 ( .A1(n11343), .A2(n11363), .ZN(n9635) );
  AND2_X1 U12307 ( .A1(n9630), .A2(n14311), .ZN(n9636) );
  INV_X1 U12308 ( .A(n15817), .ZN(n18811) );
  NAND2_X1 U12309 ( .A1(n13310), .A2(n15770), .ZN(n9637) );
  AND2_X1 U12310 ( .A1(n10013), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9638) );
  AND2_X1 U12311 ( .A1(n10002), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9639) );
  AND2_X1 U12312 ( .A1(n9707), .A2(n9974), .ZN(n9640) );
  AND2_X1 U12313 ( .A1(n14617), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9641) );
  AND2_X1 U12314 ( .A1(n9641), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9642) );
  AND2_X1 U12315 ( .A1(n10121), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9643) );
  AND2_X1 U12316 ( .A1(n9774), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9644) );
  OR2_X1 U12317 ( .A1(n18913), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9645) );
  AND2_X2 U12318 ( .A1(n9607), .A2(n15934), .ZN(n10404) );
  AND2_X2 U12319 ( .A1(n10754), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10444) );
  AND2_X2 U12320 ( .A1(n10753), .A2(n15934), .ZN(n10499) );
  OR2_X1 U12321 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n13371), .ZN(n9649) );
  NOR3_X1 U12322 ( .A1(n17691), .A2(n17329), .A3(n9758), .ZN(n9650) );
  AOI21_X1 U12323 ( .B1(n13116), .B2(n11514), .A(n11381), .ZN(n13011) );
  AND3_X1 U12324 ( .A1(n15258), .A2(n15257), .A3(n9920), .ZN(n9651) );
  NOR2_X1 U12325 ( .A1(n17419), .A2(n17747), .ZN(n17418) );
  NAND2_X1 U12326 ( .A1(n10313), .A2(n10312), .ZN(n10346) );
  INV_X2 U12327 ( .A(n11946), .ZN(n11933) );
  AND2_X1 U12328 ( .A1(n10385), .A2(n10083), .ZN(n12394) );
  AND2_X1 U12329 ( .A1(n13303), .A2(n9619), .ZN(n9652) );
  OR2_X1 U12330 ( .A1(n14628), .A2(n15816), .ZN(n9653) );
  INV_X1 U12331 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10773) );
  AND4_X1 U12332 ( .A1(n14510), .A2(n14557), .A3(n14564), .A4(n13341), .ZN(
        n9655) );
  OR2_X1 U12333 ( .A1(n14299), .A2(n14293), .ZN(n9656) );
  AND2_X1 U12334 ( .A1(n10062), .A2(n14881), .ZN(n9657) );
  INV_X1 U12335 ( .A(n9842), .ZN(n9841) );
  OAI21_X1 U12336 ( .B1(n10124), .B2(n9613), .A(n9843), .ZN(n9842) );
  OR2_X1 U12337 ( .A1(n9615), .A2(n13930), .ZN(n9658) );
  INV_X2 U12338 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15934) );
  AND3_X1 U12339 ( .A1(n9931), .A2(n9929), .A3(n9928), .ZN(n9659) );
  OR2_X1 U12340 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n13301), .ZN(n9660) );
  NAND2_X1 U12341 ( .A1(n14496), .A2(n9643), .ZN(n10122) );
  AND2_X1 U12342 ( .A1(n9614), .A2(n9804), .ZN(n9661) );
  OR2_X1 U12343 ( .A1(n9993), .A2(n9990), .ZN(n9662) );
  NOR2_X1 U12344 ( .A1(n13668), .A2(n13669), .ZN(n13569) );
  NOR2_X1 U12345 ( .A1(n9863), .A2(n9862), .ZN(n13532) );
  INV_X1 U12346 ( .A(n13532), .ZN(n9861) );
  AND3_X1 U12347 ( .A1(n14512), .A2(n13354), .A3(n14765), .ZN(n9663) );
  AND2_X1 U12348 ( .A1(n9987), .A2(n14180), .ZN(n9664) );
  AND2_X1 U12349 ( .A1(n15550), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9665) );
  OR2_X1 U12350 ( .A1(n13668), .A2(n10051), .ZN(n9666) );
  AND2_X1 U12351 ( .A1(n9615), .A2(n13930), .ZN(n9667) );
  NAND2_X1 U12352 ( .A1(n11488), .A2(n11487), .ZN(n13638) );
  NAND2_X1 U12353 ( .A1(n13327), .A2(n9630), .ZN(n9972) );
  NOR2_X1 U12354 ( .A1(n13668), .A2(n10048), .ZN(n13555) );
  NOR2_X1 U12355 ( .A1(n13530), .A2(n13519), .ZN(n13507) );
  INV_X1 U12356 ( .A(n13910), .ZN(n13889) );
  AND2_X1 U12357 ( .A1(n10032), .A2(n10031), .ZN(n9668) );
  NAND2_X1 U12358 ( .A1(n10088), .A2(n9905), .ZN(n9669) );
  AND3_X1 U12359 ( .A1(n19887), .A2(n12469), .A3(n10095), .ZN(n9670) );
  AND2_X1 U12360 ( .A1(n9612), .A2(n9746), .ZN(n9671) );
  INV_X1 U12361 ( .A(n12779), .ZN(n10271) );
  AND2_X1 U12362 ( .A1(n11846), .A2(n11843), .ZN(n9672) );
  OR2_X1 U12363 ( .A1(n10099), .A2(n9879), .ZN(n9673) );
  OR2_X1 U12364 ( .A1(n17141), .A2(n16004), .ZN(n9674) );
  NAND4_X1 U12365 ( .A1(n9832), .A2(n9831), .A3(n19992), .A4(n9635), .ZN(n9675) );
  AND2_X1 U12366 ( .A1(n11023), .A2(n12484), .ZN(n11298) );
  INV_X1 U12367 ( .A(n11278), .ZN(n11394) );
  INV_X1 U12368 ( .A(n11394), .ZN(n13203) );
  OR2_X1 U12369 ( .A1(n13592), .A2(n13591), .ZN(n9676) );
  INV_X1 U12370 ( .A(n10360), .ZN(n13037) );
  AND2_X1 U12371 ( .A1(n12850), .A2(n12864), .ZN(n12858) );
  INV_X1 U12372 ( .A(n15299), .ZN(n9927) );
  NAND2_X1 U12373 ( .A1(n19592), .A2(n19571), .ZN(n10861) );
  INV_X1 U12374 ( .A(n10861), .ZN(n14161) );
  INV_X1 U12375 ( .A(n12954), .ZN(n10010) );
  AND3_X1 U12376 ( .A1(n11396), .A2(n11397), .A3(n10043), .ZN(n13061) );
  NOR2_X1 U12377 ( .A1(n14325), .A2(n10092), .ZN(n14313) );
  AND2_X1 U12378 ( .A1(n14809), .A2(n9632), .ZN(n9677) );
  AND2_X1 U12379 ( .A1(n12962), .A2(n10006), .ZN(n9678) );
  NOR3_X1 U12380 ( .A1(n15705), .A2(n13420), .A3(n14727), .ZN(n9679) );
  AND2_X1 U12381 ( .A1(n9937), .A2(n12865), .ZN(n9680) );
  AND2_X1 U12382 ( .A1(n10067), .A2(n14852), .ZN(n9681) );
  AND2_X1 U12383 ( .A1(n10484), .A2(n9915), .ZN(n14305) );
  AND3_X1 U12384 ( .A1(n11396), .A2(n11397), .A3(n10042), .ZN(n9682) );
  OR2_X1 U12385 ( .A1(n10963), .A2(n10962), .ZN(n13426) );
  INV_X1 U12386 ( .A(n13426), .ZN(n13420) );
  INV_X1 U12387 ( .A(n13250), .ZN(n14870) );
  NOR2_X1 U12388 ( .A1(n18472), .A2(n17619), .ZN(n18264) );
  AND2_X1 U12389 ( .A1(n12866), .A2(n9626), .ZN(n9683) );
  NAND2_X1 U12390 ( .A1(n10380), .A2(n10379), .ZN(n12343) );
  INV_X1 U12391 ( .A(n12951), .ZN(n9970) );
  NOR3_X1 U12392 ( .A1(n13387), .A2(n13420), .A3(n14612), .ZN(n9684) );
  AND2_X1 U12393 ( .A1(n9917), .A2(n10483), .ZN(n9685) );
  OR2_X1 U12394 ( .A1(n17691), .A2(n17329), .ZN(n9761) );
  AND2_X1 U12395 ( .A1(n9633), .A2(n13531), .ZN(n9686) );
  NOR2_X1 U12396 ( .A1(n14285), .A2(n14284), .ZN(n9687) );
  INV_X1 U12397 ( .A(n13914), .ZN(n9982) );
  NAND2_X1 U12398 ( .A1(n18899), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n9688) );
  AND2_X1 U12399 ( .A1(n10009), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9689) );
  AND2_X1 U12400 ( .A1(n18899), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n9690) );
  NOR2_X1 U12401 ( .A1(n14325), .A2(n14326), .ZN(n10091) );
  NOR2_X1 U12402 ( .A1(n15472), .A2(n9864), .ZN(n9869) );
  NAND2_X1 U12403 ( .A1(n13893), .A2(n13193), .ZN(n9691) );
  AND2_X1 U12404 ( .A1(n9955), .A2(n14121), .ZN(n9692) );
  AND2_X1 U12405 ( .A1(n11729), .A2(n11728), .ZN(n13545) );
  OR2_X1 U12406 ( .A1(n10046), .A2(n10044), .ZN(n9693) );
  INV_X1 U12407 ( .A(n10101), .ZN(n13453) );
  NAND2_X1 U12408 ( .A1(n11161), .A2(n11120), .ZN(n10101) );
  INV_X1 U12409 ( .A(n9965), .ZN(n13246) );
  OR2_X1 U12410 ( .A1(n12773), .A2(n12774), .ZN(n9965) );
  INV_X1 U12411 ( .A(n9956), .ZN(n9955) );
  NOR2_X1 U12412 ( .A1(n9615), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9956) );
  OR2_X1 U12413 ( .A1(n9684), .A2(n9802), .ZN(n9694) );
  NOR2_X1 U12414 ( .A1(n14504), .A2(n10132), .ZN(n9695) );
  AND2_X1 U12415 ( .A1(n10084), .A2(n10341), .ZN(n9696) );
  AND2_X1 U12416 ( .A1(n12746), .A2(n9771), .ZN(n9697) );
  AND2_X1 U12417 ( .A1(n10058), .A2(n10057), .ZN(n9698) );
  AND2_X1 U12418 ( .A1(n10090), .A2(n14314), .ZN(n9699) );
  AND2_X1 U12419 ( .A1(n9681), .A2(n10066), .ZN(n9700) );
  AND2_X1 U12420 ( .A1(n9635), .A2(n11383), .ZN(n9701) );
  AND2_X1 U12421 ( .A1(n9626), .A2(n13014), .ZN(n9702) );
  INV_X1 U12422 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14147) );
  INV_X1 U12423 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14594) );
  OR2_X1 U12424 ( .A1(n15325), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9703) );
  AND2_X1 U12425 ( .A1(n9890), .A2(n13406), .ZN(n9704) );
  INV_X1 U12426 ( .A(n12575), .ZN(n19767) );
  NAND2_X1 U12427 ( .A1(n12673), .A2(n12672), .ZN(n12476) );
  NOR2_X1 U12428 ( .A1(n13152), .A2(n13153), .ZN(n9850) );
  OR2_X1 U12429 ( .A1(n12450), .A2(n12427), .ZN(n19838) );
  INV_X1 U12430 ( .A(n19838), .ZN(n19823) );
  AND2_X1 U12431 ( .A1(n14152), .A2(n10002), .ZN(n9705) );
  AND2_X1 U12432 ( .A1(n12850), .A2(n10089), .ZN(n9706) );
  INV_X1 U12433 ( .A(n18525), .ZN(n18527) );
  AND2_X1 U12434 ( .A1(n9975), .A2(n13355), .ZN(n9707) );
  AND3_X1 U12435 ( .A1(n15348), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n13426), .ZN(n9708) );
  AND4_X1 U12436 ( .A1(n17313), .A2(n17635), .A3(n17349), .A4(n17660), .ZN(
        n9709) );
  INV_X1 U12437 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11277) );
  INV_X1 U12438 ( .A(n14464), .ZN(n9999) );
  INV_X1 U12439 ( .A(n10623), .ZN(n10087) );
  OR2_X1 U12440 ( .A1(n10772), .A2(n10771), .ZN(n13405) );
  INV_X1 U12441 ( .A(n13405), .ZN(n10134) );
  AND2_X1 U12442 ( .A1(n14438), .A2(n14439), .ZN(n9710) );
  INV_X1 U12443 ( .A(n12558), .ZN(n9906) );
  INV_X1 U12444 ( .A(n13523), .ZN(n9860) );
  INV_X1 U12445 ( .A(n14302), .ZN(n9913) );
  AND2_X1 U12446 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9711) );
  AND2_X1 U12447 ( .A1(n10065), .A2(n14405), .ZN(n9712) );
  AND2_X1 U12448 ( .A1(n12673), .A2(n9634), .ZN(n9713) );
  INV_X1 U12449 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n9978) );
  INV_X1 U12450 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n9804) );
  AND2_X1 U12451 ( .A1(n14163), .A2(n14162), .ZN(n9714) );
  INV_X1 U12452 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U12453 ( .A1(n11956), .A2(n11955), .ZN(n9715) );
  AND2_X1 U12454 ( .A1(n10070), .A2(n14183), .ZN(n9716) );
  AND2_X1 U12455 ( .A1(n10719), .A2(n10718), .ZN(n9717) );
  INV_X1 U12456 ( .A(n13966), .ZN(n9882) );
  AND2_X1 U12457 ( .A1(n15572), .A2(n14054), .ZN(n9718) );
  INV_X1 U12458 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U12459 ( .A1(n9882), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9719) );
  INV_X1 U12460 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9925) );
  INV_X1 U12461 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10008) );
  INV_X1 U12462 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n15967) );
  INV_X1 U12463 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9990) );
  INV_X1 U12464 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10004) );
  INV_X1 U12465 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10014) );
  OAI221_X1 U12466 ( .B1(n20017), .B2(n20232), .C1(n20017), .C2(n20001), .A(
        n20297), .ZN(n20019) );
  NOR3_X2 U12467 ( .A1(n18166), .A2(n18119), .A3(n18090), .ZN(n18085) );
  AOI22_X2 U12468 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18916), .ZN(n19410) );
  NOR2_X2 U12469 ( .A1(n18861), .A2(n18860), .ZN(n18916) );
  NOR3_X2 U12470 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18166), .A3(
        n18044), .ZN(n18012) );
  NOR2_X2 U12471 ( .A1(n18419), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18166) );
  CLKBUF_X1 U12472 ( .A(n16500), .Z(n9720) );
  INV_X1 U12473 ( .A(n9720), .ZN(n18330) );
  NOR4_X2 U12474 ( .A1(n9597), .A2(n18488), .A3(n9720), .A4(n18320), .ZN(
        n16529) );
  NOR4_X1 U12475 ( .A1(n18429), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_0__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n16500)
         );
  NOR2_X1 U12476 ( .A1(n19896), .A2(n10095), .ZN(n9721) );
  NOR2_X1 U12477 ( .A1(n16209), .A2(n16208), .ZN(n16207) );
  NOR2_X1 U12478 ( .A1(n17168), .A2(n16257), .ZN(n16256) );
  NOR2_X1 U12479 ( .A1(n16249), .A2(n16248), .ZN(n16247) );
  NOR2_X1 U12480 ( .A1(n16281), .A2(n16280), .ZN(n16279) );
  NOR2_X1 U12481 ( .A1(n17231), .A2(n16299), .ZN(n16298) );
  INV_X1 U12482 ( .A(n9885), .ZN(n13779) );
  NAND2_X1 U12483 ( .A1(n13808), .A2(n13981), .ZN(n13786) );
  NAND2_X1 U12484 ( .A1(n9896), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U12485 ( .A1(n10096), .A2(n11153), .ZN(n11196) );
  XNOR2_X1 U12486 ( .A(n11196), .B(n11195), .ZN(n11276) );
  XNOR2_X2 U12487 ( .A(n12047), .B(n12050), .ZN(n12713) );
  NAND2_X2 U12488 ( .A1(n10369), .A2(n10328), .ZN(n12047) );
  NAND3_X2 U12489 ( .A1(n10364), .A2(n10365), .A3(n10363), .ZN(n10369) );
  AND2_X2 U12490 ( .A1(n10328), .A2(n10307), .ZN(n10365) );
  NAND2_X1 U12491 ( .A1(n10327), .A2(n10349), .ZN(n10364) );
  NAND3_X1 U12492 ( .A1(n9723), .A2(n10816), .A3(n18913), .ZN(n12807) );
  NAND3_X1 U12493 ( .A1(n10823), .A2(n10822), .A3(n9722), .ZN(n12786) );
  AND2_X1 U12494 ( .A1(n12808), .A2(n9723), .ZN(n9722) );
  NAND2_X1 U12495 ( .A1(n10821), .A2(n18892), .ZN(n9723) );
  AND2_X2 U12496 ( .A1(n9728), .A2(n9726), .ZN(n14876) );
  NAND2_X1 U12497 ( .A1(n9727), .A2(n14895), .ZN(n9726) );
  NAND2_X1 U12498 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9727) );
  NAND2_X1 U12499 ( .A1(n9729), .A2(n14894), .ZN(n9728) );
  INV_X1 U12500 ( .A(n14896), .ZN(n9729) );
  NOR2_X2 U12501 ( .A1(n9730), .A2(n12719), .ZN(n13233) );
  NOR2_X2 U12502 ( .A1(n9730), .A2(n12734), .ZN(n13232) );
  NAND2_X1 U12503 ( .A1(n12714), .A2(n13001), .ZN(n9730) );
  NOR2_X4 U12504 ( .A1(n14519), .A2(n14739), .ZN(n15741) );
  NAND3_X1 U12505 ( .A1(n16045), .A2(n16047), .A3(n9732), .ZN(P3_U2834) );
  NAND3_X1 U12506 ( .A1(n9740), .A2(n9736), .A3(n9733), .ZN(n15306) );
  NAND3_X1 U12507 ( .A1(n15249), .A2(n15245), .A3(n9738), .ZN(n9737) );
  NAND2_X1 U12508 ( .A1(n15337), .A2(n9742), .ZN(n9741) );
  NAND2_X1 U12509 ( .A1(n9756), .A2(n9671), .ZN(n9753) );
  INV_X1 U12510 ( .A(n17418), .ZN(n9756) );
  NAND2_X1 U12511 ( .A1(n9756), .A2(n9612), .ZN(n9747) );
  OAI21_X1 U12512 ( .B1(n9612), .B2(n15326), .A(n9703), .ZN(n9749) );
  NAND2_X1 U12513 ( .A1(n17403), .A2(n9752), .ZN(n9751) );
  INV_X1 U12514 ( .A(n15326), .ZN(n9755) );
  INV_X2 U12515 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18443) );
  INV_X1 U12516 ( .A(n9761), .ZN(n17665) );
  NAND3_X1 U12517 ( .A1(n15283), .A2(n15282), .A3(n9766), .ZN(n9765) );
  NAND2_X1 U12518 ( .A1(n15801), .A2(n15799), .ZN(n13429) );
  NAND2_X1 U12519 ( .A1(n14588), .A2(n13421), .ZN(n9767) );
  NAND3_X1 U12520 ( .A1(n9772), .A2(n9697), .A3(n9770), .ZN(n13408) );
  AND2_X2 U12521 ( .A1(n9768), .A2(n13239), .ZN(n13254) );
  NAND3_X1 U12522 ( .A1(n13228), .A2(n9621), .A3(n9769), .ZN(n9768) );
  INV_X1 U12523 ( .A(n12737), .ZN(n19267) );
  NAND2_X1 U12524 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n9773) );
  NAND2_X1 U12525 ( .A1(n12770), .A2(n12771), .ZN(n9890) );
  NAND3_X1 U12526 ( .A1(n9890), .A2(n13406), .A3(n13420), .ZN(n9776) );
  NOR2_X1 U12527 ( .A1(n10911), .A2(n9791), .ZN(n9790) );
  OR2_X2 U12528 ( .A1(n9845), .A2(n9801), .ZN(n9800) );
  INV_X1 U12529 ( .A(n12774), .ZN(n9807) );
  NAND2_X2 U12530 ( .A1(n14495), .A2(n10148), .ZN(n10146) );
  NAND3_X1 U12531 ( .A1(n9982), .A2(n9819), .A3(n9983), .ZN(n13902) );
  XNOR2_X1 U12532 ( .A(n13915), .B(n9819), .ZN(n14092) );
  NAND3_X1 U12533 ( .A1(n9824), .A2(n9822), .A3(n9821), .ZN(n9828) );
  NAND3_X1 U12534 ( .A1(n9832), .A2(n9831), .A3(n9829), .ZN(n13137) );
  NAND3_X1 U12535 ( .A1(n9830), .A2(n9832), .A3(n9831), .ZN(n9981) );
  OAI21_X2 U12536 ( .B1(n13786), .B2(n9834), .A(n9833), .ZN(n9885) );
  NAND2_X2 U12537 ( .A1(n9849), .A2(n9848), .ZN(n10126) );
  NAND3_X1 U12538 ( .A1(n9949), .A2(n9854), .A3(n9853), .ZN(P1_U3000) );
  NOR2_X1 U12539 ( .A1(n13561), .A2(n13547), .ZN(n13546) );
  INV_X1 U12540 ( .A(n9869), .ZN(n13671) );
  AND2_X4 U12541 ( .A1(n11024), .A2(n14110), .ZN(n11816) );
  AND2_X2 U12542 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14110) );
  NAND2_X1 U12543 ( .A1(n9871), .A2(n9870), .ZN(n15547) );
  NAND3_X1 U12544 ( .A1(n10103), .A2(n10105), .A3(n9872), .ZN(n9871) );
  NAND3_X1 U12545 ( .A1(n10103), .A2(n10105), .A3(n15556), .ZN(n15555) );
  NOR2_X1 U12546 ( .A1(n13828), .A2(n13937), .ZN(n9883) );
  NAND2_X1 U12547 ( .A1(n9875), .A2(n9874), .ZN(n13788) );
  NAND3_X1 U12548 ( .A1(n10099), .A2(n13852), .A3(n13799), .ZN(n9881) );
  NAND3_X1 U12549 ( .A1(n9877), .A2(n9876), .A3(n9673), .ZN(n9875) );
  NOR2_X1 U12550 ( .A1(n13828), .A2(n9719), .ZN(n9876) );
  NAND2_X2 U12551 ( .A1(n13852), .A2(n10099), .ZN(n13848) );
  INV_X1 U12552 ( .A(n13852), .ZN(n9878) );
  XNOR2_X2 U12553 ( .A(n11193), .B(n11192), .ZN(n11257) );
  OAI21_X1 U12554 ( .B1(n13964), .B2(n19804), .A(n13785), .ZN(P1_U2969) );
  XNOR2_X1 U12555 ( .A(n9885), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13964) );
  NAND3_X1 U12556 ( .A1(n9887), .A2(n14876), .A3(n14874), .ZN(n9886) );
  NAND2_X1 U12557 ( .A1(n9889), .A2(n14878), .ZN(n9888) );
  NAND2_X1 U12558 ( .A1(n14599), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13417) );
  NAND3_X1 U12559 ( .A1(n9890), .A2(n13406), .A3(n12835), .ZN(n15825) );
  OAI21_X2 U12560 ( .B1(n12428), .B2(n12354), .A(n12430), .ZN(n9894) );
  NAND3_X1 U12561 ( .A1(n9960), .A2(n9958), .A3(n9672), .ZN(n9896) );
  NAND2_X1 U12562 ( .A1(n11488), .A2(n9897), .ZN(n13605) );
  INV_X1 U12563 ( .A(n13605), .ZN(n11553) );
  NAND2_X1 U12564 ( .A1(n9899), .A2(n12845), .ZN(n13006) );
  NAND3_X1 U12565 ( .A1(n12470), .A2(n19883), .A3(n11155), .ZN(n12444) );
  AND2_X1 U12566 ( .A1(n13680), .A2(n9902), .ZN(n13542) );
  NAND2_X1 U12567 ( .A1(n13680), .A2(n13582), .ZN(n13668) );
  NAND3_X1 U12568 ( .A1(n10323), .A2(n9904), .A3(n10275), .ZN(n9933) );
  NAND2_X1 U12569 ( .A1(n10825), .A2(n9904), .ZN(n14912) );
  NOR2_X1 U12570 ( .A1(n12558), .A2(n9907), .ZN(n12850) );
  NAND2_X1 U12571 ( .A1(n14252), .A2(n10077), .ZN(n10072) );
  INV_X1 U12572 ( .A(n14300), .ZN(n9914) );
  INV_X1 U12573 ( .A(n9919), .ZN(n15309) );
  NOR2_X1 U12574 ( .A1(n9919), .A2(n18430), .ZN(n15284) );
  XNOR2_X1 U12575 ( .A(n9919), .B(n18430), .ZN(n17479) );
  AND2_X1 U12576 ( .A1(n16993), .A2(n9919), .ZN(n9918) );
  NAND2_X1 U12577 ( .A1(n14600), .A2(n14601), .ZN(n13284) );
  NAND2_X1 U12578 ( .A1(n13253), .A2(n13252), .ZN(n14600) );
  INV_X1 U12579 ( .A(n9932), .ZN(n10354) );
  NAND2_X1 U12580 ( .A1(n10308), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10277) );
  NAND2_X2 U12581 ( .A1(n10126), .A2(n9695), .ZN(n10130) );
  NAND2_X2 U12582 ( .A1(n9935), .A2(n18830), .ZN(n10150) );
  NAND2_X1 U12583 ( .A1(n12866), .A2(n9702), .ZN(n13085) );
  INV_X1 U12584 ( .A(n14266), .ZN(n9942) );
  INV_X1 U12585 ( .A(n14279), .ZN(n9943) );
  NAND4_X1 U12586 ( .A1(n9951), .A2(n9950), .A3(n19823), .A4(n9952), .ZN(n9949) );
  NAND3_X1 U12587 ( .A1(n9951), .A2(n9952), .A3(n9950), .ZN(n13954) );
  NAND3_X1 U12588 ( .A1(n13779), .A2(n9957), .A3(n14121), .ZN(n9951) );
  INV_X1 U12589 ( .A(n9957), .ZN(n9953) );
  NAND2_X1 U12590 ( .A1(n13200), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9957) );
  NOR2_X1 U12591 ( .A1(n11161), .A2(n12443), .ZN(n9959) );
  NAND2_X1 U12592 ( .A1(n12444), .A2(n12456), .ZN(n9960) );
  OAI21_X2 U12593 ( .B1(n13882), .B2(n9962), .A(n10117), .ZN(n13852) );
  NAND2_X1 U12594 ( .A1(n13327), .A2(n9636), .ZN(n13357) );
  INV_X1 U12595 ( .A(n9972), .ZN(n13322) );
  AND2_X1 U12596 ( .A1(n13318), .A2(n9640), .ZN(n13370) );
  NAND2_X1 U12597 ( .A1(n13318), .A2(n9973), .ZN(n13371) );
  NAND2_X1 U12598 ( .A1(n13318), .A2(n9707), .ZN(n13363) );
  NAND2_X1 U12599 ( .A1(n13287), .A2(n9976), .ZN(n13301) );
  NAND2_X1 U12600 ( .A1(n13287), .A2(n13285), .ZN(n12973) );
  NAND2_X1 U12601 ( .A1(n18669), .A2(n18528), .ZN(n9986) );
  NAND2_X1 U12602 ( .A1(n15350), .A2(n18669), .ZN(n15708) );
  INV_X1 U12603 ( .A(n9986), .ZN(n9985) );
  AOI21_X1 U12604 ( .B1(n14219), .B2(n9999), .A(n18653), .ZN(n14190) );
  NAND2_X1 U12605 ( .A1(n9997), .A2(n9995), .ZN(n14189) );
  NAND2_X1 U12606 ( .A1(n14219), .A2(n9998), .ZN(n9997) );
  INV_X1 U12607 ( .A(n10000), .ZN(n14198) );
  INV_X1 U12608 ( .A(n17451), .ZN(n10019) );
  INV_X2 U12609 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18425) );
  INV_X2 U12610 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18436) );
  OAI21_X1 U12611 ( .B1(n17428), .B2(n10024), .A(n10022), .ZN(n10021) );
  NAND2_X1 U12612 ( .A1(n17428), .A2(n17429), .ZN(n17427) );
  OR2_X1 U12613 ( .A1(n17429), .A2(n10030), .ZN(n10029) );
  INV_X1 U12614 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U12615 ( .A1(n17388), .A2(n15344), .ZN(n10031) );
  NAND3_X1 U12616 ( .A1(n16006), .A2(n9625), .A3(n9674), .ZN(n10034) );
  AND2_X2 U12617 ( .A1(n11277), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11025) );
  INV_X1 U12618 ( .A(n11849), .ZN(n11144) );
  NAND2_X2 U12619 ( .A1(n12634), .A2(n19855), .ZN(n11843) );
  NAND3_X1 U12620 ( .A1(n11396), .A2(n10041), .A3(n11397), .ZN(n13180) );
  INV_X1 U12621 ( .A(n12663), .ZN(n10060) );
  NAND2_X1 U12622 ( .A1(n10060), .A2(n9627), .ZN(n10947) );
  NAND2_X1 U12623 ( .A1(n14777), .A2(n9712), .ZN(n14407) );
  INV_X1 U12624 ( .A(n15882), .ZN(n10066) );
  NAND2_X1 U12625 ( .A1(n14213), .A2(n10069), .ZN(n10071) );
  AND2_X1 U12626 ( .A1(n14213), .A2(n14202), .ZN(n14200) );
  INV_X1 U12627 ( .A(n10071), .ZN(n14164) );
  INV_X2 U12628 ( .A(n10861), .ZN(n10993) );
  NAND2_X1 U12629 ( .A1(n14252), .A2(n10074), .ZN(n10073) );
  NAND2_X1 U12630 ( .A1(n14252), .A2(n14251), .ZN(n14253) );
  OAI211_X1 U12631 ( .C1(n14252), .C2(n10076), .A(n10073), .B(n14344), .ZN(
        n12134) );
  NAND2_X1 U12632 ( .A1(n10342), .A2(n10341), .ZN(n10345) );
  NAND2_X1 U12633 ( .A1(n12394), .A2(n12395), .ZN(n10387) );
  NAND2_X1 U12634 ( .A1(n10342), .A2(n9696), .ZN(n10083) );
  INV_X1 U12635 ( .A(n10344), .ZN(n10084) );
  OAI21_X2 U12636 ( .B1(n14290), .B2(n10085), .A(n10086), .ZN(n10652) );
  NAND2_X1 U12637 ( .A1(n10095), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U12638 ( .A1(n19931), .A2(n10095), .ZN(n11275) );
  NOR2_X1 U12639 ( .A1(n19896), .A2(n10095), .ZN(n20384) );
  AND2_X1 U12640 ( .A1(n11196), .A2(n11194), .ZN(n11243) );
  NAND2_X1 U12641 ( .A1(n11169), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10096) );
  XNOR2_X2 U12642 ( .A(n10097), .B(n11165), .ZN(n19960) );
  INV_X1 U12643 ( .A(n13198), .ZN(n10099) );
  NAND2_X1 U12644 ( .A1(n11161), .A2(n10100), .ZN(n12374) );
  OAI21_X1 U12645 ( .B1(n13098), .B2(n10104), .A(n10102), .ZN(n15557) );
  AOI21_X1 U12646 ( .B1(n10108), .B2(n19790), .A(n10107), .ZN(n10102) );
  INV_X1 U12647 ( .A(n19790), .ZN(n10104) );
  NAND2_X1 U12648 ( .A1(n13098), .A2(n10106), .ZN(n10105) );
  NOR2_X1 U12649 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  INV_X1 U12650 ( .A(n13105), .ZN(n10107) );
  INV_X1 U12651 ( .A(n13097), .ZN(n10108) );
  NAND2_X1 U12652 ( .A1(n19791), .A2(n19790), .ZN(n19789) );
  NAND2_X1 U12653 ( .A1(n10333), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10304) );
  NAND2_X1 U12654 ( .A1(n10333), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10317) );
  NAND2_X1 U12655 ( .A1(n10333), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10326) );
  NAND2_X2 U12656 ( .A1(n10302), .A2(n10301), .ZN(n10333) );
  NAND2_X2 U12657 ( .A1(n10368), .A2(n10369), .ZN(n18830) );
  INV_X1 U12658 ( .A(n10122), .ZN(n14467) );
  NAND2_X1 U12659 ( .A1(n14551), .A2(n10123), .ZN(n14533) );
  CLKBUF_X1 U12660 ( .A(n10130), .Z(n10127) );
  INV_X1 U12661 ( .A(n9637), .ZN(n10131) );
  NOR2_X1 U12662 ( .A1(n14503), .A2(n14504), .ZN(n15768) );
  CLKBUF_X1 U12663 ( .A(n10139), .Z(n10135) );
  NAND2_X1 U12664 ( .A1(n10146), .A2(n10141), .ZN(n14454) );
  INV_X1 U12665 ( .A(n14493), .ZN(n10149) );
  NOR2_X1 U12666 ( .A1(n10150), .A2(n12733), .ZN(n13216) );
  NOR2_X2 U12667 ( .A1(n10150), .A2(n12726), .ZN(n19044) );
  NOR2_X2 U12668 ( .A1(n10150), .A2(n12721), .ZN(n19070) );
  NAND2_X1 U12669 ( .A1(n12617), .A2(n12616), .ZN(n12615) );
  NAND2_X1 U12670 ( .A1(n12562), .A2(n11287), .ZN(n12617) );
  NAND2_X1 U12671 ( .A1(n11553), .A2(n11552), .ZN(n13606) );
  CLKBUF_X1 U12672 ( .A(n14300), .Z(n14306) );
  NAND2_X1 U12673 ( .A1(n14305), .A2(n14307), .ZN(n14300) );
  INV_X1 U12674 ( .A(n13005), .ZN(n11396) );
  AND2_X2 U12675 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12484) );
  AND2_X1 U12676 ( .A1(n20107), .A2(n20105), .ZN(n19964) );
  NAND2_X1 U12677 ( .A1(n11097), .A2(n11096), .ZN(n11098) );
  INV_X1 U12678 ( .A(n13569), .ZN(n13667) );
  NAND2_X1 U12679 ( .A1(n11289), .A2(n11180), .ZN(n12631) );
  INV_X1 U12680 ( .A(n13028), .ZN(n10484) );
  INV_X2 U12681 ( .A(n12443), .ZN(n19855) );
  NAND2_X1 U12682 ( .A1(n13784), .A2(n11912), .ZN(n12020) );
  NAND2_X1 U12683 ( .A1(n10699), .A2(n10700), .ZN(n10701) );
  NAND2_X1 U12684 ( .A1(n14276), .A2(n14275), .ZN(n14274) );
  NAND2_X1 U12685 ( .A1(n10294), .A2(n18913), .ZN(n11012) );
  NAND2_X1 U12686 ( .A1(n12713), .A2(n12708), .ZN(n12753) );
  NOR2_X1 U12687 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11313) );
  AND2_X1 U12688 ( .A1(n10669), .A2(n10697), .ZN(n10151) );
  NAND2_X1 U12689 ( .A1(n19728), .A2(n19895), .ZN(n13698) );
  INV_X1 U12690 ( .A(n13696), .ZN(n11912) );
  AND2_X1 U12691 ( .A1(n10167), .A2(n15934), .ZN(n10153) );
  NAND2_X1 U12692 ( .A1(n10840), .A2(n10839), .ZN(n10154) );
  AND2_X1 U12693 ( .A1(n10162), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10155) );
  OR2_X1 U12694 ( .A1(n13445), .A2(n14894), .ZN(n10156) );
  INV_X1 U12695 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19636) );
  AND2_X1 U12696 ( .A1(n15803), .A2(n15802), .ZN(n10157) );
  AND3_X1 U12697 ( .A1(n11016), .A2(n11015), .A3(n11014), .ZN(n10158) );
  INV_X1 U12698 ( .A(n14875), .ZN(n13413) );
  AND2_X1 U12699 ( .A1(n12023), .A2(n12798), .ZN(n14350) );
  OR2_X1 U12700 ( .A1(n10472), .A2(n10471), .ZN(n10159) );
  OR2_X1 U12701 ( .A1(n19599), .A2(n19550), .ZN(n15908) );
  AND2_X1 U12702 ( .A1(n12133), .A2(n12132), .ZN(n10161) );
  INV_X1 U12703 ( .A(n13418), .ZN(n13412) );
  BUF_X4 U12704 ( .A(n11918), .Z(n13469) );
  AND2_X1 U12705 ( .A1(n11879), .A2(n11864), .ZN(n11885) );
  OR2_X1 U12706 ( .A1(n11879), .A2(n11878), .ZN(n11895) );
  INV_X1 U12707 ( .A(n11895), .ZN(n11897) );
  NAND2_X1 U12708 ( .A1(n11870), .A2(n12416), .ZN(n11096) );
  NAND2_X1 U12709 ( .A1(n11274), .A2(n11273), .ZN(n11225) );
  OR2_X1 U12710 ( .A1(n12125), .A2(n10330), .ZN(n10331) );
  AND2_X1 U12711 ( .A1(n20259), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11874) );
  OR2_X1 U12712 ( .A1(n11354), .A2(n11353), .ZN(n13125) );
  OR2_X1 U12714 ( .A1(n11373), .A2(n11372), .ZN(n13124) );
  NOR2_X1 U12715 ( .A1(n11142), .A2(n12889), .ZN(n11143) );
  NAND2_X1 U12716 ( .A1(n12429), .A2(n12443), .ZN(n11296) );
  OR2_X1 U12717 ( .A1(n14983), .A2(n14984), .ZN(n14978) );
  OR2_X1 U12718 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19848), .ZN(
        n11858) );
  NOR2_X1 U12719 ( .A1(n11190), .A2(n11189), .ZN(n12690) );
  NOR2_X1 U12720 ( .A1(n12469), .A2(n11260), .ZN(n11278) );
  XNOR2_X1 U12721 ( .A(n11253), .B(n11251), .ZN(n11266) );
  AND2_X1 U12722 ( .A1(n11898), .A2(n13133), .ZN(n11893) );
  NAND2_X1 U12723 ( .A1(n10777), .A2(n10792), .ZN(n10790) );
  AND2_X1 U12724 ( .A1(n18899), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13311) );
  AOI21_X1 U12725 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n14917), .A(n10324), 
        .ZN(n10325) );
  AND2_X1 U12726 ( .A1(n10670), .A2(n10151), .ZN(n10671) );
  AND2_X1 U12727 ( .A1(n11859), .A2(n11858), .ZN(n12270) );
  INV_X1 U12728 ( .A(n11724), .ZN(n11725) );
  INV_X1 U12729 ( .A(n12012), .ZN(n11998) );
  AND3_X1 U12730 ( .A1(n12377), .A2(n12507), .A3(n12376), .ZN(n12405) );
  OR2_X1 U12731 ( .A1(n11216), .A2(n11215), .ZN(n12505) );
  INV_X1 U12732 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14112) );
  NAND2_X1 U12733 ( .A1(n20110), .A2(n20401), .ZN(n11311) );
  NOR2_X1 U12734 ( .A1(n12815), .A2(n12939), .ZN(n10261) );
  NOR2_X1 U12735 ( .A1(n10263), .A2(n12779), .ZN(n10834) );
  NOR2_X1 U12736 ( .A1(n17864), .A2(n17001), .ZN(n15146) );
  INV_X1 U12737 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n20605) );
  NOR2_X1 U12738 ( .A1(n17864), .A2(n17843), .ZN(n15202) );
  AND2_X1 U12739 ( .A1(n16901), .A2(n15411), .ZN(n15152) );
  INV_X1 U12740 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20603) );
  INV_X1 U12741 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20624) );
  NAND2_X1 U12742 ( .A1(n13633), .A2(n11457), .ZN(n11488) );
  INV_X1 U12743 ( .A(n12640), .ZN(n14113) );
  OR2_X1 U12744 ( .A1(n12881), .A2(n13782), .ZN(n12882) );
  NAND2_X1 U12745 ( .A1(n11790), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12881) );
  NAND2_X1 U12746 ( .A1(n11649), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11682) );
  INV_X1 U12747 ( .A(n13608), .ZN(n11552) );
  INV_X1 U12748 ( .A(n11438), .ZN(n11514) );
  AND2_X1 U12749 ( .A1(n14030), .A2(n13938), .ZN(n13991) );
  INV_X1 U12750 ( .A(n15626), .ZN(n14073) );
  AND2_X1 U12751 ( .A1(n11142), .A2(n12889), .ZN(n13133) );
  INV_X1 U12752 ( .A(n20260), .ZN(n20337) );
  INV_X1 U12753 ( .A(n13082), .ZN(n10483) );
  INV_X1 U12754 ( .A(n12622), .ZN(n10416) );
  INV_X1 U12755 ( .A(n12344), .ZN(n10380) );
  NOR2_X1 U12756 ( .A1(n14616), .A2(n15898), .ZN(n14850) );
  AND4_X1 U12757 ( .A1(n17848), .A2(n17843), .A3(n15146), .A4(n15143), .ZN(
        n15150) );
  NOR2_X1 U12758 ( .A1(n18277), .A2(n14945), .ZN(n15186) );
  NOR2_X1 U12759 ( .A1(n18334), .A2(n17457), .ZN(n15985) );
  AND2_X1 U12760 ( .A1(n17277), .A2(n17599), .ZN(n17219) );
  NAND2_X1 U12761 ( .A1(n9600), .A2(n15201), .ZN(n18294) );
  NAND3_X1 U12762 ( .A1(n15030), .A2(n15029), .A3(n15028), .ZN(n15177) );
  OR2_X1 U12763 ( .A1(n18445), .A2(n18331), .ZN(n17830) );
  AND2_X1 U12764 ( .A1(n11627), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11628) );
  INV_X1 U12765 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13600) );
  INV_X1 U12766 ( .A(n19710), .ZN(n19686) );
  AND2_X1 U12767 ( .A1(n13208), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12899) );
  NOR2_X1 U12768 ( .A1(n12887), .A2(n19855), .ZN(n12898) );
  NAND2_X1 U12769 ( .A1(n19646), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12887) );
  AND2_X1 U12770 ( .A1(n12001), .A2(n12000), .ZN(n13547) );
  INV_X1 U12771 ( .A(n12428), .ZN(n13463) );
  XNOR2_X1 U12772 ( .A(n12882), .B(n13482), .ZN(n13208) );
  OR2_X1 U12773 ( .A1(n11682), .A2(n11681), .ZN(n11724) );
  AND2_X1 U12774 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n11588), .ZN(
        n11627) );
  INV_X1 U12775 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15466) );
  NOR2_X1 U12776 ( .A1(n11435), .A2(n19636), .ZN(n11440) );
  AND2_X1 U12777 ( .A1(n11387), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11411) );
  OR2_X1 U12778 ( .A1(n19795), .A2(n12406), .ZN(n13917) );
  AND3_X1 U12779 ( .A1(n13788), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n9615), .ZN(n13200) );
  OR2_X1 U12780 ( .A1(n14066), .A2(n13936), .ZN(n14037) );
  AND2_X1 U12781 ( .A1(n9615), .A2(n13196), .ZN(n13914) );
  AND2_X1 U12782 ( .A1(n14058), .A2(n13933), .ZN(n15626) );
  AND2_X1 U12783 ( .A1(n15626), .A2(n19812), .ZN(n15629) );
  NAND2_X1 U12784 ( .A1(n11176), .A2(n11175), .ZN(n11289) );
  OR2_X1 U12785 ( .A1(n20105), .A2(n19992), .ZN(n20081) );
  INV_X1 U12786 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20626) );
  NOR2_X1 U12787 ( .A1(n20000), .A2(n19999), .ZN(n20297) );
  INV_X1 U12788 ( .A(n20348), .ZN(n20346) );
  AND2_X1 U12789 ( .A1(n20400), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15384) );
  OR2_X1 U12790 ( .A1(n12786), .A2(n10824), .ZN(n15948) );
  AND2_X1 U12791 ( .A1(n12160), .A2(n10831), .ZN(n12790) );
  OR2_X1 U12792 ( .A1(n14639), .A2(n14340), .ZN(n12133) );
  AND3_X1 U12793 ( .A1(n10852), .A2(n10851), .A3(n10850), .ZN(n13020) );
  NAND2_X1 U12794 ( .A1(n12779), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12254) );
  AND2_X1 U12795 ( .A1(n14696), .A2(n14610), .ZN(n14675) );
  AND3_X1 U12796 ( .A1(n10855), .A2(n10854), .A3(n10853), .ZN(n12965) );
  NAND2_X1 U12797 ( .A1(n13413), .A2(n13412), .ZN(n13414) );
  INV_X1 U12798 ( .A(n18854), .ZN(n14609) );
  NAND2_X1 U12799 ( .A1(n12834), .A2(n12801), .ZN(n18832) );
  INV_X1 U12800 ( .A(n14940), .ZN(n14904) );
  AND2_X1 U12801 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19221) );
  OR2_X1 U12802 ( .A1(n19230), .A2(n19226), .ZN(n19257) );
  OR2_X1 U12803 ( .A1(n19305), .A2(n19300), .ZN(n19346) );
  OR2_X1 U12804 ( .A1(n19555), .A2(n19565), .ZN(n19296) );
  OR2_X1 U12805 ( .A1(n19566), .A2(n19162), .ZN(n18860) );
  NAND2_X1 U12806 ( .A1(n17063), .A2(n15151), .ZN(n16169) );
  NOR2_X1 U12807 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16370), .ZN(n16354) );
  NOR2_X1 U12808 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16486), .ZN(n16470) );
  INV_X1 U12809 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16487) );
  NAND2_X1 U12810 ( .A1(n17145), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17125) );
  INV_X1 U12811 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17308) );
  INV_X1 U12812 ( .A(n17689), .ZN(n17356) );
  INV_X1 U12813 ( .A(n15985), .ZN(n17267) );
  NOR3_X1 U12814 ( .A1(n17175), .A2(n17182), .A3(n17537), .ZN(n15343) );
  NOR2_X1 U12815 ( .A1(n17173), .A2(n17631), .ZN(n17536) );
  AOI21_X2 U12816 ( .B1(n18279), .B2(n9600), .A(n18278), .ZN(n18270) );
  INV_X1 U12817 ( .A(n18270), .ZN(n18282) );
  NAND2_X1 U12818 ( .A1(n11628), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11650) );
  AND2_X1 U12819 ( .A1(n19646), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19710) );
  AND2_X1 U12820 ( .A1(n19646), .A2(n12883), .ZN(n19667) );
  AND2_X1 U12821 ( .A1(n19646), .A2(n12899), .ZN(n19641) );
  INV_X1 U12822 ( .A(n13698), .ZN(n19725) );
  NAND2_X1 U12823 ( .A1(n12381), .A2(n12461), .ZN(n11911) );
  INV_X1 U12824 ( .A(n12474), .ZN(n19773) );
  NAND2_X1 U12825 ( .A1(n11441), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11471) );
  NAND2_X1 U12826 ( .A1(n11338), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11357) );
  INV_X1 U12827 ( .A(n13917), .ZN(n19799) );
  AND2_X1 U12828 ( .A1(n20348), .A2(n12397), .ZN(n19794) );
  NOR2_X1 U12829 ( .A1(n14037), .A2(n9990), .ZN(n14030) );
  NOR2_X1 U12830 ( .A1(n13931), .A2(n15597), .ZN(n15628) );
  INV_X1 U12831 ( .A(n19812), .ZN(n19831) );
  INV_X1 U12832 ( .A(n19858), .ZN(n19999) );
  INV_X1 U12833 ( .A(n20398), .ZN(n19898) );
  INV_X1 U12834 ( .A(n19991), .ZN(n19980) );
  AND2_X1 U12835 ( .A1(n19964), .A2(n20075), .ZN(n20018) );
  INV_X1 U12836 ( .A(n20066), .ZN(n20070) );
  INV_X1 U12837 ( .A(n20104), .ZN(n20095) );
  INV_X1 U12838 ( .A(n20098), .ZN(n20133) );
  INV_X1 U12839 ( .A(n20225), .ZN(n20108) );
  OAI22_X1 U12840 ( .A1(n20172), .A2(n20171), .B1(n20170), .B2(n20288), .ZN(
        n20189) );
  INV_X1 U12841 ( .A(n20218), .ZN(n20221) );
  OR2_X1 U12842 ( .A1(n20107), .A2(n20106), .ZN(n20202) );
  OAI211_X1 U12843 ( .C1(n20328), .C2(n20298), .A(n20297), .B(n20296), .ZN(
        n20330) );
  INV_X1 U12844 ( .A(n20462), .ZN(n20465) );
  INV_X1 U12845 ( .A(n20459), .ZN(n20466) );
  INV_X1 U12846 ( .A(n18679), .ZN(n18563) );
  INV_X1 U12847 ( .A(n18681), .ZN(n18667) );
  OR2_X1 U12848 ( .A1(n10450), .A2(n10449), .ZN(n12986) );
  OR2_X1 U12849 ( .A1(n10403), .A2(n10402), .ZN(n12559) );
  NOR2_X1 U12850 ( .A1(n10389), .A2(n10388), .ZN(n12672) );
  AND2_X1 U12851 ( .A1(n14333), .A2(n18913), .ZN(n14344) );
  INV_X1 U12852 ( .A(n19458), .ZN(n12798) );
  INV_X1 U12853 ( .A(n12289), .ZN(n12324) );
  AND2_X1 U12854 ( .A1(n10314), .A2(n12928), .ZN(n12173) );
  AND2_X1 U12855 ( .A1(n15833), .A2(n12234), .ZN(n15824) );
  AND2_X1 U12856 ( .A1(n12834), .A2(n12804), .ZN(n18853) );
  AND2_X1 U12857 ( .A1(n12834), .A2(n19582), .ZN(n18844) );
  AOI21_X2 U12858 ( .B1(n15408), .B2(n15407), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19405) );
  OR2_X1 U12859 ( .A1(n15943), .A2(n19571), .ZN(n15408) );
  INV_X1 U12860 ( .A(n18906), .ZN(n18944) );
  INV_X1 U12861 ( .A(n18956), .ZN(n18973) );
  INV_X1 U12862 ( .A(n19235), .ZN(n19229) );
  AND2_X1 U12863 ( .A1(n19098), .A2(n19229), .ZN(n19035) );
  INV_X1 U12864 ( .A(n19056), .ZN(n19063) );
  AND2_X1 U12865 ( .A1(n19160), .A2(n19573), .ZN(n19068) );
  INV_X1 U12866 ( .A(n19157), .ZN(n19149) );
  AND2_X1 U12867 ( .A1(n19555), .A2(n19563), .ZN(n19158) );
  NOR2_X1 U12868 ( .A1(n19353), .A2(n19235), .ZN(n19215) );
  INV_X1 U12869 ( .A(n19420), .ZN(n19319) );
  INV_X1 U12870 ( .A(n19432), .ZN(n19378) );
  NOR2_X1 U12871 ( .A1(n19297), .A2(n19296), .ZN(n19392) );
  AND2_X1 U12872 ( .A1(n18888), .A2(n18912), .ZN(n19421) );
  OR2_X1 U12873 ( .A1(n19575), .A2(n12168), .ZN(n15961) );
  INV_X1 U12874 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19485) );
  INV_X1 U12875 ( .A(n18488), .ZN(n16488) );
  NOR2_X2 U12876 ( .A1(n18487), .A2(n15200), .ZN(n18266) );
  NOR2_X1 U12877 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16283), .ZN(n16268) );
  NOR2_X1 U12878 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16303), .ZN(n16292) );
  NOR2_X1 U12879 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16320), .ZN(n16311) );
  NOR2_X1 U12880 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16392), .ZN(n16374) );
  INV_X1 U12881 ( .A(n16530), .ZN(n16510) );
  NOR2_X1 U12882 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16456), .ZN(n16445) );
  NOR4_X1 U12883 ( .A1(n17831), .A2(n16173), .A3(n18316), .A4(n16488), .ZN(
        n16276) );
  NOR3_X2 U12884 ( .A1(n17831), .A2(n16488), .A3(n16172), .ZN(n16530) );
  NOR2_X1 U12885 ( .A1(n16637), .A2(n16641), .ZN(n16610) );
  NAND2_X1 U12886 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16746), .ZN(n16705) );
  NAND2_X1 U12887 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16816), .ZN(n16774) );
  NAND2_X1 U12888 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n16886), .ZN(n16885) );
  INV_X1 U12889 ( .A(n15176), .ZN(n17853) );
  INV_X1 U12890 ( .A(n16925), .ZN(n16921) );
  NAND4_X1 U12891 ( .A1(n16968), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n16854), .ZN(n16944) );
  NOR2_X1 U12892 ( .A1(n16995), .A2(n16941), .ZN(n16968) );
  INV_X1 U12893 ( .A(n17831), .ZN(n17001) );
  NOR2_X1 U12894 ( .A1(n17107), .A2(n17834), .ZN(n17108) );
  INV_X1 U12895 ( .A(n17346), .ZN(n17285) );
  OAI22_X1 U12896 ( .A1(n17492), .A2(n17691), .B1(n17117), .B2(n17356), .ZN(
        n17383) );
  INV_X1 U12897 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17422) );
  NOR2_X1 U12898 ( .A1(n18018), .A2(n18168), .ZN(n15986) );
  INV_X1 U12899 ( .A(n17722), .ZN(n17619) );
  NOR2_X1 U12900 ( .A1(n17677), .A2(n17804), .ZN(n17710) );
  INV_X1 U12901 ( .A(n17805), .ZN(n17761) );
  INV_X1 U12902 ( .A(n17802), .ZN(n17809) );
  NOR2_X1 U12903 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18419), .ZN(
        n18445) );
  INV_X1 U12904 ( .A(n17924), .ZN(n17928) );
  INV_X1 U12905 ( .A(n20663), .ZN(n18013) );
  INV_X1 U12906 ( .A(n18034), .ZN(n18038) );
  INV_X1 U12907 ( .A(n18153), .ZN(n18161) );
  AND2_X1 U12908 ( .A1(n18171), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18210) );
  AND2_X1 U12909 ( .A1(n18482), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18355) );
  NOR2_X1 U12910 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12149), .ZN(n16130)
         );
  INV_X1 U12911 ( .A(n20487), .ZN(n20502) );
  NAND2_X1 U12912 ( .A1(n20419), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20485) );
  INV_X1 U12913 ( .A(n19707), .ZN(n19673) );
  INV_X1 U12914 ( .A(n19698), .ZN(n19714) );
  INV_X1 U12915 ( .A(n13784), .ZN(n13707) );
  INV_X1 U12916 ( .A(n19732), .ZN(n19761) );
  NOR2_X1 U12917 ( .A1(n12371), .A2(n12370), .ZN(n12575) );
  INV_X1 U12918 ( .A(n19795), .ZN(n19804) );
  INV_X1 U12919 ( .A(n19794), .ZN(n19851) );
  NOR2_X1 U12920 ( .A1(n19831), .A2(n15628), .ZN(n15606) );
  OR2_X1 U12921 ( .A1(n12450), .A2(n12432), .ZN(n19834) );
  OAI21_X1 U12922 ( .B1(n12652), .B2(n12651), .A(n19999), .ZN(n19847) );
  NAND2_X1 U12923 ( .A1(n19964), .A2(n20108), .ZN(n19930) );
  NAND2_X1 U12924 ( .A1(n19964), .A2(n20257), .ZN(n19959) );
  NAND2_X1 U12925 ( .A1(n19964), .A2(n20162), .ZN(n19991) );
  NAND2_X1 U12926 ( .A1(n20076), .A2(n20108), .ZN(n20045) );
  NAND2_X1 U12927 ( .A1(n20076), .A2(n20257), .ZN(n20066) );
  NAND2_X1 U12928 ( .A1(n20076), .A2(n20075), .ZN(n20098) );
  NAND2_X1 U12929 ( .A1(n20076), .A2(n20162), .ZN(n20104) );
  NAND2_X1 U12930 ( .A1(n20109), .A2(n20108), .ZN(n20161) );
  OR2_X1 U12931 ( .A1(n20202), .A2(n20141), .ZN(n20193) );
  OR2_X1 U12932 ( .A1(n20202), .A2(n20289), .ZN(n20218) );
  OR2_X1 U12933 ( .A1(n20202), .A2(n20201), .ZN(n20256) );
  NAND2_X1 U12934 ( .A1(n20258), .A2(n20257), .ZN(n20333) );
  NAND2_X1 U12935 ( .A1(n20258), .A2(n20075), .ZN(n20398) );
  INV_X1 U12936 ( .A(n20475), .ZN(n20405) );
  INV_X1 U12937 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20419) );
  INV_X1 U12938 ( .A(n20485), .ZN(n20487) );
  OR2_X1 U12939 ( .A1(n20422), .A2(n20502), .ZN(n20459) );
  AND2_X1 U12940 ( .A1(n15945), .A2(n12928), .ZN(n19600) );
  NAND2_X1 U12941 ( .A1(n12793), .A2(n12172), .ZN(n12214) );
  NAND2_X1 U12942 ( .A1(n19600), .A2(n12926), .ZN(n18656) );
  INV_X1 U12943 ( .A(n18639), .ZN(n18687) );
  INV_X1 U12944 ( .A(n15763), .ZN(n15864) );
  INV_X1 U12945 ( .A(n14340), .ZN(n14333) );
  XNOR2_X1 U12946 ( .A(n12395), .B(n12394), .ZN(n19160) );
  NOR2_X1 U12947 ( .A1(n18761), .A2(n18757), .ZN(n18739) );
  AND2_X1 U12948 ( .A1(n10838), .A2(n12798), .ZN(n18755) );
  NAND2_X1 U12949 ( .A1(n18766), .A2(n12255), .ZN(n12341) );
  INV_X1 U12950 ( .A(n18766), .ZN(n18799) );
  NAND2_X1 U12951 ( .A1(n12173), .A2(n13275), .ZN(n12935) );
  NAND2_X1 U12952 ( .A1(n12209), .A2(n19592), .ZN(n15817) );
  INV_X1 U12953 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18602) );
  OR2_X1 U12954 ( .A1(n14628), .A2(n18841), .ZN(n14629) );
  INV_X1 U12955 ( .A(n18846), .ZN(n18841) );
  INV_X1 U12956 ( .A(n18844), .ZN(n15926) );
  INV_X1 U12957 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U12958 ( .A1(n19158), .A2(n19098), .ZN(n18956) );
  NAND2_X1 U12959 ( .A1(n19068), .A2(n19229), .ZN(n19007) );
  NAND2_X1 U12960 ( .A1(n19068), .A2(n19304), .ZN(n19056) );
  INV_X1 U12961 ( .A(n19094), .ZN(n19089) );
  NAND2_X1 U12962 ( .A1(n19544), .A2(n19068), .ZN(n19126) );
  NAND2_X1 U12963 ( .A1(n19098), .A2(n19544), .ZN(n19157) );
  NAND2_X1 U12964 ( .A1(n19128), .A2(n19158), .ZN(n19183) );
  INV_X1 U12965 ( .A(n19210), .ZN(n19219) );
  INV_X1 U12966 ( .A(n19215), .ZN(n19262) );
  AOI21_X1 U12967 ( .B1(n19269), .B2(n19270), .A(n19268), .ZN(n19295) );
  INV_X1 U12968 ( .A(n19392), .ZN(n19389) );
  INV_X1 U12969 ( .A(n19452), .ZN(n19439) );
  NAND2_X1 U12970 ( .A1(n19544), .A2(n18870), .ZN(n19456) );
  INV_X1 U12971 ( .A(n19542), .ZN(n19467) );
  NAND2_X1 U12972 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18347), .ZN(n18483) );
  NAND2_X1 U12973 ( .A1(n18470), .A2(n18268), .ZN(n16152) );
  INV_X1 U12974 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17226) );
  INV_X1 U12975 ( .A(n16533), .ZN(n16450) );
  NAND2_X1 U12976 ( .A1(n16901), .A2(n16841), .ZN(n16834) );
  NOR2_X1 U12977 ( .A1(n16942), .A2(n16967), .ZN(n16961) );
  NOR2_X1 U12978 ( .A1(n15231), .A2(n15230), .ZN(n16977) );
  INV_X1 U12979 ( .A(n16993), .ZN(n16989) );
  INV_X1 U12980 ( .A(n17028), .ZN(n17059) );
  INV_X1 U12981 ( .A(n17108), .ZN(n17103) );
  NAND2_X1 U12982 ( .A1(n17383), .A2(n17594), .ZN(n17292) );
  NAND2_X1 U12983 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17485), .ZN(n17346) );
  INV_X1 U12984 ( .A(n17342), .ZN(n17402) );
  INV_X1 U12985 ( .A(n17480), .ZN(n17471) );
  INV_X1 U12986 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17484) );
  NAND2_X1 U12987 ( .A1(n17811), .A2(n17644), .ZN(n17727) );
  NAND2_X1 U12988 ( .A1(n17712), .A2(n17804), .ZN(n17805) );
  INV_X1 U12989 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18091) );
  INV_X1 U12990 ( .A(n18137), .ZN(n18135) );
  INV_X1 U12991 ( .A(n18250), .ZN(n18200) );
  INV_X1 U12992 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18475) );
  INV_X1 U12993 ( .A(n18416), .ZN(n18335) );
  INV_X1 U12994 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18347) );
  INV_X1 U12995 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20544) );
  NAND2_X1 U12996 ( .A1(n12020), .A2(n12019), .ZN(P1_U2842) );
  NOR2_X4 U12997 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14902) );
  AND2_X4 U12998 ( .A1(n10776), .A2(n14902), .ZN(n10391) );
  AOI22_X1 U12999 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10391), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10162) );
  AND2_X2 U13000 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14911) );
  AND2_X4 U13001 ( .A1(n14911), .A2(n13033), .ZN(n10253) );
  AND3_X4 U13002 ( .A1(n10773), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13003 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10190), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10166) );
  NOR2_X2 U13004 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10163) );
  AND2_X4 U13005 ( .A1(n10163), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10754) );
  AND2_X4 U13006 ( .A1(n14922), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10753) );
  AOI22_X1 U13007 ( .A1(n10754), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10165) );
  AND2_X2 U13008 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14914) );
  AND2_X4 U13009 ( .A1(n14914), .A2(n10776), .ZN(n10239) );
  AOI22_X1 U13010 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10164) );
  NAND4_X1 U13011 ( .A1(n10155), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10172) );
  AOI22_X1 U13012 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13013 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13014 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13015 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10168) );
  NAND4_X1 U13016 ( .A1(n10153), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10171) );
  NAND2_X2 U13017 ( .A1(n10172), .A2(n10171), .ZN(n18892) );
  AOI22_X1 U13018 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13019 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13020 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13021 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U13022 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U13023 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13024 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13025 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10178) );
  AND4_X2 U13026 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        n10182) );
  NAND2_X2 U13027 ( .A1(n10184), .A2(n10183), .ZN(n10278) );
  AOI22_X1 U13028 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13029 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13030 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13031 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10185) );
  NAND4_X1 U13032 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10189) );
  NAND2_X1 U13033 ( .A1(n10189), .A2(n15934), .ZN(n10197) );
  AOI22_X1 U13034 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13035 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U13036 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10192) );
  NAND4_X1 U13037 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10195) );
  NAND2_X1 U13038 ( .A1(n10195), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10196) );
  NAND2_X2 U13039 ( .A1(n10197), .A2(n10196), .ZN(n18903) );
  AOI22_X1 U13040 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13041 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U13042 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U13043 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10198) );
  NAND4_X1 U13044 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n10202) );
  AOI22_X1 U13045 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13046 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U13047 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10190), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10203) );
  NAND4_X1 U13048 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10207) );
  AOI22_X1 U13049 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13050 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13051 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U13052 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10210) );
  NAND4_X1 U13053 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10219) );
  AOI22_X1 U13054 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U13055 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U13056 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10214) );
  NAND4_X1 U13057 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        n10218) );
  MUX2_X2 U13058 ( .A(n10219), .B(n10218), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n18888) );
  AOI22_X1 U13059 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13060 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U13061 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U13062 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10220) );
  AND4_X1 U13063 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10233) );
  AOI22_X1 U13064 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13065 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U13066 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10229) );
  NAND3_X1 U13067 ( .A1(n10229), .A2(n10228), .A3(n10227), .ZN(n10230) );
  NOR2_X1 U13068 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  MUX2_X2 U13069 ( .A(n10233), .B(n10232), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n18884) );
  AOI22_X1 U13070 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13071 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13072 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13073 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U13074 ( .A1(n10238), .A2(n15934), .ZN(n10246) );
  AOI22_X1 U13075 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10240) );
  AND2_X1 U13076 ( .A1(n10240), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10244) );
  AOI22_X1 U13077 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13078 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13079 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10241) );
  NAND4_X1 U13080 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10245) );
  AOI22_X1 U13081 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U13082 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U13083 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13084 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10248) );
  NAND4_X1 U13085 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10252) );
  AOI22_X1 U13086 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13087 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10253), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13088 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13089 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10254) );
  NAND4_X1 U13090 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10258) );
  NAND2_X1 U13091 ( .A1(n10258), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10259) );
  INV_X1 U13092 ( .A(n18892), .ZN(n12778) );
  NAND2_X1 U13093 ( .A1(n12778), .A2(n18913), .ZN(n10285) );
  INV_X1 U13094 ( .A(n10285), .ZN(n10262) );
  NAND2_X1 U13095 ( .A1(n10832), .A2(n10262), .ZN(n10269) );
  INV_X1 U13096 ( .A(n10278), .ZN(n10263) );
  NAND2_X1 U13097 ( .A1(n10840), .A2(n10266), .ZN(n10264) );
  NAND2_X1 U13098 ( .A1(n10264), .A2(n9594), .ZN(n10267) );
  INV_X1 U13099 ( .A(n10278), .ZN(n10265) );
  NAND2_X1 U13100 ( .A1(n12021), .A2(n10819), .ZN(n10323) );
  NOR2_X1 U13101 ( .A1(n10294), .A2(n18888), .ZN(n10270) );
  AND2_X2 U13102 ( .A1(n18913), .A2(n18903), .ZN(n10293) );
  NAND4_X1 U13103 ( .A1(n10270), .A2(n10293), .A3(n12777), .A4(n18892), .ZN(
        n10289) );
  INV_X1 U13104 ( .A(n10289), .ZN(n10272) );
  NAND2_X1 U13105 ( .A1(n10272), .A2(n18868), .ZN(n10814) );
  NAND4_X1 U13106 ( .A1(n12788), .A2(n9594), .A3(n10293), .A4(n10834), .ZN(
        n10273) );
  NOR2_X2 U13107 ( .A1(n11012), .A2(n18903), .ZN(n10274) );
  NAND2_X1 U13108 ( .A1(n10314), .A2(n10298), .ZN(n10275) );
  AND2_X4 U13109 ( .A1(n10314), .A2(n10697), .ZN(n12025) );
  AOI22_X1 U13110 ( .A1(n12025), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10276) );
  OAI211_X1 U13111 ( .C1(n12125), .C2(n12996), .A(n10277), .B(n10276), .ZN(
        n10306) );
  XNOR2_X1 U13112 ( .A(n10278), .B(n18903), .ZN(n10821) );
  NAND2_X1 U13113 ( .A1(n12807), .A2(n18888), .ZN(n10280) );
  NAND2_X1 U13114 ( .A1(n10280), .A2(n10279), .ZN(n10836) );
  NAND2_X1 U13115 ( .A1(n10281), .A2(n10298), .ZN(n12805) );
  AND2_X1 U13116 ( .A1(n18903), .A2(n10263), .ZN(n10286) );
  INV_X1 U13117 ( .A(n10283), .ZN(n10284) );
  NAND3_X1 U13118 ( .A1(n10288), .A2(n10287), .A3(n18884), .ZN(n10290) );
  NAND3_X1 U13119 ( .A1(n10290), .A2(n18868), .A3(n10289), .ZN(n12812) );
  NAND2_X1 U13120 ( .A1(n10291), .A2(n12812), .ZN(n10292) );
  NAND2_X1 U13121 ( .A1(n10292), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10302) );
  INV_X1 U13122 ( .A(n10293), .ZN(n10295) );
  NOR2_X1 U13123 ( .A1(n10298), .A2(n12777), .ZN(n10299) );
  NAND2_X1 U13124 ( .A1(n15941), .A2(n10299), .ZN(n10300) );
  NAND2_X1 U13125 ( .A1(n10300), .A2(n12787), .ZN(n12022) );
  AOI21_X1 U13126 ( .B1(n15967), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U13127 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  OR2_X2 U13128 ( .A1(n10306), .A2(n10305), .ZN(n10328) );
  NAND2_X1 U13129 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  NAND2_X1 U13130 ( .A1(n10308), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10313) );
  INV_X1 U13131 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13132 ( .A1(n12025), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10309) );
  INV_X1 U13133 ( .A(n10311), .ZN(n10312) );
  INV_X1 U13134 ( .A(n10314), .ZN(n10825) );
  NAND2_X1 U13135 ( .A1(n15967), .A2(n20564), .ZN(n19599) );
  NOR2_X1 U13136 ( .A1(n19599), .A2(n19570), .ZN(n10315) );
  INV_X1 U13138 ( .A(n10347), .ZN(n10318) );
  INV_X1 U13139 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U13140 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12210) );
  NAND2_X1 U13141 ( .A1(n19599), .A2(n12210), .ZN(n10319) );
  AOI21_X1 U13142 ( .B1(n12025), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10319), .ZN(
        n10321) );
  INV_X1 U13143 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12203) );
  OAI211_X1 U13144 ( .C1(n10329), .C2(n12207), .A(n10321), .B(n10320), .ZN(
        n10322) );
  OAI21_X1 U13145 ( .B1(n19599), .B2(n19578), .A(n9603), .ZN(n10324) );
  NAND2_X1 U13146 ( .A1(n10347), .A2(n10346), .ZN(n10363) );
  INV_X1 U13147 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14614) );
  AOI22_X1 U13148 ( .A1(n12025), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10332) );
  INV_X1 U13149 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U13150 ( .A1(n10333), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10335) );
  OR2_X1 U13151 ( .A1(n19599), .A2(n19554), .ZN(n10334) );
  NAND2_X1 U13152 ( .A1(n10335), .A2(n10334), .ZN(n10336) );
  NAND2_X1 U13153 ( .A1(n10337), .A2(n10336), .ZN(n10338) );
  NAND2_X1 U13154 ( .A1(n12728), .A2(n10370), .ZN(n10342) );
  NAND2_X1 U13155 ( .A1(n18903), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U13156 ( .A1(n10339), .A2(n19571), .ZN(n10375) );
  NAND2_X1 U13157 ( .A1(n19221), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10373) );
  AOI21_X1 U13158 ( .B1(n10373), .B2(n19554), .A(n19550), .ZN(n10340) );
  INV_X1 U13159 ( .A(n19448), .ZN(n18863) );
  AOI22_X1 U13160 ( .A1(n10375), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n10340), .B2(n18863), .ZN(n10341) );
  INV_X1 U13161 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U13162 ( .A1(n10389), .A2(n10343), .ZN(n10344) );
  NAND2_X1 U13163 ( .A1(n10345), .A2(n10344), .ZN(n10385) );
  INV_X1 U13164 ( .A(n10346), .ZN(n10348) );
  XNOR2_X2 U13165 ( .A(n10348), .B(n10347), .ZN(n12706) );
  XNOR2_X2 U13166 ( .A(n12706), .B(n10357), .ZN(n12719) );
  NAND2_X1 U13167 ( .A1(n10375), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10351) );
  NAND2_X1 U13168 ( .A1(n19578), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10350) );
  NAND2_X1 U13169 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19570), .ZN(
        n19159) );
  NAND2_X1 U13170 ( .A1(n10350), .A2(n19159), .ZN(n19008) );
  NAND2_X1 U13171 ( .A1(n19008), .A2(n19355), .ZN(n19192) );
  NAND2_X1 U13172 ( .A1(n10351), .A2(n19192), .ZN(n10352) );
  INV_X1 U13173 ( .A(n10353), .ZN(n10355) );
  NAND2_X1 U13174 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  INV_X1 U13175 ( .A(n10370), .ZN(n12233) );
  NOR2_X1 U13176 ( .A1(n19550), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10358) );
  AOI21_X1 U13177 ( .B1(n10375), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10358), .ZN(n10359) );
  NAND2_X1 U13178 ( .A1(n10697), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10361) );
  XNOR2_X1 U13179 ( .A(n10360), .B(n10361), .ZN(n12349) );
  NAND2_X1 U13180 ( .A1(n13037), .A2(n10361), .ZN(n10362) );
  NAND2_X1 U13181 ( .A1(n12350), .A2(n10362), .ZN(n12344) );
  NAND2_X1 U13182 ( .A1(n10364), .A2(n10363), .ZN(n10367) );
  INV_X1 U13183 ( .A(n10365), .ZN(n10366) );
  NAND2_X1 U13184 ( .A1(n10367), .A2(n10366), .ZN(n10368) );
  INV_X1 U13185 ( .A(n19221), .ZN(n10371) );
  NAND2_X1 U13186 ( .A1(n10371), .A2(n19560), .ZN(n10372) );
  NAND2_X1 U13187 ( .A1(n10373), .A2(n10372), .ZN(n19009) );
  NOR2_X1 U13188 ( .A1(n19009), .A2(n19550), .ZN(n10374) );
  AOI21_X1 U13189 ( .B1(n10375), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10374), .ZN(n10376) );
  NAND2_X1 U13190 ( .A1(n10377), .A2(n10376), .ZN(n10382) );
  INV_X1 U13191 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10378) );
  XNOR2_X1 U13192 ( .A(n10382), .B(n10381), .ZN(n12345) );
  NAND2_X1 U13193 ( .A1(n10382), .A2(n10381), .ZN(n10383) );
  NAND2_X1 U13194 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18903), .ZN(
        n10384) );
  INV_X1 U13195 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10388) );
  INV_X1 U13196 ( .A(n9607), .ZN(n10577) );
  AND2_X2 U13197 ( .A1(n9608), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10950) );
  AOI22_X1 U13198 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10396) );
  AND2_X2 U13199 ( .A1(n10391), .A2(n15934), .ZN(n10417) );
  AND2_X2 U13200 ( .A1(n10752), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10865) );
  AOI22_X1 U13201 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10395) );
  AND2_X2 U13202 ( .A1(n10391), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10418) );
  AND2_X2 U13203 ( .A1(n10641), .A2(n15934), .ZN(n10951) );
  AOI22_X1 U13204 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10394) );
  AND2_X2 U13205 ( .A1(n10641), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10429) );
  INV_X1 U13206 ( .A(n10392), .ZN(n10578) );
  AND2_X2 U13207 ( .A1(n9604), .A2(n15934), .ZN(n10405) );
  AOI22_X1 U13208 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10393) );
  NAND4_X1 U13209 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10403) );
  AOI22_X1 U13210 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10401) );
  AND2_X2 U13211 ( .A1(n10190), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10870) );
  AOI22_X1 U13213 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10400) );
  AND2_X2 U13214 ( .A1(n10752), .A2(n15934), .ZN(n10510) );
  AOI22_X1 U13215 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10399) );
  AND2_X2 U13216 ( .A1(n10190), .A2(n15934), .ZN(n10522) );
  NAND3_X1 U13217 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12164) );
  INV_X1 U13218 ( .A(n12164), .ZN(n10397) );
  NAND2_X1 U13219 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10397), .ZN(
        n10524) );
  AOI22_X1 U13220 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10398) );
  NAND4_X1 U13221 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10402) );
  AOI22_X1 U13222 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13223 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13224 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13225 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10406) );
  NAND4_X1 U13226 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10415) );
  AOI22_X1 U13227 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13228 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13229 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13230 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10957), .ZN(n10410) );
  NAND4_X1 U13231 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10414) );
  NOR2_X1 U13232 ( .A1(n10415), .A2(n10414), .ZN(n12622) );
  AOI22_X1 U13233 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U13234 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13235 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U13236 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10419) );
  NAND4_X1 U13237 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10428) );
  AOI22_X1 U13238 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10499), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13239 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13240 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10522), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U13241 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n10957), .ZN(n10423) );
  NAND4_X1 U13242 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n10427) );
  AOI22_X1 U13243 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13244 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13245 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13246 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10430) );
  NAND4_X1 U13247 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10439) );
  AOI22_X1 U13248 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13249 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13250 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13251 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n10957), .ZN(n10434) );
  NAND4_X1 U13252 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10438) );
  AOI22_X1 U13253 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13254 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13255 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13256 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10440) );
  NAND4_X1 U13257 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10450) );
  AOI22_X1 U13258 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13259 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13260 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13261 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n10957), .ZN(n10445) );
  NAND4_X1 U13262 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10449) );
  AOI22_X1 U13263 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U13264 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13265 ( .A1(n10951), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13266 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10451) );
  NAND4_X1 U13267 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10461) );
  AOI22_X1 U13268 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13269 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13270 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13271 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10456) );
  NAND4_X1 U13272 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10460) );
  AOI22_X1 U13273 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13274 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13275 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13276 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10463) );
  NAND4_X1 U13277 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10472) );
  AOI22_X1 U13278 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10870), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13279 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10510), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13280 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10499), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13281 ( .A1(n10546), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n10957), .ZN(n10467) );
  NAND4_X1 U13282 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10471) );
  AOI22_X1 U13283 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13284 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13285 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13286 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10429), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10473) );
  NAND4_X1 U13287 ( .A1(n10476), .A2(n10475), .A3(n10474), .A4(n10473), .ZN(
        n10482) );
  AOI22_X1 U13288 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13289 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13290 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13291 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n10957), .ZN(n10477) );
  NAND4_X1 U13292 ( .A1(n10480), .A2(n10479), .A3(n10478), .A4(n10477), .ZN(
        n10481) );
  NOR2_X1 U13293 ( .A1(n10482), .A2(n10481), .ZN(n13082) );
  AOI22_X1 U13294 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13295 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13296 ( .A1(n10951), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13297 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13298 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10494) );
  AOI22_X1 U13299 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13300 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13301 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13302 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10489) );
  NAND4_X1 U13303 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10493) );
  NOR2_X1 U13304 ( .A1(n10494), .A2(n10493), .ZN(n14343) );
  AOI22_X1 U13305 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13306 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13307 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13308 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10495) );
  NAND4_X1 U13309 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10505) );
  AOI22_X1 U13310 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13311 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13312 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13313 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n10957), .ZN(n10500) );
  NAND4_X1 U13314 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  AOI22_X1 U13315 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13316 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13317 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13318 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10506) );
  NAND4_X1 U13319 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10516) );
  AOI22_X1 U13320 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13321 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13322 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13323 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n10957), .ZN(n10511) );
  NAND4_X1 U13324 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10515) );
  NOR2_X1 U13325 ( .A1(n10516), .A2(n10515), .ZN(n14326) );
  INV_X1 U13326 ( .A(n14326), .ZN(n10517) );
  AOI22_X1 U13327 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13329 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13330 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13331 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10531) );
  AOI22_X1 U13332 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13333 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13334 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10527) );
  INV_X1 U13335 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10523) );
  NOR2_X1 U13336 ( .A1(n10524), .A2(n10523), .ZN(n10525) );
  AOI21_X1 U13337 ( .B1(n10444), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n10525), .ZN(n10526) );
  NAND4_X1 U13338 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10530) );
  NOR2_X1 U13339 ( .A1(n10531), .A2(n10530), .ZN(n14322) );
  AOI22_X1 U13340 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13341 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13342 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13343 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10532) );
  NAND4_X1 U13344 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10541) );
  AOI22_X1 U13345 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13346 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13347 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13348 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n10957), .ZN(n10536) );
  NAND4_X1 U13349 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10540) );
  OR2_X1 U13350 ( .A1(n10541), .A2(n10540), .ZN(n14314) );
  AOI22_X1 U13351 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13352 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U13353 ( .A1(n10951), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13354 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10542) );
  NAND4_X1 U13355 ( .A1(n10545), .A2(n10544), .A3(n10543), .A4(n10542), .ZN(
        n10556) );
  AOI22_X1 U13356 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13357 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13358 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10552) );
  INV_X1 U13359 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10549) );
  INV_X1 U13360 ( .A(n10870), .ZN(n10548) );
  INV_X1 U13361 ( .A(n10546), .ZN(n10547) );
  INV_X1 U13362 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13225) );
  OAI22_X1 U13363 ( .A1(n10549), .A2(n10548), .B1(n10547), .B2(n13225), .ZN(
        n10550) );
  INV_X1 U13364 ( .A(n10550), .ZN(n10551) );
  NAND4_X1 U13365 ( .A1(n10554), .A2(n10553), .A3(n10552), .A4(n10551), .ZN(
        n10555) );
  AOI22_X1 U13366 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13367 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13368 ( .A1(n10951), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13369 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10557) );
  NAND4_X1 U13370 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10566) );
  AOI22_X1 U13371 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13372 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10870), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13373 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10510), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13374 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n10957), .ZN(n10561) );
  NAND4_X1 U13375 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10565) );
  NOR2_X1 U13376 ( .A1(n10566), .A2(n10565), .ZN(n14302) );
  AOI22_X1 U13377 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10404), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13378 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13379 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13380 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10429), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10567) );
  NAND4_X1 U13381 ( .A1(n10570), .A2(n10569), .A3(n10568), .A4(n10567), .ZN(
        n10576) );
  AOI22_X1 U13382 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10455), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13383 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10510), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13384 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10499), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13385 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n10957), .ZN(n10571) );
  NAND4_X1 U13386 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10575) );
  NOR2_X1 U13387 ( .A1(n10576), .A2(n10575), .ZN(n10616) );
  INV_X1 U13388 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12284) );
  OR2_X1 U13389 ( .A1(n10577), .A2(n12284), .ZN(n10582) );
  NAND2_X1 U13390 ( .A1(n10641), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10581) );
  NAND2_X1 U13391 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13392 ( .A1(n10752), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10579) );
  AND4_X1 U13393 ( .A1(n10582), .A2(n10581), .A3(n10580), .A4(n10579), .ZN(
        n10585) );
  AOI22_X1 U13394 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13395 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10583) );
  XNOR2_X1 U13396 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10747) );
  NAND4_X1 U13397 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10747), .ZN(
        n10595) );
  INV_X1 U13398 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10586) );
  OR2_X1 U13399 ( .A1(n10577), .A2(n10586), .ZN(n10590) );
  NAND2_X1 U13400 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10589) );
  NAND2_X1 U13401 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10588) );
  NAND2_X1 U13402 ( .A1(n10752), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10587) );
  AND4_X1 U13403 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10593) );
  INV_X1 U13404 ( .A(n10747), .ZN(n10755) );
  AOI22_X1 U13405 ( .A1(n10190), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10754), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13406 ( .A1(n10391), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10591) );
  NAND4_X1 U13407 ( .A1(n10593), .A2(n10755), .A3(n10592), .A4(n10591), .ZN(
        n10594) );
  NAND2_X1 U13408 ( .A1(n10595), .A2(n10594), .ZN(n10621) );
  NOR2_X1 U13409 ( .A1(n13275), .A2(n10621), .ZN(n10596) );
  XOR2_X1 U13410 ( .A(n10616), .B(n10596), .Z(n10622) );
  INV_X1 U13411 ( .A(n10621), .ZN(n10617) );
  NAND2_X1 U13412 ( .A1(n13275), .A2(n10617), .ZN(n14291) );
  NOR2_X2 U13413 ( .A1(n14292), .A2(n14291), .ZN(n14290) );
  INV_X1 U13414 ( .A(n10391), .ZN(n10729) );
  INV_X1 U13415 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10600) );
  INV_X1 U13416 ( .A(n10753), .ZN(n10728) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10599) );
  OAI22_X1 U13418 ( .A1(n10729), .A2(n10600), .B1(n10728), .B2(n10599), .ZN(
        n10604) );
  INV_X1 U13419 ( .A(n10754), .ZN(n10731) );
  INV_X1 U13420 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10602) );
  INV_X1 U13421 ( .A(n10190), .ZN(n10730) );
  INV_X1 U13422 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10601) );
  OAI22_X1 U13423 ( .A1(n10731), .A2(n10602), .B1(n10730), .B2(n10601), .ZN(
        n10603) );
  NOR2_X1 U13424 ( .A1(n10604), .A2(n10603), .ZN(n10607) );
  AOI22_X1 U13425 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13426 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10605) );
  NAND4_X1 U13427 ( .A1(n10607), .A2(n10606), .A3(n10605), .A4(n10747), .ZN(
        n10615) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10608) );
  INV_X1 U13429 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12709) );
  OAI22_X1 U13430 ( .A1(n10729), .A2(n10608), .B1(n10728), .B2(n12709), .ZN(
        n10610) );
  INV_X1 U13431 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12724) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12729) );
  OAI22_X1 U13433 ( .A1(n10731), .A2(n12724), .B1(n10730), .B2(n12729), .ZN(
        n10609) );
  NOR2_X1 U13434 ( .A1(n10610), .A2(n10609), .ZN(n10613) );
  AOI22_X1 U13435 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13436 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10611) );
  NAND4_X1 U13437 ( .A1(n10613), .A2(n10755), .A3(n10612), .A4(n10611), .ZN(
        n10614) );
  NAND2_X1 U13438 ( .A1(n10615), .A2(n10614), .ZN(n10624) );
  INV_X1 U13439 ( .A(n10616), .ZN(n10618) );
  NAND2_X1 U13440 ( .A1(n10618), .A2(n10617), .ZN(n10625) );
  XOR2_X1 U13441 ( .A(n10624), .B(n10625), .Z(n10619) );
  NAND2_X1 U13442 ( .A1(n10619), .A2(n10697), .ZN(n14284) );
  INV_X1 U13443 ( .A(n10624), .ZN(n10620) );
  NAND2_X1 U13444 ( .A1(n13275), .A2(n10620), .ZN(n14286) );
  NOR3_X1 U13445 ( .A1(n10622), .A2(n10621), .A3(n14286), .ZN(n10623) );
  NOR2_X1 U13446 ( .A1(n10625), .A2(n10624), .ZN(n10647) );
  INV_X1 U13447 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10627) );
  INV_X1 U13448 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10626) );
  OAI22_X1 U13449 ( .A1(n10729), .A2(n10627), .B1(n10728), .B2(n10626), .ZN(
        n10631) );
  INV_X1 U13450 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10629) );
  INV_X1 U13451 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10628) );
  OAI22_X1 U13452 ( .A1(n10731), .A2(n10629), .B1(n10730), .B2(n10628), .ZN(
        n10630) );
  NOR2_X1 U13453 ( .A1(n10631), .A2(n10630), .ZN(n10634) );
  AOI22_X1 U13454 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13455 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10632) );
  NAND4_X1 U13456 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10747), .ZN(
        n10646) );
  INV_X1 U13457 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10636) );
  INV_X1 U13458 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10635) );
  OAI22_X1 U13459 ( .A1(n10729), .A2(n10636), .B1(n10728), .B2(n10635), .ZN(
        n10640) );
  INV_X1 U13460 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10638) );
  INV_X1 U13461 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10637) );
  OAI22_X1 U13462 ( .A1(n10731), .A2(n10638), .B1(n10730), .B2(n10637), .ZN(
        n10639) );
  NOR2_X1 U13463 ( .A1(n10640), .A2(n10639), .ZN(n10644) );
  AOI22_X1 U13464 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13465 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10642) );
  NAND4_X1 U13466 ( .A1(n10644), .A2(n10755), .A3(n10643), .A4(n10642), .ZN(
        n10645) );
  AND2_X1 U13467 ( .A1(n10646), .A2(n10645), .ZN(n10649) );
  NAND2_X1 U13468 ( .A1(n10647), .A2(n10649), .ZN(n10694) );
  OAI211_X1 U13469 ( .C1(n10647), .C2(n10649), .A(n10697), .B(n10694), .ZN(
        n10651) );
  INV_X1 U13470 ( .A(n10651), .ZN(n10648) );
  INV_X1 U13471 ( .A(n10649), .ZN(n10650) );
  NOR2_X1 U13472 ( .A1(n19592), .A2(n10650), .ZN(n14275) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10654) );
  INV_X1 U13474 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10653) );
  OAI22_X1 U13475 ( .A1(n10729), .A2(n10654), .B1(n10728), .B2(n10653), .ZN(
        n10658) );
  INV_X1 U13476 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10656) );
  INV_X1 U13477 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10655) );
  OAI22_X1 U13478 ( .A1(n10731), .A2(n10656), .B1(n10730), .B2(n10655), .ZN(
        n10657) );
  NOR2_X1 U13479 ( .A1(n10658), .A2(n10657), .ZN(n10661) );
  AOI22_X1 U13480 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13481 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10659) );
  NAND4_X1 U13482 ( .A1(n10661), .A2(n10660), .A3(n10659), .A4(n10747), .ZN(
        n10668) );
  INV_X1 U13483 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12758) );
  INV_X1 U13484 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12754) );
  OAI22_X1 U13485 ( .A1(n10729), .A2(n12758), .B1(n10728), .B2(n12754), .ZN(
        n10663) );
  INV_X1 U13486 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12759) );
  INV_X1 U13487 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12755) );
  OAI22_X1 U13488 ( .A1(n10731), .A2(n12759), .B1(n10730), .B2(n12755), .ZN(
        n10662) );
  NOR2_X1 U13489 ( .A1(n10663), .A2(n10662), .ZN(n10666) );
  AOI22_X1 U13490 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13491 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13492 ( .A1(n10666), .A2(n10755), .A3(n10665), .A4(n10664), .ZN(
        n10667) );
  AND2_X1 U13493 ( .A1(n10668), .A2(n10667), .ZN(n10692) );
  XNOR2_X1 U13494 ( .A(n10694), .B(n10692), .ZN(n10669) );
  XNOR2_X1 U13495 ( .A(n10670), .B(n10151), .ZN(n14271) );
  NAND2_X1 U13496 ( .A1(n13275), .A2(n10692), .ZN(n14270) );
  NOR2_X1 U13497 ( .A1(n14271), .A2(n14270), .ZN(n14269) );
  INV_X1 U13498 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10673) );
  INV_X1 U13499 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10672) );
  OAI22_X1 U13500 ( .A1(n10729), .A2(n10673), .B1(n10728), .B2(n10672), .ZN(
        n10677) );
  INV_X1 U13501 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10675) );
  INV_X1 U13502 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10674) );
  OAI22_X1 U13503 ( .A1(n10731), .A2(n10675), .B1(n10730), .B2(n10674), .ZN(
        n10676) );
  NOR2_X1 U13504 ( .A1(n10677), .A2(n10676), .ZN(n10680) );
  AOI22_X1 U13505 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13506 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10678) );
  NAND4_X1 U13507 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10747), .ZN(
        n10691) );
  INV_X1 U13508 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10682) );
  INV_X1 U13509 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10681) );
  OAI22_X1 U13510 ( .A1(n10729), .A2(n10682), .B1(n10728), .B2(n10681), .ZN(
        n10686) );
  INV_X1 U13511 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10684) );
  INV_X1 U13512 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10683) );
  OAI22_X1 U13513 ( .A1(n10731), .A2(n10684), .B1(n10730), .B2(n10683), .ZN(
        n10685) );
  NOR2_X1 U13514 ( .A1(n10686), .A2(n10685), .ZN(n10689) );
  AOI22_X1 U13515 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13516 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10687) );
  NAND4_X1 U13517 ( .A1(n10689), .A2(n10755), .A3(n10688), .A4(n10687), .ZN(
        n10690) );
  NAND2_X1 U13518 ( .A1(n10691), .A2(n10690), .ZN(n10695) );
  INV_X1 U13519 ( .A(n10695), .ZN(n10702) );
  INV_X1 U13520 ( .A(n10692), .ZN(n10693) );
  OR2_X1 U13521 ( .A1(n10694), .A2(n10693), .ZN(n10696) );
  INV_X1 U13522 ( .A(n10696), .ZN(n10698) );
  OR2_X1 U13523 ( .A1(n10696), .A2(n10695), .ZN(n10739) );
  OAI211_X1 U13524 ( .C1(n10702), .C2(n10698), .A(n10739), .B(n10697), .ZN(
        n10700) );
  NAND2_X1 U13525 ( .A1(n13275), .A2(n10702), .ZN(n14262) );
  INV_X1 U13526 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10705) );
  INV_X1 U13527 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10704) );
  OAI22_X1 U13528 ( .A1(n10729), .A2(n10705), .B1(n10728), .B2(n10704), .ZN(
        n10709) );
  INV_X1 U13529 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10707) );
  INV_X1 U13530 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10706) );
  OAI22_X1 U13531 ( .A1(n10731), .A2(n10707), .B1(n10730), .B2(n10706), .ZN(
        n10708) );
  NOR2_X1 U13532 ( .A1(n10709), .A2(n10708), .ZN(n10712) );
  AOI22_X1 U13533 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13534 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10710) );
  NAND4_X1 U13535 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10747), .ZN(
        n10719) );
  INV_X1 U13536 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13220) );
  OAI22_X1 U13537 ( .A1(n10729), .A2(n13225), .B1(n10728), .B2(n13220), .ZN(
        n10714) );
  INV_X1 U13538 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13226) );
  INV_X1 U13539 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13218) );
  OAI22_X1 U13540 ( .A1(n10731), .A2(n13226), .B1(n10730), .B2(n13218), .ZN(
        n10713) );
  NOR2_X1 U13541 ( .A1(n10714), .A2(n10713), .ZN(n10717) );
  AOI22_X1 U13542 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13543 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13544 ( .A1(n10717), .A2(n10755), .A3(n10716), .A4(n10715), .ZN(
        n10718) );
  INV_X1 U13545 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10720) );
  INV_X1 U13546 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n20579) );
  OAI22_X1 U13547 ( .A1(n10729), .A2(n10720), .B1(n10731), .B2(n20579), .ZN(
        n10724) );
  INV_X1 U13548 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10722) );
  INV_X1 U13549 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10721) );
  OAI22_X1 U13550 ( .A1(n10728), .A2(n10722), .B1(n10730), .B2(n10721), .ZN(
        n10723) );
  NOR2_X1 U13551 ( .A1(n10724), .A2(n10723), .ZN(n10727) );
  AOI22_X1 U13552 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13553 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10725) );
  NAND4_X1 U13554 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10747), .ZN(
        n10738) );
  INV_X1 U13555 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13262) );
  INV_X1 U13556 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13258) );
  OAI22_X1 U13557 ( .A1(n10729), .A2(n13262), .B1(n10728), .B2(n13258), .ZN(
        n10733) );
  INV_X1 U13558 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13263) );
  INV_X1 U13559 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13259) );
  OAI22_X1 U13560 ( .A1(n10731), .A2(n13263), .B1(n10730), .B2(n13259), .ZN(
        n10732) );
  NOR2_X1 U13561 ( .A1(n10733), .A2(n10732), .ZN(n10736) );
  AOI22_X1 U13562 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10752), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13563 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10734) );
  NAND4_X1 U13564 ( .A1(n10736), .A2(n10755), .A3(n10735), .A4(n10734), .ZN(
        n10737) );
  NAND2_X1 U13565 ( .A1(n10738), .A2(n10737), .ZN(n10742) );
  INV_X1 U13566 ( .A(n10739), .ZN(n14257) );
  AND2_X1 U13567 ( .A1(n19592), .A2(n9717), .ZN(n10740) );
  NAND2_X1 U13568 ( .A1(n14257), .A2(n10740), .ZN(n10741) );
  NOR2_X1 U13569 ( .A1(n10741), .A2(n10742), .ZN(n10743) );
  AOI21_X1 U13570 ( .B1(n10742), .B2(n10741), .A(n10743), .ZN(n14251) );
  INV_X1 U13571 ( .A(n10743), .ZN(n10744) );
  AOI22_X1 U13572 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10391), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13573 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10239), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U13574 ( .A1(n10746), .A2(n10745), .ZN(n10761) );
  AOI22_X1 U13575 ( .A1(n10752), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10190), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13576 ( .A1(n10754), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10748) );
  NAND3_X1 U13577 ( .A1(n10749), .A2(n10748), .A3(n10747), .ZN(n10760) );
  AOI22_X1 U13578 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10391), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13579 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13580 ( .A1(n10751), .A2(n10750), .ZN(n10759) );
  AOI22_X1 U13581 ( .A1(n10752), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10190), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13582 ( .A1(n10754), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10756) );
  NAND3_X1 U13583 ( .A1(n10757), .A2(n10756), .A3(n10755), .ZN(n10758) );
  OAI22_X1 U13584 ( .A1(n10761), .A2(n10760), .B1(n10759), .B2(n10758), .ZN(
        n10762) );
  AOI22_X1 U13585 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10417), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13586 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13587 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10951), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13588 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10763) );
  NAND4_X1 U13589 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n10772) );
  AOI22_X1 U13590 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10522), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13591 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13592 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10499), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13593 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n10957), .ZN(n10767) );
  NAND4_X1 U13594 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(
        n10771) );
  NAND2_X1 U13595 ( .A1(n19570), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10775) );
  NAND2_X1 U13596 ( .A1(n10773), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10774) );
  NAND2_X1 U13597 ( .A1(n10775), .A2(n10774), .ZN(n10796) );
  NAND2_X1 U13598 ( .A1(n19578), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10795) );
  NAND2_X1 U13599 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19560), .ZN(
        n10791) );
  NAND2_X1 U13600 ( .A1(n10794), .A2(n10791), .ZN(n10777) );
  NAND2_X1 U13601 ( .A1(n10776), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10792) );
  XNOR2_X1 U13602 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10789) );
  INV_X1 U13603 ( .A(n10789), .ZN(n10778) );
  NAND2_X1 U13604 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15174), .ZN(
        n10807) );
  OR2_X1 U13605 ( .A1(n10806), .A2(n10807), .ZN(n10828) );
  MUX2_X1 U13606 ( .A(n13405), .B(n10828), .S(n12939), .Z(n12949) );
  AOI22_X1 U13607 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U13608 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U13609 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13610 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10779) );
  NAND4_X1 U13611 ( .A1(n10782), .A2(n10781), .A3(n10780), .A4(n10779), .ZN(
        n10788) );
  AOI22_X1 U13612 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10522), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10786) );
  AOI22_X1 U13613 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13614 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10455), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13615 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n10957), .ZN(n10783) );
  NAND4_X1 U13616 ( .A1(n10786), .A2(n10785), .A3(n10784), .A4(n10783), .ZN(
        n10787) );
  XNOR2_X1 U13617 ( .A(n10790), .B(n10789), .ZN(n10826) );
  MUX2_X1 U13618 ( .A(n12765), .B(n10826), .S(n12939), .Z(n12772) );
  NAND2_X1 U13619 ( .A1(n12949), .A2(n12772), .ZN(n12161) );
  NAND2_X1 U13620 ( .A1(n12161), .A2(n12939), .ZN(n10811) );
  AND2_X1 U13621 ( .A1(n10792), .A2(n10791), .ZN(n10793) );
  XNOR2_X1 U13622 ( .A(n10794), .B(n10793), .ZN(n10827) );
  AND2_X1 U13623 ( .A1(n12939), .A2(n10827), .ZN(n12155) );
  AOI21_X1 U13624 ( .B1(n12254), .B2(n19592), .A(n10827), .ZN(n10803) );
  INV_X1 U13625 ( .A(n10827), .ZN(n10800) );
  OAI21_X1 U13626 ( .B1(n19578), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10795), .ZN(n12201) );
  INV_X1 U13627 ( .A(n12939), .ZN(n12200) );
  OAI21_X1 U13628 ( .B1(n12201), .B2(n10796), .A(n12200), .ZN(n10799) );
  INV_X1 U13629 ( .A(n12201), .ZN(n12157) );
  NAND2_X1 U13630 ( .A1(n10796), .A2(n10795), .ZN(n12158) );
  AND2_X1 U13631 ( .A1(n10797), .A2(n12158), .ZN(n10830) );
  OAI211_X1 U13632 ( .C1(n19592), .C2(n12157), .A(n18868), .B(n10830), .ZN(
        n10798) );
  OAI211_X1 U13633 ( .C1(n10801), .C2(n10800), .A(n10799), .B(n10798), .ZN(
        n10802) );
  OAI21_X1 U13634 ( .B1(n12155), .B2(n10803), .A(n10802), .ZN(n10804) );
  NAND2_X1 U13635 ( .A1(n10804), .A2(n10826), .ZN(n10810) );
  INV_X1 U13636 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15409) );
  AND2_X1 U13637 ( .A1(n15409), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10805) );
  OAI21_X1 U13638 ( .B1(n10828), .B2(n12939), .A(n12160), .ZN(n10809) );
  AOI21_X1 U13639 ( .B1(n10811), .B2(n10810), .A(n10809), .ZN(n10812) );
  MUX2_X1 U13640 ( .A(n10812), .B(n15174), .S(n15967), .Z(n12780) );
  NAND2_X1 U13641 ( .A1(n10816), .A2(n18884), .ZN(n10817) );
  NAND2_X1 U13642 ( .A1(n10815), .A2(n10817), .ZN(n10823) );
  NAND2_X1 U13643 ( .A1(n12778), .A2(n13275), .ZN(n10824) );
  NAND2_X1 U13644 ( .A1(n10824), .A2(n18868), .ZN(n10818) );
  NAND2_X1 U13645 ( .A1(n10818), .A2(n18913), .ZN(n10820) );
  AOI21_X1 U13646 ( .B1(n10820), .B2(n18884), .A(n10819), .ZN(n10822) );
  AND2_X1 U13647 ( .A1(n12779), .A2(n13275), .ZN(n12163) );
  OAI21_X1 U13648 ( .B1(n10821), .B2(n11000), .A(n12163), .ZN(n12808) );
  NAND2_X1 U13649 ( .A1(n10825), .A2(n10815), .ZN(n15945) );
  NAND3_X1 U13650 ( .A1(n10828), .A2(n10827), .A3(n10826), .ZN(n12166) );
  INV_X1 U13651 ( .A(n12166), .ZN(n10829) );
  NAND2_X1 U13652 ( .A1(n10830), .A2(n10829), .ZN(n10831) );
  NAND2_X1 U13653 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19602) );
  NAND4_X1 U13654 ( .A1(n15945), .A2(n12790), .A3(n10832), .A4(n19602), .ZN(
        n10833) );
  OAI21_X1 U13655 ( .B1(n15943), .B2(n15948), .A(n10833), .ZN(n13041) );
  NAND3_X1 U13656 ( .A1(n12788), .A2(n10834), .A3(n18903), .ZN(n10835) );
  NOR2_X1 U13657 ( .A1(n10836), .A2(n10835), .ZN(n12818) );
  OR2_X1 U13658 ( .A1(n13041), .A2(n12818), .ZN(n10838) );
  NAND2_X1 U13659 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20564), .ZN(n12930) );
  INV_X1 U13660 ( .A(n12930), .ZN(n10837) );
  INV_X1 U13661 ( .A(n10281), .ZN(n10877) );
  NAND2_X1 U13662 ( .A1(n12024), .A2(n18761), .ZN(n11017) );
  AOI22_X1 U13663 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n10842) );
  AND2_X1 U13664 ( .A1(n18913), .A2(n19571), .ZN(n10839) );
  INV_X2 U13665 ( .A(n10154), .ZN(n10996) );
  NAND2_X1 U13666 ( .A1(n10996), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10841) );
  AND2_X1 U13667 ( .A1(n10842), .A2(n10841), .ZN(n10999) );
  AOI22_X1 U13668 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U13669 ( .A1(n10996), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10843) );
  NAND2_X1 U13670 ( .A1(n10844), .A2(n10843), .ZN(n14742) );
  INV_X1 U13671 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U13672 ( .A1(n10996), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10846) );
  NAND2_X1 U13673 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10845) );
  OAI211_X1 U13674 ( .C1(n9645), .C2(n12342), .A(n10846), .B(n10845), .ZN(
        n14415) );
  AOI22_X1 U13675 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n10848) );
  NAND2_X1 U13676 ( .A1(n10996), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10847) );
  AOI222_X1 U13677 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n10996), .B1(n14161), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n14160), .C2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14798) );
  AOI22_X1 U13678 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U13679 ( .A1(n10964), .A2(n10159), .ZN(n10851) );
  NAND2_X1 U13680 ( .A1(n10996), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13681 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U13682 ( .A1(n10964), .A2(n12986), .ZN(n10854) );
  NAND2_X1 U13683 ( .A1(n10996), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13684 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n10856) );
  OAI21_X1 U13685 ( .B1(n12851), .B2(n10976), .A(n10856), .ZN(n10857) );
  AOI21_X1 U13686 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n10996), .A(n10857), 
        .ZN(n15882) );
  INV_X1 U13687 ( .A(n12559), .ZN(n10859) );
  AOI22_X1 U13688 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n10858) );
  OAI21_X1 U13689 ( .B1(n10859), .B2(n10976), .A(n10858), .ZN(n10860) );
  AOI21_X1 U13690 ( .B1(n10996), .B2(P2_REIP_REG_8__SCAN_IN), .A(n10860), .ZN(
        n12978) );
  INV_X1 U13691 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15911) );
  INV_X1 U13692 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18783) );
  INV_X1 U13693 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19497) );
  OAI222_X1 U13694 ( .A1(n15911), .A2(n10861), .B1(n9645), .B2(n18783), .C1(
        n10154), .C2(n19497), .ZN(n15906) );
  AOI22_X1 U13695 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U13696 ( .A1(n10964), .A2(n13405), .ZN(n10863) );
  NAND2_X1 U13697 ( .A1(n10996), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13698 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13699 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13700 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13701 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10866) );
  NAND4_X1 U13702 ( .A1(n10869), .A2(n10868), .A3(n10867), .A4(n10866), .ZN(
        n10876) );
  AOI22_X1 U13703 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U13704 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13705 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13706 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10871) );
  NAND4_X1 U13707 ( .A1(n10874), .A2(n10873), .A3(n10872), .A4(n10871), .ZN(
        n10875) );
  NOR2_X1 U13708 ( .A1(n10876), .A2(n10875), .ZN(n12230) );
  OR2_X1 U13709 ( .A1(n12230), .A2(n10976), .ZN(n10880) );
  MUX2_X1 U13710 ( .A(n18913), .B(n19578), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10878) );
  NAND2_X1 U13711 ( .A1(n10993), .A2(n10877), .ZN(n10912) );
  AND2_X1 U13712 ( .A1(n10878), .A2(n10912), .ZN(n10879) );
  NAND2_X1 U13713 ( .A1(n10880), .A2(n10879), .ZN(n12280) );
  INV_X1 U13714 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18680) );
  NAND2_X1 U13715 ( .A1(n10996), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10884) );
  NAND2_X1 U13716 ( .A1(n11000), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10881) );
  OAI211_X1 U13717 ( .C1(n13275), .C2(n12207), .A(n10881), .B(n19571), .ZN(
        n10882) );
  INV_X1 U13718 ( .A(n10882), .ZN(n10883) );
  NAND2_X1 U13719 ( .A1(n10884), .A2(n10883), .ZN(n12279) );
  INV_X1 U13720 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18795) );
  INV_X1 U13721 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19486) );
  NAND2_X1 U13722 ( .A1(n10996), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10886) );
  INV_X1 U13723 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18850) );
  NAND2_X1 U13724 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10885) );
  OAI211_X1 U13725 ( .C1(n9645), .C2(n18795), .A(n10886), .B(n10885), .ZN(
        n10887) );
  NOR2_X1 U13726 ( .A1(n12282), .A2(n10887), .ZN(n10902) );
  XNOR2_X1 U13727 ( .A(n12282), .B(n10887), .ZN(n12666) );
  AOI22_X1 U13728 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10957), .ZN(n10891) );
  AOI22_X1 U13729 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13730 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10429), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13731 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10522), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10888) );
  NAND4_X1 U13732 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n10897) );
  AOI22_X1 U13733 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13734 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13735 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10405), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13736 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10865), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10892) );
  NAND4_X1 U13737 ( .A1(n10895), .A2(n10894), .A3(n10893), .A4(n10892), .ZN(
        n10896) );
  NOR2_X1 U13738 ( .A1(n10897), .A2(n10896), .ZN(n12236) );
  OR2_X1 U13739 ( .A1(n12236), .A2(n10976), .ZN(n10900) );
  NAND2_X1 U13740 ( .A1(n10281), .A2(n18913), .ZN(n10898) );
  MUX2_X1 U13741 ( .A(n10898), .B(n19570), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10899) );
  NAND2_X1 U13742 ( .A1(n10900), .A2(n10899), .ZN(n12665) );
  NOR2_X1 U13743 ( .A1(n12666), .A2(n12665), .ZN(n10901) );
  AOI22_X1 U13744 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13745 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13746 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13747 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13748 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10499), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13749 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13750 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10522), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U13751 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n10957), .ZN(n10907) );
  NAND4_X1 U13752 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n10911) );
  INV_X1 U13753 ( .A(n12232), .ZN(n12744) );
  NAND2_X1 U13754 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10913) );
  OAI211_X1 U13755 ( .C1(n10976), .C2(n12744), .A(n10913), .B(n10912), .ZN(
        n10915) );
  NOR2_X1 U13756 ( .A1(n10914), .A2(n10915), .ZN(n10918) );
  XNOR2_X1 U13757 ( .A(n10915), .B(n10914), .ZN(n12662) );
  INV_X1 U13758 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18793) );
  INV_X1 U13759 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19488) );
  NAND2_X1 U13760 ( .A1(n10996), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U13761 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10916) );
  OAI211_X1 U13762 ( .C1(n9645), .C2(n18793), .A(n10917), .B(n10916), .ZN(
        n12661) );
  NOR2_X1 U13763 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  AOI22_X1 U13764 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10922) );
  NAND2_X1 U13765 ( .A1(n10964), .A2(n12765), .ZN(n10921) );
  NAND2_X1 U13766 ( .A1(n10996), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U13767 ( .A1(n14160), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10919) );
  NAND4_X1 U13768 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(
        n12658) );
  AOI22_X1 U13769 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13770 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13771 ( .A1(n10951), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13772 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10923) );
  NAND4_X1 U13773 ( .A1(n10926), .A2(n10925), .A3(n10924), .A4(n10923), .ZN(
        n10932) );
  AOI22_X1 U13774 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13775 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13776 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13777 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U13778 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n10931) );
  AOI22_X1 U13779 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U13780 ( .A1(n10996), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10933) );
  OAI211_X1 U13781 ( .C1(n13238), .C2(n10976), .A(n10934), .B(n10933), .ZN(
        n14881) );
  AOI22_X1 U13782 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13783 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13784 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13785 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10935) );
  NAND4_X1 U13786 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(
        n10944) );
  AOI22_X1 U13787 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13788 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13789 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10870), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13790 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n10957), .ZN(n10939) );
  NAND4_X1 U13791 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10943) );
  INV_X1 U13792 ( .A(n13276), .ZN(n10945) );
  NAND2_X1 U13793 ( .A1(n10964), .A2(n10945), .ZN(n10946) );
  INV_X1 U13794 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18785) );
  NAND2_X1 U13795 ( .A1(n10996), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U13796 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10948) );
  OAI211_X1 U13797 ( .C1(n9645), .C2(n18785), .A(n10949), .B(n10948), .ZN(
        n14859) );
  AOI22_X1 U13798 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13799 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10951), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U13800 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10405), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U13801 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10952) );
  NAND4_X1 U13802 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n10963) );
  AOI22_X1 U13803 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10870), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13804 ( .A1(n10404), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13805 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10522), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13806 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n10957), .ZN(n10958) );
  NAND4_X1 U13807 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10962) );
  AOI22_X1 U13808 ( .A1(n14860), .A2(n14859), .B1(n10964), .B2(n13426), .ZN(
        n10965) );
  INV_X1 U13809 ( .A(n10965), .ZN(n15907) );
  AOI22_X1 U13810 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U13811 ( .A1(n10996), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10966) );
  OAI211_X1 U13812 ( .C1(n12622), .C2(n10976), .A(n10967), .B(n10966), .ZN(
        n14852) );
  INV_X1 U13813 ( .A(n12864), .ZN(n10970) );
  AOI22_X1 U13814 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n10969) );
  NAND2_X1 U13815 ( .A1(n10996), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10968) );
  OAI211_X1 U13816 ( .C1(n10970), .C2(n10976), .A(n10969), .B(n10968), .ZN(
        n14835) );
  NAND2_X1 U13817 ( .A1(n14834), .A2(n14835), .ZN(n14836) );
  NOR2_X2 U13818 ( .A1(n12965), .A2(n14836), .ZN(n14809) );
  INV_X1 U13819 ( .A(n12985), .ZN(n10973) );
  AOI22_X1 U13820 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n10972) );
  NAND2_X1 U13821 ( .A1(n10996), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10971) );
  OAI211_X1 U13822 ( .C1(n10973), .C2(n10976), .A(n10972), .B(n10971), .ZN(
        n14810) );
  AOI22_X1 U13823 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U13824 ( .A1(n10996), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10974) );
  OAI211_X1 U13825 ( .C1(n13082), .C2(n10976), .A(n10975), .B(n10974), .ZN(
        n15846) );
  INV_X1 U13826 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U13827 ( .A1(n10996), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U13828 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10977) );
  OAI211_X1 U13829 ( .C1(n9645), .C2(n12328), .A(n10978), .B(n10977), .ZN(
        n14424) );
  NAND2_X1 U13830 ( .A1(n14797), .A2(n14424), .ZN(n14775) );
  NOR2_X2 U13831 ( .A1(n14776), .A2(n14775), .ZN(n14777) );
  AOI22_X1 U13832 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U13833 ( .A1(n10996), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10979) );
  NAND2_X1 U13834 ( .A1(n10980), .A2(n10979), .ZN(n14228) );
  INV_X1 U13835 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U13836 ( .A1(n10996), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U13837 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10981) );
  OAI211_X1 U13838 ( .C1(n9645), .C2(n12332), .A(n10982), .B(n10981), .ZN(
        n14405) );
  NAND2_X1 U13839 ( .A1(n14742), .A2(n14741), .ZN(n14744) );
  AOI22_X1 U13840 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n10984) );
  NAND2_X1 U13841 ( .A1(n10996), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10983) );
  AND2_X1 U13842 ( .A1(n10984), .A2(n10983), .ZN(n14396) );
  AOI22_X1 U13843 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U13844 ( .A1(n10996), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U13845 ( .A1(n10986), .A2(n10985), .ZN(n14387) );
  AOI22_X1 U13846 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13847 ( .A1(n10996), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10987) );
  AND2_X1 U13848 ( .A1(n10988), .A2(n10987), .ZN(n14378) );
  AOI22_X1 U13849 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n10990) );
  NAND2_X1 U13850 ( .A1(n10996), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10989) );
  AND2_X1 U13851 ( .A1(n10990), .A2(n10989), .ZN(n14371) );
  AOI22_X1 U13852 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U13853 ( .A1(n10996), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10991) );
  AND2_X1 U13854 ( .A1(n10992), .A2(n10991), .ZN(n14212) );
  NOR2_X2 U13855 ( .A1(n14373), .A2(n14212), .ZN(n14213) );
  AOI22_X1 U13856 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n10995) );
  NAND2_X1 U13857 ( .A1(n10996), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U13858 ( .A1(n10995), .A2(n10994), .ZN(n14202) );
  AOI22_X1 U13859 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n10998) );
  NAND2_X1 U13860 ( .A1(n10996), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U13861 ( .A1(n10998), .A2(n10997), .ZN(n14183) );
  NAND2_X1 U13862 ( .A1(n14635), .A2(n18757), .ZN(n11016) );
  NAND2_X1 U13863 ( .A1(n18755), .A2(n10293), .ZN(n12277) );
  NOR4_X1 U13864 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n11004) );
  NOR4_X1 U13865 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_20__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n11003) );
  NOR4_X1 U13866 ( .A1(P2_ADDRESS_REG_9__SCAN_IN), .A2(
        P2_ADDRESS_REG_8__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n11002) );
  NOR4_X1 U13867 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_12__SCAN_IN), .A3(P2_ADDRESS_REG_11__SCAN_IN), .A4(
        P2_ADDRESS_REG_10__SCAN_IN), .ZN(n11001) );
  NAND4_X1 U13868 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11010) );
  NAND2_X1 U13869 ( .A1(n20544), .A2(n20527), .ZN(n20642) );
  INV_X1 U13870 ( .A(n20642), .ZN(n11008) );
  NOR3_X1 U13871 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_2__SCAN_IN), .A3(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n11007) );
  NOR4_X1 U13872 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n11006) );
  NOR4_X1 U13873 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n11005) );
  NAND4_X1 U13874 ( .A1(n11008), .A2(n11007), .A3(n11006), .A4(n11005), .ZN(
        n11009) );
  NOR2_X2 U13875 ( .A1(n12277), .A2(n18859), .ZN(n18703) );
  NOR2_X2 U13876 ( .A1(n12277), .A2(n18861), .ZN(n18702) );
  AOI22_X1 U13877 ( .A1(n18703), .A2(BUF1_REG_30__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n11015) );
  INV_X1 U13878 ( .A(n11012), .ZN(n11013) );
  MUX2_X1 U13879 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n18859), .Z(n18711) );
  AOI22_X1 U13880 ( .A1(n18701), .A2(n18711), .B1(n18756), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n11014) );
  NAND2_X1 U13881 ( .A1(n11017), .A2(n10158), .ZN(P2_U2889) );
  BUF_X2 U13882 ( .A(n11688), .Z(n11815) );
  AOI22_X1 U13883 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11021) );
  NOR2_X4 U13884 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14111) );
  AND2_X2 U13885 ( .A1(n11024), .A2(n14111), .ZN(n11227) );
  AOI22_X1 U13886 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11020) );
  AND2_X2 U13887 ( .A1(n11025), .A2(n12484), .ZN(n11228) );
  AOI22_X1 U13888 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11297), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11019) );
  BUF_X4 U13889 ( .A(n11707), .Z(n11826) );
  AOI22_X1 U13890 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11018) );
  NAND4_X1 U13891 ( .A1(n11021), .A2(n11020), .A3(n11019), .A4(n11018), .ZN(
        n11031) );
  AOI22_X1 U13892 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11570), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11029) );
  AND2_X4 U13893 ( .A1(n12483), .A2(n14110), .ZN(n11819) );
  AOI22_X1 U13894 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11028) );
  AND2_X2 U13895 ( .A1(n11024), .A2(n11025), .ZN(n11827) );
  BUF_X4 U13896 ( .A(n11827), .Z(n11800) );
  AND2_X4 U13897 ( .A1(n14111), .A2(n12483), .ZN(n11825) );
  AOI22_X1 U13898 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11027) );
  AND2_X2 U13899 ( .A1(n11025), .A2(n12483), .ZN(n11073) );
  AND2_X2 U13900 ( .A1(n12484), .A2(n14110), .ZN(n11303) );
  AOI22_X1 U13901 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11026) );
  NAND4_X1 U13902 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n11030) );
  OR2_X2 U13903 ( .A1(n11031), .A2(n11030), .ZN(n11907) );
  NAND2_X1 U13904 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U13905 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U13906 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11033) );
  BUF_X4 U13907 ( .A(n11707), .Z(n11616) );
  NAND2_X1 U13908 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11032) );
  BUF_X2 U13909 ( .A(n11688), .Z(n11571) );
  NAND2_X1 U13910 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11039) );
  NAND2_X1 U13911 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11038) );
  NAND2_X1 U13912 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11037) );
  NAND2_X1 U13913 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11036) );
  NAND2_X1 U13914 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U13915 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U13916 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11042) );
  NAND2_X1 U13917 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11041) );
  NAND2_X1 U13918 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11048) );
  NAND2_X1 U13919 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11047) );
  NAND2_X1 U13920 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11046) );
  NAND2_X1 U13921 ( .A1(n11303), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11045) );
  NAND4_X4 U13922 ( .A1(n11052), .A2(n11051), .A3(n11050), .A4(n11049), .ZN(
        n11142) );
  AOI22_X1 U13923 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U13924 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U13925 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U13926 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11053) );
  NAND4_X1 U13927 ( .A1(n11056), .A2(n11055), .A3(n11054), .A4(n11053), .ZN(
        n11062) );
  AOI22_X1 U13928 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11073), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U13929 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U13930 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U13931 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11057) );
  NAND4_X1 U13932 ( .A1(n11060), .A2(n11059), .A3(n11058), .A4(n11057), .ZN(
        n11061) );
  OR2_X2 U13933 ( .A1(n11062), .A2(n11061), .ZN(n12408) );
  NAND2_X1 U13934 ( .A1(n11148), .A2(n12408), .ZN(n11157) );
  AOI22_X1 U13935 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U13936 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U13937 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U13938 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11063) );
  NAND4_X1 U13939 ( .A1(n11066), .A2(n11065), .A3(n11064), .A4(n11063), .ZN(
        n11072) );
  AOI22_X1 U13940 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U13941 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U13942 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U13943 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11067) );
  NAND4_X1 U13944 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11071) );
  OR2_X2 U13945 ( .A1(n11072), .A2(n11071), .ZN(n12469) );
  AOI22_X1 U13946 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U13947 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U13948 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U13949 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11074) );
  NAND4_X1 U13950 ( .A1(n11077), .A2(n11076), .A3(n11075), .A4(n11074), .ZN(
        n11083) );
  AOI22_X1 U13951 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U13952 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U13953 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U13954 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11078) );
  NAND4_X1 U13955 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11082) );
  OR2_X2 U13956 ( .A1(n11083), .A2(n11082), .ZN(n12429) );
  NAND2_X1 U13957 ( .A1(n12429), .A2(n12469), .ZN(n11149) );
  NAND2_X1 U13958 ( .A1(n13702), .A2(n11149), .ZN(n11084) );
  NAND2_X1 U13959 ( .A1(n11157), .A2(n11084), .ZN(n11099) );
  AND2_X1 U13960 ( .A1(n11907), .A2(n11142), .ZN(n11095) );
  AOI22_X1 U13961 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U13962 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U13963 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U13964 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11085) );
  NAND4_X1 U13965 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11094) );
  AOI22_X1 U13966 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U13967 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U13968 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U13969 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11089) );
  NAND4_X1 U13970 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n11093) );
  OR2_X2 U13971 ( .A1(n11094), .A2(n11093), .ZN(n12416) );
  NAND2_X2 U13972 ( .A1(n11141), .A2(n11142), .ZN(n11870) );
  NOR2_X2 U13973 ( .A1(n11099), .A2(n11098), .ZN(n11161) );
  NAND2_X1 U13974 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11103) );
  NAND2_X1 U13975 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11102) );
  NAND2_X1 U13976 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11101) );
  NAND2_X1 U13977 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11100) );
  NAND2_X1 U13978 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11107) );
  NAND2_X1 U13979 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11106) );
  NAND2_X1 U13980 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11105) );
  NAND2_X1 U13981 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11104) );
  NAND2_X1 U13982 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11111) );
  NAND2_X1 U13983 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11110) );
  NAND2_X1 U13984 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U13985 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11108) );
  NAND2_X1 U13986 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U13987 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11114) );
  NAND2_X1 U13988 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11113) );
  NAND2_X1 U13989 ( .A1(n11303), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11112) );
  NAND4_X4 U13990 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        n12443) );
  NOR2_X1 U13991 ( .A1(n11870), .A2(n12443), .ZN(n11120) );
  NAND2_X1 U13992 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U13993 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U13994 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U13995 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U13996 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11128) );
  NAND2_X1 U13997 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U13998 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11126) );
  NAND2_X1 U13999 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14000 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14001 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11131) );
  NAND2_X1 U14002 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U14003 ( .A1(n11303), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14004 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11136) );
  NAND2_X1 U14005 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11135) );
  NAND2_X1 U14006 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14007 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11133) );
  NAND4_X4 U14008 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n12889) );
  AND2_X2 U14009 ( .A1(n19875), .A2(n12408), .ZN(n12507) );
  INV_X2 U14010 ( .A(n11142), .ZN(n19887) );
  NAND3_X1 U14011 ( .A1(n19883), .A2(n12507), .A3(n9670), .ZN(n12421) );
  NAND2_X1 U14012 ( .A1(n12443), .A2(n12889), .ZN(n11921) );
  OR2_X2 U14013 ( .A1(n12421), .A2(n19855), .ZN(n12428) );
  NAND2_X1 U14014 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20411) );
  OAI21_X1 U14015 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20411), .ZN(n12354) );
  NOR2_X2 U14016 ( .A1(n12416), .A2(n12408), .ZN(n12634) );
  NAND2_X2 U14017 ( .A1(n11144), .A2(n11259), .ZN(n12430) );
  INV_X1 U14018 ( .A(n12408), .ZN(n19879) );
  NAND2_X1 U14019 ( .A1(n19879), .A2(n12443), .ZN(n11914) );
  NAND2_X2 U14020 ( .A1(n12408), .A2(n12889), .ZN(n11918) );
  INV_X1 U14021 ( .A(n12507), .ZN(n11145) );
  NAND2_X1 U14022 ( .A1(n13472), .A2(n11145), .ZN(n11846) );
  NAND2_X1 U14023 ( .A1(n19855), .A2(n12889), .ZN(n12886) );
  NAND2_X1 U14024 ( .A1(n12416), .A2(n12443), .ZN(n11845) );
  AND2_X1 U14025 ( .A1(n12886), .A2(n11845), .ZN(n11146) );
  OAI211_X1 U14026 ( .C1(n19883), .C2(n20489), .A(n12439), .B(n11146), .ZN(
        n11154) );
  NAND2_X1 U14027 ( .A1(n19887), .A2(n11907), .ZN(n11147) );
  AND2_X1 U14028 ( .A1(n11147), .A2(n12469), .ZN(n11155) );
  NAND2_X1 U14029 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11172) );
  OAI21_X1 U14030 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11172), .ZN(n20165) );
  OR2_X1 U14031 ( .A1(n15384), .A2(n20163), .ZN(n11166) );
  OAI21_X1 U14032 ( .B1(n12407), .B2(n20165), .A(n11166), .ZN(n11151) );
  INV_X1 U14033 ( .A(n11151), .ZN(n11152) );
  MUX2_X1 U14034 ( .A(n12407), .B(n15384), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11153) );
  INV_X1 U14035 ( .A(n11154), .ZN(n11160) );
  INV_X1 U14036 ( .A(n11155), .ZN(n11156) );
  NAND2_X1 U14037 ( .A1(n14128), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19613) );
  AOI21_X1 U14038 ( .B1(n11156), .B2(n13140), .A(n19613), .ZN(n11159) );
  NAND2_X1 U14039 ( .A1(n19855), .A2(n19871), .ZN(n13465) );
  AND2_X1 U14040 ( .A1(n13465), .A2(n13469), .ZN(n12276) );
  NAND2_X1 U14041 ( .A1(n12276), .A2(n11157), .ZN(n11158) );
  OR2_X1 U14042 ( .A1(n11843), .A2(n11907), .ZN(n12438) );
  NAND3_X1 U14043 ( .A1(n12444), .A2(n12456), .A3(n12889), .ZN(n11163) );
  INV_X1 U14044 ( .A(n11161), .ZN(n11162) );
  NAND2_X1 U14045 ( .A1(n11162), .A2(n13462), .ZN(n12445) );
  NAND3_X1 U14046 ( .A1(n11164), .A2(n11163), .A3(n12445), .ZN(n11194) );
  INV_X1 U14047 ( .A(n11165), .ZN(n11168) );
  NAND2_X1 U14048 ( .A1(n11166), .A2(n14112), .ZN(n11167) );
  NAND2_X1 U14049 ( .A1(n11168), .A2(n11167), .ZN(n11178) );
  NAND2_X1 U14050 ( .A1(n11246), .A2(n11178), .ZN(n11176) );
  NOR2_X1 U14051 ( .A1(n15384), .A2(n20226), .ZN(n11170) );
  INV_X1 U14052 ( .A(n12407), .ZN(n11174) );
  INV_X1 U14053 ( .A(n11172), .ZN(n11171) );
  NAND2_X1 U14054 ( .A1(n11171), .A2(n20226), .ZN(n20194) );
  NAND2_X1 U14055 ( .A1(n11172), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11173) );
  NAND2_X1 U14056 ( .A1(n20194), .A2(n11173), .ZN(n19865) );
  NAND2_X1 U14057 ( .A1(n11174), .A2(n19865), .ZN(n11177) );
  NAND2_X1 U14058 ( .A1(n11179), .A2(n11177), .ZN(n11175) );
  NAND4_X1 U14059 ( .A1(n11246), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(
        n11180) );
  AOI22_X1 U14060 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14061 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14062 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14063 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11181) );
  NAND4_X1 U14064 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .ZN(
        n11190) );
  AOI22_X1 U14065 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14066 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14067 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14068 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11185) );
  NAND4_X1 U14069 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(
        n11189) );
  OAI22_X2 U14070 ( .A1(n12631), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12690), 
        .B2(n13134), .ZN(n11193) );
  INV_X1 U14071 ( .A(n11898), .ZN(n11890) );
  INV_X1 U14072 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U14073 ( .A1(n19855), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11226) );
  OAI22_X1 U14074 ( .A1(n11890), .A2(n11191), .B1(n12690), .B2(n11226), .ZN(
        n11192) );
  INV_X1 U14075 ( .A(n11194), .ZN(n11195) );
  NAND2_X1 U14076 ( .A1(n11276), .A2(n20401), .ZN(n11219) );
  AOI22_X1 U14077 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11200) );
  AOI22_X1 U14078 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11576), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14079 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14080 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11197) );
  NAND4_X1 U14081 ( .A1(n11200), .A2(n11199), .A3(n11198), .A4(n11197), .ZN(
        n11206) );
  AOI22_X1 U14082 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14083 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14084 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14085 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11201) );
  NAND4_X1 U14086 ( .A1(n11204), .A2(n11203), .A3(n11202), .A4(n11201), .ZN(
        n11205) );
  AOI22_X1 U14087 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14088 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14089 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14090 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11207) );
  NAND4_X1 U14091 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n11216) );
  AOI22_X1 U14092 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14093 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14094 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14095 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11211) );
  NAND4_X1 U14096 ( .A1(n11214), .A2(n11213), .A3(n11212), .A4(n11211), .ZN(
        n11215) );
  XNOR2_X1 U14097 ( .A(n11240), .B(n12505), .ZN(n11217) );
  NAND2_X1 U14098 ( .A1(n11217), .A2(n11248), .ZN(n11218) );
  NAND2_X1 U14099 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14100 ( .A1(n19855), .A2(n12505), .ZN(n11220) );
  OAI211_X1 U14101 ( .C1(n11240), .C2(n12429), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n11220), .ZN(n11221) );
  INV_X1 U14102 ( .A(n11221), .ZN(n11222) );
  NAND2_X1 U14103 ( .A1(n11248), .A2(n13139), .ZN(n11224) );
  INV_X1 U14104 ( .A(n11226), .ZN(n11239) );
  AOI22_X1 U14105 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11232) );
  BUF_X1 U14106 ( .A(n11227), .Z(n11576) );
  AOI22_X1 U14107 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14108 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14109 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11229) );
  NAND4_X1 U14110 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n11238) );
  AOI22_X1 U14111 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14112 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14113 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14114 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11233) );
  NAND4_X1 U14115 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11237) );
  AOI22_X1 U14116 ( .A1(n11248), .A2(n11240), .B1(n11239), .B2(n12506), .ZN(
        n11242) );
  NAND2_X1 U14117 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11241) );
  INV_X1 U14118 ( .A(n19960), .ZN(n11245) );
  INV_X1 U14119 ( .A(n11243), .ZN(n11244) );
  NAND2_X1 U14120 ( .A1(n11245), .A2(n11244), .ZN(n19904) );
  NAND2_X1 U14121 ( .A1(n19904), .A2(n11246), .ZN(n12871) );
  INV_X1 U14122 ( .A(n12871), .ZN(n11247) );
  NAND2_X1 U14123 ( .A1(n11247), .A2(n20401), .ZN(n11250) );
  NAND2_X1 U14124 ( .A1(n11248), .A2(n12506), .ZN(n11249) );
  NAND2_X1 U14125 ( .A1(n11266), .A2(n12504), .ZN(n11255) );
  INV_X1 U14126 ( .A(n11251), .ZN(n11252) );
  NAND2_X1 U14127 ( .A1(n11257), .A2(n11256), .ZN(n11258) );
  NAND2_X1 U14128 ( .A1(n11260), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11443) );
  AND2_X1 U14129 ( .A1(n11259), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U14130 ( .A1(n11336), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11265) );
  INV_X1 U14131 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11262) );
  OAI21_X1 U14132 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11315), .ZN(n19809) );
  NAND2_X1 U14133 ( .A1(n11313), .A2(n19809), .ZN(n11261) );
  OAI21_X1 U14134 ( .B1(n11443), .B2(n11262), .A(n11261), .ZN(n11263) );
  AOI21_X1 U14135 ( .B1(n13203), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11263), .ZN(
        n11264) );
  AND2_X1 U14136 ( .A1(n11265), .A2(n11264), .ZN(n11284) );
  XNOR2_X2 U14137 ( .A(n11268), .B(n11267), .ZN(n19932) );
  NAND2_X1 U14138 ( .A1(n19932), .A2(n11514), .ZN(n11272) );
  AOI22_X1 U14139 ( .A1(n13203), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11260), .ZN(n11270) );
  NAND2_X1 U14140 ( .A1(n11336), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11269) );
  AND2_X1 U14141 ( .A1(n11270), .A2(n11269), .ZN(n11271) );
  NAND2_X1 U14142 ( .A1(n11272), .A2(n11271), .ZN(n12498) );
  NAND2_X1 U14143 ( .A1(n11275), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12398) );
  INV_X1 U14144 ( .A(n11336), .ZN(n11320) );
  NAND2_X1 U14145 ( .A1(n11278), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11280) );
  NAND2_X1 U14146 ( .A1(n11260), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11279) );
  OAI211_X1 U14147 ( .C1(n11320), .C2(n11277), .A(n11280), .B(n11279), .ZN(
        n11281) );
  AOI21_X1 U14148 ( .B1(n19961), .B2(n11514), .A(n11281), .ZN(n11282) );
  OR2_X1 U14149 ( .A1(n12398), .A2(n11282), .ZN(n12399) );
  INV_X1 U14150 ( .A(n11282), .ZN(n12400) );
  OR2_X1 U14151 ( .A1(n12400), .A2(n11812), .ZN(n11283) );
  NAND2_X1 U14152 ( .A1(n12399), .A2(n11283), .ZN(n12499) );
  NAND2_X1 U14153 ( .A1(n12564), .A2(n12563), .ZN(n12562) );
  INV_X1 U14154 ( .A(n11284), .ZN(n11285) );
  NAND2_X1 U14155 ( .A1(n11286), .A2(n11285), .ZN(n11287) );
  NAND2_X1 U14156 ( .A1(n11290), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11295) );
  NAND3_X1 U14157 ( .A1(n20626), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20079) );
  INV_X1 U14158 ( .A(n20079), .ZN(n11291) );
  NAND2_X1 U14159 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11291), .ZN(
        n20077) );
  NAND2_X1 U14160 ( .A1(n20626), .A2(n20077), .ZN(n11292) );
  NOR3_X1 U14161 ( .A1(n20626), .A2(n20226), .A3(n20163), .ZN(n20347) );
  NAND2_X1 U14162 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20347), .ZN(
        n20335) );
  NAND2_X1 U14163 ( .A1(n11292), .A2(n20335), .ZN(n19856) );
  OAI22_X1 U14164 ( .A1(n12407), .A2(n19856), .B1(n15384), .B2(n20626), .ZN(
        n11293) );
  INV_X1 U14165 ( .A(n11293), .ZN(n11294) );
  XNOR2_X2 U14166 ( .A(n11289), .B(n19993), .ZN(n20110) );
  AOI22_X1 U14167 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14168 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14169 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14170 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11299) );
  NAND4_X1 U14171 ( .A1(n11302), .A2(n11301), .A3(n11300), .A4(n11299), .ZN(
        n11309) );
  AOI22_X1 U14172 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14173 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14174 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14175 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11304) );
  NAND4_X1 U14176 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(
        n11308) );
  AOI22_X1 U14177 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11879), .B2(n13107), .ZN(n11310) );
  INV_X1 U14178 ( .A(n19992), .ZN(n12839) );
  INV_X1 U14179 ( .A(n11315), .ZN(n11317) );
  INV_X1 U14180 ( .A(n11338), .ZN(n11316) );
  OAI21_X1 U14181 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11317), .A(
        n11316), .ZN(n12912) );
  AOI22_X1 U14182 ( .A1(n12878), .A2(n12912), .B1(n13202), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11319) );
  NAND2_X1 U14183 ( .A1(n13203), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11318) );
  OAI211_X1 U14184 ( .C1(n11320), .C2(n12495), .A(n11319), .B(n11318), .ZN(
        n11321) );
  INV_X1 U14185 ( .A(n11321), .ZN(n11322) );
  NAND2_X1 U14186 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11335) );
  AOI22_X1 U14187 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9598), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14188 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14189 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14190 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11324) );
  NAND4_X1 U14191 ( .A1(n11327), .A2(n11326), .A3(n11325), .A4(n11324), .ZN(
        n11333) );
  AOI22_X1 U14192 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14193 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14194 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14195 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11328) );
  NAND4_X1 U14196 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11332) );
  NAND2_X1 U14197 ( .A1(n11879), .A2(n13108), .ZN(n11334) );
  NAND2_X1 U14198 ( .A1(n11335), .A2(n11334), .ZN(n11343) );
  XNOR2_X1 U14199 ( .A(n11344), .B(n11343), .ZN(n13099) );
  NAND2_X1 U14200 ( .A1(n11336), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11341) );
  INV_X1 U14201 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19687) );
  AOI21_X1 U14202 ( .B1(n19687), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11337) );
  AOI21_X1 U14203 ( .B1(n13203), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11337), .ZN(
        n11340) );
  OAI21_X1 U14204 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11338), .A(
        n11357), .ZN(n19798) );
  NOR2_X1 U14205 ( .A1(n19798), .A2(n11812), .ZN(n11339) );
  AOI21_X1 U14206 ( .B1(n11341), .B2(n11340), .A(n11339), .ZN(n11342) );
  AOI21_X1 U14207 ( .B1(n13099), .B2(n11514), .A(n11342), .ZN(n12855) );
  NAND2_X1 U14208 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11356) );
  AOI22_X1 U14209 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14210 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14211 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14212 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11345) );
  NAND4_X1 U14213 ( .A1(n11348), .A2(n11347), .A3(n11346), .A4(n11345), .ZN(
        n11354) );
  AOI22_X1 U14214 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14215 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14216 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14217 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11349) );
  NAND4_X1 U14218 ( .A1(n11352), .A2(n11351), .A3(n11350), .A4(n11349), .ZN(
        n11353) );
  NAND2_X1 U14219 ( .A1(n11879), .A2(n13125), .ZN(n11355) );
  NAND2_X1 U14220 ( .A1(n11356), .A2(n11355), .ZN(n11363) );
  NAND2_X1 U14221 ( .A1(n13106), .A2(n11514), .ZN(n11362) );
  INV_X1 U14222 ( .A(n11357), .ZN(n11358) );
  INV_X1 U14223 ( .A(n11376), .ZN(n11377) );
  OAI21_X1 U14224 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11358), .A(
        n11377), .ZN(n19683) );
  NAND2_X1 U14225 ( .A1(n19683), .A2(n12878), .ZN(n11359) );
  OAI21_X1 U14226 ( .B1(n19670), .B2(n11443), .A(n11359), .ZN(n11360) );
  AOI21_X1 U14227 ( .B1(n13203), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11360), .ZN(
        n11361) );
  NAND2_X1 U14228 ( .A1(n11362), .A2(n11361), .ZN(n12844) );
  NAND2_X1 U14229 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11375) );
  AOI22_X1 U14230 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14231 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14232 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14233 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11364) );
  NAND4_X1 U14234 ( .A1(n11367), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(
        n11373) );
  AOI22_X1 U14235 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14236 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14237 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14238 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U14239 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11372) );
  NAND2_X1 U14240 ( .A1(n11879), .A2(n13124), .ZN(n11374) );
  NAND2_X1 U14241 ( .A1(n9675), .A2(n11382), .ZN(n13116) );
  INV_X1 U14242 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19747) );
  INV_X1 U14243 ( .A(n11387), .ZN(n11389) );
  INV_X1 U14244 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U14245 ( .A1(n11378), .A2(n11377), .ZN(n11379) );
  NAND2_X1 U14246 ( .A1(n11389), .A2(n11379), .ZN(n19669) );
  AOI22_X1 U14247 ( .A1(n19669), .A2(n11313), .B1(n13202), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11380) );
  OAI21_X1 U14248 ( .B1(n11394), .B2(n19747), .A(n11380), .ZN(n11381) );
  INV_X1 U14249 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U14250 ( .A1(n11879), .A2(n13139), .ZN(n11384) );
  OAI21_X1 U14251 ( .B1(n11890), .B2(n11385), .A(n11384), .ZN(n11386) );
  INV_X1 U14252 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11393) );
  INV_X1 U14253 ( .A(n11411), .ZN(n11391) );
  INV_X1 U14254 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U14255 ( .A1(n11389), .A2(n11388), .ZN(n11390) );
  NAND2_X1 U14256 ( .A1(n11391), .A2(n11390), .ZN(n19651) );
  AOI22_X1 U14257 ( .A1(n19651), .A2(n12878), .B1(n13202), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11392) );
  OAI21_X1 U14258 ( .B1(n11394), .B2(n11393), .A(n11392), .ZN(n11395) );
  AOI21_X1 U14259 ( .B1(n13123), .B2(n11514), .A(n11395), .ZN(n13005) );
  AOI22_X1 U14260 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14261 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14262 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14263 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14264 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11407) );
  AOI22_X1 U14265 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14266 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14267 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14268 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11402) );
  NAND4_X1 U14269 ( .A1(n11405), .A2(n11404), .A3(n11403), .A4(n11402), .ZN(
        n11406) );
  OAI21_X1 U14270 ( .B1(n11407), .B2(n11406), .A(n11514), .ZN(n11410) );
  XNOR2_X1 U14271 ( .A(n11411), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13145) );
  AOI22_X1 U14272 ( .A1(n13145), .A2(n11313), .B1(n13202), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11409) );
  NAND2_X1 U14273 ( .A1(n13203), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11408) );
  XOR2_X1 U14274 ( .A(n19636), .B(n11435), .Z(n19640) );
  AOI22_X1 U14275 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14276 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11571), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14277 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14278 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11412) );
  NAND4_X1 U14279 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11421) );
  AOI22_X1 U14280 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14281 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14282 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14283 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14284 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11420) );
  OR2_X1 U14285 ( .A1(n11421), .A2(n11420), .ZN(n11422) );
  AOI22_X1 U14286 ( .A1(n11514), .A2(n11422), .B1(n13202), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U14287 ( .A1(n13203), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11423) );
  OAI211_X1 U14288 ( .C1(n19640), .C2(n11812), .A(n11424), .B(n11423), .ZN(
        n13089) );
  AOI22_X1 U14289 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14290 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14291 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14292 ( .A1(n11706), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11425) );
  NAND4_X1 U14293 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11434) );
  AOI22_X1 U14294 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14295 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14296 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14297 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11429) );
  NAND4_X1 U14298 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n11433) );
  NOR2_X1 U14299 ( .A1(n11434), .A2(n11433), .ZN(n11439) );
  XNOR2_X1 U14300 ( .A(n11440), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13924) );
  NAND2_X1 U14301 ( .A1(n13924), .A2(n11313), .ZN(n11437) );
  AOI22_X1 U14302 ( .A1(n13203), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13202), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11436) );
  OAI211_X1 U14303 ( .C1(n11439), .C2(n11438), .A(n11437), .B(n11436), .ZN(
        n13150) );
  INV_X1 U14304 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11444) );
  OAI21_X1 U14305 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11441), .A(
        n11471), .ZN(n15543) );
  NAND2_X1 U14306 ( .A1(n15543), .A2(n12878), .ZN(n11442) );
  OAI21_X1 U14307 ( .B1(n11444), .B2(n11443), .A(n11442), .ZN(n11445) );
  AOI21_X1 U14308 ( .B1(n13203), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11445), .ZN(
        n13179) );
  AOI22_X1 U14309 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9598), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14310 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14311 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14312 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11446) );
  NAND4_X1 U14313 ( .A1(n11449), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11455) );
  AOI22_X1 U14314 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11571), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14315 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14316 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14317 ( .A1(n11706), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11450) );
  NAND4_X1 U14318 ( .A1(n11453), .A2(n11452), .A3(n11451), .A4(n11450), .ZN(
        n11454) );
  OR2_X1 U14319 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  NAND2_X1 U14320 ( .A1(n11514), .A2(n11456), .ZN(n13632) );
  XOR2_X1 U14321 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11489), .Z(
        n13921) );
  AOI22_X1 U14322 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11571), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14323 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14324 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14325 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11458) );
  NAND4_X1 U14326 ( .A1(n11461), .A2(n11460), .A3(n11459), .A4(n11458), .ZN(
        n11467) );
  AOI22_X1 U14327 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14328 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14329 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14330 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11462) );
  NAND4_X1 U14331 ( .A1(n11465), .A2(n11464), .A3(n11463), .A4(n11462), .ZN(
        n11466) );
  OR2_X1 U14332 ( .A1(n11467), .A2(n11466), .ZN(n11468) );
  AOI22_X1 U14333 ( .A1(n11514), .A2(n11468), .B1(n13202), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14334 ( .A1(n13203), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11469) );
  OAI211_X1 U14335 ( .C1(n13921), .C2(n11812), .A(n11470), .B(n11469), .ZN(
        n13639) );
  XOR2_X1 U14336 ( .A(n11472), .B(n11471), .Z(n15535) );
  AOI22_X1 U14337 ( .A1(n11571), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14338 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14339 ( .A1(n11706), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14340 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11473) );
  NAND4_X1 U14341 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(
        n11482) );
  AOI22_X1 U14342 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14343 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14344 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14345 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11477) );
  NAND4_X1 U14346 ( .A1(n11480), .A2(n11479), .A3(n11478), .A4(n11477), .ZN(
        n11481) );
  OAI21_X1 U14347 ( .B1(n11482), .B2(n11481), .A(n11514), .ZN(n11485) );
  NAND2_X1 U14348 ( .A1(n13203), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11484) );
  NAND2_X1 U14349 ( .A1(n13202), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11483) );
  AND3_X1 U14350 ( .A1(n11485), .A2(n11484), .A3(n11483), .ZN(n11486) );
  OAI21_X1 U14351 ( .B1(n15535), .B2(n11812), .A(n11486), .ZN(n13637) );
  AND2_X1 U14352 ( .A1(n13639), .A2(n13637), .ZN(n11487) );
  NAND2_X1 U14353 ( .A1(n11489), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11505) );
  XNOR2_X1 U14354 ( .A(n11505), .B(n15476), .ZN(n15479) );
  AOI22_X1 U14355 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n9593), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14356 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14357 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14358 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11633), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11490) );
  NAND4_X1 U14359 ( .A1(n11493), .A2(n11492), .A3(n11491), .A4(n11490), .ZN(
        n11499) );
  AOI22_X1 U14360 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14361 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11659), .B1(
        n11576), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14362 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14363 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n9598), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11494) );
  NAND4_X1 U14364 ( .A1(n11497), .A2(n11496), .A3(n11495), .A4(n11494), .ZN(
        n11498) );
  OAI21_X1 U14365 ( .B1(n11499), .B2(n11498), .A(n11514), .ZN(n11502) );
  NAND2_X1 U14366 ( .A1(n13203), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11501) );
  NAND2_X1 U14367 ( .A1(n13202), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11500) );
  NAND3_X1 U14368 ( .A1(n11502), .A2(n11501), .A3(n11500), .ZN(n11503) );
  AOI21_X1 U14369 ( .B1(n15479), .B2(n12878), .A(n11503), .ZN(n13689) );
  INV_X1 U14370 ( .A(n13689), .ZN(n11504) );
  XOR2_X1 U14371 ( .A(n15466), .B(n11522), .Z(n15527) );
  INV_X1 U14372 ( .A(n15527), .ZN(n11521) );
  AOI22_X1 U14373 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14374 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14375 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14376 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11506) );
  NAND4_X1 U14377 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11516) );
  AOI22_X1 U14378 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14379 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14380 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14381 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11510) );
  NAND4_X1 U14382 ( .A1(n11513), .A2(n11512), .A3(n11511), .A4(n11510), .ZN(
        n11515) );
  OAI21_X1 U14383 ( .B1(n11516), .B2(n11515), .A(n11514), .ZN(n11519) );
  NAND2_X1 U14384 ( .A1(n13203), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U14385 ( .A1(n13202), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11517) );
  NAND3_X1 U14386 ( .A1(n11519), .A2(n11518), .A3(n11517), .ZN(n11520) );
  AOI21_X1 U14387 ( .B1(n11521), .B2(n12878), .A(n11520), .ZN(n13762) );
  INV_X1 U14388 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13895) );
  XNOR2_X1 U14389 ( .A(n11536), .B(n13895), .ZN(n13899) );
  AOI21_X1 U14390 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13895), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11523) );
  AOI21_X1 U14391 ( .B1(n13203), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11523), .ZN(
        n11535) );
  AOI22_X1 U14392 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14393 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14394 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14395 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11524) );
  NAND4_X1 U14396 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11533) );
  AOI22_X1 U14397 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14398 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11571), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14399 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14400 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11528) );
  NAND4_X1 U14401 ( .A1(n11531), .A2(n11530), .A3(n11529), .A4(n11528), .ZN(
        n11532) );
  OAI21_X1 U14402 ( .B1(n11533), .B2(n11532), .A(n11836), .ZN(n11534) );
  AOI22_X1 U14403 ( .A1(n13899), .A2(n12878), .B1(n11535), .B2(n11534), .ZN(
        n13619) );
  XOR2_X1 U14404 ( .A(n11554), .B(n11555), .Z(n15519) );
  INV_X1 U14405 ( .A(n15519), .ZN(n11551) );
  AOI22_X1 U14406 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14407 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14408 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14409 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11538) );
  NAND4_X1 U14410 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n11547) );
  AOI22_X1 U14411 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14412 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14413 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14414 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11542) );
  NAND4_X1 U14415 ( .A1(n11545), .A2(n11544), .A3(n11543), .A4(n11542), .ZN(
        n11546) );
  NOR2_X1 U14416 ( .A1(n11547), .A2(n11546), .ZN(n11549) );
  AOI22_X1 U14417 ( .A1(n13203), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13202), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11548) );
  OAI21_X1 U14418 ( .B1(n11809), .B2(n11549), .A(n11548), .ZN(n11550) );
  AOI21_X1 U14419 ( .B1(n11551), .B2(n12878), .A(n11550), .ZN(n13608) );
  XNOR2_X1 U14420 ( .A(n11587), .B(n13600), .ZN(n13884) );
  AOI22_X1 U14421 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14422 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14423 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14424 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11556) );
  NAND4_X1 U14425 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n11565) );
  AOI22_X1 U14426 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14427 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14428 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14429 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U14430 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11564) );
  NOR2_X1 U14431 ( .A1(n11565), .A2(n11564), .ZN(n11568) );
  OAI21_X1 U14432 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n13600), .A(n11812), 
        .ZN(n11566) );
  AOI21_X1 U14433 ( .B1(n13203), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11566), .ZN(
        n11567) );
  OAI21_X1 U14434 ( .B1(n11809), .B2(n11568), .A(n11567), .ZN(n11569) );
  OAI21_X1 U14435 ( .B1(n13884), .B2(n11812), .A(n11569), .ZN(n13590) );
  NOR2_X2 U14436 ( .A1(n13606), .A2(n13590), .ZN(n13678) );
  AOI22_X1 U14437 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14438 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14439 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11571), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14440 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11572) );
  NAND4_X1 U14441 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11582) );
  AOI22_X1 U14442 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14443 ( .A1(n11706), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14444 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14445 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11577) );
  NAND4_X1 U14446 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11581) );
  NOR2_X1 U14447 ( .A1(n11582), .A2(n11581), .ZN(n11586) );
  NAND2_X1 U14448 ( .A1(n11260), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11583) );
  NAND2_X1 U14449 ( .A1(n11812), .A2(n11583), .ZN(n11584) );
  AOI21_X1 U14450 ( .B1(n11278), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11584), .ZN(
        n11585) );
  OAI21_X1 U14451 ( .B1(n11809), .B2(n11586), .A(n11585), .ZN(n11594) );
  INV_X1 U14452 ( .A(n11627), .ZN(n11592) );
  INV_X1 U14453 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11590) );
  INV_X1 U14454 ( .A(n11588), .ZN(n11589) );
  NAND2_X1 U14455 ( .A1(n11590), .A2(n11589), .ZN(n11591) );
  NAND2_X1 U14456 ( .A1(n11592), .A2(n11591), .ZN(n15514) );
  OR2_X1 U14457 ( .A1(n15514), .A2(n11812), .ZN(n11593) );
  AOI22_X1 U14458 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14459 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14460 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14461 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11595) );
  NAND4_X1 U14462 ( .A1(n11598), .A2(n11597), .A3(n11596), .A4(n11595), .ZN(
        n11604) );
  AOI22_X1 U14463 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14464 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14465 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14466 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11599) );
  NAND4_X1 U14467 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11603) );
  NOR2_X1 U14468 ( .A1(n11604), .A2(n11603), .ZN(n11608) );
  NAND2_X1 U14469 ( .A1(n11260), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14470 ( .A1(n11812), .A2(n11605), .ZN(n11606) );
  AOI21_X1 U14471 ( .B1(n11278), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11606), .ZN(
        n11607) );
  OAI21_X1 U14472 ( .B1(n11809), .B2(n11608), .A(n11607), .ZN(n11610) );
  INV_X1 U14473 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13873) );
  XNOR2_X1 U14474 ( .A(n11627), .B(n13873), .ZN(n13875) );
  NAND2_X1 U14475 ( .A1(n13875), .A2(n12878), .ZN(n11609) );
  AOI22_X1 U14476 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14477 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14478 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14479 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11611) );
  NAND4_X1 U14480 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n11622) );
  AOI22_X1 U14481 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14482 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14483 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14484 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14485 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11621) );
  NOR2_X1 U14486 ( .A1(n11622), .A2(n11621), .ZN(n11626) );
  INV_X1 U14487 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20291) );
  OAI21_X1 U14488 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20291), .A(
        n11260), .ZN(n11623) );
  INV_X1 U14489 ( .A(n11623), .ZN(n11624) );
  AOI21_X1 U14490 ( .B1(n11278), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11624), .ZN(
        n11625) );
  OAI21_X1 U14491 ( .B1(n11809), .B2(n11626), .A(n11625), .ZN(n11632) );
  INV_X1 U14492 ( .A(n11628), .ZN(n11629) );
  INV_X1 U14493 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15439) );
  NAND2_X1 U14494 ( .A1(n11629), .A2(n15439), .ZN(n11630) );
  NAND2_X1 U14495 ( .A1(n11650), .A2(n11630), .ZN(n15450) );
  OR2_X1 U14496 ( .A1(n15450), .A2(n11812), .ZN(n11631) );
  NAND2_X1 U14497 ( .A1(n11632), .A2(n11631), .ZN(n13669) );
  AOI22_X1 U14498 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n9593), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14499 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11633), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14500 ( .A1(n11634), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14501 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11635) );
  NAND4_X1 U14502 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11645) );
  AOI22_X1 U14503 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n9598), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14504 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11818), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14505 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11639), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14506 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11640) );
  NAND4_X1 U14507 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n11644) );
  NOR2_X1 U14508 ( .A1(n11645), .A2(n11644), .ZN(n11648) );
  INV_X1 U14509 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20631) );
  AOI21_X1 U14510 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20631), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11646) );
  AOI21_X1 U14511 ( .B1(n11278), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11646), .ZN(
        n11647) );
  OAI21_X1 U14512 ( .B1(n11809), .B2(n11648), .A(n11647), .ZN(n11653) );
  NAND2_X1 U14513 ( .A1(n11650), .A2(n20631), .ZN(n11651) );
  NAND2_X1 U14514 ( .A1(n11682), .A2(n11651), .ZN(n13857) );
  OR2_X1 U14515 ( .A1(n13857), .A2(n11812), .ZN(n11652) );
  NAND2_X1 U14516 ( .A1(n11653), .A2(n11652), .ZN(n13571) );
  INV_X1 U14517 ( .A(n13571), .ZN(n11654) );
  AOI22_X1 U14518 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14519 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14520 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14521 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11655) );
  NAND4_X1 U14522 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11666) );
  AOI22_X1 U14523 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14524 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14525 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14526 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11661) );
  NAND4_X1 U14527 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n11665) );
  NOR2_X1 U14528 ( .A1(n11666), .A2(n11665), .ZN(n11687) );
  AOI22_X1 U14529 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14530 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14531 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14532 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11667) );
  NAND4_X1 U14533 ( .A1(n11670), .A2(n11669), .A3(n11668), .A4(n11667), .ZN(
        n11676) );
  AOI22_X1 U14534 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14535 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14536 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14537 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11671) );
  NAND4_X1 U14538 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11675) );
  NOR2_X1 U14539 ( .A1(n11676), .A2(n11675), .ZN(n11686) );
  XNOR2_X1 U14540 ( .A(n11687), .B(n11686), .ZN(n11680) );
  NAND2_X1 U14541 ( .A1(n11260), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11677) );
  NAND2_X1 U14542 ( .A1(n11812), .A2(n11677), .ZN(n11678) );
  AOI21_X1 U14543 ( .B1(n11278), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11678), .ZN(
        n11679) );
  OAI21_X1 U14544 ( .B1(n11809), .B2(n11680), .A(n11679), .ZN(n11685) );
  INV_X1 U14545 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11681) );
  NAND2_X1 U14546 ( .A1(n11682), .A2(n11681), .ZN(n11683) );
  NAND2_X1 U14547 ( .A1(n11724), .A2(n11683), .ZN(n15427) );
  NAND2_X1 U14548 ( .A1(n11685), .A2(n11684), .ZN(n13664) );
  NOR2_X1 U14549 ( .A1(n11687), .A2(n11686), .ZN(n11719) );
  AOI22_X1 U14550 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11760), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11692) );
  INV_X1 U14551 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n20609) );
  AOI22_X1 U14552 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14553 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14554 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14555 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11698) );
  AOI22_X1 U14556 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14557 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14558 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14559 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14560 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11697) );
  OR2_X1 U14561 ( .A1(n11698), .A2(n11697), .ZN(n11718) );
  INV_X1 U14562 ( .A(n11718), .ZN(n11699) );
  XNOR2_X1 U14563 ( .A(n11719), .B(n11699), .ZN(n11700) );
  NAND2_X1 U14564 ( .A1(n11700), .A2(n11836), .ZN(n11705) );
  NAND2_X1 U14565 ( .A1(n11260), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11701) );
  NAND2_X1 U14566 ( .A1(n11812), .A2(n11701), .ZN(n11702) );
  AOI21_X1 U14567 ( .B1(n11278), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11702), .ZN(
        n11704) );
  XNOR2_X1 U14568 ( .A(n11724), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13845) );
  AOI21_X1 U14569 ( .B1(n11705), .B2(n11704), .A(n11703), .ZN(n13557) );
  AOI22_X1 U14570 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14571 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11706), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14572 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14573 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14574 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11717) );
  AOI22_X1 U14575 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14576 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14577 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14578 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11712) );
  NAND4_X1 U14579 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11716) );
  NOR2_X1 U14580 ( .A1(n11717), .A2(n11716), .ZN(n11731) );
  NAND2_X1 U14581 ( .A1(n11719), .A2(n11718), .ZN(n11730) );
  XNOR2_X1 U14582 ( .A(n11731), .B(n11730), .ZN(n11723) );
  NAND2_X1 U14583 ( .A1(n11260), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11720) );
  NAND2_X1 U14584 ( .A1(n11812), .A2(n11720), .ZN(n11721) );
  AOI21_X1 U14585 ( .B1(n11278), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11721), .ZN(
        n11722) );
  OAI21_X1 U14586 ( .B1(n11723), .B2(n11809), .A(n11722), .ZN(n11729) );
  INV_X1 U14587 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U14588 ( .A1(n11726), .A2(n13832), .ZN(n11727) );
  AND2_X1 U14589 ( .A1(n11750), .A2(n11727), .ZN(n13836) );
  NAND2_X1 U14590 ( .A1(n13836), .A2(n12878), .ZN(n11728) );
  NOR2_X1 U14591 ( .A1(n11731), .A2(n11730), .ZN(n11755) );
  AOI22_X1 U14592 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11760), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14593 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14594 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14595 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11732) );
  NAND4_X1 U14596 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11742) );
  AOI22_X1 U14597 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14598 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14599 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14600 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U14601 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11741) );
  OR2_X1 U14602 ( .A1(n11742), .A2(n11741), .ZN(n11754) );
  INV_X1 U14603 ( .A(n11754), .ZN(n11743) );
  XNOR2_X1 U14604 ( .A(n11755), .B(n11743), .ZN(n11744) );
  NAND2_X1 U14605 ( .A1(n11744), .A2(n11836), .ZN(n11749) );
  NAND2_X1 U14606 ( .A1(n11260), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14607 ( .A1(n11812), .A2(n11745), .ZN(n11746) );
  AOI21_X1 U14608 ( .B1(n11278), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11746), .ZN(
        n11748) );
  XNOR2_X1 U14609 ( .A(n11750), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13824) );
  INV_X1 U14610 ( .A(n11750), .ZN(n11751) );
  NAND2_X1 U14611 ( .A1(n11751), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11752) );
  INV_X1 U14612 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13520) );
  NAND2_X1 U14613 ( .A1(n11752), .A2(n13520), .ZN(n11753) );
  NAND2_X1 U14614 ( .A1(n11789), .A2(n11753), .ZN(n13812) );
  NAND2_X1 U14615 ( .A1(n11755), .A2(n11754), .ZN(n11782) );
  AOI22_X1 U14616 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14617 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14618 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14619 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U14620 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11766) );
  AOI22_X1 U14621 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14622 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14623 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14624 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11761) );
  NAND4_X1 U14625 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11765) );
  NOR2_X1 U14626 ( .A1(n11766), .A2(n11765), .ZN(n11783) );
  XNOR2_X1 U14627 ( .A(n11782), .B(n11783), .ZN(n11769) );
  AOI21_X1 U14628 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n11260), .A(
        n11313), .ZN(n11768) );
  NAND2_X1 U14629 ( .A1(n11278), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11767) );
  OAI211_X1 U14630 ( .C1(n11769), .C2(n11809), .A(n11768), .B(n11767), .ZN(
        n11770) );
  OAI21_X1 U14631 ( .B1(n11812), .B2(n13812), .A(n11770), .ZN(n13519) );
  AOI22_X1 U14632 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11760), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14633 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14634 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U14635 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11771) );
  NAND4_X1 U14636 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11781) );
  AOI22_X1 U14637 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14638 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14639 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14640 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11776) );
  NAND4_X1 U14641 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11780) );
  OR2_X1 U14642 ( .A1(n11781), .A2(n11780), .ZN(n11794) );
  NOR2_X1 U14643 ( .A1(n11783), .A2(n11782), .ZN(n11795) );
  XOR2_X1 U14644 ( .A(n11794), .B(n11795), .Z(n11784) );
  NAND2_X1 U14645 ( .A1(n11784), .A2(n11836), .ZN(n11788) );
  INV_X1 U14646 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13796) );
  AOI21_X1 U14647 ( .B1(n13796), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11785) );
  AOI21_X1 U14648 ( .B1(n13203), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11785), .ZN(
        n11787) );
  INV_X1 U14649 ( .A(n11789), .ZN(n11786) );
  XOR2_X1 U14650 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n11786), .Z(
        n13798) );
  AOI22_X1 U14651 ( .A1(n11788), .A2(n11787), .B1(n12878), .B2(n13798), .ZN(
        n13509) );
  INV_X1 U14652 ( .A(n11790), .ZN(n11792) );
  INV_X1 U14653 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11791) );
  NAND2_X1 U14654 ( .A1(n11792), .A2(n11791), .ZN(n11793) );
  NAND2_X1 U14655 ( .A1(n12881), .A2(n11793), .ZN(n13791) );
  NAND2_X1 U14656 ( .A1(n11795), .A2(n11794), .ZN(n11813) );
  AOI22_X1 U14657 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n9593), .B1(
        n11816), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14658 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11760), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14659 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14660 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U14661 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11806) );
  AOI22_X1 U14662 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11576), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U14663 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11818), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14664 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14665 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11801) );
  NAND4_X1 U14666 ( .A1(n11804), .A2(n11803), .A3(n11802), .A4(n11801), .ZN(
        n11805) );
  NOR2_X1 U14667 ( .A1(n11806), .A2(n11805), .ZN(n11814) );
  XNOR2_X1 U14668 ( .A(n11813), .B(n11814), .ZN(n11810) );
  AOI21_X1 U14669 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n11260), .A(
        n12878), .ZN(n11808) );
  NAND2_X1 U14670 ( .A1(n13203), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11807) );
  OAI211_X1 U14671 ( .C1(n11810), .C2(n11809), .A(n11808), .B(n11807), .ZN(
        n11811) );
  OAI21_X1 U14672 ( .B1(n11812), .B2(n13791), .A(n11811), .ZN(n13498) );
  NOR2_X1 U14673 ( .A1(n11814), .A2(n11813), .ZN(n11835) );
  AOI22_X1 U14674 ( .A1(n11816), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11815), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14675 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14676 ( .A1(n11818), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U14677 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11821) );
  NAND4_X1 U14678 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .ZN(
        n11833) );
  AOI22_X1 U14679 ( .A1(n11639), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14680 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14681 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11826), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14682 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11828) );
  NAND4_X1 U14683 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n11832) );
  NOR2_X1 U14684 ( .A1(n11833), .A2(n11832), .ZN(n11834) );
  XNOR2_X1 U14685 ( .A(n11835), .B(n11834), .ZN(n11837) );
  NAND2_X1 U14686 ( .A1(n11837), .A2(n11836), .ZN(n11840) );
  INV_X1 U14687 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13782) );
  NOR2_X1 U14688 ( .A1(n13782), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11838) );
  AOI211_X1 U14689 ( .C1(n13203), .C2(P1_EAX_REG_30__SCAN_IN), .A(n11838), .B(
        n12878), .ZN(n11839) );
  XNOR2_X1 U14690 ( .A(n12881), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13780) );
  AOI22_X1 U14691 ( .A1(n11840), .A2(n11839), .B1(n13780), .B2(n12878), .ZN(
        n13201) );
  INV_X1 U14692 ( .A(n11870), .ZN(n12404) );
  OAI211_X1 U14693 ( .C1(n12404), .C2(n12443), .A(n12377), .B(n11843), .ZN(
        n11844) );
  NAND2_X1 U14694 ( .A1(n11844), .A2(n12889), .ZN(n11848) );
  AND2_X1 U14695 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  NAND2_X1 U14696 ( .A1(n11848), .A2(n11847), .ZN(n12441) );
  NAND3_X1 U14697 ( .A1(n11849), .A2(n12439), .A3(n12421), .ZN(n11850) );
  OR2_X1 U14698 ( .A1(n12470), .A2(n19871), .ZN(n12442) );
  XNOR2_X1 U14699 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11873) );
  NAND2_X1 U14700 ( .A1(n11874), .A2(n11873), .ZN(n11852) );
  NAND2_X1 U14701 ( .A1(n20163), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11851) );
  NAND2_X1 U14702 ( .A1(n11852), .A2(n11851), .ZN(n11863) );
  XNOR2_X1 U14703 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U14704 ( .A1(n11863), .A2(n11862), .ZN(n11854) );
  NAND2_X1 U14705 ( .A1(n20226), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11853) );
  NAND2_X1 U14706 ( .A1(n11854), .A2(n11853), .ZN(n11861) );
  XNOR2_X1 U14707 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U14708 ( .A1(n11861), .A2(n11860), .ZN(n11856) );
  NAND2_X1 U14709 ( .A1(n20626), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U14710 ( .A1(n11856), .A2(n11855), .ZN(n11894) );
  INV_X1 U14711 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12648) );
  NOR2_X1 U14712 ( .A1(n12648), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11857) );
  OR2_X1 U14713 ( .A1(n11894), .A2(n11857), .ZN(n11859) );
  NAND2_X1 U14714 ( .A1(n11893), .A2(n12270), .ZN(n11906) );
  NAND2_X1 U14715 ( .A1(n12270), .A2(n11879), .ZN(n11904) );
  XNOR2_X1 U14716 ( .A(n11861), .B(n11860), .ZN(n12267) );
  XNOR2_X1 U14717 ( .A(n11863), .B(n11862), .ZN(n12265) );
  INV_X1 U14718 ( .A(n12265), .ZN(n11864) );
  NAND2_X1 U14719 ( .A1(n19887), .A2(n12443), .ZN(n11865) );
  NAND2_X1 U14720 ( .A1(n11865), .A2(n19871), .ZN(n11886) );
  INV_X1 U14721 ( .A(n11886), .ZN(n11866) );
  AOI211_X1 U14722 ( .C1(n11898), .C2(n12265), .A(n11885), .B(n11866), .ZN(
        n11889) );
  INV_X1 U14723 ( .A(n11879), .ZN(n11875) );
  INV_X1 U14724 ( .A(n11874), .ZN(n11867) );
  OAI21_X1 U14725 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20259), .A(
        n11867), .ZN(n11868) );
  NOR2_X1 U14726 ( .A1(n11875), .A2(n11868), .ZN(n11872) );
  INV_X1 U14727 ( .A(n11868), .ZN(n11869) );
  OAI211_X1 U14728 ( .C1(n19855), .C2(n11870), .A(n11869), .B(n11886), .ZN(
        n11871) );
  OAI21_X1 U14729 ( .B1(n11893), .B2(n11872), .A(n11871), .ZN(n11880) );
  INV_X1 U14730 ( .A(n11880), .ZN(n11884) );
  XNOR2_X1 U14731 ( .A(n11874), .B(n11873), .ZN(n12266) );
  NAND2_X1 U14732 ( .A1(n19887), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11877) );
  OAI21_X1 U14733 ( .B1(n19871), .B2(n11875), .A(n11877), .ZN(n11876) );
  AOI21_X1 U14734 ( .B1(n11898), .B2(n12266), .A(n11876), .ZN(n11881) );
  INV_X1 U14735 ( .A(n11881), .ZN(n11883) );
  NAND2_X1 U14736 ( .A1(n11877), .A2(n12889), .ZN(n11878) );
  AOI22_X1 U14737 ( .A1(n12266), .A2(n11895), .B1(n11881), .B2(n11880), .ZN(
        n11882) );
  AOI21_X1 U14738 ( .B1(n11884), .B2(n11883), .A(n11882), .ZN(n11888) );
  INV_X1 U14739 ( .A(n11885), .ZN(n11887) );
  OAI22_X1 U14740 ( .A1(n11889), .A2(n11888), .B1(n11887), .B2(n11886), .ZN(
        n11892) );
  NAND2_X1 U14741 ( .A1(n11890), .A2(n12267), .ZN(n11891) );
  AOI22_X1 U14742 ( .A1(n11893), .A2(n12267), .B1(n11892), .B2(n11891), .ZN(
        n11901) );
  NOR2_X1 U14743 ( .A1(n11898), .A2(n11896), .ZN(n11900) );
  INV_X1 U14744 ( .A(n11896), .ZN(n12268) );
  NAND3_X1 U14745 ( .A1(n11898), .A2(n11897), .A3(n12268), .ZN(n11899) );
  OAI21_X1 U14746 ( .B1(n11901), .B2(n11900), .A(n11899), .ZN(n11902) );
  AOI21_X1 U14747 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20401), .A(
        n11902), .ZN(n11903) );
  NAND2_X1 U14748 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  NOR2_X1 U14749 ( .A1(n11142), .A2(n19610), .ZN(n11909) );
  NOR2_X1 U14750 ( .A1(n12429), .A2(n12469), .ZN(n11908) );
  NAND4_X1 U14751 ( .A1(n12634), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n12463) );
  OR2_X1 U14752 ( .A1(n12463), .A2(n13471), .ZN(n11910) );
  INV_X1 U14753 ( .A(n11921), .ZN(n11985) );
  NAND2_X2 U14754 ( .A1(n11985), .A2(n13469), .ZN(n12006) );
  OR2_X1 U14755 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11913) );
  INV_X1 U14756 ( .A(n11914), .ZN(n11946) );
  INV_X1 U14757 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11915) );
  OR2_X1 U14758 ( .A1(n11933), .A2(n11915), .ZN(n11917) );
  INV_X1 U14759 ( .A(n11918), .ZN(n12013) );
  NAND2_X1 U14760 ( .A1(n12013), .A2(n11915), .ZN(n11916) );
  NAND2_X1 U14761 ( .A1(n11917), .A2(n11916), .ZN(n12433) );
  MUX2_X1 U14762 ( .A(n12006), .B(n13469), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11920) );
  OR2_X1 U14763 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11919) );
  AND2_X1 U14764 ( .A1(n11920), .A2(n11919), .ZN(n12611) );
  INV_X1 U14765 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19828) );
  NAND2_X1 U14766 ( .A1(n11933), .A2(n19828), .ZN(n11924) );
  INV_X1 U14767 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n11922) );
  NAND2_X1 U14768 ( .A1(n11985), .A2(n11922), .ZN(n11923) );
  NAND3_X1 U14769 ( .A1(n11924), .A2(n11923), .A3(n13469), .ZN(n11925) );
  OAI21_X1 U14770 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(n12012), .A(n11925), .ZN(
        n12618) );
  NAND2_X1 U14771 ( .A1(n12619), .A2(n12618), .ZN(n19690) );
  OR2_X1 U14772 ( .A1(n12006), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U14773 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11926) );
  OAI211_X1 U14774 ( .C1(n13471), .C2(P1_EBX_REG_4__SCAN_IN), .A(n11933), .B(
        n11926), .ZN(n11927) );
  NAND2_X1 U14775 ( .A1(n11928), .A2(n11927), .ZN(n19689) );
  OR2_X1 U14776 ( .A1(n12006), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n11931) );
  NAND2_X1 U14777 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11929) );
  OAI211_X1 U14778 ( .C1(n13471), .C2(P1_EBX_REG_6__SCAN_IN), .A(n11933), .B(
        n11929), .ZN(n11930) );
  AND2_X1 U14779 ( .A1(n11931), .A2(n11930), .ZN(n15639) );
  NAND2_X1 U14780 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U14781 ( .A1(n11933), .A2(n11932), .ZN(n11935) );
  OR2_X1 U14782 ( .A1(n13471), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U14783 ( .A1(n11935), .A2(n11934), .ZN(n11936) );
  OAI21_X1 U14784 ( .B1(n12012), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11936), .ZN(
        n15640) );
  NAND2_X1 U14785 ( .A1(n15639), .A2(n15640), .ZN(n11937) );
  OR2_X1 U14786 ( .A1(n12006), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n11940) );
  NAND2_X1 U14787 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11938) );
  OAI211_X1 U14788 ( .C1(n13471), .C2(P1_EBX_REG_8__SCAN_IN), .A(n11933), .B(
        n11938), .ZN(n11939) );
  AND2_X1 U14789 ( .A1(n11940), .A2(n11939), .ZN(n13064) );
  NAND2_X1 U14790 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U14791 ( .A1(n11933), .A2(n11941), .ZN(n11943) );
  OR2_X1 U14792 ( .A1(n13471), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U14793 ( .A1(n11943), .A2(n11942), .ZN(n11944) );
  OAI21_X1 U14794 ( .B1(n12012), .B2(P1_EBX_REG_7__SCAN_IN), .A(n11944), .ZN(
        n13065) );
  AND2_X1 U14795 ( .A1(n13064), .A2(n13065), .ZN(n11945) );
  AND2_X2 U14796 ( .A1(n15642), .A2(n11945), .ZN(n13093) );
  NAND2_X1 U14797 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11947) );
  NAND2_X1 U14798 ( .A1(n11933), .A2(n11947), .ZN(n11949) );
  OR2_X1 U14799 ( .A1(n13471), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14800 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  OAI21_X1 U14801 ( .B1(n12012), .B2(P1_EBX_REG_9__SCAN_IN), .A(n11950), .ZN(
        n13092) );
  NAND2_X1 U14802 ( .A1(n13093), .A2(n13092), .ZN(n13152) );
  MUX2_X1 U14803 ( .A(n12006), .B(n13469), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11952) );
  OR2_X1 U14804 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U14805 ( .A1(n11952), .A2(n11951), .ZN(n13153) );
  INV_X1 U14806 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15498) );
  NAND2_X1 U14807 ( .A1(n11998), .A2(n15498), .ZN(n11956) );
  INV_X1 U14808 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14097) );
  NAND2_X1 U14809 ( .A1(n11933), .A2(n14097), .ZN(n11954) );
  NAND2_X1 U14810 ( .A1(n11985), .A2(n15498), .ZN(n11953) );
  NAND3_X1 U14811 ( .A1(n11954), .A2(n11953), .A3(n13469), .ZN(n11955) );
  OR2_X1 U14812 ( .A1(n12006), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U14813 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11957) );
  OAI211_X1 U14814 ( .C1(n13471), .C2(P1_EBX_REG_12__SCAN_IN), .A(n11933), .B(
        n11957), .ZN(n11958) );
  NAND2_X1 U14815 ( .A1(n11959), .A2(n11958), .ZN(n15487) );
  NAND2_X1 U14816 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11960) );
  NAND2_X1 U14817 ( .A1(n11933), .A2(n11960), .ZN(n11962) );
  OR2_X1 U14818 ( .A1(n13471), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U14819 ( .A1(n11962), .A2(n11961), .ZN(n11963) );
  OAI21_X1 U14820 ( .B1(n12012), .B2(P1_EBX_REG_13__SCAN_IN), .A(n11963), .ZN(
        n13645) );
  OR2_X1 U14821 ( .A1(n12006), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U14822 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11964) );
  OAI211_X1 U14823 ( .C1(n13471), .C2(P1_EBX_REG_14__SCAN_IN), .A(n11933), .B(
        n11964), .ZN(n11965) );
  NAND2_X1 U14824 ( .A1(n11966), .A2(n11965), .ZN(n13693) );
  MUX2_X1 U14825 ( .A(n12006), .B(n13469), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11968) );
  OR2_X1 U14826 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11967) );
  AND2_X1 U14827 ( .A1(n11968), .A2(n11967), .ZN(n13620) );
  INV_X1 U14828 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U14829 ( .A1(n11998), .A2(n15507), .ZN(n11972) );
  INV_X1 U14830 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13192) );
  NAND2_X1 U14831 ( .A1(n11933), .A2(n13192), .ZN(n11970) );
  NAND2_X1 U14832 ( .A1(n11985), .A2(n15507), .ZN(n11969) );
  NAND3_X1 U14833 ( .A1(n11970), .A2(n11969), .A3(n13469), .ZN(n11971) );
  NAND2_X1 U14834 ( .A1(n11972), .A2(n11971), .ZN(n15471) );
  NAND2_X1 U14835 ( .A1(n13620), .A2(n15471), .ZN(n11973) );
  MUX2_X1 U14836 ( .A(n12006), .B(n13469), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n11975) );
  OR2_X1 U14837 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11974) );
  NAND2_X1 U14838 ( .A1(n11975), .A2(n11974), .ZN(n13592) );
  INV_X1 U14839 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n13612) );
  NAND2_X1 U14840 ( .A1(n11998), .A2(n13612), .ZN(n11978) );
  INV_X1 U14841 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15574) );
  NAND2_X1 U14842 ( .A1(n11933), .A2(n15574), .ZN(n11976) );
  OAI211_X1 U14843 ( .C1(n13471), .C2(P1_EBX_REG_17__SCAN_IN), .A(n11976), .B(
        n13469), .ZN(n11977) );
  AND2_X1 U14844 ( .A1(n11978), .A2(n11977), .ZN(n13591) );
  INV_X1 U14845 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14054) );
  NAND2_X1 U14846 ( .A1(n11933), .A2(n14054), .ZN(n11980) );
  INV_X1 U14847 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U14848 ( .A1(n11985), .A2(n15459), .ZN(n11979) );
  NAND3_X1 U14849 ( .A1(n11980), .A2(n11979), .A3(n13469), .ZN(n11981) );
  OAI21_X1 U14850 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(n12012), .A(n11981), .ZN(
        n13681) );
  OR2_X1 U14851 ( .A1(n12006), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U14852 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11982) );
  OAI211_X1 U14853 ( .C1(n13471), .C2(P1_EBX_REG_20__SCAN_IN), .A(n11933), .B(
        n11982), .ZN(n11983) );
  NAND2_X1 U14854 ( .A1(n11984), .A2(n11983), .ZN(n13583) );
  INV_X1 U14855 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15440) );
  NAND2_X1 U14856 ( .A1(n11998), .A2(n15440), .ZN(n11989) );
  INV_X1 U14857 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14041) );
  NAND2_X1 U14858 ( .A1(n11933), .A2(n14041), .ZN(n11987) );
  NAND2_X1 U14859 ( .A1(n11985), .A2(n15440), .ZN(n11986) );
  NAND3_X1 U14860 ( .A1(n11987), .A2(n11986), .A3(n13469), .ZN(n11988) );
  AND2_X1 U14861 ( .A1(n11989), .A2(n11988), .ZN(n13670) );
  MUX2_X1 U14862 ( .A(n12006), .B(n13469), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11991) );
  OR2_X1 U14863 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11990) );
  NAND2_X1 U14864 ( .A1(n11991), .A2(n11990), .ZN(n13572) );
  NAND2_X1 U14865 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11992) );
  NAND2_X1 U14866 ( .A1(n11933), .A2(n11992), .ZN(n11994) );
  OR2_X1 U14867 ( .A1(n13471), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n11993) );
  NAND2_X1 U14868 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  OAI21_X1 U14869 ( .B1(n12012), .B2(P1_EBX_REG_23__SCAN_IN), .A(n11995), .ZN(
        n13660) );
  NAND2_X1 U14870 ( .A1(n13661), .A2(n13660), .ZN(n13663) );
  MUX2_X1 U14871 ( .A(n12006), .B(n13469), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11997) );
  OR2_X1 U14872 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11996) );
  NAND2_X1 U14873 ( .A1(n11997), .A2(n11996), .ZN(n13559) );
  INV_X1 U14874 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U14875 ( .A1(n11998), .A2(n13658), .ZN(n12001) );
  INV_X1 U14876 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14004) );
  NAND2_X1 U14877 ( .A1(n11933), .A2(n14004), .ZN(n11999) );
  OAI211_X1 U14878 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n13471), .A(n11999), .B(
        n13469), .ZN(n12000) );
  MUX2_X1 U14879 ( .A(n12006), .B(n13469), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12003) );
  OR2_X1 U14880 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12002) );
  AND2_X1 U14881 ( .A1(n12003), .A2(n12002), .ZN(n13533) );
  INV_X1 U14882 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13990) );
  NAND2_X1 U14883 ( .A1(n11933), .A2(n13990), .ZN(n12004) );
  OAI211_X1 U14884 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n13471), .A(n12004), .B(
        n13469), .ZN(n12005) );
  OAI21_X1 U14885 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(n12012), .A(n12005), .ZN(
        n13523) );
  OR2_X1 U14886 ( .A1(n12006), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12009) );
  NAND2_X1 U14887 ( .A1(n13469), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12007) );
  OAI211_X1 U14888 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n13471), .A(n11933), .B(
        n12007), .ZN(n12008) );
  AND2_X1 U14889 ( .A1(n12009), .A2(n12008), .ZN(n13510) );
  OR2_X1 U14890 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12011) );
  OR2_X1 U14891 ( .A1(n13471), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12010) );
  NAND2_X1 U14892 ( .A1(n12011), .A2(n12010), .ZN(n12015) );
  OAI22_X1 U14893 ( .A1(n12015), .A2(n12013), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12012), .ZN(n13497) );
  NAND2_X1 U14894 ( .A1(n13512), .A2(n13497), .ZN(n13468) );
  NAND2_X1 U14895 ( .A1(n13468), .A2(n12013), .ZN(n12016) );
  INV_X1 U14896 ( .A(n13512), .ZN(n12014) );
  AOI22_X1 U14897 ( .A1(n12016), .A2(n12015), .B1(n12014), .B2(n13469), .ZN(
        n12017) );
  AOI22_X1 U14898 ( .A1(n13472), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13471), .ZN(n13470) );
  XNOR2_X1 U14899 ( .A(n12017), .B(n13470), .ZN(n13962) );
  INV_X1 U14900 ( .A(n12469), .ZN(n19895) );
  INV_X1 U14901 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13494) );
  NOR2_X1 U14902 ( .A1(n19728), .A2(n13494), .ZN(n12018) );
  AOI21_X1 U14903 ( .B1(n13962), .B2(n19725), .A(n12018), .ZN(n12019) );
  AND2_X1 U14904 ( .A1(n12021), .A2(n12022), .ZN(n15946) );
  NAND2_X1 U14905 ( .A1(n15943), .A2(n15946), .ZN(n13039) );
  INV_X1 U14906 ( .A(n14916), .ZN(n12819) );
  NAND2_X1 U14907 ( .A1(n13039), .A2(n12819), .ZN(n12023) );
  INV_X1 U14908 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15787) );
  OR2_X1 U14909 ( .A1(n13398), .A2(n15787), .ZN(n12032) );
  INV_X1 U14910 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12029) );
  INV_X1 U14911 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12026) );
  OR2_X1 U14912 ( .A1(n12119), .A2(n12026), .ZN(n12028) );
  NAND2_X1 U14913 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12027) );
  OAI211_X1 U14914 ( .C1(n12126), .C2(n12029), .A(n12028), .B(n12027), .ZN(
        n12030) );
  INV_X1 U14915 ( .A(n12030), .ZN(n12031) );
  NAND2_X1 U14916 ( .A1(n12032), .A2(n12031), .ZN(n12848) );
  INV_X1 U14917 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14849) );
  OR2_X1 U14918 ( .A1(n13398), .A2(n14849), .ZN(n12037) );
  NAND2_X1 U14919 ( .A1(n12025), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U14920 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12033) );
  OAI211_X1 U14921 ( .C1(n9978), .C2(n12119), .A(n12034), .B(n12033), .ZN(
        n12035) );
  INV_X1 U14922 ( .A(n12035), .ZN(n12036) );
  INV_X1 U14923 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15899) );
  OR2_X1 U14924 ( .A1(n13398), .A2(n15899), .ZN(n12042) );
  INV_X1 U14925 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18650) );
  NAND2_X1 U14926 ( .A1(n12025), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12039) );
  NAND2_X1 U14927 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12038) );
  OAI211_X1 U14928 ( .C1(n18650), .C2(n12119), .A(n12039), .B(n12038), .ZN(
        n12040) );
  INV_X1 U14929 ( .A(n12040), .ZN(n12041) );
  NAND2_X1 U14930 ( .A1(n12042), .A2(n12041), .ZN(n12527) );
  INV_X1 U14931 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12045) );
  NAND2_X1 U14932 ( .A1(n12124), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12044) );
  AOI22_X1 U14933 ( .A1(n12025), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12043) );
  OAI211_X1 U14934 ( .C1(n12045), .C2(n12119), .A(n12044), .B(n12043), .ZN(
        n12046) );
  INV_X1 U14935 ( .A(n12046), .ZN(n12477) );
  INV_X1 U14936 ( .A(n12048), .ZN(n12049) );
  INV_X1 U14937 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12948) );
  INV_X1 U14938 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14894) );
  OR2_X1 U14939 ( .A1(n13398), .A2(n14894), .ZN(n12052) );
  AOI22_X1 U14940 ( .A1(n12025), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12051) );
  OAI211_X1 U14941 ( .C1(n12948), .C2(n12119), .A(n12052), .B(n12051), .ZN(
        n13432) );
  NAND2_X1 U14942 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  INV_X1 U14943 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12950) );
  OR2_X1 U14944 ( .A1(n13398), .A2(n15911), .ZN(n12054) );
  AOI22_X1 U14945 ( .A1(n12025), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12053) );
  OAI211_X1 U14946 ( .C1(n12950), .C2(n12119), .A(n12054), .B(n12053), .ZN(
        n12533) );
  INV_X1 U14947 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12980) );
  OR2_X1 U14948 ( .A1(n13398), .A2(n15900), .ZN(n12056) );
  AOI22_X1 U14949 ( .A1(n12025), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12055) );
  OAI211_X1 U14950 ( .C1(n12980), .C2(n12119), .A(n12056), .B(n12055), .ZN(
        n12555) );
  INV_X1 U14951 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12059) );
  INV_X1 U14952 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14831) );
  OR2_X1 U14953 ( .A1(n13398), .A2(n14831), .ZN(n12058) );
  AOI22_X1 U14954 ( .A1(n12025), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12057) );
  OAI211_X1 U14955 ( .C1(n12119), .C2(n12059), .A(n12058), .B(n12057), .ZN(
        n12865) );
  INV_X1 U14956 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12062) );
  INV_X1 U14957 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12967) );
  OR2_X1 U14958 ( .A1(n12119), .A2(n12967), .ZN(n12061) );
  NAND2_X1 U14959 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12060) );
  OAI211_X1 U14960 ( .C1(n12126), .C2(n12062), .A(n12061), .B(n12060), .ZN(
        n12063) );
  AOI21_X1 U14961 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12063), .ZN(n12859) );
  INV_X1 U14962 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12067) );
  INV_X1 U14963 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12064) );
  OR2_X1 U14964 ( .A1(n12119), .A2(n12064), .ZN(n12066) );
  NAND2_X1 U14965 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12065) );
  OAI211_X1 U14966 ( .C1(n12126), .C2(n12067), .A(n12066), .B(n12065), .ZN(
        n12068) );
  AOI21_X1 U14967 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12068), .ZN(n12988) );
  INV_X1 U14968 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13024) );
  INV_X1 U14969 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15870) );
  OR2_X1 U14970 ( .A1(n13398), .A2(n15870), .ZN(n12070) );
  AOI22_X1 U14971 ( .A1(n12025), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12069) );
  OAI211_X1 U14972 ( .C1(n12119), .C2(n13024), .A(n12070), .B(n12069), .ZN(
        n13014) );
  INV_X1 U14973 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n12074) );
  INV_X1 U14974 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12071) );
  OR2_X1 U14975 ( .A1(n12119), .A2(n12071), .ZN(n12073) );
  NAND2_X1 U14976 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12072) );
  OAI211_X1 U14977 ( .C1(n12126), .C2(n12074), .A(n12073), .B(n12072), .ZN(
        n12075) );
  AOI21_X1 U14978 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12075), .ZN(n13084) );
  INV_X1 U14979 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n12078) );
  OR2_X1 U14980 ( .A1(n12119), .A2(n9804), .ZN(n12077) );
  NAND2_X1 U14981 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12076) );
  OAI211_X1 U14982 ( .C1(n12126), .C2(n12078), .A(n12077), .B(n12076), .ZN(
        n12079) );
  AOI21_X1 U14983 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12079), .ZN(n14347) );
  NOR2_X2 U14984 ( .A1(n14346), .A2(n14347), .ZN(n14345) );
  INV_X1 U14985 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12082) );
  INV_X1 U14986 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14553) );
  OR2_X1 U14987 ( .A1(n13398), .A2(n14553), .ZN(n12081) );
  AOI22_X1 U14988 ( .A1(n12025), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12080) );
  OAI211_X1 U14989 ( .C1(n12119), .C2(n12082), .A(n12081), .B(n12080), .ZN(
        n14336) );
  INV_X1 U14990 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14332) );
  INV_X1 U14991 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14773) );
  OR2_X1 U14992 ( .A1(n13398), .A2(n14773), .ZN(n12084) );
  AOI22_X1 U14993 ( .A1(n12025), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12083) );
  OAI211_X1 U14994 ( .C1(n12119), .C2(n14332), .A(n12084), .B(n12083), .ZN(
        n14327) );
  INV_X1 U14995 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n12088) );
  INV_X1 U14996 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12085) );
  OR2_X1 U14997 ( .A1(n12119), .A2(n12085), .ZN(n12087) );
  NAND2_X1 U14998 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12086) );
  OAI211_X1 U14999 ( .C1(n12126), .C2(n12088), .A(n12087), .B(n12086), .ZN(
        n12089) );
  AOI21_X1 U15000 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12089), .ZN(n14318) );
  INV_X1 U15001 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19515) );
  INV_X1 U15002 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12090) );
  OR2_X1 U15003 ( .A1(n12119), .A2(n12090), .ZN(n12092) );
  NAND2_X1 U15004 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12091) );
  OAI211_X1 U15005 ( .C1(n12126), .C2(n19515), .A(n12092), .B(n12091), .ZN(
        n12093) );
  AOI21_X1 U15006 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12093), .ZN(n14226) );
  INV_X1 U15007 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14311) );
  INV_X1 U15008 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14618) );
  OR2_X1 U15009 ( .A1(n13398), .A2(n14618), .ZN(n12095) );
  AOI22_X1 U15010 ( .A1(n12025), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12094) );
  OAI211_X1 U15011 ( .C1(n12119), .C2(n14311), .A(n12095), .B(n12094), .ZN(
        n14309) );
  INV_X1 U15012 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12099) );
  INV_X1 U15013 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12096) );
  OR2_X1 U15014 ( .A1(n12119), .A2(n12096), .ZN(n12098) );
  NAND2_X1 U15015 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12097) );
  OAI211_X1 U15016 ( .C1(n12126), .C2(n12099), .A(n12098), .B(n12097), .ZN(
        n12100) );
  AOI21_X1 U15017 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12100), .ZN(n14297) );
  INV_X1 U15018 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n12104) );
  INV_X1 U15019 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12101) );
  OR2_X1 U15020 ( .A1(n12119), .A2(n12101), .ZN(n12103) );
  NAND2_X1 U15021 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12102) );
  OAI211_X1 U15022 ( .C1(n12126), .C2(n12104), .A(n12103), .B(n12102), .ZN(
        n12105) );
  AOI21_X1 U15023 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12105), .ZN(n14293) );
  INV_X1 U15024 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n12108) );
  OR2_X1 U15025 ( .A1(n12119), .A2(n9974), .ZN(n12107) );
  NAND2_X1 U15026 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12106) );
  OAI211_X1 U15027 ( .C1(n12126), .C2(n12108), .A(n12107), .B(n12106), .ZN(
        n12109) );
  AOI21_X1 U15028 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12109), .ZN(n14281) );
  INV_X1 U15029 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n20558) );
  INV_X1 U15030 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14697) );
  OR2_X1 U15031 ( .A1(n13398), .A2(n14697), .ZN(n12111) );
  AOI22_X1 U15032 ( .A1(n12025), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12110) );
  OAI211_X1 U15033 ( .C1(n12119), .C2(n20558), .A(n12111), .B(n12110), .ZN(
        n14279) );
  INV_X1 U15034 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12114) );
  INV_X1 U15035 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14690) );
  OR2_X1 U15036 ( .A1(n13398), .A2(n14690), .ZN(n12113) );
  AOI22_X1 U15037 ( .A1(n12025), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12112) );
  OAI211_X1 U15038 ( .C1(n12119), .C2(n12114), .A(n12113), .B(n12112), .ZN(
        n14266) );
  INV_X1 U15039 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12117) );
  INV_X1 U15040 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14674) );
  OR2_X1 U15041 ( .A1(n13398), .A2(n14674), .ZN(n12116) );
  AOI22_X1 U15042 ( .A1(n12025), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12115) );
  OAI211_X1 U15043 ( .C1(n12119), .C2(n12117), .A(n12116), .B(n12115), .ZN(
        n14209) );
  INV_X1 U15044 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12122) );
  INV_X1 U15045 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12118) );
  OR2_X1 U15046 ( .A1(n12119), .A2(n12118), .ZN(n12121) );
  NAND2_X1 U15047 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12120) );
  OAI211_X1 U15048 ( .C1(n12126), .C2(n12122), .A(n12121), .B(n12120), .ZN(
        n12123) );
  AOI21_X1 U15049 ( .B1(n12124), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12123), .ZN(n14194) );
  INV_X1 U15050 ( .A(n12125), .ZN(n13395) );
  INV_X1 U15051 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19529) );
  INV_X1 U15052 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14446) );
  OAI22_X1 U15053 ( .A1(n12126), .A2(n19529), .B1(n20564), .B2(n14446), .ZN(
        n12128) );
  INV_X1 U15054 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14652) );
  NOR2_X1 U15055 ( .A1(n13398), .A2(n14652), .ZN(n12127) );
  AOI211_X1 U15056 ( .C1(n13395), .C2(P2_EBX_REG_29__SCAN_IN), .A(n12128), .B(
        n12127), .ZN(n14182) );
  INV_X1 U15057 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14612) );
  AOI22_X1 U15058 ( .A1(n12025), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12130) );
  NAND2_X1 U15059 ( .A1(n13395), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12129) );
  OAI211_X1 U15060 ( .C1(n13398), .C2(n14612), .A(n12130), .B(n12129), .ZN(
        n12131) );
  NAND2_X1 U15061 ( .A1(n14181), .A2(n12131), .ZN(n13400) );
  INV_X2 U15062 ( .A(n14350), .ZN(n14340) );
  NAND2_X1 U15063 ( .A1(n14340), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U15064 ( .A1(n12134), .A2(n10161), .ZN(P2_U2857) );
  NOR2_X1 U15065 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12136) );
  NOR4_X1 U15066 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12135) );
  NAND4_X1 U15067 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12136), .A4(n12135), .ZN(n12149) );
  NOR4_X1 U15068 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12140) );
  NOR4_X1 U15069 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12139) );
  NOR4_X1 U15070 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12138) );
  NOR4_X1 U15071 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12137) );
  AND4_X1 U15072 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12145) );
  NOR4_X1 U15073 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12143) );
  NOR4_X1 U15074 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12142) );
  NOR4_X1 U15075 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12141) );
  INV_X1 U15076 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20425) );
  AND4_X1 U15077 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n20425), .ZN(
        n12144) );
  NAND2_X1 U15078 ( .A1(n12145), .A2(n12144), .ZN(n12146) );
  INV_X1 U15079 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20486) );
  NOR3_X1 U15080 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20486), .ZN(n12148) );
  NOR4_X1 U15081 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15082 ( .A1(n19852), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12148), .A4(
        n12147), .ZN(U214) );
  NOR2_X1 U15083 ( .A1(n18859), .A2(n12149), .ZN(n16051) );
  NAND2_X1 U15084 ( .A1(n16051), .A2(U214), .ZN(U212) );
  INV_X1 U15085 ( .A(n10815), .ZN(n15171) );
  AND2_X1 U15086 ( .A1(n15171), .A2(n12928), .ZN(n18691) );
  INV_X1 U15087 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12150) );
  INV_X1 U15088 ( .A(n12173), .ZN(n12933) );
  NAND2_X1 U15089 ( .A1(n19355), .A2(n20564), .ZN(n12151) );
  OAI211_X1 U15090 ( .C1(n18691), .C2(n12150), .A(n12933), .B(n12151), .ZN(
        P2_U2814) );
  NOR2_X1 U15091 ( .A1(n19600), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12152)
         );
  INV_X1 U15092 ( .A(n10832), .ZN(n19594) );
  AOI22_X1 U15093 ( .A1(n12152), .A2(n12151), .B1(n19594), .B2(n19600), .ZN(
        P2_U3612) );
  INV_X1 U15094 ( .A(n15945), .ZN(n12154) );
  INV_X1 U15095 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18493) );
  NOR2_X1 U15096 ( .A1(n18493), .A2(n19485), .ZN(n19478) );
  NOR2_X1 U15097 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19468) );
  NOR3_X1 U15098 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19478), .A3(n19468), 
        .ZN(n19591) );
  NAND2_X1 U15099 ( .A1(n19602), .A2(n19591), .ZN(n13043) );
  INV_X1 U15100 ( .A(n13043), .ZN(n12783) );
  AND2_X1 U15101 ( .A1(n10832), .A2(n19602), .ZN(n12153) );
  INV_X1 U15102 ( .A(n12790), .ZN(n15944) );
  NOR4_X1 U15103 ( .A1(n12154), .A2(n12783), .A3(n12153), .A4(n15944), .ZN(
        n15952) );
  NOR2_X1 U15104 ( .A1(n15952), .A2(n19458), .ZN(n19581) );
  INV_X1 U15105 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13048) );
  INV_X1 U15106 ( .A(n12155), .ZN(n12156) );
  AND2_X1 U15107 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  NOR2_X1 U15108 ( .A1(n12243), .A2(n12159), .ZN(n12162) );
  OAI21_X1 U15109 ( .B1(n12162), .B2(n12161), .A(n12160), .ZN(n19585) );
  INV_X1 U15110 ( .A(n15941), .ZN(n12169) );
  NAND2_X1 U15111 ( .A1(n12169), .A2(n12163), .ZN(n12833) );
  OR2_X1 U15112 ( .A1(n19585), .A2(n12833), .ZN(n12171) );
  NAND2_X1 U15113 ( .A1(n15174), .A2(n12164), .ZN(n15940) );
  OAI21_X1 U15114 ( .B1(n10870), .B2(n15940), .A(n13048), .ZN(n12165) );
  AND2_X1 U15115 ( .A1(n12165), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19575) );
  OAI211_X1 U15116 ( .C1(n12201), .C2(n12166), .A(n20564), .B(n12790), .ZN(
        n12167) );
  INV_X1 U15117 ( .A(n12167), .ZN(n12168) );
  NAND3_X1 U15118 ( .A1(n12169), .A2(n19592), .A3(n15961), .ZN(n12170) );
  NAND2_X1 U15119 ( .A1(n12171), .A2(n12170), .ZN(n12793) );
  NOR2_X1 U15120 ( .A1(n18868), .A2(n19458), .ZN(n12172) );
  OAI21_X1 U15121 ( .B1(n19581), .B2(n13048), .A(n12214), .ZN(P2_U2819) );
  AND2_X1 U15122 ( .A1(n12173), .A2(n19602), .ZN(n12174) );
  NOR2_X2 U15123 ( .A1(n12310), .A2(n12174), .ZN(n12220) );
  AOI22_X1 U15124 ( .A1(n12220), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12179) );
  INV_X1 U15125 ( .A(n12174), .ZN(n12175) );
  NOR2_X2 U15126 ( .A1(n12175), .A2(n13275), .ZN(n12320) );
  INV_X1 U15127 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12176) );
  OR2_X1 U15128 ( .A1(n18859), .A2(n12176), .ZN(n12178) );
  NAND2_X1 U15129 ( .A1(n18859), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12177) );
  AND2_X1 U15130 ( .A1(n12178), .A2(n12177), .ZN(n18720) );
  INV_X1 U15131 ( .A(n18720), .ZN(n14364) );
  NAND2_X1 U15132 ( .A1(n12320), .A2(n14364), .ZN(n12300) );
  NAND2_X1 U15133 ( .A1(n12179), .A2(n12300), .ZN(P2_U2978) );
  AOI22_X1 U15134 ( .A1(n12220), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12184) );
  INV_X1 U15135 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n12180) );
  OR2_X1 U15136 ( .A1(n18859), .A2(n12180), .ZN(n12182) );
  NAND2_X1 U15137 ( .A1(n18859), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12181) );
  AND2_X1 U15138 ( .A1(n12182), .A2(n12181), .ZN(n18714) );
  INV_X1 U15139 ( .A(n18714), .ZN(n12183) );
  NAND2_X1 U15140 ( .A1(n12320), .A2(n12183), .ZN(n12189) );
  NAND2_X1 U15141 ( .A1(n12184), .A2(n12189), .ZN(P2_U2980) );
  AOI22_X1 U15142 ( .A1(n12220), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12188) );
  INV_X1 U15143 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12185) );
  OR2_X1 U15144 ( .A1(n18859), .A2(n12185), .ZN(n12187) );
  NAND2_X1 U15145 ( .A1(n18859), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12186) );
  AND2_X1 U15146 ( .A1(n12187), .A2(n12186), .ZN(n18725) );
  INV_X1 U15147 ( .A(n18725), .ZN(n14381) );
  NAND2_X1 U15148 ( .A1(n12320), .A2(n14381), .ZN(n12296) );
  NAND2_X1 U15149 ( .A1(n12188), .A2(n12296), .ZN(P2_U2976) );
  AOI22_X1 U15150 ( .A1(n12220), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n12310), .ZN(n12190) );
  NAND2_X1 U15151 ( .A1(n12190), .A2(n12189), .ZN(P2_U2965) );
  AOI22_X1 U15152 ( .A1(n12220), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12191) );
  OAI22_X1 U15153 ( .A1(n18859), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n18861), .ZN(n18891) );
  INV_X1 U15154 ( .A(n18891), .ZN(n15720) );
  NAND2_X1 U15155 ( .A1(n12320), .A2(n15720), .ZN(n12298) );
  NAND2_X1 U15156 ( .A1(n12191), .A2(n12298), .ZN(P2_U2971) );
  AOI22_X1 U15157 ( .A1(n12220), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12192) );
  OAI22_X1 U15158 ( .A1(n18859), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n18861), .ZN(n18882) );
  INV_X1 U15159 ( .A(n18882), .ZN(n18748) );
  NAND2_X1 U15160 ( .A1(n12320), .A2(n18748), .ZN(n12308) );
  NAND2_X1 U15161 ( .A1(n12192), .A2(n12308), .ZN(P2_U2969) );
  AOI22_X1 U15162 ( .A1(n12220), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15163 ( .A1(n18861), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n18859), .ZN(n18887) );
  INV_X1 U15164 ( .A(n18887), .ZN(n14418) );
  NAND2_X1 U15165 ( .A1(n12320), .A2(n14418), .ZN(n12311) );
  NAND2_X1 U15166 ( .A1(n12193), .A2(n12311), .ZN(P2_U2970) );
  AOI22_X1 U15167 ( .A1(n12220), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15168 ( .A1(n18861), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18859), .ZN(n18911) );
  INV_X1 U15169 ( .A(n18911), .ZN(n14399) );
  NAND2_X1 U15170 ( .A1(n12320), .A2(n14399), .ZN(n12304) );
  NAND2_X1 U15171 ( .A1(n12194), .A2(n12304), .ZN(P2_U2974) );
  AOI22_X1 U15172 ( .A1(n12220), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12195) );
  OAI22_X1 U15173 ( .A1(n18859), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n18861), .ZN(n18902) );
  INV_X1 U15174 ( .A(n18902), .ZN(n15713) );
  NAND2_X1 U15175 ( .A1(n12320), .A2(n15713), .ZN(n12294) );
  NAND2_X1 U15176 ( .A1(n12195), .A2(n12294), .ZN(P2_U2973) );
  AOI22_X1 U15177 ( .A1(n12220), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15178 ( .A1(n18861), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n18859), .ZN(n18897) );
  INV_X1 U15179 ( .A(n18897), .ZN(n14409) );
  NAND2_X1 U15180 ( .A1(n12320), .A2(n14409), .ZN(n12306) );
  NAND2_X1 U15181 ( .A1(n12196), .A2(n12306), .ZN(P2_U2972) );
  AOI22_X1 U15182 ( .A1(n12220), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15183 ( .A1(n18861), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18859), .ZN(n18878) );
  INV_X1 U15184 ( .A(n18878), .ZN(n14426) );
  NAND2_X1 U15185 ( .A1(n12320), .A2(n14426), .ZN(n12198) );
  NAND2_X1 U15186 ( .A1(n12197), .A2(n12198), .ZN(P2_U2968) );
  AOI22_X1 U15187 ( .A1(n12220), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U15188 ( .A1(n12199), .A2(n12198), .ZN(P2_U2953) );
  INV_X1 U15189 ( .A(n12214), .ZN(n12209) );
  MUX2_X1 U15190 ( .A(n12201), .B(n12230), .S(n12200), .Z(n12202) );
  NAND2_X1 U15191 ( .A1(n12202), .A2(n10263), .ZN(n12205) );
  AND2_X1 U15192 ( .A1(n10294), .A2(n12203), .ZN(n12237) );
  INV_X1 U15193 ( .A(n12237), .ZN(n12204) );
  NAND2_X1 U15194 ( .A1(n12205), .A2(n12204), .ZN(n18686) );
  INV_X1 U15195 ( .A(n18686), .ZN(n12206) );
  NAND2_X1 U15196 ( .A1(n12206), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18807) );
  NAND2_X1 U15197 ( .A1(n18686), .A2(n12207), .ZN(n12208) );
  NAND2_X1 U15198 ( .A1(n18807), .A2(n12208), .ZN(n15925) );
  NAND2_X1 U15199 ( .A1(n12209), .A2(n13275), .ZN(n15816) );
  NAND2_X1 U15200 ( .A1(n12230), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12227) );
  OAI21_X1 U15201 ( .B1(n12230), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12227), .ZN(n15920) );
  INV_X1 U15202 ( .A(n15920), .ZN(n12212) );
  INV_X2 U15203 ( .A(n15908), .ZN(n18815) );
  NAND2_X1 U15204 ( .A1(n18815), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n15923) );
  NAND2_X1 U15205 ( .A1(n15923), .A2(n12210), .ZN(n12211) );
  AOI21_X1 U15206 ( .B1(n18814), .B2(n12212), .A(n12211), .ZN(n12217) );
  NOR2_X1 U15207 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18495) );
  INV_X1 U15208 ( .A(n18495), .ZN(n19543) );
  NAND2_X1 U15209 ( .A1(n19550), .A2(n19543), .ZN(n19561) );
  NAND2_X1 U15210 ( .A1(n19561), .A2(n15967), .ZN(n12213) );
  NAND2_X1 U15211 ( .A1(n15833), .A2(n12233), .ZN(n12215) );
  NAND2_X1 U15212 ( .A1(n12215), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12216) );
  OAI211_X1 U15213 ( .C1(n15817), .C2(n15925), .A(n12217), .B(n12216), .ZN(
        P2_U3014) );
  INV_X1 U15214 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18769) );
  NAND2_X1 U15215 ( .A1(n12220), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12219) );
  NAND2_X1 U15216 ( .A1(n12320), .A2(n18711), .ZN(n12315) );
  OAI211_X1 U15217 ( .C1(n18769), .C2(n12935), .A(n12219), .B(n12315), .ZN(
        P2_U2981) );
  INV_X1 U15218 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12222) );
  INV_X1 U15219 ( .A(n12220), .ZN(n12289) );
  INV_X1 U15220 ( .A(n12320), .ZN(n12225) );
  OAI22_X1 U15221 ( .A1(n18859), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n18861), .ZN(n18866) );
  INV_X1 U15222 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12221) );
  OAI222_X1 U15223 ( .A1(n12222), .A2(n12289), .B1(n12225), .B2(n18866), .C1(
        n12935), .C2(n12221), .ZN(P2_U2967) );
  INV_X1 U15224 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12223) );
  INV_X1 U15225 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12330) );
  OAI222_X1 U15226 ( .A1(n12223), .A2(n12289), .B1(n12935), .B2(n12330), .C1(
        n12225), .C2(n18866), .ZN(P2_U2952) );
  INV_X1 U15227 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15228 ( .A1(n18861), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18859), .ZN(n18709) );
  INV_X1 U15229 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12224) );
  OAI222_X1 U15230 ( .A1(n12226), .A2(n12289), .B1(n12225), .B2(n18709), .C1(
        n12935), .C2(n12224), .ZN(P2_U2982) );
  AND2_X1 U15231 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19562) );
  NOR2_X1 U15232 ( .A1(n12236), .A2(n12227), .ZN(n12229) );
  AND2_X1 U15233 ( .A1(n12230), .A2(n12207), .ZN(n12228) );
  XNOR2_X1 U15234 ( .A(n12228), .B(n12236), .ZN(n18813) );
  NOR2_X1 U15235 ( .A1(n18850), .A2(n18813), .ZN(n18812) );
  NOR2_X1 U15236 ( .A1(n12229), .A2(n18812), .ZN(n12829) );
  XOR2_X1 U15237 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12829), .Z(
        n12832) );
  NOR2_X1 U15238 ( .A1(n12230), .A2(n12236), .ZN(n12231) );
  NAND2_X1 U15239 ( .A1(n13275), .A2(n12231), .ZN(n12745) );
  XNOR2_X1 U15240 ( .A(n12745), .B(n12232), .ZN(n12831) );
  XNOR2_X1 U15241 ( .A(n12832), .B(n12831), .ZN(n18842) );
  INV_X1 U15242 ( .A(n18842), .ZN(n12250) );
  OAI21_X1 U15243 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20564), .A(n12233), 
        .ZN(n12234) );
  OAI21_X1 U15244 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12922), .ZN(n12994) );
  NAND2_X1 U15245 ( .A1(n18815), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n18827) );
  NAND2_X1 U15246 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12235) );
  OAI211_X1 U15247 ( .C1(n18817), .C2(n12994), .A(n18827), .B(n12235), .ZN(
        n12249) );
  OR2_X1 U15248 ( .A1(n12236), .A2(n10294), .ZN(n12239) );
  NAND2_X1 U15249 ( .A1(n12237), .A2(n10310), .ZN(n12238) );
  NAND2_X1 U15250 ( .A1(n12239), .A2(n12238), .ZN(n12245) );
  INV_X1 U15251 ( .A(n12245), .ZN(n12241) );
  NAND3_X1 U15252 ( .A1(n18899), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U15253 ( .A1(n12241), .A2(n12240), .ZN(n18808) );
  NOR2_X1 U15254 ( .A1(n18807), .A2(n18808), .ZN(n12242) );
  NAND2_X1 U15255 ( .A1(n18807), .A2(n18808), .ZN(n18806) );
  OAI21_X1 U15256 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12242), .A(
        n18806), .ZN(n12247) );
  INV_X1 U15257 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12996) );
  MUX2_X1 U15258 ( .A(n12243), .B(n12996), .S(n10294), .Z(n12244) );
  OAI21_X1 U15259 ( .B1(n12245), .B2(n12244), .A(n12773), .ZN(n12997) );
  INV_X1 U15260 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12828) );
  XNOR2_X1 U15261 ( .A(n12997), .B(n12828), .ZN(n12246) );
  OR2_X1 U15262 ( .A1(n12247), .A2(n12246), .ZN(n18825) );
  NAND2_X1 U15263 ( .A1(n12247), .A2(n12246), .ZN(n18824) );
  AND3_X1 U15264 ( .A1(n18825), .A2(n18811), .A3(n18824), .ZN(n12248) );
  AOI211_X1 U15265 ( .C1(n18814), .C2(n12250), .A(n12249), .B(n12248), .ZN(
        n12251) );
  OAI21_X1 U15266 ( .B1(n13001), .B2(n15828), .A(n12251), .ZN(P2_U3012) );
  INV_X1 U15267 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14353) );
  OR2_X1 U15268 ( .A1(n15943), .A2(n13275), .ZN(n13042) );
  OR2_X1 U15269 ( .A1(n10815), .A2(n19458), .ZN(n12252) );
  OAI21_X1 U15270 ( .B1(n13042), .B2(n12252), .A(n12935), .ZN(n12253) );
  AND2_X1 U15271 ( .A1(n12253), .A2(n19591), .ZN(n18766) );
  INV_X1 U15272 ( .A(n12254), .ZN(n12255) );
  NAND2_X1 U15273 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n15405) );
  NOR2_X1 U15274 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15405), .ZN(n18797) );
  CLKBUF_X2 U15275 ( .A(n18797), .Z(n19603) );
  NOR2_X4 U15276 ( .A1(n18766), .A2(n19603), .ZN(n18796) );
  AOI22_X1 U15277 ( .A1(n19603), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12256) );
  OAI21_X1 U15278 ( .B1(n14353), .B2(n12341), .A(n12256), .ZN(P2_U2922) );
  INV_X1 U15279 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15280 ( .A1(n19603), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12257) );
  OAI21_X1 U15281 ( .B1(n12317), .B2(n12341), .A(n12257), .ZN(P2_U2921) );
  INV_X1 U15282 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n20521) );
  AOI22_X1 U15283 ( .A1(n19603), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12258) );
  OAI21_X1 U15284 ( .B1(n20521), .B2(n12341), .A(n12258), .ZN(P2_U2927) );
  INV_X1 U15285 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15286 ( .A1(n19603), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12259) );
  OAI21_X1 U15287 ( .B1(n12260), .B2(n12341), .A(n12259), .ZN(P2_U2926) );
  INV_X1 U15288 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n20640) );
  AOI22_X1 U15289 ( .A1(n19603), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12261) );
  OAI21_X1 U15290 ( .B1(n20640), .B2(n12341), .A(n12261), .ZN(P2_U2925) );
  INV_X1 U15291 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15292 ( .A1(n19603), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12262) );
  OAI21_X1 U15293 ( .B1(n12263), .B2(n12341), .A(n12262), .ZN(P2_U2924) );
  INV_X1 U15294 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15295 ( .A1(n19603), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12264) );
  OAI21_X1 U15296 ( .B1(n12314), .B2(n12341), .A(n12264), .ZN(P2_U2923) );
  NOR4_X1 U15297 ( .A1(n12268), .A2(n12267), .A3(n12266), .A4(n12265), .ZN(
        n12269) );
  NOR2_X1 U15298 ( .A1(n12270), .A2(n12269), .ZN(n13451) );
  AND2_X1 U15299 ( .A1(n13453), .A2(n13451), .ZN(n13464) );
  NAND2_X1 U15300 ( .A1(n13464), .A2(n12461), .ZN(n12273) );
  NOR2_X2 U15301 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20348) );
  AND2_X1 U15302 ( .A1(n20348), .A2(n20400), .ZN(n13071) );
  INV_X1 U15303 ( .A(n12371), .ZN(n12271) );
  AOI211_X1 U15304 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n12273), .A(n13071), 
        .B(n12271), .ZN(n12272) );
  INV_X1 U15305 ( .A(n12272), .ZN(P1_U2801) );
  INV_X1 U15306 ( .A(n20496), .ZN(n12275) );
  OAI21_X1 U15307 ( .B1(n13071), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12275), 
        .ZN(n12274) );
  OAI21_X1 U15308 ( .B1(n12276), .B2(n12275), .A(n12274), .ZN(P1_U3487) );
  INV_X1 U15309 ( .A(n12277), .ZN(n12278) );
  OR2_X1 U15310 ( .A1(n18701), .A2(n12278), .ZN(n18747) );
  INV_X1 U15311 ( .A(n18747), .ZN(n18765) );
  NOR2_X1 U15312 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  NOR2_X1 U15313 ( .A1(n12282), .A2(n12281), .ZN(n18683) );
  AOI22_X1 U15314 ( .A1(n18757), .A2(n18683), .B1(n18756), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n12288) );
  AND2_X1 U15315 ( .A1(n19571), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12283) );
  OAI211_X1 U15316 ( .C1(n13275), .C2(n12284), .A(n10266), .B(n12283), .ZN(
        n12285) );
  INV_X1 U15317 ( .A(n12285), .ZN(n12286) );
  NAND2_X1 U15318 ( .A1(n19127), .A2(n18683), .ZN(n18759) );
  OAI211_X1 U15319 ( .C1(n19127), .C2(n18683), .A(n18759), .B(n18761), .ZN(
        n12287) );
  OAI211_X1 U15320 ( .C1(n18765), .C2(n18866), .A(n12288), .B(n12287), .ZN(
        P2_U2919) );
  AOI22_X1 U15321 ( .A1(n12324), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n12310), .ZN(n12293) );
  INV_X1 U15322 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n12290) );
  OR2_X1 U15323 ( .A1(n18859), .A2(n12290), .ZN(n12292) );
  NAND2_X1 U15324 ( .A1(n18859), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12291) );
  AND2_X1 U15325 ( .A1(n12292), .A2(n12291), .ZN(n18728) );
  INV_X1 U15326 ( .A(n18728), .ZN(n14390) );
  NAND2_X1 U15327 ( .A1(n12320), .A2(n14390), .ZN(n12302) );
  NAND2_X1 U15328 ( .A1(n12293), .A2(n12302), .ZN(P2_U2960) );
  AOI22_X1 U15329 ( .A1(n12324), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n12310), .ZN(n12295) );
  NAND2_X1 U15330 ( .A1(n12295), .A2(n12294), .ZN(P2_U2958) );
  AOI22_X1 U15331 ( .A1(n12324), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n12310), .ZN(n12297) );
  NAND2_X1 U15332 ( .A1(n12297), .A2(n12296), .ZN(P2_U2961) );
  AOI22_X1 U15333 ( .A1(n12324), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n12310), .ZN(n12299) );
  NAND2_X1 U15334 ( .A1(n12299), .A2(n12298), .ZN(P2_U2956) );
  AOI22_X1 U15335 ( .A1(n12324), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n12310), .ZN(n12301) );
  NAND2_X1 U15336 ( .A1(n12301), .A2(n12300), .ZN(P2_U2963) );
  AOI22_X1 U15337 ( .A1(n12324), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U15338 ( .A1(n12303), .A2(n12302), .ZN(P2_U2975) );
  AOI22_X1 U15339 ( .A1(n12324), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12305) );
  NAND2_X1 U15340 ( .A1(n12305), .A2(n12304), .ZN(P2_U2959) );
  AOI22_X1 U15341 ( .A1(n12324), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U15342 ( .A1(n12307), .A2(n12306), .ZN(P2_U2957) );
  AOI22_X1 U15343 ( .A1(n12324), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n12310), .ZN(n12309) );
  NAND2_X1 U15344 ( .A1(n12309), .A2(n12308), .ZN(P2_U2954) );
  AOI22_X1 U15345 ( .A1(n12324), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n12310), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15346 ( .A1(n12312), .A2(n12311), .ZN(P2_U2955) );
  NAND2_X1 U15347 ( .A1(n12324), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12313) );
  MUX2_X1 U15348 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n18859), .Z(n18717) );
  NAND2_X1 U15349 ( .A1(n12320), .A2(n18717), .ZN(n12325) );
  OAI211_X1 U15350 ( .C1(n12314), .C2(n12935), .A(n12313), .B(n12325), .ZN(
        P2_U2964) );
  NAND2_X1 U15351 ( .A1(n12324), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12316) );
  OAI211_X1 U15352 ( .C1(n12317), .C2(n12935), .A(n12316), .B(n12315), .ZN(
        P2_U2966) );
  INV_X1 U15353 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18777) );
  NAND2_X1 U15354 ( .A1(n12324), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12321) );
  NAND2_X1 U15355 ( .A1(n18859), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12319) );
  INV_X1 U15356 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16085) );
  OR2_X1 U15357 ( .A1(n18859), .A2(n16085), .ZN(n12318) );
  NAND2_X1 U15358 ( .A1(n12319), .A2(n12318), .ZN(n18722) );
  NAND2_X1 U15359 ( .A1(n12320), .A2(n18722), .ZN(n12322) );
  OAI211_X1 U15360 ( .C1(n18777), .C2(n12935), .A(n12321), .B(n12322), .ZN(
        P2_U2977) );
  NAND2_X1 U15361 ( .A1(n12324), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12323) );
  OAI211_X1 U15362 ( .C1(n20640), .C2(n12935), .A(n12323), .B(n12322), .ZN(
        P2_U2962) );
  INV_X1 U15363 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18773) );
  NAND2_X1 U15364 ( .A1(n12324), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12326) );
  OAI211_X1 U15365 ( .C1(n18773), .C2(n12935), .A(n12326), .B(n12325), .ZN(
        P2_U2979) );
  AOI22_X1 U15366 ( .A1(n18797), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12327) );
  OAI21_X1 U15367 ( .B1(n12328), .B2(n12341), .A(n12327), .ZN(P2_U2934) );
  AOI22_X1 U15368 ( .A1(n18797), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12329) );
  OAI21_X1 U15369 ( .B1(n12330), .B2(n12341), .A(n12329), .ZN(P2_U2935) );
  AOI22_X1 U15370 ( .A1(n19603), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12331) );
  OAI21_X1 U15371 ( .B1(n12332), .B2(n12341), .A(n12331), .ZN(P2_U2930) );
  INV_X1 U15372 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15373 ( .A1(n19603), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12333) );
  OAI21_X1 U15374 ( .B1(n12334), .B2(n12341), .A(n12333), .ZN(P2_U2933) );
  INV_X1 U15375 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15376 ( .A1(n19603), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12335) );
  OAI21_X1 U15377 ( .B1(n12336), .B2(n12341), .A(n12335), .ZN(P2_U2929) );
  INV_X1 U15378 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15379 ( .A1(n19603), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12337) );
  OAI21_X1 U15380 ( .B1(n12338), .B2(n12341), .A(n12337), .ZN(P2_U2928) );
  INV_X1 U15381 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n20627) );
  AOI22_X1 U15382 ( .A1(n19603), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12339) );
  OAI21_X1 U15383 ( .B1(n20627), .B2(n12341), .A(n12339), .ZN(P2_U2931) );
  AOI22_X1 U15384 ( .A1(n19603), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12340) );
  OAI21_X1 U15385 ( .B1(n12342), .B2(n12341), .A(n12340), .ZN(P2_U2932) );
  NAND2_X1 U15386 ( .A1(n12345), .A2(n12344), .ZN(n12346) );
  MUX2_X1 U15387 ( .A(n12996), .B(n13001), .S(n14333), .Z(n12347) );
  OAI21_X1 U15388 ( .B1(n19555), .B2(n14342), .A(n12347), .ZN(P2_U2885) );
  OR2_X1 U15389 ( .A1(n12349), .A2(n12348), .ZN(n12351) );
  MUX2_X1 U15390 ( .A(n10310), .B(n12734), .S(n14333), .Z(n12352) );
  OAI21_X1 U15391 ( .B1(n19563), .B2(n14342), .A(n12352), .ZN(P2_U2886) );
  MUX2_X1 U15392 ( .A(n12203), .B(n13035), .S(n14333), .Z(n12353) );
  OAI21_X1 U15393 ( .B1(n19573), .B2(n14342), .A(n12353), .ZN(P2_U2887) );
  INV_X1 U15394 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12358) );
  OR2_X1 U15395 ( .A1(n12354), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15401) );
  INV_X1 U15396 ( .A(n15401), .ZN(n20488) );
  NAND3_X1 U15397 ( .A1(n13463), .A2(n19871), .A3(n20488), .ZN(n15380) );
  NAND2_X1 U15398 ( .A1(n13453), .A2(n12889), .ZN(n12640) );
  NAND2_X1 U15399 ( .A1(n14113), .A2(n20488), .ZN(n12356) );
  INV_X1 U15400 ( .A(n12466), .ZN(n12355) );
  NAND2_X1 U15401 ( .A1(n19732), .A2(n12443), .ZN(n12552) );
  NAND2_X1 U15402 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15664) );
  INV_X1 U15403 ( .A(n15664), .ZN(n15660) );
  NAND2_X1 U15404 ( .A1(n20401), .A2(n15660), .ZN(n19730) );
  NOR2_X4 U15405 ( .A1(n19732), .A2(n19759), .ZN(n19758) );
  AOI22_X1 U15406 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12357) );
  OAI21_X1 U15407 ( .B1(n12358), .B2(n12552), .A(n12357), .ZN(P1_U2911) );
  INV_X1 U15408 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15409 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12359) );
  OAI21_X1 U15410 ( .B1(n12360), .B2(n12552), .A(n12359), .ZN(P1_U2912) );
  INV_X1 U15411 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15412 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12361) );
  OAI21_X1 U15413 ( .B1(n12362), .B2(n12552), .A(n12361), .ZN(P1_U2908) );
  INV_X1 U15414 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15415 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12363) );
  OAI21_X1 U15416 ( .B1(n12364), .B2(n12552), .A(n12363), .ZN(P1_U2906) );
  INV_X1 U15417 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n20585) );
  AOI22_X1 U15418 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12365) );
  OAI21_X1 U15419 ( .B1(n20585), .B2(n12552), .A(n12365), .ZN(P1_U2907) );
  INV_X1 U15420 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15421 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12366) );
  OAI21_X1 U15422 ( .B1(n12367), .B2(n12552), .A(n12366), .ZN(P1_U2909) );
  INV_X1 U15423 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15424 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12368) );
  OAI21_X1 U15425 ( .B1(n12369), .B2(n12552), .A(n12368), .ZN(P1_U2910) );
  NAND2_X1 U15426 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20415) );
  INV_X1 U15427 ( .A(n20415), .ZN(n20491) );
  AND2_X1 U15428 ( .A1(n20489), .A2(n20491), .ZN(n12370) );
  OR2_X1 U15429 ( .A1(n19767), .A2(n12889), .ZN(n12567) );
  INV_X1 U15430 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13763) );
  OR2_X1 U15431 ( .A1(n19767), .A2(n19871), .ZN(n12474) );
  INV_X1 U15432 ( .A(DATAI_15_), .ZN(n12373) );
  INV_X1 U15433 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12372) );
  MUX2_X1 U15434 ( .A(n12373), .B(n12372), .S(n19852), .Z(n13765) );
  INV_X1 U15435 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19731) );
  OAI222_X1 U15436 ( .A1(n12567), .A2(n13763), .B1(n12474), .B2(n13765), .C1(
        n12575), .C2(n19731), .ZN(P1_U2967) );
  NAND2_X1 U15437 ( .A1(n13451), .A2(n20415), .ZN(n12375) );
  NOR2_X1 U15438 ( .A1(n12374), .A2(n12375), .ZN(n12462) );
  NAND2_X1 U15439 ( .A1(n12456), .A2(n19855), .ZN(n12376) );
  OAI21_X1 U15440 ( .B1(n13140), .B2(n12470), .A(n12444), .ZN(n12378) );
  NAND2_X1 U15441 ( .A1(n12405), .A2(n12378), .ZN(n12379) );
  NAND2_X1 U15442 ( .A1(n10101), .A2(n12379), .ZN(n12419) );
  OAI21_X1 U15443 ( .B1(n12886), .B2(n12416), .A(n12419), .ZN(n12380) );
  OR3_X1 U15444 ( .A1(n12381), .A2(n12462), .A3(n12380), .ZN(n12389) );
  NAND2_X1 U15445 ( .A1(n12640), .A2(n12421), .ZN(n12382) );
  NAND3_X1 U15446 ( .A1(n12382), .A2(n20488), .A3(n20415), .ZN(n12387) );
  NAND2_X1 U15447 ( .A1(n12405), .A2(n13462), .ZN(n13455) );
  INV_X1 U15448 ( .A(n12383), .ZN(n12384) );
  NAND2_X1 U15449 ( .A1(n12384), .A2(n20415), .ZN(n12385) );
  NAND2_X1 U15450 ( .A1(n13455), .A2(n12385), .ZN(n12465) );
  INV_X1 U15451 ( .A(n12465), .ZN(n12386) );
  AOI21_X1 U15452 ( .B1(n12387), .B2(n12386), .A(n13456), .ZN(n12388) );
  NAND2_X1 U15453 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15660), .ZN(n12651) );
  INV_X1 U15454 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19617) );
  OAI22_X1 U15455 ( .A1(n15360), .A2(n19610), .B1(n12651), .B2(n19617), .ZN(
        n12392) );
  AOI21_X1 U15456 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20401), .A(n12392), 
        .ZN(n12390) );
  INV_X1 U15457 ( .A(n12390), .ZN(n14133) );
  INV_X1 U15458 ( .A(n19993), .ZN(n20229) );
  OR2_X1 U15459 ( .A1(n11289), .A2(n20229), .ZN(n12391) );
  XNOR2_X1 U15460 ( .A(n12391), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19697) );
  INV_X1 U15461 ( .A(n12374), .ZN(n12646) );
  NAND4_X1 U15462 ( .A1(n19697), .A2(n14128), .A3(n12646), .A4(n12392), .ZN(
        n12393) );
  OAI21_X1 U15463 ( .B1(n14133), .B2(n12648), .A(n12393), .ZN(P1_U3468) );
  MUX2_X1 U15464 ( .A(n10330), .B(n9935), .S(n14333), .Z(n12396) );
  OAI21_X1 U15465 ( .B1(n19160), .B2(n14342), .A(n12396), .ZN(P2_U2884) );
  NOR2_X1 U15466 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20400), .ZN(n20499) );
  NAND2_X1 U15467 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20499), .ZN(n15658) );
  INV_X1 U15468 ( .A(n15658), .ZN(n12397) );
  INV_X1 U15469 ( .A(n12398), .ZN(n12401) );
  OAI21_X1 U15470 ( .B1(n12401), .B2(n12400), .A(n12399), .ZN(n13060) );
  NAND2_X1 U15471 ( .A1(n20401), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U15472 ( .A1(n20291), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12402) );
  AND2_X1 U15473 ( .A1(n12403), .A2(n12402), .ZN(n12500) );
  NAND2_X1 U15474 ( .A1(n12405), .A2(n12404), .ZN(n13454) );
  NAND2_X1 U15475 ( .A1(n20346), .A2(n12407), .ZN(n20497) );
  AND2_X1 U15476 ( .A1(n20497), .A2(n20401), .ZN(n12406) );
  NAND2_X1 U15477 ( .A1(n12500), .A2(n13917), .ZN(n12413) );
  INV_X1 U15478 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20482) );
  NOR2_X1 U15479 ( .A1(n15601), .A2(n20482), .ZN(n12437) );
  INV_X1 U15480 ( .A(n13133), .ZN(n12689) );
  NAND2_X1 U15481 ( .A1(n19855), .A2(n12408), .ZN(n12682) );
  OAI21_X1 U15482 ( .B1(n20489), .B2(n12505), .A(n12682), .ZN(n12409) );
  INV_X1 U15483 ( .A(n12409), .ZN(n12410) );
  OAI21_X1 U15484 ( .B1(n12411), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12679), .ZN(n12452) );
  NOR2_X1 U15485 ( .A1(n12452), .A2(n19804), .ZN(n12412) );
  AOI211_X1 U15486 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n12413), .A(
        n12437), .B(n12412), .ZN(n12414) );
  OAI21_X1 U15487 ( .B1(n19851), .B2(n13060), .A(n12414), .ZN(P1_U2999) );
  INV_X1 U15488 ( .A(n12456), .ZN(n14115) );
  NAND3_X1 U15489 ( .A1(n13456), .A2(n14115), .A3(n12889), .ZN(n12418) );
  NAND2_X1 U15490 ( .A1(n12889), .A2(n15401), .ZN(n12415) );
  NAND4_X1 U15491 ( .A1(n13451), .A2(n12416), .A3(n20415), .A4(n12415), .ZN(
        n12417) );
  NAND3_X1 U15492 ( .A1(n12419), .A2(n12418), .A3(n12417), .ZN(n12420) );
  NAND2_X1 U15493 ( .A1(n12420), .A2(n12461), .ZN(n12424) );
  OAI21_X1 U15494 ( .B1(n12889), .B2(n20488), .A(n20415), .ZN(n12888) );
  OAI211_X1 U15495 ( .C1(n12421), .C2(n12888), .A(n12443), .B(n13702), .ZN(
        n12422) );
  NAND3_X1 U15496 ( .A1(n12466), .A2(n19875), .A3(n12422), .ZN(n12423) );
  OAI211_X1 U15497 ( .C1(n19883), .C2(n12430), .A(n13455), .B(n13454), .ZN(
        n12425) );
  NOR2_X1 U15498 ( .A1(n12426), .A2(n12425), .ZN(n12427) );
  OAI22_X1 U15499 ( .A1(n12430), .A2(n12429), .B1(n12889), .B2(n12428), .ZN(
        n12431) );
  INV_X1 U15500 ( .A(n12431), .ZN(n12432) );
  INV_X1 U15501 ( .A(n12433), .ZN(n12435) );
  OR2_X1 U15502 ( .A1(n13472), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12434) );
  AND2_X1 U15503 ( .A1(n12435), .A2(n12434), .ZN(n13056) );
  NAND2_X1 U15504 ( .A1(n12450), .A2(n15601), .ZN(n13172) );
  INV_X1 U15505 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14119) );
  AOI21_X1 U15506 ( .B1(n14058), .B2(n13172), .A(n14119), .ZN(n12436) );
  AOI211_X1 U15507 ( .C1(n19825), .C2(n13056), .A(n12437), .B(n12436), .ZN(
        n12451) );
  OAI21_X1 U15508 ( .B1(n12439), .B2(n12443), .A(n12438), .ZN(n12440) );
  OR2_X1 U15509 ( .A1(n12441), .A2(n12440), .ZN(n12447) );
  NAND3_X1 U15510 ( .A1(n12444), .A2(n12443), .A3(n12442), .ZN(n12446) );
  NAND2_X1 U15511 ( .A1(n12446), .A2(n12445), .ZN(n12453) );
  NOR2_X1 U15512 ( .A1(n12447), .A2(n12453), .ZN(n12448) );
  INV_X1 U15513 ( .A(n13450), .ZN(n12449) );
  OAI21_X1 U15514 ( .B1(n13170), .B2(n19831), .A(n14119), .ZN(n12518) );
  OAI211_X1 U15515 ( .C1(n12452), .C2(n19838), .A(n12451), .B(n12518), .ZN(
        P1_U3031) );
  INV_X1 U15516 ( .A(n15388), .ZN(n14132) );
  INV_X1 U15517 ( .A(n19961), .ZN(n12655) );
  NOR2_X1 U15518 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  AND2_X1 U15519 ( .A1(n12374), .A2(n12455), .ZN(n14118) );
  OAI22_X1 U15520 ( .A1(n12655), .A2(n14118), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12456), .ZN(n15357) );
  AOI22_X1 U15521 ( .A1(n15357), .A2(n14128), .B1(P1_STATE2_REG_1__SCAN_IN), 
        .B2(n14119), .ZN(n12457) );
  OAI21_X1 U15522 ( .B1(n14132), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12457), .ZN(n12458) );
  NAND2_X1 U15523 ( .A1(n12458), .A2(n14133), .ZN(n12460) );
  NOR2_X1 U15524 ( .A1(n12640), .A2(n11277), .ZN(n15356) );
  NAND2_X1 U15525 ( .A1(n15356), .A2(n14128), .ZN(n12459) );
  OAI211_X1 U15526 ( .C1(n14133), .C2(n11277), .A(n12460), .B(n12459), .ZN(
        P1_U3474) );
  NAND2_X1 U15527 ( .A1(n12462), .A2(n12461), .ZN(n12468) );
  NOR2_X1 U15528 ( .A1(n12463), .A2(n13465), .ZN(n12464) );
  NAND2_X1 U15529 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  NAND2_X2 U15530 ( .A1(n13764), .A2(n12471), .ZN(n13777) );
  INV_X1 U15531 ( .A(n19852), .ZN(n19849) );
  NAND2_X1 U15532 ( .A1(n19849), .A2(DATAI_0_), .ZN(n12473) );
  NAND2_X1 U15533 ( .A1(n19852), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12472) );
  AND2_X1 U15534 ( .A1(n12473), .A2(n12472), .ZN(n19863) );
  INV_X1 U15535 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19762) );
  OAI222_X1 U15536 ( .A1(n13060), .A2(n13777), .B1(n13766), .B2(n19863), .C1(
        n13764), .C2(n19762), .ZN(P1_U2904) );
  MUX2_X1 U15537 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n19852), .Z(
        n13769) );
  NAND2_X1 U15538 ( .A1(n19773), .A2(n13769), .ZN(n19783) );
  NAND2_X1 U15539 ( .A1(n19767), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n12475) );
  OAI211_X1 U15540 ( .C1(n20585), .C2(n12567), .A(n19783), .B(n12475), .ZN(
        P1_U2950) );
  XOR2_X1 U15541 ( .A(n12476), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n12480)
         );
  AOI21_X1 U15542 ( .B1(n12477), .B2(n13434), .A(n12526), .ZN(n18672) );
  NOR2_X1 U15543 ( .A1(n14350), .A2(n12045), .ZN(n12478) );
  AOI21_X1 U15544 ( .B1(n18672), .B2(n14350), .A(n12478), .ZN(n12479) );
  OAI21_X1 U15545 ( .B1(n12480), .B2(n14342), .A(n12479), .ZN(P2_U2882) );
  AOI21_X1 U15546 ( .B1(n14110), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12481) );
  NOR2_X1 U15547 ( .A1(n11736), .A2(n12481), .ZN(n12493) );
  INV_X1 U15548 ( .A(n14118), .ZN(n12636) );
  NAND2_X1 U15549 ( .A1(n12634), .A2(n12493), .ZN(n12492) );
  NAND2_X1 U15550 ( .A1(n20110), .A2(n12636), .ZN(n12491) );
  INV_X1 U15551 ( .A(n13455), .ZN(n12482) );
  OR2_X1 U15552 ( .A1(n13450), .A2(n12482), .ZN(n12632) );
  MUX2_X1 U15553 ( .A(n12483), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14110), .Z(n12485) );
  NOR2_X1 U15554 ( .A1(n12485), .A2(n12484), .ZN(n12489) );
  NAND2_X1 U15555 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12486) );
  INV_X1 U15556 ( .A(n12486), .ZN(n12487) );
  MUX2_X1 U15557 ( .A(n12487), .B(n12486), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12488) );
  AOI22_X1 U15558 ( .A1(n12632), .A2(n12489), .B1(n14113), .B2(n12488), .ZN(
        n12490) );
  OAI211_X1 U15559 ( .C1(n12636), .C2(n12492), .A(n12491), .B(n12490), .ZN(
        n12630) );
  AOI22_X1 U15560 ( .A1(n15388), .A2(n12493), .B1(n14128), .B2(n12630), .ZN(
        n12494) );
  MUX2_X1 U15561 ( .A(n12495), .B(n12494), .S(n14133), .Z(n12496) );
  INV_X1 U15562 ( .A(n12496), .ZN(P1_U3469) );
  INV_X1 U15563 ( .A(n12563), .ZN(n12497) );
  OAI21_X1 U15564 ( .B1(n12499), .B2(n12498), .A(n12497), .ZN(n12910) );
  INV_X1 U15565 ( .A(n12500), .ZN(n12501) );
  INV_X1 U15566 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12900) );
  NAND2_X1 U15567 ( .A1(n12502), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n12517) );
  OAI21_X1 U15568 ( .B1(n13917), .B2(n12900), .A(n12517), .ZN(n12503) );
  AOI21_X1 U15569 ( .B1(n15536), .B2(n12900), .A(n12503), .ZN(n12514) );
  NAND2_X1 U15570 ( .A1(n12504), .A2(n12889), .ZN(n12511) );
  NAND2_X1 U15571 ( .A1(n12506), .A2(n12505), .ZN(n12691) );
  OAI21_X1 U15572 ( .B1(n12506), .B2(n12505), .A(n12691), .ZN(n12508) );
  OAI211_X1 U15573 ( .C1(n12508), .C2(n20489), .A(n12507), .B(n11142), .ZN(
        n12509) );
  INV_X1 U15574 ( .A(n12509), .ZN(n12510) );
  NAND2_X1 U15575 ( .A1(n12511), .A2(n12510), .ZN(n12677) );
  XNOR2_X1 U15576 ( .A(n12679), .B(n12677), .ZN(n12512) );
  OR2_X1 U15577 ( .A1(n12512), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12516) );
  NAND2_X1 U15578 ( .A1(n12512), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12681) );
  NAND3_X1 U15579 ( .A1(n12516), .A2(n12681), .A3(n19795), .ZN(n12513) );
  OAI211_X1 U15580 ( .C1(n12910), .C2(n19851), .A(n12514), .B(n12513), .ZN(
        P1_U2998) );
  XNOR2_X1 U15581 ( .A(n12515), .B(n13471), .ZN(n12892) );
  NAND3_X1 U15582 ( .A1(n12516), .A2(n12681), .A3(n19823), .ZN(n12523) );
  AOI211_X1 U15583 ( .C1(n14119), .C2(n14058), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n15629), .ZN(n12521) );
  INV_X1 U15584 ( .A(n12517), .ZN(n12520) );
  INV_X1 U15585 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14120) );
  AOI21_X1 U15586 ( .B1(n12518), .B2(n13172), .A(n14120), .ZN(n12519) );
  NOR3_X1 U15587 ( .A1(n12521), .A2(n12520), .A3(n12519), .ZN(n12522) );
  OAI211_X1 U15588 ( .C1(n12892), .C2(n19834), .A(n12523), .B(n12522), .ZN(
        P1_U3030) );
  NAND2_X1 U15589 ( .A1(n19849), .A2(DATAI_1_), .ZN(n12525) );
  NAND2_X1 U15590 ( .A1(n19852), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12524) );
  AND2_X1 U15591 ( .A1(n12525), .A2(n12524), .ZN(n19872) );
  INV_X1 U15592 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19757) );
  OAI222_X1 U15593 ( .A1(n12910), .A2(n13777), .B1(n13766), .B2(n19872), .C1(
        n13764), .C2(n19757), .ZN(P1_U2903) );
  NOR2_X1 U15594 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  OR2_X1 U15595 ( .A1(n12534), .A2(n12528), .ZN(n18657) );
  NOR2_X1 U15596 ( .A1(n12476), .A2(n10549), .ZN(n12529) );
  OAI211_X1 U15597 ( .C1(n12529), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14344), .B(n12532), .ZN(n12531) );
  NAND2_X1 U15598 ( .A1(n14340), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12530) );
  OAI211_X1 U15599 ( .C1(n18657), .C2(n14340), .A(n12531), .B(n12530), .ZN(
        P2_U2881) );
  INV_X1 U15600 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12903) );
  OAI222_X1 U15601 ( .A1(n12892), .A2(n13698), .B1(n12903), .B2(n19728), .C1(
        n13696), .C2(n12910), .ZN(P1_U2871) );
  XOR2_X1 U15602 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n12532), .Z(n12537)
         );
  NOR2_X1 U15603 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  OR2_X1 U15604 ( .A1(n12556), .A2(n12535), .ZN(n18642) );
  MUX2_X1 U15605 ( .A(n18642), .B(n12950), .S(n14340), .Z(n12536) );
  OAI21_X1 U15606 ( .B1(n12537), .B2(n14342), .A(n12536), .ZN(P2_U2880) );
  INV_X1 U15607 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15608 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12538) );
  OAI21_X1 U15609 ( .B1(n12539), .B2(n12552), .A(n12538), .ZN(P1_U2916) );
  INV_X1 U15610 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U15611 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12540) );
  OAI21_X1 U15612 ( .B1(n12541), .B2(n12552), .A(n12540), .ZN(P1_U2919) );
  INV_X1 U15613 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15614 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12542) );
  OAI21_X1 U15615 ( .B1(n12543), .B2(n12552), .A(n12542), .ZN(P1_U2913) );
  AOI22_X1 U15616 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12544) );
  OAI21_X1 U15617 ( .B1(n13744), .B2(n12552), .A(n12544), .ZN(P1_U2918) );
  INV_X1 U15618 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15619 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12545) );
  OAI21_X1 U15620 ( .B1(n12546), .B2(n12552), .A(n12545), .ZN(P1_U2914) );
  INV_X1 U15621 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15622 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12547) );
  OAI21_X1 U15623 ( .B1(n12548), .B2(n12552), .A(n12547), .ZN(P1_U2920) );
  INV_X1 U15624 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15625 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12549) );
  OAI21_X1 U15626 ( .B1(n12550), .B2(n12552), .A(n12549), .ZN(P1_U2917) );
  INV_X1 U15627 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15628 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12551) );
  OAI21_X1 U15629 ( .B1(n12553), .B2(n12552), .A(n12551), .ZN(P1_U2915) );
  INV_X1 U15630 ( .A(n13056), .ZN(n12554) );
  OAI222_X1 U15631 ( .A1(n12554), .A2(n13698), .B1(n19728), .B2(n11915), .C1(
        n13060), .C2(n13696), .ZN(P1_U2872) );
  OR2_X1 U15632 ( .A1(n12556), .A2(n12555), .ZN(n12557) );
  NAND2_X1 U15633 ( .A1(n12557), .A2(n12624), .ZN(n15893) );
  OAI211_X1 U15634 ( .C1(n9713), .C2(n12559), .A(n12558), .B(n14344), .ZN(
        n12561) );
  NAND2_X1 U15635 ( .A1(n14340), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12560) );
  OAI211_X1 U15636 ( .C1(n15893), .C2(n14340), .A(n12561), .B(n12560), .ZN(
        P2_U2879) );
  OAI21_X1 U15637 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n19805) );
  NAND2_X1 U15638 ( .A1(n19849), .A2(DATAI_2_), .ZN(n12566) );
  NAND2_X1 U15639 ( .A1(n19852), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12565) );
  AND2_X1 U15640 ( .A1(n12566), .A2(n12565), .ZN(n19876) );
  INV_X1 U15641 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19755) );
  OAI222_X1 U15642 ( .A1(n19805), .A2(n13777), .B1(n13766), .B2(n19876), .C1(
        n13764), .C2(n19755), .ZN(P1_U2902) );
  AOI22_X1 U15643 ( .A1(n19786), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19785), .ZN(n12571) );
  NAND2_X1 U15644 ( .A1(n19849), .A2(DATAI_4_), .ZN(n12569) );
  NAND2_X1 U15645 ( .A1(n19852), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12568) );
  AND2_X1 U15646 ( .A1(n12569), .A2(n12568), .ZN(n19884) );
  INV_X1 U15647 ( .A(n19884), .ZN(n12570) );
  NAND2_X1 U15648 ( .A1(n19773), .A2(n12570), .ZN(n12605) );
  NAND2_X1 U15649 ( .A1(n12571), .A2(n12605), .ZN(P1_U2941) );
  AOI22_X1 U15650 ( .A1(n19786), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19785), .ZN(n12574) );
  NAND2_X1 U15651 ( .A1(n19849), .A2(DATAI_5_), .ZN(n12573) );
  NAND2_X1 U15652 ( .A1(n19852), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12572) );
  AND2_X1 U15653 ( .A1(n12573), .A2(n12572), .ZN(n19888) );
  INV_X1 U15654 ( .A(n19888), .ZN(n13734) );
  NAND2_X1 U15655 ( .A1(n19773), .A2(n13734), .ZN(n12576) );
  NAND2_X1 U15656 ( .A1(n12574), .A2(n12576), .ZN(P1_U2942) );
  INV_X1 U15657 ( .A(n12575), .ZN(n19785) );
  AOI22_X1 U15658 ( .A1(n19786), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19785), .ZN(n12577) );
  NAND2_X1 U15659 ( .A1(n12577), .A2(n12576), .ZN(P1_U2957) );
  AOI22_X1 U15660 ( .A1(n19786), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19785), .ZN(n12581) );
  NAND2_X1 U15661 ( .A1(n19849), .A2(DATAI_6_), .ZN(n12579) );
  NAND2_X1 U15662 ( .A1(n19852), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12578) );
  AND2_X1 U15663 ( .A1(n12579), .A2(n12578), .ZN(n19891) );
  INV_X1 U15664 ( .A(n19891), .ZN(n12580) );
  NAND2_X1 U15665 ( .A1(n19773), .A2(n12580), .ZN(n12609) );
  NAND2_X1 U15666 ( .A1(n12581), .A2(n12609), .ZN(P1_U2943) );
  AOI22_X1 U15667 ( .A1(n19786), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19785), .ZN(n12584) );
  NAND2_X1 U15668 ( .A1(n19849), .A2(DATAI_3_), .ZN(n12583) );
  NAND2_X1 U15669 ( .A1(n19852), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12582) );
  AND2_X1 U15670 ( .A1(n12583), .A2(n12582), .ZN(n19880) );
  INV_X1 U15671 ( .A(n19880), .ZN(n13741) );
  NAND2_X1 U15672 ( .A1(n19773), .A2(n13741), .ZN(n12603) );
  NAND2_X1 U15673 ( .A1(n12584), .A2(n12603), .ZN(P1_U2940) );
  AOI22_X1 U15674 ( .A1(n19786), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19785), .ZN(n12588) );
  NAND2_X1 U15675 ( .A1(n19849), .A2(DATAI_7_), .ZN(n12586) );
  NAND2_X1 U15676 ( .A1(n19852), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12585) );
  AND2_X1 U15677 ( .A1(n12586), .A2(n12585), .ZN(n19899) );
  INV_X1 U15678 ( .A(n19899), .ZN(n12587) );
  NAND2_X1 U15679 ( .A1(n19773), .A2(n12587), .ZN(n12594) );
  NAND2_X1 U15680 ( .A1(n12588), .A2(n12594), .ZN(P1_U2944) );
  AOI22_X1 U15681 ( .A1(n19786), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19785), .ZN(n12589) );
  MUX2_X1 U15682 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n19852), .Z(
        n13717) );
  NAND2_X1 U15683 ( .A1(n19773), .A2(n13717), .ZN(n12607) );
  NAND2_X1 U15684 ( .A1(n12589), .A2(n12607), .ZN(P1_U2947) );
  AOI22_X1 U15685 ( .A1(n19786), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19785), .ZN(n12591) );
  INV_X1 U15686 ( .A(n19863), .ZN(n12590) );
  NAND2_X1 U15687 ( .A1(n19773), .A2(n12590), .ZN(n12599) );
  NAND2_X1 U15688 ( .A1(n12591), .A2(n12599), .ZN(P1_U2937) );
  AOI22_X1 U15689 ( .A1(n19786), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19785), .ZN(n12593) );
  INV_X1 U15690 ( .A(n19876), .ZN(n12592) );
  NAND2_X1 U15691 ( .A1(n19773), .A2(n12592), .ZN(n12597) );
  NAND2_X1 U15692 ( .A1(n12593), .A2(n12597), .ZN(P1_U2954) );
  AOI22_X1 U15693 ( .A1(n19786), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19785), .ZN(n12595) );
  NAND2_X1 U15694 ( .A1(n12595), .A2(n12594), .ZN(P1_U2959) );
  AOI22_X1 U15695 ( .A1(n19786), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19785), .ZN(n12596) );
  INV_X1 U15696 ( .A(n19872), .ZN(n13751) );
  NAND2_X1 U15697 ( .A1(n19773), .A2(n13751), .ZN(n12601) );
  NAND2_X1 U15698 ( .A1(n12596), .A2(n12601), .ZN(P1_U2938) );
  AOI22_X1 U15699 ( .A1(n19786), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19785), .ZN(n12598) );
  NAND2_X1 U15700 ( .A1(n12598), .A2(n12597), .ZN(P1_U2939) );
  AOI22_X1 U15701 ( .A1(n19786), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19785), .ZN(n12600) );
  NAND2_X1 U15702 ( .A1(n12600), .A2(n12599), .ZN(P1_U2952) );
  AOI22_X1 U15703 ( .A1(n19786), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19785), .ZN(n12602) );
  NAND2_X1 U15704 ( .A1(n12602), .A2(n12601), .ZN(P1_U2953) );
  AOI22_X1 U15705 ( .A1(n19786), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19785), .ZN(n12604) );
  NAND2_X1 U15706 ( .A1(n12604), .A2(n12603), .ZN(P1_U2955) );
  AOI22_X1 U15707 ( .A1(n19786), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19785), .ZN(n12606) );
  NAND2_X1 U15708 ( .A1(n12606), .A2(n12605), .ZN(P1_U2956) );
  AOI22_X1 U15709 ( .A1(n19786), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19785), .ZN(n12608) );
  NAND2_X1 U15710 ( .A1(n12608), .A2(n12607), .ZN(P1_U2962) );
  AOI22_X1 U15711 ( .A1(n19786), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19785), .ZN(n12610) );
  NAND2_X1 U15712 ( .A1(n12610), .A2(n12609), .ZN(P1_U2958) );
  NOR2_X1 U15713 ( .A1(n12612), .A2(n12611), .ZN(n12613) );
  OR2_X1 U15714 ( .A1(n12619), .A2(n12613), .ZN(n19835) );
  INV_X1 U15715 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12614) );
  OAI222_X1 U15716 ( .A1(n19835), .A2(n13698), .B1(n12614), .B2(n19728), .C1(
        n13696), .C2(n19805), .ZN(P1_U2870) );
  OAI21_X1 U15717 ( .B1(n12617), .B2(n12616), .A(n12615), .ZN(n12921) );
  OR2_X1 U15718 ( .A1(n12619), .A2(n12618), .ZN(n12620) );
  AND2_X1 U15719 ( .A1(n19690), .A2(n12620), .ZN(n19824) );
  INV_X1 U15720 ( .A(n19728), .ZN(n13694) );
  AOI22_X1 U15721 ( .A1(n19725), .A2(n19824), .B1(n13694), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n12621) );
  OAI21_X1 U15722 ( .B1(n12921), .B2(n13696), .A(n12621), .ZN(P1_U2869) );
  OAI211_X1 U15723 ( .C1(n9906), .C2(n10416), .A(n14344), .B(n12623), .ZN(
        n12629) );
  NAND2_X1 U15724 ( .A1(n12625), .A2(n12624), .ZN(n12627) );
  INV_X1 U15725 ( .A(n12847), .ZN(n12626) );
  AND2_X1 U15726 ( .A1(n12627), .A2(n12626), .ZN(n18632) );
  NAND2_X1 U15727 ( .A1(n14350), .A2(n18632), .ZN(n12628) );
  OAI211_X1 U15728 ( .C1(n14333), .C2(n9978), .A(n12629), .B(n12628), .ZN(
        P2_U2878) );
  NOR2_X1 U15729 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20400), .ZN(n12650) );
  MUX2_X1 U15730 ( .A(n12630), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15360), .Z(n15368) );
  AOI22_X1 U15731 ( .A1(n12650), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20400), .B2(n15368), .ZN(n12645) );
  OR2_X1 U15732 ( .A1(n20230), .A2(n14118), .ZN(n12643) );
  XNOR2_X1 U15733 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12639) );
  XNOR2_X1 U15734 ( .A(n14110), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14131) );
  NAND2_X1 U15735 ( .A1(n12632), .A2(n14131), .ZN(n12638) );
  INV_X1 U15736 ( .A(n14131), .ZN(n12633) );
  NAND2_X1 U15737 ( .A1(n12634), .A2(n12633), .ZN(n12635) );
  OR2_X1 U15738 ( .A1(n12636), .A2(n12635), .ZN(n12637) );
  OAI211_X1 U15739 ( .C1(n12640), .C2(n12639), .A(n12638), .B(n12637), .ZN(
        n12641) );
  INV_X1 U15740 ( .A(n12641), .ZN(n12642) );
  NAND2_X1 U15741 ( .A1(n12643), .A2(n12642), .ZN(n14129) );
  MUX2_X1 U15742 ( .A(n14129), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15360), .Z(n15364) );
  AOI22_X1 U15743 ( .A1(n15364), .A2(n20400), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n12650), .ZN(n12644) );
  OR2_X1 U15744 ( .A1(n12645), .A2(n12644), .ZN(n15375) );
  OR2_X1 U15745 ( .A1(n15375), .A2(n14111), .ZN(n12653) );
  AOI21_X1 U15746 ( .B1(n19697), .B2(n12646), .A(n15360), .ZN(n12647) );
  AOI211_X1 U15747 ( .C1(n15360), .C2(n12648), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n12647), .ZN(n12649) );
  AOI21_X1 U15748 ( .B1(n12650), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n12649), .ZN(n15377) );
  AND3_X1 U15749 ( .A1(n12653), .A2(n15377), .A3(n19617), .ZN(n12652) );
  NAND2_X1 U15750 ( .A1(n11260), .A2(n20400), .ZN(n20494) );
  AND3_X1 U15751 ( .A1(n12653), .A2(n15377), .A3(n15660), .ZN(n15382) );
  NAND2_X1 U15752 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20232), .ZN(n12702) );
  INV_X1 U15753 ( .A(n12702), .ZN(n12654) );
  OAI22_X1 U15754 ( .A1(n19931), .A2(n20346), .B1(n12655), .B2(n12654), .ZN(
        n12656) );
  OAI21_X1 U15755 ( .B1(n15382), .B2(n12656), .A(n19847), .ZN(n12657) );
  OAI21_X1 U15756 ( .B1(n19847), .B2(n20259), .A(n12657), .ZN(P1_U3478) );
  INV_X1 U15757 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19753) );
  OAI222_X1 U15758 ( .A1(n12921), .A2(n13777), .B1(n13766), .B2(n19880), .C1(
        n13764), .C2(n19753), .ZN(P1_U2901) );
  OR2_X1 U15759 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  NAND2_X1 U15760 ( .A1(n12660), .A2(n12668), .ZN(n19546) );
  XOR2_X1 U15761 ( .A(n19546), .B(n19160), .Z(n18743) );
  INV_X1 U15762 ( .A(n19555), .ZN(n12667) );
  NAND2_X1 U15763 ( .A1(n12662), .A2(n12661), .ZN(n12664) );
  NAND2_X1 U15764 ( .A1(n12664), .A2(n10060), .ZN(n19558) );
  XNOR2_X1 U15765 ( .A(n12666), .B(n12665), .ZN(n19568) );
  XNOR2_X1 U15766 ( .A(n19563), .B(n19568), .ZN(n18760) );
  NAND2_X1 U15767 ( .A1(n18760), .A2(n18759), .ZN(n18758) );
  OAI21_X1 U15768 ( .B1(n19568), .B2(n19565), .A(n18758), .ZN(n18750) );
  XNOR2_X1 U15769 ( .A(n19555), .B(n19558), .ZN(n18751) );
  NAND2_X1 U15770 ( .A1(n18750), .A2(n18751), .ZN(n18749) );
  OAI21_X1 U15771 ( .B1(n12667), .B2(n19558), .A(n18749), .ZN(n18742) );
  NAND2_X1 U15772 ( .A1(n18743), .A2(n18742), .ZN(n18741) );
  NAND2_X1 U15773 ( .A1(n19160), .A2(n19546), .ZN(n12671) );
  INV_X1 U15774 ( .A(n12668), .ZN(n12669) );
  XNOR2_X1 U15775 ( .A(n12670), .B(n12669), .ZN(n14893) );
  AOI21_X1 U15776 ( .B1(n18741), .B2(n12671), .A(n14893), .ZN(n18735) );
  OAI21_X1 U15777 ( .B1(n12673), .B2(n12672), .A(n12476), .ZN(n18734) );
  XNOR2_X1 U15778 ( .A(n18735), .B(n18734), .ZN(n12676) );
  INV_X1 U15779 ( .A(n18761), .ZN(n18733) );
  AOI22_X1 U15780 ( .A1(n18757), .A2(n14893), .B1(n18756), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U15781 ( .A1(n18747), .A2(n15720), .ZN(n12674) );
  OAI211_X1 U15782 ( .C1(n12676), .C2(n18733), .A(n12675), .B(n12674), .ZN(
        P2_U2915) );
  INV_X1 U15783 ( .A(n12677), .ZN(n12678) );
  OR2_X1 U15784 ( .A1(n12679), .A2(n12678), .ZN(n12680) );
  INV_X1 U15785 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19841) );
  XNOR2_X1 U15786 ( .A(n12687), .B(n19841), .ZN(n19801) );
  XNOR2_X1 U15787 ( .A(n12691), .B(n12690), .ZN(n12684) );
  INV_X1 U15788 ( .A(n12682), .ZN(n12683) );
  AOI21_X1 U15789 ( .B1(n12684), .B2(n13140), .A(n12683), .ZN(n12685) );
  NAND2_X1 U15790 ( .A1(n12686), .A2(n12685), .ZN(n19800) );
  NAND2_X1 U15791 ( .A1(n19801), .A2(n19800), .ZN(n19803) );
  NAND2_X1 U15792 ( .A1(n12687), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12688) );
  XNOR2_X1 U15793 ( .A(n13096), .B(n19828), .ZN(n12697) );
  OR2_X1 U15794 ( .A1(n20107), .A2(n12689), .ZN(n12695) );
  NAND2_X1 U15795 ( .A1(n12691), .A2(n12690), .ZN(n13110) );
  INV_X1 U15796 ( .A(n13107), .ZN(n12692) );
  XNOR2_X1 U15797 ( .A(n13110), .B(n12692), .ZN(n12693) );
  NAND2_X1 U15798 ( .A1(n12693), .A2(n13140), .ZN(n12694) );
  NAND2_X1 U15799 ( .A1(n12695), .A2(n12694), .ZN(n12696) );
  OAI21_X1 U15800 ( .B1(n12697), .B2(n12696), .A(n13098), .ZN(n19821) );
  INV_X1 U15801 ( .A(n12921), .ZN(n12700) );
  AOI22_X1 U15802 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n12698) );
  OAI21_X1 U15803 ( .B1(n19810), .B2(n12912), .A(n12698), .ZN(n12699) );
  AOI21_X1 U15804 ( .B1(n12700), .B2(n19794), .A(n12699), .ZN(n12701) );
  OAI21_X1 U15805 ( .B1(n19821), .B2(n19804), .A(n12701), .ZN(P1_U2996) );
  NAND2_X1 U15806 ( .A1(n19847), .A2(n12702), .ZN(n12877) );
  NAND2_X1 U15807 ( .A1(n19847), .A2(n20348), .ZN(n12872) );
  NAND2_X1 U15808 ( .A1(n19932), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20198) );
  XNOR2_X1 U15809 ( .A(n20105), .B(n20198), .ZN(n12703) );
  OAI222_X1 U15810 ( .A1(n12877), .A2(n20230), .B1(n19847), .B2(n20226), .C1(
        n12872), .C2(n12703), .ZN(P1_U3476) );
  NAND2_X1 U15811 ( .A1(n12719), .A2(n13035), .ZN(n12721) );
  NOR2_X2 U15812 ( .A1(n12720), .A2(n12721), .ZN(n18950) );
  INV_X1 U15813 ( .A(n13035), .ZN(n18690) );
  INV_X1 U15814 ( .A(n12733), .ZN(n12704) );
  AND2_X1 U15815 ( .A1(n18830), .A2(n12704), .ZN(n12705) );
  INV_X1 U15817 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12711) );
  INV_X1 U15818 ( .A(n12726), .ZN(n12707) );
  AND2_X1 U15819 ( .A1(n18830), .A2(n12707), .ZN(n12708) );
  OAI211_X1 U15820 ( .C1(n19404), .C2(n12711), .A(n12710), .B(n19592), .ZN(
        n12712) );
  AOI21_X1 U15821 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18950), .A(
        n12712), .ZN(n12718) );
  NOR2_X2 U15822 ( .A1(n12720), .A2(n12726), .ZN(n18922) );
  AOI22_X1 U15823 ( .A1(n19044), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18922), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15824 ( .A1(n12713), .A2(n13035), .ZN(n12736) );
  INV_X1 U15825 ( .A(n12736), .ZN(n12714) );
  INV_X1 U15826 ( .A(n18830), .ZN(n13001) );
  NAND2_X1 U15827 ( .A1(n13232), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12716) );
  NAND2_X1 U15828 ( .A1(n13233), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12715) );
  OR2_X1 U15829 ( .A1(n12719), .A2(n18690), .ZN(n12722) );
  NOR2_X2 U15830 ( .A1(n12720), .A2(n12722), .ZN(n18869) );
  NOR2_X2 U15831 ( .A1(n12720), .A2(n12733), .ZN(n18983) );
  AOI22_X1 U15832 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18869), .B1(
        n18983), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15833 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19070), .B1(
        n19010), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U15834 ( .A1(n18830), .A2(n12719), .ZN(n12723) );
  NOR2_X1 U15835 ( .A1(n13224), .A2(n12724), .ZN(n12732) );
  INV_X1 U15836 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12730) );
  NOR2_X1 U15837 ( .A1(n18830), .A2(n12733), .ZN(n12725) );
  NAND2_X1 U15838 ( .A1(n12728), .A2(n12725), .ZN(n19223) );
  NOR2_X1 U15839 ( .A1(n18830), .A2(n12726), .ZN(n12727) );
  NAND2_X1 U15840 ( .A1(n12728), .A2(n12727), .ZN(n13217) );
  OAI22_X1 U15841 ( .A1(n12730), .A2(n19223), .B1(n13217), .B2(n12729), .ZN(
        n12731) );
  NOR2_X1 U15842 ( .A1(n12732), .A2(n12731), .ZN(n12739) );
  NAND2_X1 U15843 ( .A1(n12734), .A2(n18830), .ZN(n12735) );
  AOI22_X1 U15844 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13216), .B1(
        n12737), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12738) );
  NAND2_X1 U15845 ( .A1(n12745), .A2(n12744), .ZN(n12746) );
  AOI22_X1 U15846 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18869), .B1(
        n19044), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15847 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18983), .B1(
        n19070), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U15848 ( .A1(n13232), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12748) );
  NAND2_X1 U15849 ( .A1(n13233), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12747) );
  AOI22_X1 U15850 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13216), .B1(
        n19010), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15851 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18950), .B1(
        n18922), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12763) );
  INV_X1 U15852 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12752) );
  INV_X1 U15853 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12751) );
  OAI22_X1 U15854 ( .A1(n12752), .A2(n19404), .B1(n19223), .B2(n12751), .ZN(
        n12757) );
  OAI22_X1 U15855 ( .A1(n12755), .A2(n13217), .B1(n12753), .B2(n12754), .ZN(
        n12756) );
  NOR2_X1 U15856 ( .A1(n12757), .A2(n12756), .ZN(n12762) );
  INV_X1 U15857 ( .A(n12760), .ZN(n12761) );
  INV_X1 U15858 ( .A(n12765), .ZN(n12766) );
  NAND2_X1 U15859 ( .A1(n12766), .A2(n13275), .ZN(n12767) );
  INV_X1 U15860 ( .A(n12768), .ZN(n12771) );
  INV_X1 U15861 ( .A(n12769), .ZN(n12770) );
  NAND2_X1 U15862 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  NAND2_X1 U15863 ( .A1(n9965), .A2(n12775), .ZN(n12941) );
  OAI21_X1 U15864 ( .B1(n12997), .B2(n12828), .A(n18825), .ZN(n13241) );
  XNOR2_X1 U15865 ( .A(n13241), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12776) );
  XNOR2_X1 U15866 ( .A(n13242), .B(n12776), .ZN(n15830) );
  INV_X1 U15867 ( .A(n15830), .ZN(n12838) );
  NAND2_X1 U15868 ( .A1(n12777), .A2(n12783), .ZN(n12797) );
  OAI21_X1 U15869 ( .B1(n12780), .B2(n12779), .A(n12778), .ZN(n12781) );
  INV_X1 U15870 ( .A(n12781), .ZN(n12782) );
  NAND2_X1 U15871 ( .A1(n13042), .A2(n12782), .ZN(n12796) );
  NAND2_X1 U15872 ( .A1(n12790), .A2(n12783), .ZN(n12784) );
  NOR2_X1 U15873 ( .A1(n12784), .A2(n12787), .ZN(n12785) );
  NOR2_X1 U15874 ( .A1(n12786), .A2(n12785), .ZN(n13038) );
  NAND2_X1 U15875 ( .A1(n12787), .A2(n19592), .ZN(n12791) );
  INV_X1 U15876 ( .A(n12788), .ZN(n12789) );
  NAND4_X1 U15877 ( .A1(n12791), .A2(n12790), .A3(n19602), .A4(n12789), .ZN(
        n12792) );
  NAND2_X1 U15878 ( .A1(n13038), .A2(n12792), .ZN(n12794) );
  NOR2_X1 U15879 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  OAI211_X1 U15880 ( .C1(n12797), .C2(n13042), .A(n12796), .B(n12795), .ZN(
        n12799) );
  NOR2_X1 U15881 ( .A1(n15941), .A2(n12939), .ZN(n19582) );
  INV_X1 U15882 ( .A(n15946), .ZN(n14913) );
  NAND2_X1 U15883 ( .A1(n15945), .A2(n19592), .ZN(n12800) );
  NAND2_X1 U15884 ( .A1(n14913), .A2(n12800), .ZN(n12801) );
  NAND2_X1 U15885 ( .A1(n14912), .A2(n13275), .ZN(n12802) );
  NAND2_X1 U15886 ( .A1(n12803), .A2(n12802), .ZN(n12804) );
  OAI22_X1 U15887 ( .A1(n19546), .A2(n18832), .B1(n9935), .B2(n15894), .ZN(
        n12827) );
  INV_X1 U15888 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19489) );
  AOI21_X1 U15889 ( .B1(n12806), .B2(n12805), .A(n19594), .ZN(n12816) );
  NAND2_X1 U15890 ( .A1(n12807), .A2(n19592), .ZN(n13031) );
  NAND2_X1 U15891 ( .A1(n13031), .A2(n12808), .ZN(n12809) );
  NAND2_X1 U15892 ( .A1(n12809), .A2(n18888), .ZN(n12814) );
  OAI22_X1 U15893 ( .A1(n10832), .A2(n18892), .B1(n18884), .B2(n18868), .ZN(
        n12810) );
  INV_X1 U15894 ( .A(n12810), .ZN(n12811) );
  AND2_X1 U15895 ( .A1(n12812), .A2(n12811), .ZN(n12813) );
  OAI211_X1 U15896 ( .C1(n12816), .C2(n12815), .A(n12814), .B(n12813), .ZN(
        n12817) );
  OR2_X1 U15897 ( .A1(n12818), .A2(n12817), .ZN(n14940) );
  NAND2_X1 U15898 ( .A1(n14904), .A2(n12819), .ZN(n12820) );
  NAND2_X1 U15899 ( .A1(n12834), .A2(n12820), .ZN(n14789) );
  INV_X1 U15900 ( .A(n14789), .ZN(n12822) );
  NAND2_X1 U15901 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18855) );
  NOR2_X1 U15902 ( .A1(n12828), .A2(n18855), .ZN(n18837) );
  INV_X1 U15903 ( .A(n15948), .ZN(n12821) );
  NAND2_X1 U15904 ( .A1(n12828), .A2(n18855), .ZN(n12823) );
  AOI22_X1 U15905 ( .A1(n12822), .A2(n18837), .B1(n18836), .B2(n12823), .ZN(
        n14615) );
  INV_X1 U15906 ( .A(n12823), .ZN(n18838) );
  NOR2_X1 U15907 ( .A1(n14789), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18823) );
  INV_X1 U15908 ( .A(n18855), .ZN(n18822) );
  INV_X1 U15909 ( .A(n12834), .ZN(n12824) );
  NAND2_X1 U15910 ( .A1(n12824), .A2(n15908), .ZN(n18851) );
  OAI21_X1 U15911 ( .B1(n14789), .B2(n18822), .A(n18851), .ZN(n18835) );
  AOI211_X1 U15912 ( .C1(n18836), .C2(n18838), .A(n18823), .B(n18835), .ZN(
        n14606) );
  MUX2_X1 U15913 ( .A(n14615), .B(n14606), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n12825) );
  OAI21_X1 U15914 ( .B1(n19489), .B2(n15908), .A(n12825), .ZN(n12826) );
  NOR2_X1 U15915 ( .A1(n12827), .A2(n12826), .ZN(n12837) );
  OR2_X1 U15916 ( .A1(n12829), .A2(n12828), .ZN(n12830) );
  OAI21_X1 U15917 ( .B1(n12832), .B2(n12831), .A(n12830), .ZN(n13403) );
  XNOR2_X1 U15918 ( .A(n13403), .B(n14614), .ZN(n12835) );
  OR2_X1 U15919 ( .A1(n9704), .A2(n12835), .ZN(n15826) );
  INV_X1 U15920 ( .A(n12833), .ZN(n19584) );
  NAND3_X1 U15921 ( .A1(n15826), .A2(n18846), .A3(n15825), .ZN(n12836) );
  OAI211_X1 U15922 ( .C1(n12838), .C2(n15926), .A(n12837), .B(n12836), .ZN(
        P2_U3043) );
  INV_X1 U15923 ( .A(n20110), .ZN(n12843) );
  INV_X1 U15924 ( .A(n12872), .ZN(n12841) );
  NOR2_X1 U15925 ( .A1(n20290), .A2(n20198), .ZN(n20341) );
  AOI211_X1 U15926 ( .C1(n20107), .C2(n20198), .A(n20341), .B(n19964), .ZN(
        n12840) );
  INV_X1 U15927 ( .A(n19847), .ZN(n12875) );
  AOI22_X1 U15928 ( .A1(n12841), .A2(n12840), .B1(n12875), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12842) );
  OAI21_X1 U15929 ( .B1(n12843), .B2(n12877), .A(n12842), .ZN(P1_U3475) );
  OAI21_X1 U15930 ( .B1(n12845), .B2(n12844), .A(n13012), .ZN(n15559) );
  INV_X1 U15931 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19749) );
  OAI222_X1 U15932 ( .A1(n15559), .A2(n13777), .B1(n13766), .B2(n19888), .C1(
        n13764), .C2(n19749), .ZN(P1_U2899) );
  INV_X1 U15933 ( .A(n19692), .ZN(n15641) );
  XNOR2_X1 U15934 ( .A(n15641), .B(n15640), .ZN(n19674) );
  INV_X1 U15935 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12846) );
  OAI222_X1 U15936 ( .A1(n15559), .A2(n13696), .B1(n13698), .B2(n19674), .C1(
        n19728), .C2(n12846), .ZN(P1_U2867) );
  NOR2_X1 U15937 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  NOR2_X1 U15938 ( .A1(n12866), .A2(n12849), .ZN(n18618) );
  NOR2_X1 U15939 ( .A1(n14333), .A2(n12026), .ZN(n12853) );
  AOI211_X1 U15940 ( .C1(n12851), .C2(n12623), .A(n14342), .B(n12850), .ZN(
        n12852) );
  AOI211_X1 U15941 ( .C1(n18618), .C2(n14350), .A(n12853), .B(n12852), .ZN(
        n12854) );
  INV_X1 U15942 ( .A(n12854), .ZN(P2_U2877) );
  INV_X1 U15943 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19751) );
  INV_X1 U15944 ( .A(n12855), .ZN(n12856) );
  XNOR2_X1 U15945 ( .A(n12615), .B(n12856), .ZN(n19793) );
  INV_X1 U15946 ( .A(n19793), .ZN(n12857) );
  OAI222_X1 U15947 ( .A1(n13764), .A2(n19751), .B1(n13766), .B2(n19884), .C1(
        n13777), .C2(n12857), .ZN(P1_U2900) );
  XNOR2_X1 U15948 ( .A(n12858), .B(n12986), .ZN(n12862) );
  NAND2_X1 U15949 ( .A1(n12867), .A2(n12859), .ZN(n12860) );
  NAND2_X1 U15950 ( .A1(n12989), .A2(n12860), .ZN(n15875) );
  MUX2_X1 U15951 ( .A(n15875), .B(n12967), .S(n14340), .Z(n12861) );
  OAI21_X1 U15952 ( .B1(n12862), .B2(n14342), .A(n12861), .ZN(P2_U2875) );
  INV_X1 U15953 ( .A(n12858), .ZN(n12863) );
  OAI211_X1 U15954 ( .C1(n12850), .C2(n12864), .A(n12863), .B(n14344), .ZN(
        n12870) );
  OR2_X1 U15955 ( .A1(n12866), .A2(n12865), .ZN(n12868) );
  AND2_X1 U15956 ( .A1(n12868), .A2(n12867), .ZN(n18609) );
  NAND2_X1 U15957 ( .A1(n18609), .A2(n14350), .ZN(n12869) );
  OAI211_X1 U15958 ( .C1(n14333), .C2(n12059), .A(n12870), .B(n12869), .ZN(
        P2_U2876) );
  INV_X1 U15959 ( .A(n19932), .ZN(n12873) );
  INV_X1 U15960 ( .A(n20198), .ZN(n19963) );
  AOI211_X1 U15961 ( .C1(n12873), .C2(n20291), .A(n19963), .B(n12872), .ZN(
        n12874) );
  AOI21_X1 U15962 ( .B1(n12875), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n12874), .ZN(n12876) );
  OAI21_X1 U15963 ( .B1(n20111), .B2(n12877), .A(n12876), .ZN(P1_U3477) );
  INV_X1 U15964 ( .A(n20494), .ZN(n15389) );
  NAND2_X1 U15965 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15389), .ZN(n15385) );
  NAND2_X1 U15966 ( .A1(n12878), .A2(n20499), .ZN(n12879) );
  OAI211_X1 U15967 ( .C1(n15385), .C2(n20401), .A(n15601), .B(n12879), .ZN(
        n12880) );
  INV_X1 U15968 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13482) );
  NOR2_X1 U15969 ( .A1(n13208), .A2(n20400), .ZN(n12883) );
  INV_X1 U15970 ( .A(n12887), .ZN(n12884) );
  NAND2_X1 U15971 ( .A1(n12884), .A2(n13462), .ZN(n12885) );
  NAND2_X1 U15972 ( .A1(n15480), .A2(n12885), .ZN(n19698) );
  NOR2_X1 U15973 ( .A1(n12887), .A2(n12886), .ZN(n19717) );
  INV_X1 U15974 ( .A(n19717), .ZN(n12907) );
  NOR2_X1 U15975 ( .A1(n12888), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12896) );
  INV_X1 U15976 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20476) );
  NAND2_X1 U15977 ( .A1(n12889), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12894) );
  AND2_X1 U15978 ( .A1(n20415), .A2(n20291), .ZN(n12890) );
  NOR2_X1 U15979 ( .A1(n12894), .A2(n12890), .ZN(n12891) );
  INV_X1 U15980 ( .A(n12892), .ZN(n12893) );
  AOI22_X1 U15981 ( .A1(n19709), .A2(n20476), .B1(n19707), .B2(n12893), .ZN(
        n12906) );
  INV_X1 U15982 ( .A(n12894), .ZN(n12895) );
  NOR2_X1 U15983 ( .A1(n12896), .A2(n12895), .ZN(n12897) );
  INV_X1 U15984 ( .A(n19646), .ZN(n19705) );
  AOI22_X1 U15985 ( .A1(n19641), .A2(n12900), .B1(n19705), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n12902) );
  NAND2_X1 U15986 ( .A1(n19710), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12901) );
  OAI211_X1 U15987 ( .C1(n19695), .C2(n12903), .A(n12902), .B(n12901), .ZN(
        n12904) );
  INV_X1 U15988 ( .A(n12904), .ZN(n12905) );
  OAI211_X1 U15989 ( .C1(n20111), .C2(n12907), .A(n12906), .B(n12905), .ZN(
        n12908) );
  INV_X1 U15990 ( .A(n12908), .ZN(n12909) );
  OAI21_X1 U15991 ( .B1(n12910), .B2(n19714), .A(n12909), .ZN(P1_U2839) );
  OAI221_X1 U15992 ( .B1(n19678), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n19678), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n19646), .ZN(n12911) );
  AOI22_X1 U15993 ( .A1(n19710), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n12911), .ZN(n12915) );
  INV_X1 U15994 ( .A(n12912), .ZN(n12913) );
  NAND2_X1 U15995 ( .A1(n19641), .A2(n12913), .ZN(n12914) );
  OAI211_X1 U15996 ( .C1(n19695), .C2(n11922), .A(n12915), .B(n12914), .ZN(
        n12918) );
  INV_X1 U15997 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n12916) );
  NOR4_X1 U15998 ( .A1(n19678), .A2(P1_REIP_REG_3__SCAN_IN), .A3(n12916), .A4(
        n20476), .ZN(n12917) );
  AOI211_X1 U15999 ( .C1(n19824), .C2(n19707), .A(n12918), .B(n12917), .ZN(
        n12920) );
  NAND2_X1 U16000 ( .A1(n20110), .A2(n19717), .ZN(n12919) );
  OAI211_X1 U16001 ( .C1(n12921), .C2(n19714), .A(n12920), .B(n12919), .ZN(
        P1_U2837) );
  INV_X1 U16002 ( .A(n18691), .ZN(n13449) );
  AOI21_X1 U16003 ( .B1(n15834), .B2(n12922), .A(n12955), .ZN(n15823) );
  INV_X1 U16004 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14622) );
  INV_X1 U16005 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18522) );
  INV_X1 U16006 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14543) );
  INV_X1 U16007 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14145) );
  INV_X1 U16008 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20563) );
  INV_X1 U16009 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14487) );
  INV_X1 U16010 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14155) );
  INV_X1 U16011 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14469) );
  INV_X1 U16012 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20511) );
  OAI22_X4 U16013 ( .A1(n15967), .A2(n14622), .B1(n13402), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n18669) );
  OAI22_X1 U16014 ( .A1(n15967), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n14245) );
  INV_X1 U16015 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14237) );
  OAI22_X1 U16016 ( .A1(n15967), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14237), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14244) );
  AND2_X1 U16017 ( .A1(n14245), .A2(n14244), .ZN(n12993) );
  NAND2_X1 U16018 ( .A1(n12993), .A2(n12994), .ZN(n12953) );
  NAND2_X1 U16019 ( .A1(n18669), .A2(n12953), .ZN(n12924) );
  XNOR2_X1 U16020 ( .A(n15823), .B(n12924), .ZN(n12925) );
  INV_X1 U16021 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n18921) );
  INV_X1 U16022 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19072) );
  NAND4_X1 U16023 ( .A1(n18921), .A2(n15967), .A3(n19072), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19465) );
  NAND2_X1 U16024 ( .A1(n12925), .A2(n18678), .ZN(n12947) );
  NAND2_X1 U16025 ( .A1(n19072), .A2(n19602), .ZN(n12937) );
  NOR2_X1 U16026 ( .A1(n12939), .A2(n12937), .ZN(n12926) );
  NOR2_X1 U16027 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13043), .ZN(n12934) );
  AND2_X1 U16028 ( .A1(n13275), .A2(n12934), .ZN(n12927) );
  AND2_X1 U16029 ( .A1(n10314), .A2(n12927), .ZN(n15964) );
  NOR2_X1 U16030 ( .A1(n19571), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19011) );
  INV_X1 U16031 ( .A(n19011), .ZN(n12929) );
  NOR2_X1 U16032 ( .A1(n12930), .A2(n12929), .ZN(n15959) );
  INV_X1 U16033 ( .A(n15959), .ZN(n12931) );
  INV_X2 U16034 ( .A(n18815), .ZN(n18662) );
  NAND3_X1 U16035 ( .A1(n12931), .A2(n18662), .A3(n19465), .ZN(n12932) );
  NAND2_X1 U16036 ( .A1(n18681), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18663) );
  NOR2_X1 U16037 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12933), .ZN(n12936) );
  NOR2_X1 U16038 ( .A1(n12935), .A2(n12934), .ZN(n14165) );
  AOI21_X2 U16039 ( .B1(n12937), .B2(n12936), .A(n14165), .ZN(n18679) );
  OAI22_X1 U16040 ( .A1(n18679), .A2(n10330), .B1(n19489), .B2(n18681), .ZN(
        n12943) );
  NAND2_X1 U16041 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12937), .ZN(n12938) );
  NOR2_X1 U16042 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  NOR2_X1 U16043 ( .A1(n12941), .A2(n18687), .ZN(n12942) );
  AOI211_X1 U16044 ( .C1(n18677), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n12943), .B(n12942), .ZN(n12944) );
  OAI21_X1 U16045 ( .B1(n19546), .B2(n18676), .A(n12944), .ZN(n12945) );
  AOI21_X1 U16046 ( .B1(n12728), .B2(n18689), .A(n12945), .ZN(n12946) );
  OAI211_X1 U16047 ( .C1(n19160), .C2(n13449), .A(n12947), .B(n12946), .ZN(
        P2_U2852) );
  MUX2_X1 U16048 ( .A(n12949), .B(n12948), .S(n18899), .Z(n13245) );
  MUX2_X1 U16049 ( .A(n13238), .B(P2_EBX_REG_5__SCAN_IN), .S(n18899), .Z(
        n13240) );
  MUX2_X1 U16050 ( .A(n13276), .B(P2_EBX_REG_6__SCAN_IN), .S(n18899), .Z(
        n13279) );
  MUX2_X1 U16051 ( .A(n13426), .B(n12950), .S(n18899), .Z(n13285) );
  NAND2_X1 U16052 ( .A1(n18899), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U16053 ( .A1(n9970), .A2(n9660), .ZN(n12952) );
  NAND2_X1 U16054 ( .A1(n13312), .A2(n12952), .ZN(n13309) );
  AOI21_X1 U16055 ( .B1(n18602), .B2(n12960), .A(n12962), .ZN(n18608) );
  AOI21_X1 U16056 ( .B1(n18625), .B2(n12958), .A(n12961), .ZN(n18631) );
  AOI21_X1 U16057 ( .B1(n14594), .B2(n12956), .A(n12959), .ZN(n18637) );
  AOI21_X1 U16058 ( .B1(n15822), .B2(n12954), .A(n12957), .ZN(n18671) );
  NOR2_X1 U16059 ( .A1(n15823), .A2(n12953), .ZN(n13438) );
  OAI21_X1 U16060 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12955), .A(
        n12954), .ZN(n18805) );
  NAND2_X1 U16061 ( .A1(n13438), .A2(n18805), .ZN(n18668) );
  NOR2_X1 U16062 ( .A1(n18671), .A2(n18668), .ZN(n18652) );
  OAI21_X1 U16063 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12957), .A(
        n12956), .ZN(n18655) );
  NAND2_X1 U16064 ( .A1(n18652), .A2(n18655), .ZN(n18636) );
  NOR2_X1 U16065 ( .A1(n18637), .A2(n18636), .ZN(n12975) );
  OAI21_X1 U16066 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12959), .A(
        n12958), .ZN(n15813) );
  NAND2_X1 U16067 ( .A1(n12975), .A2(n15813), .ZN(n18629) );
  NOR2_X1 U16068 ( .A1(n18631), .A2(n18629), .ZN(n18613) );
  OAI21_X1 U16069 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12961), .A(
        n12960), .ZN(n18615) );
  NAND2_X1 U16070 ( .A1(n18613), .A2(n18615), .ZN(n18606) );
  NOR2_X1 U16071 ( .A1(n18608), .A2(n18606), .ZN(n13017) );
  NOR2_X1 U16072 ( .A1(n18653), .A2(n13017), .ZN(n12963) );
  OAI21_X1 U16073 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12962), .A(
        n13016), .ZN(n15775) );
  XNOR2_X1 U16074 ( .A(n12963), .B(n15775), .ZN(n12964) );
  NAND2_X1 U16075 ( .A1(n12964), .A2(n18678), .ZN(n12971) );
  INV_X1 U16076 ( .A(n18676), .ZN(n18684) );
  AOI21_X1 U16077 ( .B1(n12965), .B2(n14836), .A(n14809), .ZN(n18716) );
  AOI22_X1 U16078 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18667), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18677), .ZN(n12966) );
  OAI211_X1 U16079 ( .C1(n18679), .C2(n12967), .A(n15908), .B(n12966), .ZN(
        n12969) );
  NOR2_X1 U16080 ( .A1(n15875), .A2(n18656), .ZN(n12968) );
  AOI211_X1 U16081 ( .C1(n18684), .C2(n18716), .A(n12969), .B(n12968), .ZN(
        n12970) );
  OAI211_X1 U16082 ( .C1(n18687), .C2(n13309), .A(n12971), .B(n12970), .ZN(
        P2_U2843) );
  NAND2_X1 U16083 ( .A1(n12973), .A2(n12972), .ZN(n12974) );
  NAND2_X1 U16084 ( .A1(n13294), .A2(n12974), .ZN(n13290) );
  NOR2_X1 U16085 ( .A1(n18653), .A2(n12975), .ZN(n12976) );
  XNOR2_X1 U16086 ( .A(n12976), .B(n15813), .ZN(n12977) );
  NAND2_X1 U16087 ( .A1(n12977), .A2(n18678), .ZN(n12984) );
  AOI21_X1 U16088 ( .B1(n12978), .B2(n15905), .A(n14851), .ZN(n18727) );
  AOI22_X1 U16089 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18677), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18667), .ZN(n12979) );
  OAI211_X1 U16090 ( .C1(n18679), .C2(n12980), .A(n15908), .B(n12979), .ZN(
        n12982) );
  NOR2_X1 U16091 ( .A1(n15893), .A2(n18656), .ZN(n12981) );
  AOI211_X1 U16092 ( .C1(n18684), .C2(n18727), .A(n12982), .B(n12981), .ZN(
        n12983) );
  OAI211_X1 U16093 ( .C1(n18687), .C2(n13290), .A(n12984), .B(n12983), .ZN(
        P2_U2847) );
  AOI21_X1 U16094 ( .B1(n12858), .B2(n12986), .A(n12985), .ZN(n12987) );
  OR3_X1 U16095 ( .A1(n9706), .A2(n12987), .A3(n14342), .ZN(n12992) );
  AND2_X1 U16096 ( .A1(n12989), .A2(n12988), .ZN(n12990) );
  OR2_X1 U16097 ( .A1(n12990), .A2(n9683), .ZN(n14814) );
  INV_X1 U16098 ( .A(n14814), .ZN(n18598) );
  NAND2_X1 U16099 ( .A1(n18598), .A2(n14350), .ZN(n12991) );
  OAI211_X1 U16100 ( .C1(n14350), .C2(n12064), .A(n12992), .B(n12991), .ZN(
        P2_U2874) );
  NOR2_X1 U16101 ( .A1(n18653), .A2(n12993), .ZN(n14243) );
  XNOR2_X1 U16102 ( .A(n14243), .B(n12994), .ZN(n12995) );
  NAND2_X1 U16103 ( .A1(n12995), .A2(n18678), .ZN(n13004) );
  OAI22_X1 U16104 ( .A1(n18679), .A2(n12996), .B1(n19488), .B2(n18681), .ZN(
        n12999) );
  NOR2_X1 U16105 ( .A1(n18687), .A2(n12997), .ZN(n12998) );
  AOI211_X1 U16106 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n18677), .A(
        n12999), .B(n12998), .ZN(n13000) );
  OAI21_X1 U16107 ( .B1(n13001), .B2(n18656), .A(n13000), .ZN(n13002) );
  AOI21_X1 U16108 ( .B1(n19558), .B2(n18684), .A(n13002), .ZN(n13003) );
  OAI211_X1 U16109 ( .C1(n13449), .C2(n19555), .A(n13004), .B(n13003), .ZN(
        P2_U2853) );
  NAND2_X1 U16110 ( .A1(n13006), .A2(n13005), .ZN(n13007) );
  AND2_X1 U16111 ( .A1(n13062), .A2(n13007), .ZN(n19647) );
  INV_X1 U16112 ( .A(n19647), .ZN(n13010) );
  INV_X1 U16113 ( .A(n13065), .ZN(n13008) );
  XNOR2_X1 U16114 ( .A(n15642), .B(n13008), .ZN(n19654) );
  INV_X1 U16115 ( .A(n19654), .ZN(n13009) );
  INV_X1 U16116 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19652) );
  OAI222_X1 U16117 ( .A1(n13010), .A2(n13696), .B1(n13698), .B2(n13009), .C1(
        n19728), .C2(n19652), .ZN(P1_U2865) );
  OAI222_X1 U16118 ( .A1(n13010), .A2(n13777), .B1(n13766), .B2(n19899), .C1(
        n13764), .C2(n11393), .ZN(P1_U2897) );
  XOR2_X1 U16119 ( .A(n13012), .B(n13011), .Z(n19722) );
  INV_X1 U16120 ( .A(n19722), .ZN(n13013) );
  OAI222_X1 U16121 ( .A1(n13764), .A2(n19747), .B1(n13766), .B2(n19891), .C1(
        n13777), .C2(n13013), .ZN(P1_U2898) );
  OR2_X1 U16122 ( .A1(n9683), .A2(n13014), .ZN(n13015) );
  AND2_X1 U16123 ( .A1(n13015), .A2(n13085), .ZN(n15763) );
  AOI21_X1 U16124 ( .B1(n18591), .B2(n13016), .A(n9678), .ZN(n18597) );
  NAND2_X1 U16125 ( .A1(n13017), .A2(n15775), .ZN(n18595) );
  NOR2_X1 U16126 ( .A1(n18597), .A2(n18595), .ZN(n14148) );
  NOR2_X1 U16127 ( .A1(n18653), .A2(n14148), .ZN(n13018) );
  OAI21_X1 U16128 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9678), .A(
        n14146), .ZN(n15766) );
  XNOR2_X1 U16129 ( .A(n13018), .B(n15766), .ZN(n13019) );
  NAND2_X1 U16130 ( .A1(n13019), .A2(n18678), .ZN(n13027) );
  AOI21_X1 U16131 ( .B1(n13020), .B2(n14811), .A(n9677), .ZN(n15860) );
  INV_X1 U16132 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19506) );
  XNOR2_X1 U16133 ( .A(n13314), .B(n9688), .ZN(n13349) );
  AOI22_X1 U16134 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18677), .B1(
        n18639), .B2(n13349), .ZN(n13021) );
  OAI21_X1 U16135 ( .B1(n19506), .B2(n18681), .A(n13021), .ZN(n13022) );
  INV_X1 U16136 ( .A(n13022), .ZN(n13023) );
  OAI211_X1 U16137 ( .C1(n18679), .C2(n13024), .A(n15908), .B(n13023), .ZN(
        n13025) );
  AOI21_X1 U16138 ( .B1(n18684), .B2(n15860), .A(n13025), .ZN(n13026) );
  OAI211_X1 U16139 ( .C1(n15864), .C2(n18656), .A(n13027), .B(n13026), .ZN(
        P2_U2841) );
  OAI211_X1 U16140 ( .C1(n9706), .C2(n10159), .A(n14344), .B(n13028), .ZN(
        n13030) );
  NAND2_X1 U16141 ( .A1(n14340), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13029) );
  OAI211_X1 U16142 ( .C1(n15864), .C2(n14340), .A(n13030), .B(n13029), .ZN(
        P2_U2873) );
  INV_X1 U16143 ( .A(n14912), .ZN(n14936) );
  INV_X1 U16144 ( .A(n13031), .ZN(n13032) );
  NOR2_X1 U16145 ( .A1(n13032), .A2(n12021), .ZN(n14903) );
  MUX2_X1 U16146 ( .A(n14936), .B(n14903), .S(n13033), .Z(n13034) );
  OAI21_X1 U16147 ( .B1(n13035), .B2(n14904), .A(n13034), .ZN(n15927) );
  INV_X1 U16148 ( .A(n15408), .ZN(n15965) );
  INV_X1 U16149 ( .A(n14245), .ZN(n13036) );
  AOI22_X1 U16150 ( .A1(n18653), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13036), .B2(n18669), .ZN(n14907) );
  AOI222_X1 U16151 ( .A1(n15927), .A2(n18495), .B1(n13037), .B2(n15965), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n14907), .ZN(n13053) );
  NAND2_X1 U16152 ( .A1(n13039), .A2(n13038), .ZN(n13040) );
  NOR2_X1 U16153 ( .A1(n13041), .A2(n13040), .ZN(n13047) );
  INV_X1 U16154 ( .A(n13042), .ZN(n13045) );
  NOR2_X1 U16155 ( .A1(n10815), .A2(n13043), .ZN(n13044) );
  NAND2_X1 U16156 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  AND2_X1 U16157 ( .A1(n13047), .A2(n13046), .ZN(n15958) );
  NOR2_X1 U16158 ( .A1(n15958), .A2(n19458), .ZN(n13050) );
  NOR2_X1 U16159 ( .A1(n15967), .A2(n15405), .ZN(n15962) );
  AOI21_X1 U16160 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n15967), .A(n15962), 
        .ZN(n15973) );
  AOI21_X1 U16161 ( .B1(n13048), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15973), 
        .ZN(n13049) );
  OR2_X1 U16162 ( .A1(n13050), .A2(n13049), .ZN(n15175) );
  INV_X1 U16163 ( .A(n15175), .ZN(n13052) );
  NAND2_X1 U16164 ( .A1(n13052), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13051) );
  OAI21_X1 U16165 ( .B1(n13053), .B2(n13052), .A(n13051), .ZN(P2_U3601) );
  OAI21_X1 U16166 ( .B1(n19710), .B2(n19641), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13054) );
  OAI21_X1 U16167 ( .B1(n19695), .B2(n11915), .A(n13054), .ZN(n13055) );
  AOI21_X1 U16168 ( .B1(n19707), .B2(n13056), .A(n13055), .ZN(n13057) );
  OAI21_X1 U16169 ( .B1(n13640), .B2(n20482), .A(n13057), .ZN(n13058) );
  AOI21_X1 U16170 ( .B1(n19961), .B2(n19717), .A(n13058), .ZN(n13059) );
  OAI21_X1 U16171 ( .B1(n13060), .B2(n19714), .A(n13059), .ZN(P1_U2840) );
  AOI21_X1 U16172 ( .B1(n13063), .B2(n13062), .A(n13061), .ZN(n13070) );
  AOI21_X1 U16173 ( .B1(n15642), .B2(n13065), .A(n13064), .ZN(n13066) );
  OR2_X1 U16174 ( .A1(n13093), .A2(n13066), .ZN(n13074) );
  INV_X1 U16175 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13067) );
  OAI22_X1 U16176 ( .A1(n13074), .A2(n13698), .B1(n13067), .B2(n19728), .ZN(
        n13068) );
  AOI21_X1 U16177 ( .B1(n13070), .B2(n11912), .A(n13068), .ZN(n13069) );
  INV_X1 U16178 ( .A(n13069), .ZN(P1_U2864) );
  INV_X1 U16179 ( .A(n13070), .ZN(n13149) );
  INV_X1 U16180 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20433) );
  NAND4_X1 U16181 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19677)
         );
  NAND2_X1 U16182 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19648) );
  NOR3_X1 U16183 ( .A1(n20433), .A2(n19677), .A3(n19648), .ZN(n13073) );
  NAND2_X1 U16184 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13073), .ZN(n13475) );
  NOR2_X1 U16185 ( .A1(n19705), .A2(n13475), .ZN(n13641) );
  NOR2_X1 U16186 ( .A1(n13640), .A2(n13641), .ZN(n19638) );
  NAND2_X1 U16187 ( .A1(n19646), .A2(n13071), .ZN(n19693) );
  AOI21_X1 U16188 ( .B1(n19710), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19650), .ZN(n13072) );
  OAI21_X1 U16189 ( .B1(n13145), .B2(n19713), .A(n13072), .ZN(n13078) );
  NAND2_X1 U16190 ( .A1(n19709), .A2(n13073), .ZN(n13076) );
  INV_X1 U16191 ( .A(n13074), .ZN(n15623) );
  AOI22_X1 U16192 ( .A1(n15623), .A2(n19707), .B1(n19708), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n13075) );
  OAI21_X1 U16193 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n13076), .A(n13075), .ZN(
        n13077) );
  AOI211_X1 U16194 ( .C1(n19638), .C2(P1_REIP_REG_8__SCAN_IN), .A(n13078), .B(
        n13077), .ZN(n13079) );
  OAI21_X1 U16195 ( .B1(n13149), .B2(n15480), .A(n13079), .ZN(P1_U2832) );
  INV_X1 U16196 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U16197 ( .A1(n19852), .A2(n12290), .ZN(n13080) );
  OAI21_X1 U16198 ( .B1(n19852), .B2(DATAI_8_), .A(n13080), .ZN(n13722) );
  OAI222_X1 U16199 ( .A1(n13149), .A2(n13777), .B1(n13764), .B2(n13081), .C1(
        n13722), .C2(n13766), .ZN(P1_U2896) );
  OAI211_X1 U16200 ( .C1(n10484), .C2(n10483), .A(n14344), .B(n13083), .ZN(
        n13088) );
  NAND2_X1 U16201 ( .A1(n13085), .A2(n13084), .ZN(n13086) );
  AND2_X1 U16202 ( .A1(n14346), .A2(n13086), .ZN(n15852) );
  NAND2_X1 U16203 ( .A1(n15852), .A2(n14350), .ZN(n13087) );
  OAI211_X1 U16204 ( .C1(n14350), .C2(n12071), .A(n13088), .B(n13087), .ZN(
        P2_U2872) );
  NOR2_X1 U16205 ( .A1(n13061), .A2(n13089), .ZN(n13090) );
  OR2_X1 U16206 ( .A1(n9682), .A2(n13090), .ZN(n19639) );
  INV_X1 U16207 ( .A(n13766), .ZN(n13775) );
  MUX2_X1 U16208 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n19852), .Z(
        n19765) );
  AOI22_X1 U16209 ( .A1(n13775), .A2(n19765), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n13774), .ZN(n13091) );
  OAI21_X1 U16210 ( .B1(n19639), .B2(n13777), .A(n13091), .ZN(P1_U2895) );
  OR2_X1 U16211 ( .A1(n13093), .A2(n13092), .ZN(n13094) );
  NAND2_X1 U16212 ( .A1(n13152), .A2(n13094), .ZN(n19635) );
  INV_X1 U16213 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13095) );
  OAI222_X1 U16214 ( .A1(n19635), .A2(n13698), .B1(n13095), .B2(n19728), .C1(
        n19639), .C2(n13696), .ZN(P1_U2863) );
  NAND2_X1 U16215 ( .A1(n13096), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13097) );
  NAND2_X1 U16216 ( .A1(n13099), .A2(n13133), .ZN(n13103) );
  NAND2_X1 U16217 ( .A1(n13110), .A2(n13107), .ZN(n13100) );
  XNOR2_X1 U16218 ( .A(n13100), .B(n13108), .ZN(n13101) );
  NAND2_X1 U16219 ( .A1(n13101), .A2(n13140), .ZN(n13102) );
  NAND2_X1 U16220 ( .A1(n13103), .A2(n13102), .ZN(n13104) );
  INV_X1 U16221 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19820) );
  XNOR2_X1 U16222 ( .A(n13104), .B(n19820), .ZN(n19790) );
  NAND2_X1 U16223 ( .A1(n13104), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13105) );
  NAND2_X1 U16224 ( .A1(n13106), .A2(n13133), .ZN(n13113) );
  AND2_X1 U16225 ( .A1(n13108), .A2(n13107), .ZN(n13109) );
  NAND2_X1 U16226 ( .A1(n13110), .A2(n13109), .ZN(n13127) );
  XNOR2_X1 U16227 ( .A(n13127), .B(n13125), .ZN(n13111) );
  NAND2_X1 U16228 ( .A1(n13111), .A2(n13140), .ZN(n13112) );
  NAND2_X1 U16229 ( .A1(n13113), .A2(n13112), .ZN(n13114) );
  INV_X1 U16230 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15624) );
  XNOR2_X1 U16231 ( .A(n13114), .B(n15624), .ZN(n15556) );
  NAND2_X1 U16232 ( .A1(n13114), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13115) );
  NAND3_X1 U16233 ( .A1(n13137), .A2(n13133), .A3(n13116), .ZN(n13121) );
  INV_X1 U16234 ( .A(n13127), .ZN(n13117) );
  NAND2_X1 U16235 ( .A1(n13117), .A2(n13125), .ZN(n13118) );
  XNOR2_X1 U16236 ( .A(n13118), .B(n13124), .ZN(n13119) );
  NAND2_X1 U16237 ( .A1(n13119), .A2(n13140), .ZN(n13120) );
  NAND2_X1 U16238 ( .A1(n13121), .A2(n13120), .ZN(n15550) );
  OR2_X1 U16239 ( .A1(n15550), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13122) );
  NAND2_X1 U16240 ( .A1(n13123), .A2(n13133), .ZN(n13130) );
  NAND2_X1 U16241 ( .A1(n13125), .A2(n13124), .ZN(n13126) );
  OR2_X1 U16242 ( .A1(n13127), .A2(n13126), .ZN(n13138) );
  XNOR2_X1 U16243 ( .A(n13138), .B(n13139), .ZN(n13128) );
  NAND2_X1 U16244 ( .A1(n13128), .A2(n13140), .ZN(n13129) );
  NAND2_X1 U16245 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  OR2_X1 U16246 ( .A1(n13131), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15545) );
  NAND2_X1 U16247 ( .A1(n15547), .A2(n15545), .ZN(n13132) );
  NAND2_X1 U16248 ( .A1(n13131), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15544) );
  NAND2_X1 U16249 ( .A1(n13133), .A2(n13139), .ZN(n13135) );
  NOR2_X1 U16250 ( .A1(n13135), .A2(n13134), .ZN(n13136) );
  INV_X1 U16251 ( .A(n13138), .ZN(n13141) );
  NAND3_X1 U16252 ( .A1(n13141), .A2(n13140), .A3(n13139), .ZN(n13142) );
  NAND2_X1 U16253 ( .A1(n9615), .A2(n13142), .ZN(n13163) );
  XNOR2_X1 U16254 ( .A(n13163), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13143) );
  XNOR2_X1 U16255 ( .A(n13162), .B(n13143), .ZN(n15630) );
  NAND2_X1 U16256 ( .A1(n15630), .A2(n19795), .ZN(n13148) );
  INV_X1 U16257 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13144) );
  NOR2_X1 U16258 ( .A1(n15601), .A2(n13144), .ZN(n15622) );
  NOR2_X1 U16259 ( .A1(n19810), .A2(n13145), .ZN(n13146) );
  AOI211_X1 U16260 ( .C1(n19799), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15622), .B(n13146), .ZN(n13147) );
  OAI211_X1 U16261 ( .C1(n19851), .C2(n13149), .A(n13148), .B(n13147), .ZN(
        P1_U2991) );
  OAI21_X1 U16262 ( .B1(n9682), .B2(n13150), .A(n13180), .ZN(n13928) );
  INV_X1 U16263 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20570) );
  INV_X1 U16264 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20435) );
  NOR2_X1 U16265 ( .A1(n20570), .A2(n20435), .ZN(n15491) );
  AOI21_X1 U16266 ( .B1(n15491), .B2(n13641), .A(n13640), .ZN(n15503) );
  AOI21_X1 U16267 ( .B1(n19710), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19650), .ZN(n13151) );
  OAI21_X1 U16268 ( .B1(n13924), .B2(n19713), .A(n13151), .ZN(n13157) );
  AOI21_X1 U16269 ( .B1(n13153), .B2(n13152), .A(n9850), .ZN(n15613) );
  AOI22_X1 U16270 ( .A1(n15613), .A2(n19707), .B1(n19708), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n13155) );
  NOR2_X1 U16271 ( .A1(n19678), .A2(n13475), .ZN(n19634) );
  NAND3_X1 U16272 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20570), .A3(n19634), 
        .ZN(n13154) );
  NAND2_X1 U16273 ( .A1(n13155), .A2(n13154), .ZN(n13156) );
  AOI211_X1 U16274 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15503), .A(n13157), 
        .B(n13156), .ZN(n13158) );
  OAI21_X1 U16275 ( .B1(n13928), .B2(n15480), .A(n13158), .ZN(P1_U2830) );
  AOI22_X1 U16276 ( .A1(n15613), .A2(n19725), .B1(n13694), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n13159) );
  OAI21_X1 U16277 ( .B1(n13928), .B2(n13696), .A(n13159), .ZN(P1_U2862) );
  INV_X1 U16278 ( .A(n13717), .ZN(n13160) );
  INV_X1 U16279 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20639) );
  OAI222_X1 U16280 ( .A1(n13928), .A2(n13777), .B1(n13766), .B2(n13160), .C1(
        n13764), .C2(n20639), .ZN(P1_U2894) );
  INV_X1 U16281 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13930) );
  MUX2_X1 U16282 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n13930), .S(n9615), .Z(n13165) );
  OR2_X1 U16283 ( .A1(n13163), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13161) );
  NAND2_X1 U16284 ( .A1(n13163), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13164) );
  XOR2_X1 U16285 ( .A(n13165), .B(n13186), .Z(n13178) );
  NAND2_X1 U16286 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13931) );
  NAND2_X1 U16287 ( .A1(n13170), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13166) );
  AND2_X1 U16288 ( .A1(n13166), .A2(n14058), .ZN(n15597) );
  INV_X1 U16289 ( .A(n15606), .ZN(n15650) );
  NOR2_X1 U16290 ( .A1(n19820), .A2(n19828), .ZN(n19815) );
  OAI21_X1 U16291 ( .B1(n14119), .B2(n14120), .A(n19841), .ZN(n19811) );
  NAND3_X1 U16292 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19815), .A3(
        n19811), .ZN(n15605) );
  NAND3_X1 U16293 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13167) );
  NOR2_X1 U16294 ( .A1(n15605), .A2(n13167), .ZN(n15611) );
  AND2_X1 U16295 ( .A1(n15650), .A2(n15611), .ZN(n13169) );
  OAI22_X1 U16296 ( .A1(n19635), .A2(n19834), .B1(n20435), .B2(n15601), .ZN(
        n13168) );
  AOI21_X1 U16297 ( .B1(n13169), .B2(n13930), .A(n13168), .ZN(n13174) );
  NAND2_X1 U16298 ( .A1(n13170), .A2(n14119), .ZN(n13171) );
  NAND2_X1 U16299 ( .A1(n13172), .A2(n13171), .ZN(n14103) );
  AOI21_X1 U16300 ( .B1(n14073), .B2(n13931), .A(n14103), .ZN(n19839) );
  INV_X1 U16301 ( .A(n19839), .ZN(n19813) );
  AOI21_X1 U16302 ( .B1(n19831), .B2(n15605), .A(n19813), .ZN(n15625) );
  OAI21_X1 U16303 ( .B1(n15629), .B2(n15611), .A(n15625), .ZN(n15615) );
  NAND2_X1 U16304 ( .A1(n15615), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13173) );
  OAI211_X1 U16305 ( .C1(n13178), .C2(n19838), .A(n13174), .B(n13173), .ZN(
        P1_U3022) );
  OAI22_X1 U16306 ( .A1(n13917), .A2(n19636), .B1(n15601), .B2(n20435), .ZN(
        n13176) );
  NOR2_X1 U16307 ( .A1(n19639), .A2(n19851), .ZN(n13175) );
  AOI211_X1 U16308 ( .C1(n15536), .C2(n19640), .A(n13176), .B(n13175), .ZN(
        n13177) );
  OAI21_X1 U16309 ( .B1(n13178), .B2(n19804), .A(n13177), .ZN(P1_U2990) );
  NAND2_X1 U16310 ( .A1(n13180), .A2(n13179), .ZN(n13181) );
  AND2_X1 U16311 ( .A1(n13633), .A2(n13181), .ZN(n13636) );
  XNOR2_X1 U16312 ( .A(n13636), .B(n13632), .ZN(n15539) );
  INV_X1 U16313 ( .A(n15539), .ZN(n13185) );
  OAI21_X1 U16314 ( .B1(n9850), .B2(n9715), .A(n15488), .ZN(n15499) );
  INV_X1 U16315 ( .A(n15499), .ZN(n13182) );
  AOI22_X1 U16316 ( .A1(n13182), .A2(n19725), .B1(n13694), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n13183) );
  OAI21_X1 U16317 ( .B1(n13185), .B2(n13696), .A(n13183), .ZN(P1_U2861) );
  MUX2_X1 U16318 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n19852), .Z(
        n19768) );
  AOI22_X1 U16319 ( .A1(n13775), .A2(n19768), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n13774), .ZN(n13184) );
  OAI21_X1 U16320 ( .B1(n13185), .B2(n13777), .A(n13184), .ZN(P1_U2893) );
  INV_X1 U16321 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14089) );
  NAND2_X1 U16322 ( .A1(n9615), .A2(n14089), .ZN(n13187) );
  NAND2_X1 U16323 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13188) );
  AND2_X1 U16324 ( .A1(n9615), .A2(n13188), .ZN(n13912) );
  INV_X1 U16325 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13196) );
  INV_X1 U16326 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15589) );
  NAND2_X1 U16327 ( .A1(n9615), .A2(n15589), .ZN(n13189) );
  OR2_X1 U16328 ( .A1(n9615), .A2(n15589), .ZN(n13190) );
  NAND2_X1 U16329 ( .A1(n13901), .A2(n13190), .ZN(n15523) );
  NOR2_X1 U16330 ( .A1(n9615), .A2(n13192), .ZN(n13191) );
  NOR2_X1 U16331 ( .A1(n15523), .A2(n13191), .ZN(n13195) );
  XNOR2_X1 U16332 ( .A(n9615), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13893) );
  NAND2_X1 U16333 ( .A1(n9615), .A2(n13192), .ZN(n13193) );
  INV_X1 U16334 ( .A(n13195), .ZN(n13891) );
  NOR2_X1 U16335 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13197) );
  NAND2_X1 U16336 ( .A1(n13913), .A2(n13911), .ZN(n13888) );
  AND2_X1 U16337 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14042) );
  NAND2_X1 U16338 ( .A1(n14042), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13936) );
  INV_X1 U16339 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15572) );
  AND2_X1 U16340 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14022) );
  NAND2_X1 U16341 ( .A1(n14022), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13999) );
  INV_X1 U16342 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13937) );
  NOR2_X1 U16343 ( .A1(n13198), .A2(n10117), .ZN(n13828) );
  INV_X1 U16344 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13199) );
  INV_X1 U16345 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14029) );
  NAND2_X1 U16346 ( .A1(n13199), .A2(n14029), .ZN(n14023) );
  NOR2_X1 U16347 ( .A1(n14023), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13799) );
  NAND2_X1 U16348 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13966) );
  NOR2_X1 U16349 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13981) );
  NAND2_X1 U16350 ( .A1(n11842), .A2(n13201), .ZN(n13206) );
  AOI22_X1 U16351 ( .A1(n13203), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n13202), .ZN(n13204) );
  INV_X1 U16352 ( .A(n13204), .ZN(n13205) );
  NAND2_X1 U16353 ( .A1(n12502), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U16354 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13207) );
  OAI211_X1 U16355 ( .C1(n19810), .C2(n13208), .A(n13950), .B(n13207), .ZN(
        n13209) );
  OAI21_X1 U16356 ( .B1(n13954), .B2(n19804), .A(n13210), .ZN(P1_U2968) );
  NAND2_X1 U16357 ( .A1(n18899), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13328) );
  OAI21_X1 U16358 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n18899), .ZN(n13211) );
  NAND2_X1 U16359 ( .A1(n18899), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n13355) );
  AND2_X1 U16360 ( .A1(n18899), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n13359) );
  INV_X1 U16361 ( .A(n13391), .ZN(n13212) );
  NAND2_X1 U16362 ( .A1(n18899), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13213) );
  INV_X1 U16363 ( .A(n13213), .ZN(n13214) );
  NAND2_X1 U16364 ( .A1(n13214), .A2(n9649), .ZN(n13215) );
  NAND2_X1 U16365 ( .A1(n13376), .A2(n13215), .ZN(n14215) );
  AOI22_X1 U16366 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19102), .B1(
        n19044), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U16367 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18869), .B1(
        n18922), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13230) );
  INV_X1 U16368 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13219) );
  OAI22_X1 U16369 ( .A1(n13219), .A2(n19404), .B1(n13217), .B2(n13218), .ZN(
        n13223) );
  INV_X1 U16370 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13221) );
  OAI22_X1 U16371 ( .A1(n13221), .A2(n19223), .B1(n12753), .B2(n13220), .ZN(
        n13222) );
  NOR2_X1 U16372 ( .A1(n13223), .A2(n13222), .ZN(n13229) );
  OAI22_X1 U16373 ( .A1(n13226), .A2(n13224), .B1(n19267), .B2(n13225), .ZN(
        n13227) );
  INV_X1 U16374 ( .A(n13227), .ZN(n13228) );
  AOI22_X1 U16375 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18950), .B1(
        n18983), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13237) );
  AOI22_X1 U16376 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19070), .B1(
        n19010), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U16377 ( .A1(n13232), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U16378 ( .A1(n13233), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n13234) );
  NAND2_X1 U16379 ( .A1(n13238), .A2(n13275), .ZN(n13239) );
  XNOR2_X1 U16380 ( .A(n13248), .B(n13240), .ZN(n18664) );
  NAND2_X1 U16381 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13243) );
  NAND2_X1 U16382 ( .A1(n13244), .A2(n13243), .ZN(n14889) );
  OR2_X1 U16383 ( .A1(n13246), .A2(n13245), .ZN(n13247) );
  NAND2_X1 U16384 ( .A1(n13248), .A2(n13247), .ZN(n13445) );
  XNOR2_X1 U16385 ( .A(n13445), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14888) );
  NAND2_X1 U16386 ( .A1(n14889), .A2(n14888), .ZN(n13249) );
  NAND2_X1 U16387 ( .A1(n13249), .A2(n10156), .ZN(n14871) );
  NAND2_X1 U16388 ( .A1(n13250), .A2(n14871), .ZN(n13253) );
  NAND2_X1 U16389 ( .A1(n13251), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13252) );
  AOI22_X1 U16390 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19102), .B1(
        n19010), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U16391 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18983), .B1(
        n19070), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13267) );
  INV_X1 U16392 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13257) );
  INV_X1 U16393 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13256) );
  OAI22_X1 U16394 ( .A1(n13257), .A2(n19404), .B1(n19223), .B2(n13256), .ZN(
        n13261) );
  OAI22_X1 U16395 ( .A1(n13259), .A2(n13217), .B1(n12753), .B2(n13258), .ZN(
        n13260) );
  NOR2_X1 U16396 ( .A1(n13261), .A2(n13260), .ZN(n13266) );
  OAI22_X1 U16397 ( .A1(n13263), .A2(n13224), .B1(n19267), .B2(n13262), .ZN(
        n13264) );
  INV_X1 U16398 ( .A(n13264), .ZN(n13265) );
  NAND4_X1 U16399 ( .A1(n13268), .A2(n13267), .A3(n13266), .A4(n13265), .ZN(
        n13274) );
  AOI22_X1 U16400 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18950), .B1(
        n18922), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U16401 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18869), .B1(
        n19044), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U16402 ( .A1(n13232), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13270) );
  NAND2_X1 U16403 ( .A1(n13233), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13269) );
  NAND4_X1 U16404 ( .A1(n13272), .A2(n13271), .A3(n13270), .A4(n13269), .ZN(
        n13273) );
  NAND2_X1 U16405 ( .A1(n13276), .A2(n13275), .ZN(n13277) );
  NAND2_X1 U16406 ( .A1(n13411), .A2(n13420), .ZN(n13281) );
  XNOR2_X1 U16407 ( .A(n13280), .B(n13279), .ZN(n18647) );
  NAND2_X1 U16408 ( .A1(n13281), .A2(n18647), .ZN(n13282) );
  XNOR2_X1 U16409 ( .A(n13282), .B(n15899), .ZN(n14601) );
  NAND2_X1 U16410 ( .A1(n13282), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13283) );
  NAND2_X1 U16411 ( .A1(n13284), .A2(n13283), .ZN(n14590) );
  INV_X1 U16412 ( .A(n13285), .ZN(n13286) );
  XNOR2_X1 U16413 ( .A(n13287), .B(n13286), .ZN(n18640) );
  AND2_X1 U16414 ( .A1(n18640), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14591) );
  INV_X1 U16415 ( .A(n14591), .ZN(n13288) );
  NOR2_X1 U16416 ( .A1(n13290), .A2(n13420), .ZN(n13291) );
  AND2_X1 U16417 ( .A1(n13291), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15805) );
  INV_X1 U16418 ( .A(n13291), .ZN(n13292) );
  NAND2_X1 U16419 ( .A1(n13292), .A2(n15900), .ZN(n15803) );
  INV_X1 U16420 ( .A(n18640), .ZN(n13293) );
  NAND2_X1 U16421 ( .A1(n13293), .A2(n15911), .ZN(n15802) );
  AND2_X1 U16422 ( .A1(n18899), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13295) );
  MUX2_X1 U16423 ( .A(n10263), .B(n13295), .S(n13294), .Z(n13296) );
  NOR2_X1 U16424 ( .A1(n13296), .A2(n13300), .ZN(n18624) );
  AOI21_X1 U16425 ( .B1(n18624), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14844) );
  NOR2_X1 U16426 ( .A1(n13300), .A2(n12026), .ZN(n13297) );
  NAND2_X1 U16427 ( .A1(n18899), .A2(n13297), .ZN(n13298) );
  NAND2_X1 U16428 ( .A1(n13368), .A2(n13298), .ZN(n13299) );
  AOI21_X1 U16429 ( .B1(n13300), .B2(n12026), .A(n13299), .ZN(n18616) );
  NAND2_X1 U16430 ( .A1(n18616), .A2(n13426), .ZN(n13307) );
  NAND2_X1 U16431 ( .A1(n13307), .A2(n15787), .ZN(n15784) );
  AND3_X1 U16432 ( .A1(n18899), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n13301), .ZN(
        n13302) );
  NOR2_X1 U16433 ( .A1(n13303), .A2(n13302), .ZN(n13304) );
  AOI21_X1 U16434 ( .B1(n13304), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14827) );
  INV_X1 U16435 ( .A(n13304), .ZN(n18603) );
  NAND2_X1 U16436 ( .A1(n13386), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13305) );
  AND2_X1 U16437 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13306) );
  NAND2_X1 U16438 ( .A1(n18624), .A2(n13306), .ZN(n14843) );
  OR2_X1 U16439 ( .A1(n15787), .A2(n13307), .ZN(n15783) );
  AND2_X1 U16440 ( .A1(n14843), .A2(n15783), .ZN(n14823) );
  NAND2_X1 U16441 ( .A1(n14825), .A2(n14823), .ZN(n14504) );
  NAND2_X1 U16442 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13308) );
  OR2_X1 U16443 ( .A1(n13309), .A2(n13308), .ZN(n15767) );
  OR2_X1 U16444 ( .A1(n13309), .A2(n13420), .ZN(n13310) );
  INV_X1 U16445 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15770) );
  NAND2_X1 U16446 ( .A1(n13312), .A2(n13311), .ZN(n13313) );
  AND2_X1 U16447 ( .A1(n13314), .A2(n13313), .ZN(n18590) );
  NAND2_X1 U16448 ( .A1(n18590), .A2(n13426), .ZN(n13351) );
  INV_X1 U16449 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U16450 ( .A1(n13351), .A2(n13315), .ZN(n14574) );
  NAND2_X1 U16451 ( .A1(n18899), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n13316) );
  NOR2_X1 U16452 ( .A1(n13322), .A2(n13316), .ZN(n13317) );
  NOR2_X1 U16453 ( .A1(n13318), .A2(n13317), .ZN(n18524) );
  AOI21_X1 U16454 ( .B1(n18524), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14516) );
  NAND2_X1 U16455 ( .A1(n13326), .A2(n14332), .ZN(n13321) );
  NAND3_X1 U16456 ( .A1(n13321), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n18899), 
        .ZN(n13319) );
  NAND2_X1 U16457 ( .A1(n13319), .A2(n13323), .ZN(n18536) );
  NOR2_X1 U16458 ( .A1(n18536), .A2(n13420), .ZN(n13345) );
  NOR2_X1 U16459 ( .A1(n13345), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14538) );
  NAND2_X1 U16460 ( .A1(n18899), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13320) );
  NOR2_X1 U16461 ( .A1(n14538), .A2(n14539), .ZN(n14525) );
  NAND2_X1 U16462 ( .A1(n18899), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13324) );
  MUX2_X1 U16463 ( .A(n18899), .B(n13324), .S(n13323), .Z(n13325) );
  NAND2_X1 U16464 ( .A1(n9972), .A2(n13325), .ZN(n14236) );
  INV_X1 U16465 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14757) );
  OAI21_X1 U16466 ( .B1(n14236), .B2(n13420), .A(n14757), .ZN(n14527) );
  NAND2_X1 U16467 ( .A1(n14525), .A2(n14527), .ZN(n14514) );
  INV_X1 U16468 ( .A(n13326), .ZN(n13332) );
  INV_X1 U16469 ( .A(n13327), .ZN(n13330) );
  INV_X1 U16470 ( .A(n13328), .ZN(n13329) );
  NAND2_X1 U16471 ( .A1(n13330), .A2(n13329), .ZN(n13331) );
  NAND2_X1 U16472 ( .A1(n13332), .A2(n13331), .ZN(n18561) );
  OR2_X1 U16473 ( .A1(n18561), .A2(n13420), .ZN(n13333) );
  NAND2_X1 U16474 ( .A1(n13333), .A2(n14553), .ZN(n14510) );
  AND2_X1 U16475 ( .A1(n18899), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13335) );
  INV_X1 U16476 ( .A(n13368), .ZN(n13334) );
  AOI21_X1 U16477 ( .B1(n13336), .B2(n13335), .A(n13334), .ZN(n13338) );
  AND2_X1 U16478 ( .A1(n13338), .A2(n13337), .ZN(n18573) );
  NAND2_X1 U16479 ( .A1(n18573), .A2(n13426), .ZN(n13339) );
  XNOR2_X1 U16480 ( .A(n13339), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14557) );
  NAND2_X1 U16481 ( .A1(n13349), .A2(n13426), .ZN(n13340) );
  NAND2_X1 U16482 ( .A1(n13340), .A2(n15870), .ZN(n14564) );
  XNOR2_X1 U16483 ( .A(n9652), .B(n9690), .ZN(n18583) );
  AOI21_X1 U16484 ( .B1(n18583), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14566) );
  INV_X1 U16485 ( .A(n14566), .ZN(n13341) );
  NAND2_X1 U16486 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13342) );
  NOR2_X1 U16487 ( .A1(n14236), .A2(n13342), .ZN(n14513) );
  INV_X1 U16488 ( .A(n18524), .ZN(n13344) );
  NAND2_X1 U16489 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13343) );
  NOR2_X1 U16490 ( .A1(n13344), .A2(n13343), .ZN(n14515) );
  NAND2_X1 U16491 ( .A1(n13345), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14512) );
  NAND2_X1 U16492 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13346) );
  OR2_X1 U16493 ( .A1(n18561), .A2(n13346), .ZN(n14509) );
  AND2_X1 U16494 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13347) );
  AND2_X1 U16495 ( .A1(n18583), .A2(n13347), .ZN(n14565) );
  AND2_X1 U16496 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13348) );
  NOR2_X1 U16497 ( .A1(n14565), .A2(n15756), .ZN(n14505) );
  AND2_X1 U16498 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13350) );
  NAND2_X1 U16499 ( .A1(n18573), .A2(n13350), .ZN(n14507) );
  INV_X1 U16500 ( .A(n13351), .ZN(n13352) );
  NAND2_X1 U16501 ( .A1(n13352), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14575) );
  AND4_X1 U16502 ( .A1(n14509), .A2(n14505), .A3(n14507), .A4(n14575), .ZN(
        n13354) );
  AND2_X1 U16503 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13353) );
  NAND2_X1 U16504 ( .A1(n18547), .A2(n13353), .ZN(n14765) );
  INV_X1 U16505 ( .A(n13355), .ZN(n13356) );
  NAND2_X1 U16506 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  AND2_X1 U16507 ( .A1(n13360), .A2(n13358), .ZN(n15348) );
  AOI21_X1 U16508 ( .B1(n15348), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14732) );
  NAND2_X1 U16509 ( .A1(n13360), .A2(n13359), .ZN(n13361) );
  NAND2_X1 U16510 ( .A1(n13363), .A2(n13361), .ZN(n15705) );
  NOR2_X1 U16511 ( .A1(n15705), .A2(n13420), .ZN(n13362) );
  XOR2_X1 U16512 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n13362), .Z(
        n14719) );
  INV_X1 U16513 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14727) );
  INV_X1 U16514 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14709) );
  NAND2_X1 U16515 ( .A1(n18899), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13364) );
  MUX2_X1 U16516 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n13364), .S(n13363), .Z(
        n13365) );
  NAND2_X1 U16517 ( .A1(n13365), .A2(n13368), .ZN(n15690) );
  NOR2_X1 U16518 ( .A1(n15690), .A2(n13420), .ZN(n14493) );
  NOR2_X1 U16519 ( .A1(n13370), .A2(n20558), .ZN(n13366) );
  NAND2_X1 U16520 ( .A1(n18899), .A2(n13366), .ZN(n13367) );
  NAND2_X1 U16521 ( .A1(n13368), .A2(n13367), .ZN(n13369) );
  AOI21_X1 U16522 ( .B1(n13370), .B2(n20558), .A(n13369), .ZN(n15687) );
  AOI21_X1 U16523 ( .B1(n15687), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14484) );
  NAND3_X1 U16524 ( .A1(n18899), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n13371), 
        .ZN(n13372) );
  NAND2_X1 U16525 ( .A1(n18899), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13374) );
  INV_X1 U16526 ( .A(n13374), .ZN(n13375) );
  NAND2_X1 U16527 ( .A1(n13376), .A2(n13375), .ZN(n13377) );
  NAND2_X1 U16528 ( .A1(n14206), .A2(n13426), .ZN(n14458) );
  INV_X1 U16529 ( .A(n15687), .ZN(n13378) );
  INV_X1 U16530 ( .A(n13379), .ZN(n13380) );
  NAND2_X1 U16531 ( .A1(n14475), .A2(n13381), .ZN(n14452) );
  NAND2_X1 U16532 ( .A1(n18899), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13383) );
  XOR2_X1 U16533 ( .A(n13383), .B(n13382), .Z(n13388) );
  OAI21_X1 U16534 ( .B1(n13388), .B2(n13420), .A(n14652), .ZN(n14441) );
  INV_X1 U16535 ( .A(n13382), .ZN(n13384) );
  NAND2_X1 U16536 ( .A1(n13384), .A2(n13383), .ZN(n13389) );
  NAND2_X1 U16537 ( .A1(n18899), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13385) );
  XNOR2_X1 U16538 ( .A(n13389), .B(n13385), .ZN(n14179) );
  AOI21_X1 U16539 ( .B1(n14179), .B2(n13386), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14433) );
  INV_X1 U16540 ( .A(n14179), .ZN(n13387) );
  INV_X1 U16541 ( .A(n13388), .ZN(n14186) );
  NAND3_X1 U16542 ( .A1(n14186), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13426), .ZN(n14440) );
  NOR2_X1 U16543 ( .A1(n13389), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13390) );
  MUX2_X1 U16544 ( .A(n13391), .B(n13390), .S(n18899), .Z(n14169) );
  NAND2_X1 U16545 ( .A1(n14169), .A2(n13426), .ZN(n13392) );
  XNOR2_X1 U16546 ( .A(n13392), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13393) );
  XNOR2_X1 U16547 ( .A(n13394), .B(n13393), .ZN(n14631) );
  AOI22_X1 U16548 ( .A1(n12025), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13397) );
  NAND2_X1 U16549 ( .A1(n13395), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13396) );
  OAI211_X1 U16550 ( .C1(n13398), .C2(n14622), .A(n13397), .B(n13396), .ZN(
        n13399) );
  XNOR2_X1 U16551 ( .A(n13400), .B(n13399), .ZN(n14627) );
  NAND2_X1 U16552 ( .A1(n18815), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14624) );
  NAND2_X1 U16553 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13401) );
  OAI211_X1 U16554 ( .C1(n13402), .C2(n18817), .A(n14624), .B(n13401), .ZN(
        n13431) );
  NAND2_X1 U16555 ( .A1(n13403), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13404) );
  NAND2_X1 U16556 ( .A1(n13406), .A2(n10134), .ZN(n13407) );
  NAND2_X1 U16557 ( .A1(n13408), .A2(n13407), .ZN(n14895) );
  NAND2_X1 U16558 ( .A1(n13410), .A2(n9934), .ZN(n14874) );
  NAND2_X1 U16559 ( .A1(n13415), .A2(n13411), .ZN(n13416) );
  NAND2_X1 U16560 ( .A1(n14586), .A2(n15911), .ZN(n13421) );
  INV_X1 U16561 ( .A(n14586), .ZN(n13422) );
  NAND2_X1 U16562 ( .A1(n13422), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13423) );
  INV_X1 U16563 ( .A(n13424), .ZN(n13427) );
  NAND2_X1 U16564 ( .A1(n13427), .A2(n13426), .ZN(n13425) );
  XNOR2_X1 U16565 ( .A(n13425), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15799) );
  NAND3_X1 U16566 ( .A1(n13427), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n13426), .ZN(n13428) );
  NAND2_X2 U16567 ( .A1(n13429), .A2(n13428), .ZN(n14551) );
  NAND3_X1 U16568 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14808) );
  INV_X1 U16569 ( .A(n14808), .ZN(n14783) );
  NAND2_X1 U16570 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15859) );
  NOR2_X1 U16571 ( .A1(n15870), .A2(n15859), .ZN(n15858) );
  NAND2_X1 U16572 ( .A1(n14783), .A2(n15858), .ZN(n14786) );
  INV_X1 U16573 ( .A(n14786), .ZN(n13430) );
  AND4_X1 U16574 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n13430), .ZN(n14617) );
  INV_X1 U16575 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15838) );
  OR2_X2 U16576 ( .A1(n14533), .A2(n14618), .ZN(n14519) );
  INV_X1 U16577 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U16578 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14620) );
  NAND2_X1 U16579 ( .A1(n14340), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13437) );
  OR2_X1 U16580 ( .A1(n13433), .A2(n13432), .ZN(n13435) );
  AND2_X1 U16581 ( .A1(n13435), .A2(n13434), .ZN(n18801) );
  NAND2_X1 U16582 ( .A1(n18801), .A2(n14350), .ZN(n13436) );
  OAI211_X1 U16583 ( .C1(n18734), .C2(n14342), .A(n13437), .B(n13436), .ZN(
        P2_U2883) );
  INV_X1 U16584 ( .A(n18805), .ZN(n13441) );
  NOR2_X1 U16585 ( .A1(n18653), .A2(n13438), .ZN(n13440) );
  AOI21_X1 U16586 ( .B1(n13441), .B2(n13440), .A(n19465), .ZN(n13439) );
  OAI21_X1 U16587 ( .B1(n13441), .B2(n13440), .A(n13439), .ZN(n13448) );
  INV_X1 U16588 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19491) );
  AOI22_X1 U16589 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18677), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n18563), .ZN(n13442) );
  OAI211_X1 U16590 ( .C1(n18681), .C2(n19491), .A(n13442), .B(n15908), .ZN(
        n13443) );
  AOI21_X1 U16591 ( .B1(n18684), .B2(n14893), .A(n13443), .ZN(n13444) );
  OAI21_X1 U16592 ( .B1(n13445), .B2(n18687), .A(n13444), .ZN(n13446) );
  AOI21_X1 U16593 ( .B1(n18801), .B2(n18689), .A(n13446), .ZN(n13447) );
  OAI211_X1 U16594 ( .C1(n18734), .C2(n13449), .A(n13448), .B(n13447), .ZN(
        P2_U2851) );
  INV_X1 U16595 ( .A(n13456), .ZN(n13461) );
  NAND2_X1 U16596 ( .A1(n13450), .A2(n13461), .ZN(n13460) );
  INV_X1 U16597 ( .A(n13451), .ZN(n13452) );
  AOI22_X1 U16598 ( .A1(n13453), .A2(n13452), .B1(n13456), .B2(n13463), .ZN(
        n13459) );
  NAND2_X1 U16599 ( .A1(n13455), .A2(n13454), .ZN(n13457) );
  NAND2_X1 U16600 ( .A1(n13457), .A2(n13456), .ZN(n13458) );
  AND3_X1 U16601 ( .A1(n13460), .A2(n13459), .A3(n13458), .ZN(n15374) );
  INV_X1 U16602 ( .A(n15374), .ZN(n13467) );
  OAI22_X1 U16603 ( .A1(n13464), .A2(n13463), .B1(n13462), .B2(n13461), .ZN(
        n19611) );
  NAND3_X1 U16604 ( .A1(n13465), .A2(n13471), .A3(n15401), .ZN(n20490) );
  AND2_X1 U16605 ( .A1(n20490), .A2(n20415), .ZN(n13466) );
  NOR2_X1 U16606 ( .A1(n19611), .A2(n13466), .ZN(n15371) );
  NOR2_X1 U16607 ( .A1(n15371), .A2(n19610), .ZN(n19618) );
  MUX2_X1 U16608 ( .A(P1_MORE_REG_SCAN_IN), .B(n13467), .S(n19618), .Z(
        P1_U3484) );
  MUX2_X1 U16609 ( .A(n13470), .B(n13469), .S(n13468), .Z(n13474) );
  AOI22_X1 U16610 ( .A1(n13472), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13471), .ZN(n13473) );
  NAND2_X1 U16611 ( .A1(n13700), .A2(n19667), .ZN(n13489) );
  AND2_X1 U16612 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n13481) );
  INV_X1 U16613 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n13537) );
  INV_X1 U16614 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n13476) );
  INV_X1 U16615 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n13649) );
  NAND4_X1 U16616 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_10__SCAN_IN), .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n13644)
         );
  NOR4_X1 U16617 ( .A1(n13476), .A2(n13649), .A3(n13475), .A4(n13644), .ZN(
        n13596) );
  INV_X1 U16618 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n13477) );
  NAND3_X1 U16619 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n13595) );
  NOR2_X1 U16620 ( .A1(n13477), .A2(n13595), .ZN(n15454) );
  NAND3_X1 U16621 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n13596), .A3(n15454), 
        .ZN(n13576) );
  NAND4_X1 U16622 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .A4(P1_REIP_REG_20__SCAN_IN), .ZN(n13483) );
  NOR3_X1 U16623 ( .A1(n19705), .A2(n13576), .A3(n13483), .ZN(n13566) );
  NAND2_X1 U16624 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n13566), .ZN(n13548) );
  NOR2_X1 U16625 ( .A1(n13537), .A2(n13548), .ZN(n13478) );
  AND2_X1 U16626 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n13478), .ZN(n13479) );
  OR2_X1 U16627 ( .A1(n13640), .A2(n13479), .ZN(n13538) );
  NAND2_X1 U16628 ( .A1(n13538), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n13526) );
  INV_X1 U16629 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n13795) );
  OR2_X1 U16630 ( .A1(n13526), .A2(n13795), .ZN(n13480) );
  INV_X1 U16631 ( .A(n13640), .ZN(n13578) );
  NAND2_X1 U16632 ( .A1(n13480), .A2(n13578), .ZN(n13513) );
  OAI21_X1 U16633 ( .B1(n13640), .B2(n13481), .A(n13513), .ZN(n13490) );
  INV_X1 U16634 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n13652) );
  OAI22_X1 U16635 ( .A1(n19695), .A2(n13652), .B1(n13482), .B2(n19686), .ZN(
        n13487) );
  NOR2_X1 U16636 ( .A1(n19678), .A2(n13576), .ZN(n13584) );
  INV_X1 U16637 ( .A(n13584), .ZN(n13484) );
  NOR2_X1 U16638 ( .A1(n13484), .A2(n13483), .ZN(n13564) );
  NAND3_X1 U16639 ( .A1(n13564), .A2(P1_REIP_REG_24__SCAN_IN), .A3(
        P1_REIP_REG_25__SCAN_IN), .ZN(n13534) );
  NOR2_X1 U16640 ( .A1(n13534), .A2(n13537), .ZN(n13527) );
  NAND3_X1 U16641 ( .A1(n13527), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n13501) );
  INV_X1 U16642 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20463) );
  INV_X1 U16643 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13485) );
  NOR4_X1 U16644 ( .A1(n13501), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n20463), 
        .A4(n13485), .ZN(n13486) );
  AOI211_X1 U16645 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n13490), .A(n13487), 
        .B(n13486), .ZN(n13488) );
  OAI211_X1 U16646 ( .C1(n13929), .C2(n19673), .A(n13489), .B(n13488), .ZN(
        P1_U2809) );
  NOR2_X1 U16647 ( .A1(n13501), .A2(n20463), .ZN(n13491) );
  OAI21_X1 U16648 ( .B1(n13491), .B2(P1_REIP_REG_30__SCAN_IN), .A(n13490), 
        .ZN(n13493) );
  AOI22_X1 U16649 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19710), .B1(
        n19641), .B2(n13780), .ZN(n13492) );
  OAI211_X1 U16650 ( .C1(n19695), .C2(n13494), .A(n13493), .B(n13492), .ZN(
        n13495) );
  AOI21_X1 U16651 ( .B1(n13962), .B2(n19707), .A(n13495), .ZN(n13496) );
  OAI21_X1 U16652 ( .B1(n13707), .B2(n15480), .A(n13496), .ZN(P1_U2810) );
  XNOR2_X1 U16653 ( .A(n13512), .B(n13497), .ZN(n13965) );
  AOI21_X1 U16654 ( .B1(n13498), .B2(n13508), .A(n11842), .ZN(n13793) );
  NAND2_X1 U16655 ( .A1(n13793), .A2(n19667), .ZN(n13506) );
  INV_X1 U16656 ( .A(n13513), .ZN(n13504) );
  INV_X1 U16657 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n13653) );
  INV_X1 U16658 ( .A(n13791), .ZN(n13499) );
  AOI22_X1 U16659 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19710), .B1(
        n19641), .B2(n13499), .ZN(n13500) );
  OAI21_X1 U16660 ( .B1(n19695), .B2(n13653), .A(n13500), .ZN(n13503) );
  NOR2_X1 U16661 ( .A1(n13501), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n13502) );
  AOI211_X1 U16662 ( .C1(n13504), .C2(P1_REIP_REG_29__SCAN_IN), .A(n13503), 
        .B(n13502), .ZN(n13505) );
  OAI211_X1 U16663 ( .C1(n13965), .C2(n19673), .A(n13506), .B(n13505), .ZN(
        P1_U2811) );
  OAI21_X1 U16664 ( .B1(n13507), .B2(n13509), .A(n13508), .ZN(n13807) );
  NOR2_X1 U16665 ( .A1(n13521), .A2(n13510), .ZN(n13511) );
  OR2_X1 U16666 ( .A1(n13512), .A2(n13511), .ZN(n13985) );
  INV_X1 U16667 ( .A(n13985), .ZN(n13517) );
  AOI21_X1 U16668 ( .B1(n13795), .B2(n13526), .A(n13513), .ZN(n13516) );
  INV_X1 U16669 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n20638) );
  AOI22_X1 U16670 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19710), .B1(
        n19641), .B2(n13798), .ZN(n13514) );
  OAI21_X1 U16671 ( .B1(n19695), .B2(n20638), .A(n13514), .ZN(n13515) );
  AOI211_X1 U16672 ( .C1(n13517), .C2(n19707), .A(n13516), .B(n13515), .ZN(
        n13518) );
  OAI21_X1 U16673 ( .B1(n13807), .B2(n15480), .A(n13518), .ZN(P1_U2812) );
  AOI21_X1 U16674 ( .B1(n13519), .B2(n13530), .A(n13507), .ZN(n13814) );
  INV_X1 U16675 ( .A(n13814), .ZN(n13716) );
  OAI22_X1 U16676 ( .A1(n13520), .A2(n19686), .B1(n19713), .B2(n13812), .ZN(
        n13525) );
  INV_X1 U16677 ( .A(n13521), .ZN(n13522) );
  OAI21_X1 U16678 ( .B1(n13532), .B2(n13523), .A(n13522), .ZN(n13993) );
  NOR2_X1 U16679 ( .A1(n13993), .A2(n19673), .ZN(n13524) );
  AOI211_X1 U16680 ( .C1(n19708), .C2(P1_EBX_REG_27__SCAN_IN), .A(n13525), .B(
        n13524), .ZN(n13529) );
  OAI21_X1 U16681 ( .B1(n13527), .B2(P1_REIP_REG_27__SCAN_IN), .A(n13526), 
        .ZN(n13528) );
  OAI211_X1 U16682 ( .C1(n13716), .C2(n15480), .A(n13529), .B(n13528), .ZN(
        P1_U2813) );
  OAI21_X1 U16683 ( .B1(n13543), .B2(n13531), .A(n13530), .ZN(n13821) );
  OAI21_X1 U16684 ( .B1(n13533), .B2(n13546), .A(n9861), .ZN(n13655) );
  INV_X1 U16685 ( .A(n13655), .ZN(n14003) );
  NOR2_X1 U16686 ( .A1(n13534), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U16687 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19710), .B1(
        n19641), .B2(n13824), .ZN(n13536) );
  NAND2_X1 U16688 ( .A1(n19708), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n13535) );
  OAI211_X1 U16689 ( .C1(n13538), .C2(n13537), .A(n13536), .B(n13535), .ZN(
        n13539) );
  AOI211_X1 U16690 ( .C1(n14003), .C2(n19707), .A(n13540), .B(n13539), .ZN(
        n13541) );
  OAI21_X1 U16691 ( .B1(n13821), .B2(n15480), .A(n13541), .ZN(P1_U2814) );
  INV_X1 U16692 ( .A(n13543), .ZN(n13544) );
  OAI21_X1 U16693 ( .B1(n13545), .B2(n13542), .A(n13544), .ZN(n13833) );
  AOI21_X1 U16694 ( .B1(n13547), .B2(n13561), .A(n13546), .ZN(n13657) );
  NAND3_X1 U16695 ( .A1(n13548), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n13578), 
        .ZN(n13550) );
  AOI22_X1 U16696 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19710), .B1(
        n19641), .B2(n13836), .ZN(n13549) );
  OAI211_X1 U16697 ( .C1(n13658), .C2(n19695), .A(n13550), .B(n13549), .ZN(
        n13551) );
  AOI21_X1 U16698 ( .B1(n13657), .B2(n19707), .A(n13551), .ZN(n13554) );
  INV_X1 U16699 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n13552) );
  NAND3_X1 U16700 ( .A1(n13564), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n13552), 
        .ZN(n13553) );
  OAI211_X1 U16701 ( .C1(n13833), .C2(n15480), .A(n13554), .B(n13553), .ZN(
        P1_U2815) );
  INV_X1 U16702 ( .A(n13542), .ZN(n13556) );
  OAI21_X1 U16703 ( .B1(n13557), .B2(n13555), .A(n13556), .ZN(n13842) );
  INV_X1 U16704 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n13565) );
  INV_X1 U16705 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U16706 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19710), .B1(
        n19641), .B2(n13845), .ZN(n13558) );
  OAI21_X1 U16707 ( .B1(n19695), .B2(n13659), .A(n13558), .ZN(n13563) );
  NAND2_X1 U16708 ( .A1(n13663), .A2(n13559), .ZN(n13560) );
  NAND2_X1 U16709 ( .A1(n13561), .A2(n13560), .ZN(n14017) );
  NOR2_X1 U16710 ( .A1(n14017), .A2(n19673), .ZN(n13562) );
  AOI211_X1 U16711 ( .C1(n13565), .C2(n13564), .A(n13563), .B(n13562), .ZN(
        n13568) );
  NOR2_X1 U16712 ( .A1(n13640), .A2(n13566), .ZN(n15434) );
  NAND2_X1 U16713 ( .A1(n15434), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n13567) );
  OAI211_X1 U16714 ( .C1(n13842), .C2(n15480), .A(n13568), .B(n13567), .ZN(
        P1_U2816) );
  INV_X1 U16715 ( .A(n9666), .ZN(n13570) );
  AOI21_X1 U16716 ( .B1(n13571), .B2(n13667), .A(n13570), .ZN(n13859) );
  INV_X1 U16717 ( .A(n13859), .ZN(n13733) );
  AOI21_X1 U16718 ( .B1(n13572), .B2(n13673), .A(n13661), .ZN(n14040) );
  NAND2_X1 U16719 ( .A1(n19708), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13575) );
  INV_X1 U16720 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n13855) );
  NAND3_X1 U16721 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n13584), .A3(
        P1_REIP_REG_20__SCAN_IN), .ZN(n15432) );
  INV_X1 U16722 ( .A(n15432), .ZN(n13573) );
  AOI22_X1 U16723 ( .A1(n19710), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n13855), .B2(n13573), .ZN(n13574) );
  OAI211_X1 U16724 ( .C1(n19713), .C2(n13857), .A(n13575), .B(n13574), .ZN(
        n13580) );
  INV_X1 U16725 ( .A(n13576), .ZN(n13577) );
  NAND2_X1 U16726 ( .A1(n13577), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15442) );
  OAI21_X1 U16727 ( .B1(n19705), .B2(n15442), .A(n13578), .ZN(n15443) );
  INV_X1 U16728 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20451) );
  NAND2_X1 U16729 ( .A1(n19709), .A2(n20451), .ZN(n15441) );
  AOI21_X1 U16730 ( .B1(n15443), .B2(n15441), .A(n13855), .ZN(n13579) );
  AOI211_X1 U16731 ( .C1(n14040), .C2(n19707), .A(n13580), .B(n13579), .ZN(
        n13581) );
  OAI21_X1 U16732 ( .B1(n13733), .B2(n15480), .A(n13581), .ZN(P1_U2818) );
  OAI21_X1 U16733 ( .B1(n13680), .B2(n13582), .A(n13668), .ZN(n13876) );
  AOI21_X1 U16734 ( .B1(n13583), .B2(n9631), .A(n9869), .ZN(n14057) );
  NOR2_X1 U16735 ( .A1(n13584), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n13587) );
  AOI22_X1 U16736 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19710), .B1(
        n19641), .B2(n13875), .ZN(n13586) );
  NAND2_X1 U16737 ( .A1(n19708), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n13585) );
  OAI211_X1 U16738 ( .C1(n15443), .C2(n13587), .A(n13586), .B(n13585), .ZN(
        n13588) );
  AOI21_X1 U16739 ( .B1(n14057), .B2(n19707), .A(n13588), .ZN(n13589) );
  OAI21_X1 U16740 ( .B1(n13876), .B2(n15480), .A(n13589), .ZN(P1_U2820) );
  AOI21_X1 U16741 ( .B1(n13590), .B2(n13606), .A(n13678), .ZN(n13886) );
  INV_X1 U16742 ( .A(n13886), .ZN(n13749) );
  NAND2_X1 U16743 ( .A1(n19709), .A2(n13596), .ZN(n15452) );
  NOR3_X1 U16744 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n13595), .A3(n15452), 
        .ZN(n15462) );
  INV_X1 U16745 ( .A(n13591), .ZN(n13610) );
  INV_X1 U16746 ( .A(n13592), .ZN(n13593) );
  AOI21_X1 U16747 ( .B1(n13621), .B2(n13610), .A(n13593), .ZN(n13594) );
  OR2_X1 U16748 ( .A1(n13682), .A2(n13594), .ZN(n15567) );
  NOR2_X1 U16749 ( .A1(n15567), .A2(n19673), .ZN(n13603) );
  INV_X1 U16750 ( .A(n13595), .ZN(n13598) );
  OR2_X1 U16751 ( .A1(n19678), .A2(n13596), .ZN(n13597) );
  NAND2_X1 U16752 ( .A1(n13597), .A2(n19646), .ZN(n13623) );
  INV_X1 U16753 ( .A(n13623), .ZN(n15486) );
  OAI21_X1 U16754 ( .B1(n19678), .B2(n13598), .A(n15486), .ZN(n15461) );
  AOI22_X1 U16755 ( .A1(n19708), .A2(P1_EBX_REG_18__SCAN_IN), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n15461), .ZN(n13599) );
  OAI211_X1 U16756 ( .C1(n19686), .C2(n13600), .A(n13599), .B(n19693), .ZN(
        n13602) );
  NOR2_X1 U16757 ( .A1(n13884), .A2(n19713), .ZN(n13601) );
  NOR4_X1 U16758 ( .A1(n15462), .A2(n13603), .A3(n13602), .A4(n13601), .ZN(
        n13604) );
  OAI21_X1 U16759 ( .B1(n13749), .B2(n15480), .A(n13604), .ZN(P1_U2822) );
  INV_X1 U16760 ( .A(n13606), .ZN(n13607) );
  AOI21_X1 U16761 ( .B1(n13608), .B2(n13605), .A(n13607), .ZN(n15520) );
  INV_X1 U16762 ( .A(n15520), .ZN(n13755) );
  NAND2_X1 U16763 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n13609) );
  INV_X1 U16764 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20445) );
  OAI21_X1 U16765 ( .B1(n13609), .B2(n15452), .A(n20445), .ZN(n13616) );
  XNOR2_X1 U16766 ( .A(n13621), .B(n13610), .ZN(n15576) );
  NAND2_X1 U16767 ( .A1(n19710), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13611) );
  OAI211_X1 U16768 ( .C1(n19695), .C2(n13612), .A(n13611), .B(n19693), .ZN(
        n13613) );
  AOI21_X1 U16769 ( .B1(n19641), .B2(n15519), .A(n13613), .ZN(n13614) );
  OAI21_X1 U16770 ( .B1(n15576), .B2(n19673), .A(n13614), .ZN(n13615) );
  AOI21_X1 U16771 ( .B1(n13616), .B2(n15461), .A(n13615), .ZN(n13617) );
  OAI21_X1 U16772 ( .B1(n13755), .B2(n15480), .A(n13617), .ZN(P1_U2823) );
  OAI21_X1 U16773 ( .B1(n13618), .B2(n13619), .A(n13605), .ZN(n13896) );
  INV_X1 U16774 ( .A(n15472), .ZN(n13691) );
  AOI21_X1 U16775 ( .B1(n13691), .B2(n15471), .A(n13620), .ZN(n13622) );
  OR2_X1 U16776 ( .A1(n13622), .A2(n13621), .ZN(n14081) );
  INV_X1 U16777 ( .A(n14081), .ZN(n13630) );
  INV_X1 U16778 ( .A(n13899), .ZN(n13627) );
  NOR2_X1 U16779 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15452), .ZN(n15470) );
  OAI21_X1 U16780 ( .B1(n15470), .B2(n13623), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n13624) );
  OAI211_X1 U16781 ( .C1(n19686), .C2(n13895), .A(n13624), .B(n19693), .ZN(
        n13625) );
  AOI21_X1 U16782 ( .B1(n19708), .B2(P1_EBX_REG_16__SCAN_IN), .A(n13625), .ZN(
        n13626) );
  OAI21_X1 U16783 ( .B1(n13627), .B2(n19713), .A(n13626), .ZN(n13629) );
  INV_X1 U16784 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20443) );
  NOR3_X1 U16785 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20443), .A3(n15452), 
        .ZN(n13628) );
  AOI211_X1 U16786 ( .C1(n13630), .C2(n19707), .A(n13629), .B(n13628), .ZN(
        n13631) );
  OAI21_X1 U16787 ( .B1(n13896), .B2(n15480), .A(n13631), .ZN(P1_U2824) );
  INV_X1 U16788 ( .A(n13632), .ZN(n13635) );
  INV_X1 U16789 ( .A(n13633), .ZN(n13634) );
  AOI21_X1 U16790 ( .B1(n13636), .B2(n13635), .A(n13634), .ZN(n13773) );
  INV_X1 U16791 ( .A(n13637), .ZN(n13772) );
  NOR2_X1 U16792 ( .A1(n13773), .A2(n13772), .ZN(n13771) );
  OAI21_X1 U16793 ( .B1(n13771), .B2(n13639), .A(n13638), .ZN(n13918) );
  INV_X1 U16794 ( .A(n13644), .ZN(n13642) );
  AOI21_X1 U16795 ( .B1(n13642), .B2(n13641), .A(n13640), .ZN(n15492) );
  INV_X1 U16796 ( .A(n19634), .ZN(n13643) );
  NOR2_X1 U16797 ( .A1(n13644), .A2(n13643), .ZN(n15475) );
  OR2_X1 U16798 ( .A1(n15490), .A2(n13645), .ZN(n13646) );
  NAND2_X1 U16799 ( .A1(n13692), .A2(n13646), .ZN(n14087) );
  AOI22_X1 U16800 ( .A1(n19708), .A2(P1_EBX_REG_13__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19710), .ZN(n13647) );
  OAI211_X1 U16801 ( .C1(n14087), .C2(n19673), .A(n13647), .B(n19693), .ZN(
        n13648) );
  AOI221_X1 U16802 ( .B1(n15492), .B2(P1_REIP_REG_13__SCAN_IN), .C1(n15475), 
        .C2(n13649), .A(n13648), .ZN(n13651) );
  NAND2_X1 U16803 ( .A1(n19641), .A2(n13921), .ZN(n13650) );
  OAI211_X1 U16804 ( .C1(n13918), .C2(n15480), .A(n13651), .B(n13650), .ZN(
        P1_U2827) );
  OAI22_X1 U16805 ( .A1(n13929), .A2(n13698), .B1(n13652), .B2(n19728), .ZN(
        P1_U2841) );
  INV_X1 U16806 ( .A(n13793), .ZN(n13711) );
  OAI222_X1 U16807 ( .A1(n13653), .A2(n19728), .B1(n13698), .B2(n13965), .C1(
        n13696), .C2(n13711), .ZN(P1_U2843) );
  OAI222_X1 U16808 ( .A1(n20638), .A2(n19728), .B1(n13698), .B2(n13985), .C1(
        n13807), .C2(n13696), .ZN(P1_U2844) );
  INV_X1 U16809 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n13654) );
  OAI222_X1 U16810 ( .A1(n13654), .A2(n19728), .B1(n13698), .B2(n13993), .C1(
        n13716), .C2(n13696), .ZN(P1_U2845) );
  INV_X1 U16811 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n13656) );
  OAI222_X1 U16812 ( .A1(n13696), .A2(n13821), .B1(n19728), .B2(n13656), .C1(
        n13655), .C2(n13698), .ZN(P1_U2846) );
  INV_X1 U16813 ( .A(n13657), .ZN(n14012) );
  OAI222_X1 U16814 ( .A1(n13658), .A2(n19728), .B1(n13698), .B2(n14012), .C1(
        n13833), .C2(n13696), .ZN(P1_U2847) );
  OAI222_X1 U16815 ( .A1(n13696), .A2(n13842), .B1(n19728), .B2(n13659), .C1(
        n14017), .C2(n13698), .ZN(P1_U2848) );
  INV_X1 U16816 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15426) );
  OR2_X1 U16817 ( .A1(n13661), .A2(n13660), .ZN(n13662) );
  NAND2_X1 U16818 ( .A1(n13663), .A2(n13662), .ZN(n15438) );
  AND2_X1 U16819 ( .A1(n9666), .A2(n13664), .ZN(n13665) );
  INV_X1 U16820 ( .A(n15435), .ZN(n13728) );
  OAI222_X1 U16821 ( .A1(n15426), .A2(n19728), .B1(n13698), .B2(n15438), .C1(
        n13728), .C2(n13696), .ZN(P1_U2849) );
  AOI22_X1 U16822 ( .A1(n14040), .A2(n19725), .B1(n13694), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n13666) );
  OAI21_X1 U16823 ( .B1(n13733), .B2(n13696), .A(n13666), .ZN(P1_U2850) );
  AOI21_X1 U16824 ( .B1(n13669), .B2(n13668), .A(n13569), .ZN(n13869) );
  INV_X1 U16825 ( .A(n13869), .ZN(n15445) );
  NAND2_X1 U16826 ( .A1(n13671), .A2(n13670), .ZN(n13672) );
  NAND2_X1 U16827 ( .A1(n13673), .A2(n13672), .ZN(n15444) );
  OAI22_X1 U16828 ( .A1(n15444), .A2(n13698), .B1(n15440), .B2(n19728), .ZN(
        n13674) );
  INV_X1 U16829 ( .A(n13674), .ZN(n13675) );
  OAI21_X1 U16830 ( .B1(n15445), .B2(n13696), .A(n13675), .ZN(P1_U2851) );
  AOI22_X1 U16831 ( .A1(n14057), .A2(n19725), .B1(n13694), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n13676) );
  OAI21_X1 U16832 ( .B1(n13876), .B2(n13696), .A(n13676), .ZN(P1_U2852) );
  NOR2_X1 U16833 ( .A1(n13678), .A2(n13677), .ZN(n13679) );
  OR2_X1 U16834 ( .A1(n13680), .A2(n13679), .ZN(n15451) );
  OR2_X1 U16835 ( .A1(n13682), .A2(n13681), .ZN(n13683) );
  NAND2_X1 U16836 ( .A1(n9631), .A2(n13683), .ZN(n15465) );
  OAI22_X1 U16837 ( .A1(n15465), .A2(n13698), .B1(n15459), .B2(n19728), .ZN(
        n13684) );
  INV_X1 U16838 ( .A(n13684), .ZN(n13685) );
  OAI21_X1 U16839 ( .B1(n15451), .B2(n13696), .A(n13685), .ZN(P1_U2853) );
  INV_X1 U16840 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n13686) );
  OAI222_X1 U16841 ( .A1(n15567), .A2(n13698), .B1(n13686), .B2(n19728), .C1(
        n13749), .C2(n13696), .ZN(P1_U2854) );
  OAI222_X1 U16842 ( .A1(n13755), .A2(n13696), .B1(n13698), .B2(n15576), .C1(
        n19728), .C2(n13612), .ZN(P1_U2855) );
  INV_X1 U16843 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n13687) );
  OAI222_X1 U16844 ( .A1(n14081), .A2(n13698), .B1(n13687), .B2(n19728), .C1(
        n13896), .C2(n13696), .ZN(P1_U2856) );
  NAND2_X1 U16845 ( .A1(n13638), .A2(n13689), .ZN(n13690) );
  NAND2_X1 U16846 ( .A1(n13688), .A2(n13690), .ZN(n15481) );
  AOI21_X1 U16847 ( .B1(n13693), .B2(n13692), .A(n13691), .ZN(n15592) );
  AOI22_X1 U16848 ( .A1(n15592), .A2(n19725), .B1(n13694), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n13695) );
  OAI21_X1 U16849 ( .B1(n15481), .B2(n13696), .A(n13695), .ZN(P1_U2858) );
  INV_X1 U16850 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13697) );
  OAI222_X1 U16851 ( .A1(n14087), .A2(n13698), .B1(n19728), .B2(n13697), .C1(
        n13696), .C2(n13918), .ZN(P1_U2859) );
  NOR2_X1 U16852 ( .A1(n13702), .A2(n19849), .ZN(n13699) );
  NAND2_X1 U16853 ( .A1(n13764), .A2(n13699), .ZN(n13756) );
  INV_X1 U16854 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n18910) );
  AND2_X1 U16855 ( .A1(n13764), .A2(n19895), .ZN(n13701) );
  NAND2_X1 U16856 ( .A1(n13701), .A2(n13700), .ZN(n13704) );
  NOR3_X4 U16857 ( .A1(n13774), .A2(n13702), .A3(n19852), .ZN(n13760) );
  AOI22_X1 U16858 ( .A1(n13760), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n13774), .ZN(n13703) );
  OAI211_X1 U16859 ( .C1(n13756), .C2(n18910), .A(n13704), .B(n13703), .ZN(
        P1_U2873) );
  AOI22_X1 U16860 ( .A1(n13750), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n13774), .ZN(n13706) );
  NOR3_X2 U16861 ( .A1(n13774), .A2(n19895), .A3(n11142), .ZN(n13752) );
  MUX2_X1 U16862 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n19852), .Z(
        n19772) );
  AOI22_X1 U16863 ( .A1(n13752), .A2(n19772), .B1(n13760), .B2(DATAI_30_), 
        .ZN(n13705) );
  OAI211_X1 U16864 ( .C1(n13707), .C2(n13777), .A(n13706), .B(n13705), .ZN(
        P1_U2874) );
  INV_X1 U16865 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n18896) );
  OAI22_X1 U16866 ( .A1(n13756), .A2(n18896), .B1(n20585), .B2(n13764), .ZN(
        n13708) );
  INV_X1 U16867 ( .A(n13708), .ZN(n13710) );
  AOI22_X1 U16868 ( .A1(n13752), .A2(n13769), .B1(n13760), .B2(DATAI_29_), 
        .ZN(n13709) );
  OAI211_X1 U16869 ( .C1(n13711), .C2(n13777), .A(n13710), .B(n13709), .ZN(
        P1_U2875) );
  AOI22_X1 U16870 ( .A1(n13750), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n13774), .ZN(n13713) );
  MUX2_X1 U16871 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n19852), .Z(
        n19770) );
  AOI22_X1 U16872 ( .A1(n13752), .A2(n19770), .B1(n13760), .B2(DATAI_28_), 
        .ZN(n13712) );
  OAI211_X1 U16873 ( .C1(n13807), .C2(n13777), .A(n13713), .B(n13712), .ZN(
        P1_U2876) );
  AOI22_X1 U16874 ( .A1(n13750), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n13774), .ZN(n13715) );
  AOI22_X1 U16875 ( .A1(n13752), .A2(n19768), .B1(n13760), .B2(DATAI_27_), 
        .ZN(n13714) );
  OAI211_X1 U16876 ( .C1(n13716), .C2(n13777), .A(n13715), .B(n13714), .ZN(
        P1_U2877) );
  AOI22_X1 U16877 ( .A1(n13750), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n13774), .ZN(n13719) );
  AOI22_X1 U16878 ( .A1(n13752), .A2(n13717), .B1(n13760), .B2(DATAI_26_), 
        .ZN(n13718) );
  OAI211_X1 U16879 ( .C1(n13821), .C2(n13777), .A(n13719), .B(n13718), .ZN(
        P1_U2878) );
  AOI22_X1 U16880 ( .A1(n13750), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n13774), .ZN(n13721) );
  AOI22_X1 U16881 ( .A1(n13752), .A2(n19765), .B1(n13760), .B2(DATAI_25_), 
        .ZN(n13720) );
  OAI211_X1 U16882 ( .C1(n13833), .C2(n13777), .A(n13721), .B(n13720), .ZN(
        P1_U2879) );
  AOI22_X1 U16883 ( .A1(n13750), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n13774), .ZN(n13724) );
  INV_X1 U16884 ( .A(n13722), .ZN(n19763) );
  AOI22_X1 U16885 ( .A1(n13752), .A2(n19763), .B1(n13760), .B2(DATAI_24_), 
        .ZN(n13723) );
  OAI211_X1 U16886 ( .C1(n13842), .C2(n13777), .A(n13724), .B(n13723), .ZN(
        P1_U2880) );
  INV_X1 U16887 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16064) );
  OAI22_X1 U16888 ( .A1(n13756), .A2(n16064), .B1(n12543), .B2(n13764), .ZN(
        n13726) );
  INV_X1 U16889 ( .A(n13752), .ZN(n13757) );
  NOR2_X1 U16890 ( .A1(n13757), .A2(n19899), .ZN(n13725) );
  AOI211_X1 U16891 ( .C1(n13760), .C2(DATAI_23_), .A(n13726), .B(n13725), .ZN(
        n13727) );
  OAI21_X1 U16892 ( .B1(n13728), .B2(n13777), .A(n13727), .ZN(P1_U2881) );
  NOR2_X1 U16893 ( .A1(n13756), .A2(n16066), .ZN(n13731) );
  INV_X1 U16894 ( .A(n13760), .ZN(n13729) );
  OAI22_X1 U16895 ( .A1(n13757), .A2(n19891), .B1(n13729), .B2(n20590), .ZN(
        n13730) );
  AOI211_X1 U16896 ( .C1(n13774), .C2(P1_EAX_REG_22__SCAN_IN), .A(n13731), .B(
        n13730), .ZN(n13732) );
  OAI21_X1 U16897 ( .B1(n13733), .B2(n13777), .A(n13732), .ZN(P1_U2882) );
  AOI22_X1 U16898 ( .A1(n13750), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n13774), .ZN(n13736) );
  AOI22_X1 U16899 ( .A1(n13752), .A2(n13734), .B1(n13760), .B2(DATAI_21_), 
        .ZN(n13735) );
  OAI211_X1 U16900 ( .C1(n15445), .C2(n13777), .A(n13736), .B(n13735), .ZN(
        P1_U2883) );
  INV_X1 U16901 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n13737) );
  OAI22_X1 U16902 ( .A1(n13756), .A2(n13737), .B1(n12539), .B2(n13764), .ZN(
        n13739) );
  NOR2_X1 U16903 ( .A1(n13757), .A2(n19884), .ZN(n13738) );
  AOI211_X1 U16904 ( .C1(n13760), .C2(DATAI_20_), .A(n13739), .B(n13738), .ZN(
        n13740) );
  OAI21_X1 U16905 ( .B1(n13876), .B2(n13777), .A(n13740), .ZN(P1_U2884) );
  AOI22_X1 U16906 ( .A1(n13750), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n13774), .ZN(n13743) );
  AOI22_X1 U16907 ( .A1(n13752), .A2(n13741), .B1(n13760), .B2(DATAI_19_), 
        .ZN(n13742) );
  OAI211_X1 U16908 ( .C1(n15451), .C2(n13777), .A(n13743), .B(n13742), .ZN(
        P1_U2885) );
  INV_X1 U16909 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n13745) );
  INV_X1 U16910 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13744) );
  OAI22_X1 U16911 ( .A1(n13756), .A2(n13745), .B1(n13744), .B2(n13764), .ZN(
        n13747) );
  NOR2_X1 U16912 ( .A1(n13757), .A2(n19876), .ZN(n13746) );
  AOI211_X1 U16913 ( .C1(n13760), .C2(DATAI_18_), .A(n13747), .B(n13746), .ZN(
        n13748) );
  OAI21_X1 U16914 ( .B1(n13749), .B2(n13777), .A(n13748), .ZN(P1_U2886) );
  AOI22_X1 U16915 ( .A1(n13750), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n13774), .ZN(n13754) );
  AOI22_X1 U16916 ( .A1(n13752), .A2(n13751), .B1(n13760), .B2(DATAI_17_), 
        .ZN(n13753) );
  OAI211_X1 U16917 ( .C1(n13755), .C2(n13777), .A(n13754), .B(n13753), .ZN(
        P1_U2887) );
  OAI22_X1 U16918 ( .A1(n13756), .A2(n16076), .B1(n12548), .B2(n13764), .ZN(
        n13759) );
  NOR2_X1 U16919 ( .A1(n13757), .A2(n19863), .ZN(n13758) );
  AOI211_X1 U16920 ( .C1(n13760), .C2(DATAI_16_), .A(n13759), .B(n13758), .ZN(
        n13761) );
  OAI21_X1 U16921 ( .B1(n13896), .B2(n13777), .A(n13761), .ZN(P1_U2888) );
  AOI21_X1 U16922 ( .B1(n13762), .B2(n13688), .A(n13618), .ZN(n15528) );
  INV_X1 U16923 ( .A(n15528), .ZN(n13767) );
  OAI222_X1 U16924 ( .A1(n13767), .A2(n13777), .B1(n13766), .B2(n13765), .C1(
        n13764), .C2(n13763), .ZN(P1_U2889) );
  AOI22_X1 U16925 ( .A1(n13775), .A2(n19772), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n13774), .ZN(n13768) );
  OAI21_X1 U16926 ( .B1(n15481), .B2(n13777), .A(n13768), .ZN(P1_U2890) );
  AOI22_X1 U16927 ( .A1(n13775), .A2(n13769), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n13774), .ZN(n13770) );
  OAI21_X1 U16928 ( .B1(n13918), .B2(n13777), .A(n13770), .ZN(P1_U2891) );
  AOI21_X1 U16929 ( .B1(n13773), .B2(n13772), .A(n13771), .ZN(n15534) );
  INV_X1 U16930 ( .A(n15534), .ZN(n13778) );
  AOI22_X1 U16931 ( .A1(n13775), .A2(n19770), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n13774), .ZN(n13776) );
  OAI21_X1 U16932 ( .B1(n13778), .B2(n13777), .A(n13776), .ZN(P1_U2892) );
  NAND2_X1 U16933 ( .A1(n15536), .A2(n13780), .ZN(n13781) );
  NAND2_X1 U16934 ( .A1(n12502), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13955) );
  OAI211_X1 U16935 ( .C1(n13917), .C2(n13782), .A(n13781), .B(n13955), .ZN(
        n13783) );
  AOI21_X1 U16936 ( .B1(n13784), .B2(n19794), .A(n13783), .ZN(n13785) );
  INV_X1 U16937 ( .A(n13786), .ZN(n13787) );
  MUX2_X1 U16938 ( .A(n13788), .B(n13787), .S(n10117), .Z(n13789) );
  XNOR2_X1 U16939 ( .A(n13789), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13975) );
  NOR2_X1 U16940 ( .A1(n15601), .A2(n20463), .ZN(n13969) );
  AOI21_X1 U16941 ( .B1(n19799), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n13969), .ZN(n13790) );
  OAI21_X1 U16942 ( .B1(n19810), .B2(n13791), .A(n13790), .ZN(n13792) );
  AOI21_X1 U16943 ( .B1(n13793), .B2(n19794), .A(n13792), .ZN(n13794) );
  OAI21_X1 U16944 ( .B1(n19804), .B2(n13975), .A(n13794), .ZN(P1_U2970) );
  NOR2_X1 U16945 ( .A1(n15601), .A2(n13795), .ZN(n13982) );
  NOR2_X1 U16946 ( .A1(n13917), .A2(n13796), .ZN(n13797) );
  AOI211_X1 U16947 ( .C1(n15536), .C2(n13798), .A(n13982), .B(n13797), .ZN(
        n13806) );
  NAND2_X1 U16948 ( .A1(n9615), .A2(n13999), .ZN(n13817) );
  NAND2_X1 U16949 ( .A1(n13848), .A2(n13817), .ZN(n13803) );
  INV_X1 U16950 ( .A(n13799), .ZN(n13800) );
  OAI21_X1 U16951 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n13800), .A(
        n13803), .ZN(n13802) );
  MUX2_X1 U16952 ( .A(n13990), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9615), .Z(n13801) );
  OAI211_X1 U16953 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n13803), .A(
        n13802), .B(n13801), .ZN(n13804) );
  XNOR2_X1 U16954 ( .A(n13804), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13976) );
  NAND2_X1 U16955 ( .A1(n13976), .A2(n19795), .ZN(n13805) );
  OAI211_X1 U16956 ( .C1(n13807), .C2(n19851), .A(n13806), .B(n13805), .ZN(
        P1_U2971) );
  MUX2_X1 U16957 ( .A(n13809), .B(n13808), .S(n10117), .Z(n13810) );
  XNOR2_X1 U16958 ( .A(n13810), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13997) );
  INV_X1 U16959 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20460) );
  NOR2_X1 U16960 ( .A1(n15601), .A2(n20460), .ZN(n13989) );
  AOI21_X1 U16961 ( .B1(n19799), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n13989), .ZN(n13811) );
  OAI21_X1 U16962 ( .B1(n19810), .B2(n13812), .A(n13811), .ZN(n13813) );
  AOI21_X1 U16963 ( .B1(n13814), .B2(n19794), .A(n13813), .ZN(n13815) );
  OAI21_X1 U16964 ( .B1(n13997), .B2(n19804), .A(n13815), .ZN(P1_U2972) );
  INV_X1 U16965 ( .A(n13816), .ZN(n13818) );
  OAI211_X1 U16966 ( .C1(n10117), .C2(n13848), .A(n13818), .B(n13817), .ZN(
        n13819) );
  XOR2_X1 U16967 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n13819), .Z(
        n14009) );
  INV_X1 U16968 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13820) );
  NAND2_X1 U16969 ( .A1(n12502), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n13998) );
  OAI21_X1 U16970 ( .B1(n13917), .B2(n13820), .A(n13998), .ZN(n13823) );
  NOR2_X1 U16971 ( .A1(n13821), .A2(n19851), .ZN(n13822) );
  AOI211_X1 U16972 ( .C1(n15536), .C2(n13824), .A(n13823), .B(n13822), .ZN(
        n13825) );
  OAI21_X1 U16973 ( .B1(n19804), .B2(n14009), .A(n13825), .ZN(P1_U2973) );
  INV_X1 U16974 ( .A(n14023), .ZN(n13826) );
  NAND2_X1 U16975 ( .A1(n13827), .A2(n13826), .ZN(n13830) );
  NAND2_X1 U16976 ( .A1(n13839), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13829) );
  MUX2_X1 U16977 ( .A(n13830), .B(n13829), .S(n9615), .Z(n13831) );
  XNOR2_X1 U16978 ( .A(n13831), .B(n14004), .ZN(n14016) );
  NAND2_X1 U16979 ( .A1(n12502), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14011) );
  OAI21_X1 U16980 ( .B1(n13917), .B2(n13832), .A(n14011), .ZN(n13835) );
  NOR2_X1 U16981 ( .A1(n13833), .A2(n19851), .ZN(n13834) );
  AOI211_X1 U16982 ( .C1(n15536), .C2(n13836), .A(n13835), .B(n13834), .ZN(
        n13837) );
  OAI21_X1 U16983 ( .B1(n19804), .B2(n14016), .A(n13837), .ZN(P1_U2974) );
  NOR2_X1 U16984 ( .A1(n13839), .A2(n13848), .ZN(n13838) );
  MUX2_X1 U16985 ( .A(n13839), .B(n13838), .S(n10117), .Z(n13840) );
  XNOR2_X1 U16986 ( .A(n13840), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14027) );
  INV_X1 U16987 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U16988 ( .A1(n12502), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14018) );
  OAI21_X1 U16989 ( .B1(n13917), .B2(n13841), .A(n14018), .ZN(n13844) );
  NOR2_X1 U16990 ( .A1(n13842), .A2(n19851), .ZN(n13843) );
  AOI211_X1 U16991 ( .C1(n15536), .C2(n13845), .A(n13844), .B(n13843), .ZN(
        n13846) );
  OAI21_X1 U16992 ( .B1(n19804), .B2(n14027), .A(n13846), .ZN(P1_U2975) );
  XNOR2_X1 U16993 ( .A(n9615), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13847) );
  XNOR2_X1 U16994 ( .A(n13848), .B(n13847), .ZN(n14036) );
  NAND2_X1 U16995 ( .A1(n12502), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14032) );
  NAND2_X1 U16996 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13849) );
  OAI211_X1 U16997 ( .C1(n19810), .C2(n15427), .A(n14032), .B(n13849), .ZN(
        n13850) );
  AOI21_X1 U16998 ( .B1(n15435), .B2(n19794), .A(n13850), .ZN(n13851) );
  OAI21_X1 U16999 ( .B1(n14036), .B2(n19804), .A(n13851), .ZN(P1_U2976) );
  NAND2_X1 U17000 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  XOR2_X1 U17001 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n13854), .Z(
        n14047) );
  NOR2_X1 U17002 ( .A1(n15601), .A2(n13855), .ZN(n14039) );
  AOI21_X1 U17003 ( .B1(n19799), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14039), .ZN(n13856) );
  OAI21_X1 U17004 ( .B1(n19810), .B2(n13857), .A(n13856), .ZN(n13858) );
  AOI21_X1 U17005 ( .B1(n13859), .B2(n19794), .A(n13858), .ZN(n13860) );
  OAI21_X1 U17006 ( .B1(n19804), .B2(n14047), .A(n13860), .ZN(P1_U2977) );
  INV_X1 U17007 ( .A(n14042), .ZN(n13946) );
  NOR2_X1 U17008 ( .A1(n13880), .A2(n13946), .ZN(n13865) );
  INV_X1 U17009 ( .A(n13880), .ZN(n13861) );
  NAND2_X1 U17010 ( .A1(n13861), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13863) );
  AOI21_X1 U17011 ( .B1(n10117), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n13861), .ZN(n14065) );
  NAND2_X1 U17012 ( .A1(n14065), .A2(n14054), .ZN(n13862) );
  MUX2_X1 U17013 ( .A(n13863), .B(n13862), .S(n10117), .Z(n13871) );
  NOR2_X1 U17014 ( .A1(n13871), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13864) );
  MUX2_X1 U17015 ( .A(n13865), .B(n13864), .S(n10117), .Z(n13866) );
  XNOR2_X1 U17016 ( .A(n13866), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14053) );
  NAND2_X1 U17017 ( .A1(n12502), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14049) );
  NAND2_X1 U17018 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13867) );
  OAI211_X1 U17019 ( .C1(n19810), .C2(n15450), .A(n14049), .B(n13867), .ZN(
        n13868) );
  AOI21_X1 U17020 ( .B1(n13869), .B2(n19794), .A(n13868), .ZN(n13870) );
  OAI21_X1 U17021 ( .B1(n14053), .B2(n19804), .A(n13870), .ZN(P1_U2978) );
  XOR2_X1 U17022 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n13871), .Z(
        n14063) );
  INV_X1 U17023 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n13872) );
  NOR2_X1 U17024 ( .A1(n15601), .A2(n13872), .ZN(n14056) );
  NOR2_X1 U17025 ( .A1(n13917), .A2(n13873), .ZN(n13874) );
  AOI211_X1 U17026 ( .C1(n15536), .C2(n13875), .A(n14056), .B(n13874), .ZN(
        n13879) );
  INV_X1 U17027 ( .A(n13876), .ZN(n13877) );
  NAND2_X1 U17028 ( .A1(n13877), .A2(n19794), .ZN(n13878) );
  OAI211_X1 U17029 ( .C1(n14063), .C2(n19804), .A(n13879), .B(n13878), .ZN(
        P1_U2979) );
  OAI21_X1 U17030 ( .B1(n13882), .B2(n13881), .A(n13880), .ZN(n15566) );
  AOI22_X1 U17031 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n13883) );
  OAI21_X1 U17032 ( .B1(n13884), .B2(n19810), .A(n13883), .ZN(n13885) );
  AOI21_X1 U17033 ( .B1(n13886), .B2(n19794), .A(n13885), .ZN(n13887) );
  OAI21_X1 U17034 ( .B1(n19804), .B2(n15566), .A(n13887), .ZN(P1_U2981) );
  NOR2_X1 U17035 ( .A1(n13889), .A2(n13888), .ZN(n13903) );
  NOR2_X1 U17036 ( .A1(n13903), .A2(n13890), .ZN(n15524) );
  NOR2_X1 U17037 ( .A1(n15524), .A2(n13891), .ZN(n13892) );
  NOR2_X1 U17038 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14076) );
  NOR2_X1 U17039 ( .A1(n13892), .A2(n14076), .ZN(n13894) );
  OAI22_X1 U17040 ( .A1(n13894), .A2(n13893), .B1(n13892), .B2(n9691), .ZN(
        n14084) );
  NAND2_X1 U17041 ( .A1(n12502), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n14080) );
  OAI21_X1 U17042 ( .B1(n13917), .B2(n13895), .A(n14080), .ZN(n13898) );
  NOR2_X1 U17043 ( .A1(n13896), .A2(n19851), .ZN(n13897) );
  AOI211_X1 U17044 ( .C1(n15536), .C2(n13899), .A(n13898), .B(n13897), .ZN(
        n13900) );
  OAI21_X1 U17045 ( .B1(n14084), .B2(n19804), .A(n13900), .ZN(P1_U2983) );
  OAI21_X1 U17046 ( .B1(n13903), .B2(n13902), .A(n13901), .ZN(n13905) );
  XNOR2_X1 U17047 ( .A(n9615), .B(n15589), .ZN(n13904) );
  XNOR2_X1 U17048 ( .A(n13905), .B(n13904), .ZN(n15593) );
  NAND2_X1 U17049 ( .A1(n15593), .A2(n19795), .ZN(n13909) );
  INV_X1 U17050 ( .A(n15479), .ZN(n13907) );
  OAI22_X1 U17051 ( .A1(n13917), .A2(n15476), .B1(n15601), .B2(n13476), .ZN(
        n13906) );
  AOI21_X1 U17052 ( .B1(n15536), .B2(n13907), .A(n13906), .ZN(n13908) );
  OAI211_X1 U17053 ( .C1(n19851), .C2(n15481), .A(n13909), .B(n13908), .ZN(
        P1_U2985) );
  OAI21_X1 U17054 ( .B1(n13910), .B2(n13912), .A(n13911), .ZN(n15533) );
  NAND2_X1 U17055 ( .A1(n9982), .A2(n13913), .ZN(n15532) );
  NOR2_X1 U17056 ( .A1(n15533), .A2(n15532), .ZN(n15531) );
  NOR2_X1 U17057 ( .A1(n15531), .A2(n13914), .ZN(n13915) );
  INV_X1 U17058 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13916) );
  NAND2_X1 U17059 ( .A1(n12502), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n14085) );
  OAI21_X1 U17060 ( .B1(n13917), .B2(n13916), .A(n14085), .ZN(n13920) );
  NOR2_X1 U17061 ( .A1(n13918), .A2(n19851), .ZN(n13919) );
  AOI211_X1 U17062 ( .C1(n15536), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        n13922) );
  OAI21_X1 U17063 ( .B1(n19804), .B2(n14092), .A(n13922), .ZN(P1_U2986) );
  MUX2_X1 U17064 ( .A(n14093), .B(n13910), .S(n9615), .Z(n13923) );
  XNOR2_X1 U17065 ( .A(n13923), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15614) );
  NAND2_X1 U17066 ( .A1(n15614), .A2(n19795), .ZN(n13927) );
  NOR2_X1 U17067 ( .A1(n15601), .A2(n20570), .ZN(n15612) );
  NOR2_X1 U17068 ( .A1(n19810), .A2(n13924), .ZN(n13925) );
  AOI211_X1 U17069 ( .C1(n19799), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15612), .B(n13925), .ZN(n13926) );
  OAI211_X1 U17070 ( .C1(n19851), .C2(n13928), .A(n13927), .B(n13926), .ZN(
        P1_U2989) );
  NAND3_X1 U17071 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15575) );
  NOR2_X1 U17072 ( .A1(n15574), .A2(n15575), .ZN(n15565) );
  INV_X1 U17073 ( .A(n15565), .ZN(n15562) );
  NOR2_X1 U17074 ( .A1(n15572), .A2(n15562), .ZN(n13939) );
  INV_X1 U17075 ( .A(n19815), .ZN(n13932) );
  INV_X1 U17076 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14094) );
  NOR2_X1 U17077 ( .A1(n14094), .A2(n13930), .ZN(n15619) );
  NAND4_X1 U17078 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n15619), .ZN(n14100) );
  NOR4_X1 U17079 ( .A1(n15624), .A2(n13932), .A3(n13931), .A4(n14100), .ZN(
        n14101) );
  NAND3_X1 U17080 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n14101), .ZN(n13940) );
  NOR2_X1 U17081 ( .A1(n13933), .A2(n13940), .ZN(n13934) );
  NAND2_X1 U17082 ( .A1(n15611), .A2(n15619), .ZN(n14099) );
  NOR3_X1 U17083 ( .A1(n13196), .A2(n14097), .A3(n14099), .ZN(n13941) );
  AOI22_X1 U17084 ( .A1(n13934), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19831), .B2(n13941), .ZN(n14059) );
  OAI21_X1 U17085 ( .B1(n14058), .B2(n13940), .A(n14059), .ZN(n14090) );
  NAND2_X1 U17086 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14090), .ZN(
        n15583) );
  INV_X1 U17087 ( .A(n15583), .ZN(n13935) );
  NAND2_X1 U17088 ( .A1(n13939), .A2(n13935), .ZN(n14066) );
  NOR2_X1 U17089 ( .A1(n13999), .A2(n13937), .ZN(n13938) );
  NAND3_X1 U17090 ( .A1(n13991), .A2(n9882), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13958) );
  INV_X1 U17091 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14121) );
  NAND2_X1 U17092 ( .A1(n14121), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13952) );
  INV_X1 U17093 ( .A(n15629), .ZN(n15563) );
  INV_X1 U17094 ( .A(n13939), .ZN(n13943) );
  OR2_X1 U17095 ( .A1(n14089), .A2(n13940), .ZN(n14072) );
  AOI221_X1 U17096 ( .B1(n13943), .B2(n14073), .C1(n14072), .C2(n14073), .A(
        n14103), .ZN(n13945) );
  AND2_X1 U17097 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n13941), .ZN(
        n15590) );
  INV_X1 U17098 ( .A(n15590), .ZN(n13942) );
  OAI21_X1 U17099 ( .B1(n13943), .B2(n13942), .A(n19831), .ZN(n13944) );
  NAND2_X1 U17100 ( .A1(n13945), .A2(n13944), .ZN(n14069) );
  AOI21_X1 U17101 ( .B1(n13946), .B2(n15563), .A(n14069), .ZN(n13947) );
  INV_X1 U17102 ( .A(n13947), .ZN(n14051) );
  NAND2_X1 U17103 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13948) );
  NAND2_X1 U17104 ( .A1(n13947), .A2(n15629), .ZN(n13977) );
  OAI21_X1 U17105 ( .B1(n14051), .B2(n13948), .A(n13977), .ZN(n14028) );
  OAI21_X1 U17106 ( .B1(n14022), .B2(n15629), .A(n14028), .ZN(n14014) );
  AND2_X1 U17107 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13979) );
  NAND2_X1 U17108 ( .A1(n9882), .A2(n13979), .ZN(n13949) );
  OAI21_X1 U17109 ( .B1(n14014), .B2(n13949), .A(n13977), .ZN(n13971) );
  OAI211_X1 U17110 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15629), .A(
        n13971), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13956) );
  NAND3_X1 U17111 ( .A1(n13956), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13977), .ZN(n13951) );
  OAI211_X1 U17112 ( .C1(n13958), .C2(n13952), .A(n13951), .B(n13950), .ZN(
        n13953) );
  INV_X1 U17113 ( .A(n13955), .ZN(n13961) );
  INV_X1 U17114 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13959) );
  INV_X1 U17115 ( .A(n13956), .ZN(n13957) );
  AOI21_X1 U17116 ( .B1(n13959), .B2(n13958), .A(n13957), .ZN(n13960) );
  AOI211_X1 U17117 ( .C1(n19825), .C2(n13962), .A(n13961), .B(n13960), .ZN(
        n13963) );
  OAI21_X1 U17118 ( .B1(n13964), .B2(n19838), .A(n13963), .ZN(P1_U3001) );
  INV_X1 U17119 ( .A(n13965), .ZN(n13970) );
  INV_X1 U17120 ( .A(n13991), .ZN(n13967) );
  NOR3_X1 U17121 ( .A1(n13967), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13966), .ZN(n13968) );
  AOI211_X1 U17122 ( .C1(n13970), .C2(n19825), .A(n13969), .B(n13968), .ZN(
        n13974) );
  INV_X1 U17123 ( .A(n13971), .ZN(n13972) );
  NAND2_X1 U17124 ( .A1(n13972), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13973) );
  OAI211_X1 U17125 ( .C1(n13975), .C2(n19838), .A(n13974), .B(n13973), .ZN(
        P1_U3002) );
  INV_X1 U17126 ( .A(n13976), .ZN(n13988) );
  INV_X1 U17127 ( .A(n14014), .ZN(n13980) );
  INV_X1 U17128 ( .A(n13977), .ZN(n13978) );
  AOI21_X1 U17129 ( .B1(n13980), .B2(n13979), .A(n13978), .ZN(n13995) );
  NOR2_X1 U17130 ( .A1(n13981), .A2(n9882), .ZN(n13983) );
  AOI21_X1 U17131 ( .B1(n13991), .B2(n13983), .A(n13982), .ZN(n13984) );
  OAI21_X1 U17132 ( .B1(n13985), .B2(n19834), .A(n13984), .ZN(n13986) );
  AOI21_X1 U17133 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n13995), .A(
        n13986), .ZN(n13987) );
  OAI21_X1 U17134 ( .B1(n13988), .B2(n19838), .A(n13987), .ZN(P1_U3003) );
  AOI21_X1 U17135 ( .B1(n13991), .B2(n13990), .A(n13989), .ZN(n13992) );
  OAI21_X1 U17136 ( .B1(n13993), .B2(n19834), .A(n13992), .ZN(n13994) );
  AOI21_X1 U17137 ( .B1(n13995), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13994), .ZN(n13996) );
  OAI21_X1 U17138 ( .B1(n13997), .B2(n19838), .A(n13996), .ZN(P1_U3004) );
  INV_X1 U17139 ( .A(n13998), .ZN(n14002) );
  INV_X1 U17140 ( .A(n14030), .ZN(n14000) );
  NOR3_X1 U17141 ( .A1(n14000), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n13999), .ZN(n14001) );
  AOI211_X1 U17142 ( .C1(n14003), .C2(n19825), .A(n14002), .B(n14001), .ZN(
        n14008) );
  AND2_X1 U17143 ( .A1(n14022), .A2(n14004), .ZN(n14005) );
  NAND2_X1 U17144 ( .A1(n14030), .A2(n14005), .ZN(n14010) );
  INV_X1 U17145 ( .A(n14010), .ZN(n14006) );
  OAI21_X1 U17146 ( .B1(n14014), .B2(n14006), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14007) );
  OAI211_X1 U17147 ( .C1(n14009), .C2(n19838), .A(n14008), .B(n14007), .ZN(
        P1_U3005) );
  OAI211_X1 U17148 ( .C1(n14012), .C2(n19834), .A(n14011), .B(n14010), .ZN(
        n14013) );
  AOI21_X1 U17149 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14014), .A(
        n14013), .ZN(n14015) );
  OAI21_X1 U17150 ( .B1(n14016), .B2(n19838), .A(n14015), .ZN(P1_U3006) );
  INV_X1 U17151 ( .A(n14017), .ZN(n14020) );
  INV_X1 U17152 ( .A(n14018), .ZN(n14019) );
  AOI21_X1 U17153 ( .B1(n14020), .B2(n19825), .A(n14019), .ZN(n14026) );
  INV_X1 U17154 ( .A(n15597), .ZN(n19842) );
  NOR2_X1 U17155 ( .A1(n19842), .A2(n19831), .ZN(n14021) );
  OAI21_X1 U17156 ( .B1(n14022), .B2(n14021), .A(n14028), .ZN(n14024) );
  OAI211_X1 U17157 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14030), .A(
        n14024), .B(n14023), .ZN(n14025) );
  OAI211_X1 U17158 ( .C1(n14027), .C2(n19838), .A(n14026), .B(n14025), .ZN(
        P1_U3007) );
  INV_X1 U17159 ( .A(n14028), .ZN(n14034) );
  NAND2_X1 U17160 ( .A1(n14030), .A2(n14029), .ZN(n14031) );
  OAI211_X1 U17161 ( .C1(n15438), .C2(n19834), .A(n14032), .B(n14031), .ZN(
        n14033) );
  AOI21_X1 U17162 ( .B1(n14034), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14033), .ZN(n14035) );
  OAI21_X1 U17163 ( .B1(n14036), .B2(n19838), .A(n14035), .ZN(P1_U3008) );
  NOR2_X1 U17164 ( .A1(n14037), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14038) );
  AOI211_X1 U17165 ( .C1(n14040), .C2(n19825), .A(n14039), .B(n14038), .ZN(
        n14046) );
  NAND2_X1 U17166 ( .A1(n14042), .A2(n14041), .ZN(n14043) );
  OR2_X1 U17167 ( .A1(n14066), .A2(n14043), .ZN(n14048) );
  INV_X1 U17168 ( .A(n14048), .ZN(n14044) );
  OAI21_X1 U17169 ( .B1(n14051), .B2(n14044), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14045) );
  OAI211_X1 U17170 ( .C1(n14047), .C2(n19838), .A(n14046), .B(n14045), .ZN(
        P1_U3009) );
  OAI211_X1 U17171 ( .C1(n15444), .C2(n19834), .A(n14049), .B(n14048), .ZN(
        n14050) );
  AOI21_X1 U17172 ( .B1(n14051), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14050), .ZN(n14052) );
  OAI21_X1 U17173 ( .B1(n14053), .B2(n19838), .A(n14052), .ZN(P1_U3010) );
  NOR3_X1 U17174 ( .A1(n14066), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n14054), .ZN(n14055) );
  AOI211_X1 U17175 ( .C1(n14057), .C2(n19825), .A(n14056), .B(n14055), .ZN(
        n14062) );
  AOI21_X1 U17176 ( .B1(n14059), .B2(n14058), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14060) );
  OAI21_X1 U17177 ( .B1(n14069), .B2(n14060), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14061) );
  OAI211_X1 U17178 ( .C1(n14063), .C2(n19838), .A(n14062), .B(n14061), .ZN(
        P1_U3011) );
  XNOR2_X1 U17179 ( .A(n9615), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14064) );
  XNOR2_X1 U17180 ( .A(n14065), .B(n14064), .ZN(n15511) );
  INV_X1 U17181 ( .A(n15511), .ZN(n14071) );
  NOR2_X1 U17182 ( .A1(n15465), .A2(n19834), .ZN(n14068) );
  OAI22_X1 U17183 ( .A1(n14066), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20449), .B2(n15601), .ZN(n14067) );
  AOI211_X1 U17184 ( .C1(n14069), .C2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14068), .B(n14067), .ZN(n14070) );
  OAI21_X1 U17185 ( .B1(n14071), .B2(n19838), .A(n14070), .ZN(P1_U3012) );
  AOI21_X1 U17186 ( .B1(n14073), .B2(n14072), .A(n14103), .ZN(n14074) );
  OAI21_X1 U17187 ( .B1(n15590), .B2(n19812), .A(n14074), .ZN(n15591) );
  INV_X1 U17188 ( .A(n15591), .ZN(n14075) );
  OAI21_X1 U17189 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15629), .A(
        n14075), .ZN(n15582) );
  NAND2_X1 U17190 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14078) );
  NOR3_X1 U17191 ( .A1(n14076), .A2(n15583), .A3(n15589), .ZN(n14077) );
  NAND2_X1 U17192 ( .A1(n14078), .A2(n14077), .ZN(n14079) );
  OAI211_X1 U17193 ( .C1(n14081), .C2(n19834), .A(n14080), .B(n14079), .ZN(
        n14082) );
  AOI21_X1 U17194 ( .B1(n15582), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14082), .ZN(n14083) );
  OAI21_X1 U17195 ( .B1(n14084), .B2(n19838), .A(n14083), .ZN(P1_U3015) );
  NAND2_X1 U17196 ( .A1(n15591), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14086) );
  OAI211_X1 U17197 ( .C1(n19834), .C2(n14087), .A(n14086), .B(n14085), .ZN(
        n14088) );
  AOI21_X1 U17198 ( .B1(n14090), .B2(n14089), .A(n14088), .ZN(n14091) );
  OAI21_X1 U17199 ( .B1(n14092), .B2(n19838), .A(n14091), .ZN(P1_U3018) );
  NOR2_X1 U17200 ( .A1(n14093), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14096) );
  NOR2_X1 U17201 ( .A1(n13910), .A2(n14094), .ZN(n14095) );
  MUX2_X1 U17202 ( .A(n14096), .B(n14095), .S(n9615), .Z(n14098) );
  XNOR2_X1 U17203 ( .A(n14098), .B(n14097), .ZN(n15540) );
  NOR2_X1 U17204 ( .A1(n15606), .A2(n14099), .ZN(n14105) );
  NOR2_X1 U17205 ( .A1(n14097), .A2(n14100), .ZN(n15607) );
  OAI22_X1 U17206 ( .A1(n15626), .A2(n14101), .B1(n15607), .B2(n19812), .ZN(
        n14102) );
  AOI211_X1 U17207 ( .C1(n19831), .C2(n15605), .A(n14103), .B(n14102), .ZN(
        n15598) );
  INV_X1 U17208 ( .A(n15598), .ZN(n14104) );
  MUX2_X1 U17209 ( .A(n14105), .B(n14104), .S(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(n14108) );
  INV_X1 U17210 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n14106) );
  OAI22_X1 U17211 ( .A1(n15499), .A2(n19834), .B1(n15601), .B2(n14106), .ZN(
        n14107) );
  AOI211_X1 U17212 ( .C1(n15540), .C2(n19823), .A(n14108), .B(n14107), .ZN(
        n14109) );
  INV_X1 U17213 ( .A(n14109), .ZN(P1_U3020) );
  NOR2_X1 U17214 ( .A1(n14111), .A2(n14110), .ZN(n14114) );
  INV_X1 U17215 ( .A(n14114), .ZN(n14123) );
  NAND2_X1 U17216 ( .A1(n14113), .A2(n14112), .ZN(n14117) );
  NAND2_X1 U17217 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  OAI211_X1 U17218 ( .C1(n20111), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        n15358) );
  NOR2_X1 U17219 ( .A1(n20400), .A2(n14119), .ZN(n14127) );
  OAI22_X1 U17220 ( .A1(n14121), .A2(n14120), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17221 ( .A1(n15358), .A2(n14128), .B1(n14127), .B2(n14125), .ZN(
        n14122) );
  OAI21_X1 U17222 ( .B1(n14132), .B2(n14123), .A(n14122), .ZN(n14124) );
  MUX2_X1 U17223 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14124), .S(
        n14133), .Z(P1_U3473) );
  INV_X1 U17224 ( .A(n14125), .ZN(n14126) );
  AOI22_X1 U17225 ( .A1(n14129), .A2(n14128), .B1(n14127), .B2(n14126), .ZN(
        n14130) );
  OAI21_X1 U17226 ( .B1(n14132), .B2(n14131), .A(n14130), .ZN(n14134) );
  MUX2_X1 U17227 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14134), .S(
        n14133), .Z(P1_U3472) );
  INV_X1 U17228 ( .A(n14627), .ZN(n14172) );
  XOR2_X1 U17229 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n14135), .Z(
        n14437) );
  INV_X1 U17230 ( .A(n14137), .ZN(n14136) );
  AOI21_X1 U17231 ( .B1(n14446), .B2(n14136), .A(n14135), .ZN(n14444) );
  INV_X1 U17232 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14461) );
  INV_X1 U17233 ( .A(n14139), .ZN(n14138) );
  AOI21_X1 U17234 ( .B1(n14461), .B2(n14138), .A(n14137), .ZN(n14464) );
  AOI21_X1 U17235 ( .B1(n14469), .B2(n14158), .A(n14139), .ZN(n14472) );
  INV_X1 U17236 ( .A(n14156), .ZN(n14140) );
  AOI21_X1 U17237 ( .B1(n14487), .B2(n14142), .A(n14140), .ZN(n15680) );
  OR2_X1 U17238 ( .A1(n14143), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14141) );
  NAND2_X1 U17239 ( .A1(n14142), .A2(n14141), .ZN(n15697) );
  AOI21_X1 U17240 ( .B1(n20563), .B2(n14153), .A(n14143), .ZN(n15734) );
  INV_X1 U17241 ( .A(n15734), .ZN(n15709) );
  AOI21_X1 U17242 ( .B1(n18522), .B2(n14144), .A(n14154), .ZN(n18528) );
  OAI21_X1 U17243 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9705), .A(
        n14144), .ZN(n14532) );
  AOI21_X1 U17244 ( .B1(n14543), .B2(n14151), .A(n9705), .ZN(n18534) );
  AOI21_X1 U17245 ( .B1(n14145), .B2(n14149), .A(n14152), .ZN(n18559) );
  AOI21_X1 U17246 ( .B1(n14147), .B2(n14146), .A(n14150), .ZN(n18581) );
  NAND2_X1 U17247 ( .A1(n14148), .A2(n15766), .ZN(n18580) );
  NOR2_X1 U17248 ( .A1(n18581), .A2(n18580), .ZN(n18570) );
  OAI21_X1 U17249 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14150), .A(
        n14149), .ZN(n18571) );
  NAND2_X1 U17250 ( .A1(n18570), .A2(n18571), .ZN(n18557) );
  NOR2_X1 U17251 ( .A1(n18559), .A2(n18557), .ZN(n18544) );
  OAI21_X1 U17252 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14152), .A(
        n14151), .ZN(n18545) );
  NAND2_X1 U17253 ( .A1(n18544), .A2(n18545), .ZN(n18532) );
  OAI21_X1 U17254 ( .B1(n18534), .B2(n18532), .A(n18669), .ZN(n14225) );
  NAND2_X1 U17255 ( .A1(n14532), .A2(n14225), .ZN(n14224) );
  NAND2_X1 U17256 ( .A1(n18669), .A2(n14224), .ZN(n18525) );
  OAI21_X1 U17257 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14154), .A(
        n14153), .ZN(n15749) );
  NAND2_X1 U17258 ( .A1(n15709), .A2(n15708), .ZN(n15707) );
  NAND2_X1 U17259 ( .A1(n18669), .A2(n15707), .ZN(n15696) );
  NAND2_X1 U17260 ( .A1(n15697), .A2(n15696), .ZN(n15695) );
  OAI21_X1 U17261 ( .B1(n15680), .B2(n15695), .A(n18669), .ZN(n15674) );
  NAND2_X1 U17262 ( .A1(n14156), .A2(n14155), .ZN(n14157) );
  NAND2_X1 U17263 ( .A1(n14158), .A2(n14157), .ZN(n15673) );
  NAND2_X1 U17264 ( .A1(n15674), .A2(n15673), .ZN(n15672) );
  AND2_X1 U17265 ( .A1(n18669), .A2(n15672), .ZN(n14220) );
  NOR2_X1 U17266 ( .A1(n14472), .A2(n14220), .ZN(n14219) );
  NOR2_X1 U17267 ( .A1(n18653), .A2(n14189), .ZN(n14174) );
  NOR2_X1 U17268 ( .A1(n18653), .A2(n19465), .ZN(n14159) );
  NAND2_X1 U17269 ( .A1(n14173), .A2(n14159), .ZN(n14171) );
  AOI22_X1 U17270 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n14160), .B2(P2_EAX_REG_31__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U17271 ( .A1(n10996), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U17272 ( .A1(n14165), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18677), .ZN(n14167) );
  NAND2_X1 U17273 ( .A1(n18667), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14166) );
  OAI211_X1 U17274 ( .C1(n18696), .C2(n18676), .A(n14167), .B(n14166), .ZN(
        n14168) );
  AOI21_X1 U17275 ( .B1(n14169), .B2(n18639), .A(n14168), .ZN(n14170) );
  OAI211_X1 U17276 ( .C1(n14172), .C2(n18656), .A(n14171), .B(n14170), .ZN(
        P2_U2824) );
  INV_X1 U17277 ( .A(n14635), .ZN(n14177) );
  NAND2_X1 U17278 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18677), .ZN(
        n14176) );
  AOI22_X1 U17279 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n18563), .ZN(n14175) );
  OAI211_X1 U17280 ( .C1(n14177), .C2(n18676), .A(n14176), .B(n14175), .ZN(
        n14178) );
  AOI21_X1 U17281 ( .B1(n14179), .B2(n18639), .A(n14178), .ZN(n14180) );
  AOI21_X1 U17282 ( .B1(n14182), .B2(n14196), .A(n14181), .ZN(n14645) );
  INV_X1 U17283 ( .A(n14645), .ZN(n14256) );
  OR2_X1 U17284 ( .A1(n14200), .A2(n14183), .ZN(n14184) );
  NAND2_X1 U17285 ( .A1(n14185), .A2(n14184), .ZN(n14352) );
  AOI22_X1 U17286 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n18563), .ZN(n14188) );
  AOI22_X1 U17287 ( .A1(n14186), .A2(n18639), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18677), .ZN(n14187) );
  OAI211_X1 U17288 ( .C1(n14352), .C2(n18676), .A(n14188), .B(n14187), .ZN(
        n14192) );
  AOI211_X1 U17289 ( .C1(n14444), .C2(n14190), .A(n14189), .B(n19465), .ZN(
        n14191) );
  NOR2_X1 U17290 ( .A1(n14192), .A2(n14191), .ZN(n14193) );
  OAI21_X1 U17291 ( .B1(n14256), .B2(n18656), .A(n14193), .ZN(P2_U2826) );
  NAND2_X1 U17292 ( .A1(n14211), .A2(n14194), .ZN(n14195) );
  NAND2_X1 U17293 ( .A1(n14196), .A2(n14195), .ZN(n14664) );
  AOI211_X1 U17294 ( .C1(n14464), .C2(n14198), .A(n14197), .B(n19465), .ZN(
        n14199) );
  INV_X1 U17295 ( .A(n14199), .ZN(n14208) );
  INV_X1 U17296 ( .A(n14200), .ZN(n14201) );
  OAI21_X1 U17297 ( .B1(n14213), .B2(n14202), .A(n14201), .ZN(n14663) );
  NAND2_X1 U17298 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18677), .ZN(
        n14204) );
  AOI22_X1 U17299 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n18563), .ZN(n14203) );
  OAI211_X1 U17300 ( .C1(n14663), .C2(n18676), .A(n14204), .B(n14203), .ZN(
        n14205) );
  AOI21_X1 U17301 ( .B1(n14206), .B2(n18639), .A(n14205), .ZN(n14207) );
  OAI211_X1 U17302 ( .C1(n18656), .C2(n14664), .A(n14208), .B(n14207), .ZN(
        P2_U2827) );
  OR2_X1 U17303 ( .A1(n14268), .A2(n14209), .ZN(n14210) );
  NAND2_X1 U17304 ( .A1(n14211), .A2(n14210), .ZN(n14673) );
  AND2_X1 U17305 ( .A1(n14373), .A2(n14212), .ZN(n14214) );
  OR2_X1 U17306 ( .A1(n14214), .A2(n14213), .ZN(n14678) );
  AOI22_X1 U17307 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n18563), .ZN(n14218) );
  OAI22_X1 U17308 ( .A1(n14215), .A2(n18687), .B1(n18663), .B2(n14469), .ZN(
        n14216) );
  INV_X1 U17309 ( .A(n14216), .ZN(n14217) );
  OAI211_X1 U17310 ( .C1(n14678), .C2(n18676), .A(n14218), .B(n14217), .ZN(
        n14222) );
  AOI211_X1 U17311 ( .C1(n14472), .C2(n14220), .A(n14219), .B(n19465), .ZN(
        n14221) );
  NOR2_X1 U17312 ( .A1(n14222), .A2(n14221), .ZN(n14223) );
  OAI21_X1 U17313 ( .B1(n14673), .B2(n18656), .A(n14223), .ZN(P2_U2828) );
  OAI211_X1 U17314 ( .C1(n14532), .C2(n14225), .A(n18678), .B(n14224), .ZN(
        n14235) );
  AND2_X1 U17315 ( .A1(n14320), .A2(n14226), .ZN(n14227) );
  NOR2_X1 U17316 ( .A1(n14310), .A2(n14227), .ZN(n14754) );
  NOR2_X1 U17317 ( .A1(n14417), .A2(n14228), .ZN(n14229) );
  NOR2_X1 U17318 ( .A1(n14406), .A2(n14229), .ZN(n15721) );
  OAI22_X1 U17319 ( .A1(n18679), .A2(n12090), .B1(n19515), .B2(n18681), .ZN(
        n14231) );
  NOR2_X1 U17320 ( .A1(n18663), .A2(n10004), .ZN(n14230) );
  AOI211_X1 U17321 ( .C1(n15721), .C2(n18684), .A(n14231), .B(n14230), .ZN(
        n14232) );
  INV_X1 U17322 ( .A(n14232), .ZN(n14233) );
  AOI21_X1 U17323 ( .B1(n14754), .B2(n18689), .A(n14233), .ZN(n14234) );
  OAI211_X1 U17324 ( .C1(n14236), .C2(n18687), .A(n14235), .B(n14234), .ZN(
        P2_U2835) );
  INV_X1 U17325 ( .A(n18808), .ZN(n14240) );
  OAI22_X1 U17326 ( .A1(n18679), .A2(n10310), .B1(n19486), .B2(n18681), .ZN(
        n14239) );
  NOR2_X1 U17327 ( .A1(n18663), .A2(n14237), .ZN(n14238) );
  AOI211_X1 U17328 ( .C1(n18639), .C2(n14240), .A(n14239), .B(n14238), .ZN(
        n14242) );
  NAND2_X1 U17329 ( .A1(n19568), .A2(n18684), .ZN(n14241) );
  OAI211_X1 U17330 ( .C1(n12734), .C2(n18656), .A(n14242), .B(n14241), .ZN(
        n14247) );
  OAI21_X1 U17331 ( .B1(n14245), .B2(n14244), .A(n14243), .ZN(n14908) );
  AOI221_X1 U17332 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n14908), .C1(
        n18669), .C2(n14908), .A(n19465), .ZN(n14246) );
  AOI211_X1 U17333 ( .C1(n18691), .C2(n19565), .A(n14247), .B(n14246), .ZN(
        n14248) );
  INV_X1 U17334 ( .A(n14248), .ZN(P2_U2854) );
  INV_X1 U17335 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U17336 ( .A1(n14627), .A2(n14350), .ZN(n14249) );
  OAI21_X1 U17337 ( .B1(n14350), .B2(n14250), .A(n14249), .ZN(P2_U2856) );
  OR2_X1 U17338 ( .A1(n14252), .A2(n14251), .ZN(n14351) );
  NAND3_X1 U17339 ( .A1(n14351), .A2(n14253), .A3(n14344), .ZN(n14255) );
  NAND2_X1 U17340 ( .A1(n14340), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14254) );
  OAI211_X1 U17341 ( .C1(n14340), .C2(n14256), .A(n14255), .B(n14254), .ZN(
        P2_U2858) );
  NOR2_X1 U17342 ( .A1(n9910), .A2(n14257), .ZN(n14258) );
  XNOR2_X1 U17343 ( .A(n14258), .B(n9717), .ZN(n14362) );
  NAND2_X1 U17344 ( .A1(n14362), .A2(n14344), .ZN(n14260) );
  NAND2_X1 U17345 ( .A1(n14340), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14259) );
  OAI211_X1 U17346 ( .C1(n14664), .C2(n14340), .A(n14260), .B(n14259), .ZN(
        P2_U2859) );
  AOI21_X1 U17347 ( .B1(n14263), .B2(n14262), .A(n14261), .ZN(n14368) );
  NAND2_X1 U17348 ( .A1(n14368), .A2(n14344), .ZN(n14265) );
  NAND2_X1 U17349 ( .A1(n14340), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14264) );
  OAI211_X1 U17350 ( .C1(n14673), .C2(n14340), .A(n14265), .B(n14264), .ZN(
        P2_U2860) );
  NOR2_X1 U17351 ( .A1(n14277), .A2(n14266), .ZN(n14267) );
  OR2_X1 U17352 ( .A1(n14268), .A2(n14267), .ZN(n15670) );
  AOI21_X1 U17353 ( .B1(n14271), .B2(n14270), .A(n14269), .ZN(n14370) );
  NAND2_X1 U17354 ( .A1(n14370), .A2(n14344), .ZN(n14273) );
  NAND2_X1 U17355 ( .A1(n14340), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14272) );
  OAI211_X1 U17356 ( .C1(n15670), .C2(n14340), .A(n14273), .B(n14272), .ZN(
        P2_U2861) );
  OAI21_X1 U17357 ( .B1(n14276), .B2(n14275), .A(n14274), .ZN(n14386) );
  INV_X1 U17358 ( .A(n14277), .ZN(n14278) );
  OAI21_X1 U17359 ( .B1(n14282), .B2(n14279), .A(n14278), .ZN(n15684) );
  MUX2_X1 U17360 ( .A(n20558), .B(n15684), .S(n14333), .Z(n14280) );
  OAI21_X1 U17361 ( .B1(n14386), .B2(n14342), .A(n14280), .ZN(P2_U2862) );
  AND2_X1 U17362 ( .A1(n9656), .A2(n14281), .ZN(n14283) );
  OR2_X1 U17363 ( .A1(n14283), .A2(n14282), .ZN(n15693) );
  AOI21_X1 U17364 ( .B1(n14285), .B2(n14284), .A(n9687), .ZN(n14287) );
  XNOR2_X1 U17365 ( .A(n14287), .B(n14286), .ZN(n14394) );
  NAND2_X1 U17366 ( .A1(n14394), .A2(n14344), .ZN(n14289) );
  NAND2_X1 U17367 ( .A1(n14340), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14288) );
  OAI211_X1 U17368 ( .C1(n15693), .C2(n14340), .A(n14289), .B(n14288), .ZN(
        P2_U2863) );
  AOI21_X1 U17369 ( .B1(n14292), .B2(n14291), .A(n14290), .ZN(n14403) );
  NAND2_X1 U17370 ( .A1(n14403), .A2(n14344), .ZN(n14296) );
  NAND2_X1 U17371 ( .A1(n14299), .A2(n14293), .ZN(n14294) );
  AND2_X1 U17372 ( .A1(n9656), .A2(n14294), .ZN(n15738) );
  NAND2_X1 U17373 ( .A1(n15738), .A2(n14350), .ZN(n14295) );
  OAI211_X1 U17374 ( .C1(n14333), .C2(n12101), .A(n14296), .B(n14295), .ZN(
        P2_U2864) );
  NAND2_X1 U17375 ( .A1(n14308), .A2(n14297), .ZN(n14298) );
  NAND2_X1 U17376 ( .A1(n14299), .A2(n14298), .ZN(n15743) );
  AOI21_X1 U17377 ( .B1(n14302), .B2(n14306), .A(n14301), .ZN(n15716) );
  NAND2_X1 U17378 ( .A1(n15716), .A2(n14344), .ZN(n14304) );
  NAND2_X1 U17379 ( .A1(n14340), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14303) );
  OAI211_X1 U17380 ( .C1(n15743), .C2(n14340), .A(n14304), .B(n14303), .ZN(
        P2_U2865) );
  OAI21_X1 U17381 ( .B1(n14305), .B2(n14307), .A(n14306), .ZN(n14414) );
  OAI21_X1 U17382 ( .B1(n14310), .B2(n14309), .A(n14308), .ZN(n15421) );
  MUX2_X1 U17383 ( .A(n14311), .B(n15421), .S(n14333), .Z(n14312) );
  OAI21_X1 U17384 ( .B1(n14414), .B2(n14342), .A(n14312), .ZN(P2_U2866) );
  NOR2_X1 U17385 ( .A1(n14313), .A2(n14314), .ZN(n14315) );
  OR2_X1 U17386 ( .A1(n14305), .A2(n14315), .ZN(n15724) );
  NOR2_X1 U17387 ( .A1(n14350), .A2(n12090), .ZN(n14316) );
  AOI21_X1 U17388 ( .B1(n14754), .B2(n14350), .A(n14316), .ZN(n14317) );
  OAI21_X1 U17389 ( .B1(n15724), .B2(n14342), .A(n14317), .ZN(P2_U2867) );
  NAND2_X1 U17390 ( .A1(n14329), .A2(n14318), .ZN(n14319) );
  NAND2_X1 U17391 ( .A1(n14320), .A2(n14319), .ZN(n18539) );
  AOI21_X1 U17392 ( .B1(n14322), .B2(n14321), .A(n14313), .ZN(n14422) );
  NAND2_X1 U17393 ( .A1(n14422), .A2(n14344), .ZN(n14324) );
  NAND2_X1 U17394 ( .A1(n14340), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14323) );
  OAI211_X1 U17395 ( .C1(n18539), .C2(n14340), .A(n14324), .B(n14323), .ZN(
        P2_U2868) );
  AOI21_X1 U17396 ( .B1(n14326), .B2(n14325), .A(n10091), .ZN(n15730) );
  NAND2_X1 U17397 ( .A1(n15730), .A2(n14344), .ZN(n14331) );
  OR2_X1 U17398 ( .A1(n14338), .A2(n14327), .ZN(n14328) );
  NAND2_X1 U17399 ( .A1(n14329), .A2(n14328), .ZN(n18552) );
  INV_X1 U17400 ( .A(n18552), .ZN(n15752) );
  NAND2_X1 U17401 ( .A1(n15752), .A2(n14350), .ZN(n14330) );
  OAI211_X1 U17402 ( .C1(n14333), .C2(n14332), .A(n14331), .B(n14330), .ZN(
        P2_U2869) );
  OAI21_X1 U17403 ( .B1(n14334), .B2(n14335), .A(n14325), .ZN(n14431) );
  NOR2_X1 U17404 ( .A1(n14345), .A2(n14336), .ZN(n14337) );
  OR2_X1 U17405 ( .A1(n14338), .A2(n14337), .ZN(n18565) );
  NOR2_X1 U17406 ( .A1(n18565), .A2(n14340), .ZN(n14339) );
  AOI21_X1 U17407 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n14340), .A(n14339), .ZN(
        n14341) );
  OAI21_X1 U17408 ( .B1(n14431), .B2(n14342), .A(n14341), .ZN(P2_U2870) );
  AOI21_X1 U17409 ( .B1(n14343), .B2(n13083), .A(n14334), .ZN(n18705) );
  NAND2_X1 U17410 ( .A1(n18705), .A2(n14344), .ZN(n14349) );
  AOI21_X1 U17411 ( .B1(n14347), .B2(n14346), .A(n14345), .ZN(n18576) );
  NAND2_X1 U17412 ( .A1(n18576), .A2(n14350), .ZN(n14348) );
  OAI211_X1 U17413 ( .C1(n14350), .C2(n9804), .A(n14349), .B(n14348), .ZN(
        P2_U2871) );
  NAND3_X1 U17414 ( .A1(n14351), .A2(n14253), .A3(n18761), .ZN(n14358) );
  INV_X1 U17415 ( .A(n14352), .ZN(n14649) );
  INV_X1 U17416 ( .A(n18701), .ZN(n14354) );
  OAI22_X1 U17417 ( .A1(n14354), .A2(n18714), .B1(n18755), .B2(n14353), .ZN(
        n14355) );
  AOI21_X1 U17418 ( .B1(n18757), .B2(n14649), .A(n14355), .ZN(n14357) );
  AOI22_X1 U17419 ( .A1(n18703), .A2(BUF1_REG_29__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14356) );
  NAND3_X1 U17420 ( .A1(n14358), .A2(n14357), .A3(n14356), .ZN(P2_U2890) );
  AOI22_X1 U17421 ( .A1(n18703), .A2(BUF1_REG_28__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U17422 ( .A1(n18701), .A2(n18717), .B1(n18756), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n14359) );
  OAI211_X1 U17423 ( .C1(n15723), .C2(n14663), .A(n14360), .B(n14359), .ZN(
        n14361) );
  AOI21_X1 U17424 ( .B1(n14362), .B2(n18761), .A(n14361), .ZN(n14363) );
  INV_X1 U17425 ( .A(n14363), .ZN(P2_U2891) );
  AOI22_X1 U17426 ( .A1(n18703), .A2(BUF1_REG_27__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U17427 ( .A1(n18701), .A2(n14364), .B1(n18756), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n14365) );
  OAI211_X1 U17428 ( .C1(n15723), .C2(n14678), .A(n14366), .B(n14365), .ZN(
        n14367) );
  AOI21_X1 U17429 ( .B1(n14368), .B2(n18761), .A(n14367), .ZN(n14369) );
  INV_X1 U17430 ( .A(n14369), .ZN(P2_U2892) );
  NAND2_X1 U17431 ( .A1(n14370), .A2(n18761), .ZN(n14377) );
  AOI22_X1 U17432 ( .A1(n18701), .A2(n18722), .B1(n18756), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U17433 ( .A1(n18703), .A2(BUF1_REG_26__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U17434 ( .A1(n14380), .A2(n14371), .ZN(n14372) );
  AND2_X1 U17435 ( .A1(n14373), .A2(n14372), .ZN(n15668) );
  NAND2_X1 U17436 ( .A1(n18757), .A2(n15668), .ZN(n14374) );
  NAND4_X1 U17437 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        P2_U2893) );
  NAND2_X1 U17438 ( .A1(n14389), .A2(n14378), .ZN(n14379) );
  NAND2_X1 U17439 ( .A1(n14380), .A2(n14379), .ZN(n15683) );
  AOI22_X1 U17440 ( .A1(n18703), .A2(BUF1_REG_25__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U17441 ( .A1(n18701), .A2(n14381), .B1(n18756), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n14382) );
  OAI211_X1 U17442 ( .C1(n15723), .C2(n15683), .A(n14383), .B(n14382), .ZN(
        n14384) );
  INV_X1 U17443 ( .A(n14384), .ZN(n14385) );
  OAI21_X1 U17444 ( .B1(n14386), .B2(n18733), .A(n14385), .ZN(P2_U2894) );
  OR2_X1 U17445 ( .A1(n14398), .A2(n14387), .ZN(n14388) );
  NAND2_X1 U17446 ( .A1(n14389), .A2(n14388), .ZN(n15692) );
  AOI22_X1 U17447 ( .A1(n18703), .A2(BUF1_REG_24__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U17448 ( .A1(n18701), .A2(n14390), .B1(n18756), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n14391) );
  OAI211_X1 U17449 ( .C1(n15723), .C2(n15692), .A(n14392), .B(n14391), .ZN(
        n14393) );
  AOI21_X1 U17450 ( .B1(n14394), .B2(n18761), .A(n14393), .ZN(n14395) );
  INV_X1 U17451 ( .A(n14395), .ZN(P2_U2895) );
  AND2_X1 U17452 ( .A1(n14744), .A2(n14396), .ZN(n14397) );
  OR2_X1 U17453 ( .A1(n14398), .A2(n14397), .ZN(n15712) );
  AOI22_X1 U17454 ( .A1(n18703), .A2(BUF1_REG_23__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U17455 ( .A1(n18701), .A2(n14399), .B1(n18756), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n14400) );
  OAI211_X1 U17456 ( .C1(n15723), .C2(n15712), .A(n14401), .B(n14400), .ZN(
        n14402) );
  AOI21_X1 U17457 ( .B1(n14403), .B2(n18761), .A(n14402), .ZN(n14404) );
  INV_X1 U17458 ( .A(n14404), .ZN(P2_U2896) );
  OR2_X1 U17459 ( .A1(n14406), .A2(n14405), .ZN(n14408) );
  NAND2_X1 U17460 ( .A1(n14408), .A2(n14407), .ZN(n18531) );
  AOI22_X1 U17461 ( .A1(n18703), .A2(BUF1_REG_21__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U17462 ( .A1(n18701), .A2(n14409), .B1(n18756), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n14410) );
  OAI211_X1 U17463 ( .C1(n15723), .C2(n18531), .A(n14411), .B(n14410), .ZN(
        n14412) );
  INV_X1 U17464 ( .A(n14412), .ZN(n14413) );
  OAI21_X1 U17465 ( .B1(n14414), .B2(n18733), .A(n14413), .ZN(P2_U2898) );
  NOR2_X1 U17466 ( .A1(n14415), .A2(n14777), .ZN(n14416) );
  OR2_X1 U17467 ( .A1(n14417), .A2(n14416), .ZN(n18538) );
  AOI22_X1 U17468 ( .A1(n18703), .A2(BUF1_REG_19__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U17469 ( .A1(n18701), .A2(n14418), .B1(n18756), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14419) );
  OAI211_X1 U17470 ( .C1(n15723), .C2(n18538), .A(n14420), .B(n14419), .ZN(
        n14421) );
  AOI21_X1 U17471 ( .B1(n14422), .B2(n18761), .A(n14421), .ZN(n14423) );
  INV_X1 U17472 ( .A(n14423), .ZN(P2_U2900) );
  OR2_X1 U17473 ( .A1(n14424), .A2(n14797), .ZN(n14425) );
  NAND2_X1 U17474 ( .A1(n14425), .A2(n14775), .ZN(n18564) );
  AOI22_X1 U17475 ( .A1(n18703), .A2(BUF1_REG_17__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U17476 ( .A1(n18701), .A2(n14426), .B1(n18756), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14427) );
  OAI211_X1 U17477 ( .C1(n15723), .C2(n18564), .A(n14428), .B(n14427), .ZN(
        n14429) );
  INV_X1 U17478 ( .A(n14429), .ZN(n14430) );
  OAI21_X1 U17479 ( .B1(n14431), .B2(n18733), .A(n14430), .ZN(P2_U2902) );
  NAND2_X1 U17480 ( .A1(n14432), .A2(n14440), .ZN(n14435) );
  NOR2_X1 U17481 ( .A1(n14433), .A2(n9684), .ZN(n14434) );
  XNOR2_X1 U17482 ( .A(n14448), .B(n14612), .ZN(n14641) );
  INV_X1 U17483 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14436) );
  NOR2_X1 U17484 ( .A1(n18662), .A2(n14436), .ZN(n14634) );
  AOI21_X1 U17485 ( .B1(n18810), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14634), .ZN(n14439) );
  NAND2_X1 U17486 ( .A1(n14437), .A2(n15824), .ZN(n14438) );
  NAND2_X1 U17487 ( .A1(n14441), .A2(n14440), .ZN(n14443) );
  XOR2_X1 U17488 ( .A(n14443), .B(n14442), .Z(n14657) );
  NAND2_X1 U17489 ( .A1(n14444), .A2(n15824), .ZN(n14445) );
  NAND2_X1 U17490 ( .A1(n18815), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14646) );
  OAI211_X1 U17491 ( .C1(n15833), .C2(n14446), .A(n14445), .B(n14646), .ZN(
        n14447) );
  AOI21_X1 U17492 ( .B1(n14645), .B2(n18819), .A(n14447), .ZN(n14450) );
  AOI21_X1 U17493 ( .B1(n14652), .B2(n14451), .A(n14448), .ZN(n14655) );
  NAND2_X1 U17494 ( .A1(n14655), .A2(n18814), .ZN(n14449) );
  OAI211_X1 U17495 ( .C1(n14657), .C2(n15817), .A(n14450), .B(n14449), .ZN(
        P2_U2985) );
  OAI21_X1 U17496 ( .B1(n14467), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14451), .ZN(n14670) );
  INV_X1 U17497 ( .A(n14452), .ZN(n14453) );
  INV_X1 U17498 ( .A(n14455), .ZN(n14457) );
  XOR2_X1 U17499 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14458), .Z(
        n14459) );
  NAND2_X1 U17500 ( .A1(n14658), .A2(n18811), .ZN(n14466) );
  NAND2_X1 U17501 ( .A1(n18815), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14662) );
  OAI21_X1 U17502 ( .B1(n15833), .B2(n14461), .A(n14662), .ZN(n14463) );
  NOR2_X1 U17503 ( .A1(n14664), .A2(n15828), .ZN(n14462) );
  AOI211_X1 U17504 ( .C1(n15824), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        n14465) );
  OAI211_X1 U17505 ( .C1(n15816), .C2(n14670), .A(n14466), .B(n14465), .ZN(
        P2_U2986) );
  OAI21_X1 U17506 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n9616), .A(
        n10122), .ZN(n14684) );
  OR2_X1 U17507 ( .A1(n14468), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14672) );
  NAND3_X1 U17508 ( .A1(n14672), .A2(n14671), .A3(n18811), .ZN(n14474) );
  NAND2_X1 U17509 ( .A1(n18815), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14676) );
  OAI21_X1 U17510 ( .B1(n15833), .B2(n14469), .A(n14676), .ZN(n14471) );
  NOR2_X1 U17511 ( .A1(n14673), .A2(n15828), .ZN(n14470) );
  AOI211_X1 U17512 ( .C1(n15824), .C2(n14472), .A(n14471), .B(n14470), .ZN(
        n14473) );
  OAI211_X1 U17513 ( .C1(n15816), .C2(n14684), .A(n14474), .B(n14473), .ZN(
        P2_U2987) );
  INV_X1 U17514 ( .A(n14475), .ZN(n14483) );
  NOR2_X1 U17515 ( .A1(n14476), .A2(n14483), .ZN(n14477) );
  XOR2_X1 U17516 ( .A(n14478), .B(n14477), .Z(n14695) );
  INV_X1 U17517 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19524) );
  NOR2_X1 U17518 ( .A1(n18662), .A2(n19524), .ZN(n14688) );
  NOR2_X1 U17519 ( .A1(n15673), .A2(n18817), .ZN(n14479) );
  AOI211_X1 U17520 ( .C1(n18810), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14688), .B(n14479), .ZN(n14480) );
  OAI21_X1 U17521 ( .B1(n15670), .B2(n15828), .A(n14480), .ZN(n14481) );
  AOI21_X1 U17522 ( .B1(n14693), .B2(n18814), .A(n14481), .ZN(n14482) );
  OAI21_X1 U17523 ( .B1(n14695), .B2(n15817), .A(n14482), .ZN(P2_U2988) );
  NOR2_X1 U17524 ( .A1(n14484), .A2(n14483), .ZN(n14486) );
  XOR2_X1 U17525 ( .A(n14486), .B(n14485), .Z(n14708) );
  NAND2_X1 U17526 ( .A1(n18815), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n14700) );
  OAI21_X1 U17527 ( .B1(n15833), .B2(n14487), .A(n14700), .ZN(n14489) );
  NOR2_X1 U17528 ( .A1(n15684), .A2(n15828), .ZN(n14488) );
  AOI211_X1 U17529 ( .C1(n15824), .C2(n15680), .A(n14489), .B(n14488), .ZN(
        n14492) );
  NAND2_X1 U17530 ( .A1(n14490), .A2(n14697), .ZN(n14704) );
  NAND3_X1 U17531 ( .A1(n14705), .A2(n18814), .A3(n14704), .ZN(n14491) );
  OAI211_X1 U17532 ( .C1(n14708), .C2(n15817), .A(n14492), .B(n14491), .ZN(
        P2_U2989) );
  XNOR2_X1 U17533 ( .A(n14493), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14494) );
  XNOR2_X1 U17534 ( .A(n14495), .B(n14494), .ZN(n14718) );
  INV_X1 U17535 ( .A(n14496), .ZN(n14498) );
  AOI21_X1 U17536 ( .B1(n14709), .B2(n14498), .A(n14497), .ZN(n14716) );
  NOR2_X1 U17537 ( .A1(n15693), .A2(n15828), .ZN(n14501) );
  AOI22_X1 U17538 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18815), .ZN(n14499) );
  OAI21_X1 U17539 ( .B1(n15697), .B2(n18817), .A(n14499), .ZN(n14500) );
  AOI211_X1 U17540 ( .C1(n14716), .C2(n18814), .A(n14501), .B(n14500), .ZN(
        n14502) );
  OAI21_X1 U17541 ( .B1(n14718), .B2(n15817), .A(n14502), .ZN(P2_U2990) );
  AOI21_X1 U17542 ( .B1(n14506), .B2(n14505), .A(n14566), .ZN(n14558) );
  INV_X1 U17543 ( .A(n14507), .ZN(n14508) );
  AOI21_X1 U17544 ( .B1(n14558), .B2(n14557), .A(n14508), .ZN(n14549) );
  INV_X1 U17545 ( .A(n14549), .ZN(n14511) );
  NAND2_X1 U17546 ( .A1(n14510), .A2(n14509), .ZN(n14548) );
  OAI21_X1 U17547 ( .B1(n14511), .B2(n14548), .A(n14510), .ZN(n14764) );
  NAND2_X1 U17548 ( .A1(n14764), .A2(n14765), .ZN(n14763) );
  INV_X1 U17549 ( .A(n14512), .ZN(n14537) );
  NOR2_X1 U17550 ( .A1(n14763), .A2(n14537), .ZN(n14524) );
  INV_X1 U17551 ( .A(n14513), .ZN(n14528) );
  OAI21_X1 U17552 ( .B1(n14524), .B2(n14514), .A(n14528), .ZN(n14518) );
  NOR2_X1 U17553 ( .A1(n14516), .A2(n14515), .ZN(n14517) );
  XNOR2_X1 U17554 ( .A(n14518), .B(n14517), .ZN(n15425) );
  INV_X1 U17555 ( .A(n14519), .ZN(n14735) );
  AOI21_X1 U17556 ( .B1(n14618), .B2(n14533), .A(n14735), .ZN(n15422) );
  INV_X1 U17557 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19517) );
  NOR2_X1 U17558 ( .A1(n19517), .A2(n18662), .ZN(n15419) );
  NOR2_X1 U17559 ( .A1(n15833), .A2(n18522), .ZN(n14520) );
  AOI211_X1 U17560 ( .C1(n18528), .C2(n15824), .A(n15419), .B(n14520), .ZN(
        n14521) );
  OAI21_X1 U17561 ( .B1(n15421), .B2(n15828), .A(n14521), .ZN(n14522) );
  AOI21_X1 U17562 ( .B1(n15422), .B2(n18814), .A(n14522), .ZN(n14523) );
  OAI21_X1 U17563 ( .B1(n15425), .B2(n15817), .A(n14523), .ZN(P2_U2993) );
  INV_X1 U17564 ( .A(n14524), .ZN(n14526) );
  NAND2_X1 U17565 ( .A1(n14526), .A2(n14525), .ZN(n14530) );
  NAND2_X1 U17566 ( .A1(n14528), .A2(n14527), .ZN(n14529) );
  XNOR2_X1 U17567 ( .A(n14530), .B(n14529), .ZN(n14762) );
  NOR2_X1 U17568 ( .A1(n18662), .A2(n19515), .ZN(n14753) );
  AOI21_X1 U17569 ( .B1(n18810), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14753), .ZN(n14531) );
  OAI21_X1 U17570 ( .B1(n14532), .B2(n18817), .A(n14531), .ZN(n14535) );
  OAI21_X1 U17571 ( .B1(n14542), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14533), .ZN(n14750) );
  NOR2_X1 U17572 ( .A1(n14750), .A2(n15816), .ZN(n14534) );
  AOI211_X1 U17573 ( .C1(n18819), .C2(n14754), .A(n14535), .B(n14534), .ZN(
        n14536) );
  OAI21_X1 U17574 ( .B1(n14762), .B2(n15817), .A(n14536), .ZN(P2_U2994) );
  NOR2_X1 U17575 ( .A1(n14538), .A2(n14537), .ZN(n14541) );
  INV_X1 U17576 ( .A(n14539), .ZN(n14767) );
  NAND2_X1 U17577 ( .A1(n14763), .A2(n14767), .ZN(n14540) );
  XOR2_X1 U17578 ( .A(n14541), .B(n14540), .Z(n15844) );
  AOI21_X1 U17579 ( .B1(n15838), .B2(n14769), .A(n14542), .ZN(n15841) );
  OAI22_X1 U17580 ( .A1(n15833), .A2(n14543), .B1(n12088), .B2(n18662), .ZN(
        n14544) );
  AOI21_X1 U17581 ( .B1(n18534), .B2(n15824), .A(n14544), .ZN(n14545) );
  OAI21_X1 U17582 ( .B1(n18539), .B2(n15828), .A(n14545), .ZN(n14546) );
  AOI21_X1 U17583 ( .B1(n15841), .B2(n18814), .A(n14546), .ZN(n14547) );
  OAI21_X1 U17584 ( .B1(n15844), .B2(n15817), .A(n14547), .ZN(P2_U2995) );
  XNOR2_X1 U17585 ( .A(n14549), .B(n14548), .ZN(n14796) );
  INV_X1 U17586 ( .A(n18565), .ZN(n14793) );
  INV_X1 U17587 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19510) );
  AOI22_X1 U17588 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n15824), .B2(n18559), .ZN(n14550) );
  OAI21_X1 U17589 ( .B1(n19510), .B2(n18662), .A(n14550), .ZN(n14555) );
  NAND2_X1 U17590 ( .A1(n14551), .A2(n14783), .ZN(n15771) );
  INV_X1 U17591 ( .A(n15858), .ZN(n14784) );
  INV_X1 U17592 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15850) );
  NOR2_X2 U17593 ( .A1(n15760), .A2(n15850), .ZN(n14785) );
  NAND2_X1 U17594 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14785), .ZN(
        n14787) );
  INV_X1 U17595 ( .A(n14771), .ZN(n14552) );
  AOI211_X1 U17596 ( .C1(n14787), .C2(n14553), .A(n15816), .B(n14552), .ZN(
        n14554) );
  AOI211_X1 U17597 ( .C1(n14793), .C2(n18819), .A(n14555), .B(n14554), .ZN(
        n14556) );
  OAI21_X1 U17598 ( .B1(n14796), .B2(n15817), .A(n14556), .ZN(P2_U2997) );
  XNOR2_X1 U17599 ( .A(n14558), .B(n14557), .ZN(n14806) );
  NOR2_X1 U17600 ( .A1(n12078), .A2(n18662), .ZN(n14561) );
  INV_X1 U17601 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14559) );
  OAI22_X1 U17602 ( .A1(n15833), .A2(n14559), .B1(n18817), .B2(n18571), .ZN(
        n14560) );
  AOI211_X1 U17603 ( .C1(n18819), .C2(n18576), .A(n14561), .B(n14560), .ZN(
        n14563) );
  OAI211_X1 U17604 ( .C1(n14785), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n18814), .B(n14787), .ZN(n14562) );
  OAI211_X1 U17605 ( .C1(n14806), .C2(n15817), .A(n14563), .B(n14562), .ZN(
        P2_U2998) );
  NAND2_X1 U17606 ( .A1(n14579), .A2(n14575), .ZN(n15755) );
  NOR2_X1 U17607 ( .A1(n15755), .A2(n15756), .ZN(n15754) );
  INV_X1 U17608 ( .A(n14564), .ZN(n15758) );
  NOR2_X1 U17609 ( .A1(n15754), .A2(n15758), .ZN(n14568) );
  NOR2_X1 U17610 ( .A1(n14566), .A2(n14565), .ZN(n14567) );
  XNOR2_X1 U17611 ( .A(n14568), .B(n14567), .ZN(n15857) );
  AND2_X1 U17612 ( .A1(n15760), .A2(n15850), .ZN(n14569) );
  OR2_X1 U17613 ( .A1(n14569), .A2(n14785), .ZN(n15853) );
  AOI22_X1 U17614 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n15824), .B2(n18581), .ZN(n14571) );
  AOI22_X1 U17615 ( .A1(n15852), .A2(n18819), .B1(P2_REIP_REG_15__SCAN_IN), 
        .B2(n18815), .ZN(n14570) );
  OAI211_X1 U17616 ( .C1(n15853), .C2(n15816), .A(n14571), .B(n14570), .ZN(
        n14572) );
  INV_X1 U17617 ( .A(n14572), .ZN(n14573) );
  OAI21_X1 U17618 ( .B1(n15857), .B2(n15817), .A(n14573), .ZN(P2_U2999) );
  INV_X1 U17619 ( .A(n14575), .ZN(n14578) );
  AND2_X1 U17620 ( .A1(n14575), .A2(n14574), .ZN(n14576) );
  OAI22_X1 U17621 ( .A1(n14579), .A2(n14578), .B1(n14577), .B2(n14576), .ZN(
        n14822) );
  INV_X1 U17622 ( .A(n15771), .ZN(n14580) );
  INV_X1 U17623 ( .A(n15859), .ZN(n14807) );
  NAND2_X1 U17624 ( .A1(n14580), .A2(n14807), .ZN(n15762) );
  INV_X1 U17625 ( .A(n15762), .ZN(n14582) );
  AOI21_X1 U17626 ( .B1(n14580), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14581) );
  NOR2_X1 U17627 ( .A1(n14582), .A2(n14581), .ZN(n14820) );
  AOI22_X1 U17628 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n15824), .B2(n18597), .ZN(n14583) );
  NAND2_X1 U17629 ( .A1(n18815), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n14813) );
  OAI211_X1 U17630 ( .C1(n15828), .C2(n14814), .A(n14583), .B(n14813), .ZN(
        n14584) );
  AOI21_X1 U17631 ( .B1(n14820), .B2(n18814), .A(n14584), .ZN(n14585) );
  OAI21_X1 U17632 ( .B1(n14822), .B2(n15817), .A(n14585), .ZN(P2_U3001) );
  XNOR2_X1 U17633 ( .A(n14586), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14587) );
  XNOR2_X1 U17634 ( .A(n14588), .B(n14587), .ZN(n15917) );
  INV_X1 U17635 ( .A(n15802), .ZN(n14593) );
  OAI21_X1 U17636 ( .B1(n14591), .B2(n14593), .A(n14590), .ZN(n14592) );
  OAI21_X1 U17637 ( .B1(n14589), .B2(n14593), .A(n14592), .ZN(n15914) );
  OAI22_X1 U17638 ( .A1(n15833), .A2(n14594), .B1(n19497), .B2(n18662), .ZN(
        n14597) );
  INV_X1 U17639 ( .A(n18637), .ZN(n14595) );
  OAI22_X1 U17640 ( .A1(n18642), .A2(n15828), .B1(n18817), .B2(n14595), .ZN(
        n14596) );
  AOI211_X1 U17641 ( .C1(n15914), .C2(n18811), .A(n14597), .B(n14596), .ZN(
        n14598) );
  OAI21_X1 U17642 ( .B1(n15816), .B2(n15917), .A(n14598), .ZN(P2_U3007) );
  XNOR2_X1 U17643 ( .A(n14599), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14869) );
  XOR2_X1 U17644 ( .A(n14601), .B(n14600), .Z(n14867) );
  INV_X1 U17645 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19495) );
  OAI22_X1 U17646 ( .A1(n19495), .A2(n18662), .B1(n18817), .B2(n18655), .ZN(
        n14603) );
  OAI22_X1 U17647 ( .A1(n15828), .A2(n18657), .B1(n15833), .B2(n10008), .ZN(
        n14602) );
  AOI211_X1 U17648 ( .C1(n14867), .C2(n18811), .A(n14603), .B(n14602), .ZN(
        n14604) );
  OAI21_X1 U17649 ( .B1(n14869), .B2(n15816), .A(n14604), .ZN(P2_U3008) );
  INV_X1 U17650 ( .A(n18836), .ZN(n14605) );
  AND2_X1 U17651 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14721) );
  NOR2_X1 U17652 ( .A1(n14757), .A2(n15838), .ZN(n14751) );
  NAND3_X1 U17653 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14616) );
  INV_X1 U17654 ( .A(n14616), .ZN(n14607) );
  NAND2_X1 U17655 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14879) );
  OAI21_X1 U17656 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14609), .A(
        n14606), .ZN(n14891) );
  AOI21_X1 U17657 ( .B1(n18854), .B2(n14879), .A(n14891), .ZN(n15891) );
  OAI21_X1 U17658 ( .B1(n14609), .B2(n14607), .A(n15891), .ZN(n14848) );
  AOI21_X1 U17659 ( .B1(n14617), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n14609), .ZN(n14608) );
  NOR2_X1 U17660 ( .A1(n14848), .A2(n14608), .ZN(n15835) );
  OAI21_X1 U17661 ( .B1(n14609), .B2(n14751), .A(n15835), .ZN(n15420) );
  AOI21_X1 U17662 ( .B1(n18854), .B2(n14618), .A(n15420), .ZN(n14738) );
  OAI21_X1 U17663 ( .B1(n14721), .B2(n14609), .A(n14738), .ZN(n14712) );
  AOI21_X1 U17664 ( .B1(n18854), .B2(n14709), .A(n14712), .ZN(n14696) );
  NAND2_X1 U17665 ( .A1(n18854), .A2(n14620), .ZN(n14610) );
  NAND2_X1 U17666 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14621) );
  OAI21_X1 U17667 ( .B1(n14652), .B2(n14621), .A(n18854), .ZN(n14611) );
  NAND2_X1 U17668 ( .A1(n14675), .A2(n14611), .ZN(n14636) );
  AOI21_X1 U17669 ( .B1(n14612), .B2(n18854), .A(n14636), .ZN(n14613) );
  NOR2_X1 U17670 ( .A1(n14613), .A2(n14622), .ZN(n14626) );
  NOR2_X1 U17671 ( .A1(n14615), .A2(n14614), .ZN(n14892) );
  NAND3_X1 U17672 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n14892), .ZN(n15898) );
  NAND2_X1 U17673 ( .A1(n14617), .A2(n14850), .ZN(n14774) );
  NOR2_X1 U17674 ( .A1(n14773), .A2(n14774), .ZN(n15839) );
  NAND3_X1 U17675 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n15839), .ZN(n15417) );
  NOR2_X1 U17676 ( .A1(n14618), .A2(n15417), .ZN(n14736) );
  AND2_X1 U17677 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14736), .ZN(
        n14619) );
  INV_X1 U17678 ( .A(n14620), .ZN(n14686) );
  NAND2_X1 U17679 ( .A1(n14698), .A2(n14686), .ZN(n14644) );
  NOR2_X1 U17680 ( .A1(n14644), .A2(n14621), .ZN(n14632) );
  NAND4_X1 U17681 ( .A1(n14632), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n14622), .ZN(n14623) );
  OAI211_X1 U17682 ( .C1(n18696), .C2(n18832), .A(n14624), .B(n14623), .ZN(
        n14625) );
  AOI211_X1 U17683 ( .C1(n14627), .C2(n18853), .A(n14626), .B(n14625), .ZN(
        n14630) );
  OAI211_X1 U17684 ( .C1(n14631), .C2(n15926), .A(n14630), .B(n14629), .ZN(
        P2_U3015) );
  INV_X1 U17685 ( .A(n14632), .ZN(n14647) );
  NOR3_X1 U17686 ( .A1(n14647), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14652), .ZN(n14633) );
  AOI211_X1 U17687 ( .C1(n14635), .C2(n18847), .A(n14634), .B(n14633), .ZN(
        n14638) );
  NAND2_X1 U17688 ( .A1(n14636), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14637) );
  OAI211_X1 U17689 ( .C1(n14639), .C2(n15894), .A(n14638), .B(n14637), .ZN(
        n14640) );
  AOI21_X1 U17690 ( .B1(n14641), .B2(n18846), .A(n14640), .ZN(n14642) );
  OAI21_X1 U17691 ( .B1(n14643), .B2(n15926), .A(n14642), .ZN(P2_U3016) );
  INV_X1 U17692 ( .A(n14644), .ZN(n14660) );
  INV_X1 U17693 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14659) );
  NAND2_X1 U17694 ( .A1(n14660), .A2(n14674), .ZN(n14677) );
  NAND2_X1 U17695 ( .A1(n14675), .A2(n14677), .ZN(n14667) );
  AOI21_X1 U17696 ( .B1(n14660), .B2(n14659), .A(n14667), .ZN(n14653) );
  NAND2_X1 U17697 ( .A1(n14645), .A2(n18853), .ZN(n14651) );
  OAI21_X1 U17698 ( .B1(n14647), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14646), .ZN(n14648) );
  AOI21_X1 U17699 ( .B1(n14649), .B2(n18847), .A(n14648), .ZN(n14650) );
  OAI211_X1 U17700 ( .C1(n14653), .C2(n14652), .A(n14651), .B(n14650), .ZN(
        n14654) );
  AOI21_X1 U17701 ( .B1(n14655), .B2(n18846), .A(n14654), .ZN(n14656) );
  OAI21_X1 U17702 ( .B1(n14657), .B2(n15926), .A(n14656), .ZN(P2_U3017) );
  NAND2_X1 U17703 ( .A1(n14658), .A2(n18844), .ZN(n14669) );
  NAND3_X1 U17704 ( .A1(n14660), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14659), .ZN(n14661) );
  OAI211_X1 U17705 ( .C1(n14663), .C2(n18832), .A(n14662), .B(n14661), .ZN(
        n14666) );
  NOR2_X1 U17706 ( .A1(n14664), .A2(n15894), .ZN(n14665) );
  AOI211_X1 U17707 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n14667), .A(
        n14666), .B(n14665), .ZN(n14668) );
  OAI211_X1 U17708 ( .C1(n14670), .C2(n18841), .A(n14669), .B(n14668), .ZN(
        P2_U3018) );
  NAND3_X1 U17709 ( .A1(n14672), .A2(n14671), .A3(n18844), .ZN(n14683) );
  INV_X1 U17710 ( .A(n14673), .ZN(n14681) );
  NOR2_X1 U17711 ( .A1(n14675), .A2(n14674), .ZN(n14680) );
  OAI211_X1 U17712 ( .C1(n18832), .C2(n14678), .A(n14677), .B(n14676), .ZN(
        n14679) );
  AOI211_X1 U17713 ( .C1(n14681), .C2(n18853), .A(n14680), .B(n14679), .ZN(
        n14682) );
  OAI211_X1 U17714 ( .C1(n14684), .C2(n18841), .A(n14683), .B(n14682), .ZN(
        P2_U3019) );
  NOR2_X1 U17715 ( .A1(n15670), .A2(n15894), .ZN(n14692) );
  INV_X1 U17716 ( .A(n14698), .ZN(n14685) );
  AOI211_X1 U17717 ( .C1(n14690), .C2(n14697), .A(n14686), .B(n14685), .ZN(
        n14687) );
  AOI211_X1 U17718 ( .C1(n18847), .C2(n15668), .A(n14688), .B(n14687), .ZN(
        n14689) );
  OAI21_X1 U17719 ( .B1(n14696), .B2(n14690), .A(n14689), .ZN(n14691) );
  AOI211_X1 U17720 ( .C1(n14693), .C2(n18846), .A(n14692), .B(n14691), .ZN(
        n14694) );
  OAI21_X1 U17721 ( .B1(n14695), .B2(n15926), .A(n14694), .ZN(P2_U3020) );
  INV_X1 U17722 ( .A(n15684), .ZN(n14703) );
  NOR2_X1 U17723 ( .A1(n14696), .A2(n14697), .ZN(n14702) );
  NAND2_X1 U17724 ( .A1(n14698), .A2(n14697), .ZN(n14699) );
  OAI211_X1 U17725 ( .C1(n18832), .C2(n15683), .A(n14700), .B(n14699), .ZN(
        n14701) );
  AOI211_X1 U17726 ( .C1(n14703), .C2(n18853), .A(n14702), .B(n14701), .ZN(
        n14707) );
  NAND3_X1 U17727 ( .A1(n14705), .A2(n18846), .A3(n14704), .ZN(n14706) );
  OAI211_X1 U17728 ( .C1(n14708), .C2(n15926), .A(n14707), .B(n14706), .ZN(
        P2_U3021) );
  NOR2_X1 U17729 ( .A1(n15693), .A2(n15894), .ZN(n14715) );
  AND3_X1 U17730 ( .A1(n14721), .A2(n14736), .A3(n14709), .ZN(n14711) );
  NOR2_X1 U17731 ( .A1(n12108), .A2(n18662), .ZN(n14710) );
  AOI211_X1 U17732 ( .C1(n14712), .C2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14711), .B(n14710), .ZN(n14713) );
  OAI21_X1 U17733 ( .B1(n18832), .B2(n15692), .A(n14713), .ZN(n14714) );
  AOI211_X1 U17734 ( .C1(n14716), .C2(n18846), .A(n14715), .B(n14714), .ZN(
        n14717) );
  OAI21_X1 U17735 ( .B1(n14718), .B2(n15926), .A(n14717), .ZN(P2_U3022) );
  XNOR2_X1 U17736 ( .A(n14720), .B(n14719), .ZN(n15736) );
  AOI21_X1 U17737 ( .B1(n14727), .B2(n14739), .A(n14721), .ZN(n14723) );
  NOR2_X1 U17738 ( .A1(n12104), .A2(n18662), .ZN(n14722) );
  AOI21_X1 U17739 ( .B1(n14736), .B2(n14723), .A(n14722), .ZN(n14726) );
  INV_X1 U17740 ( .A(n15712), .ZN(n14724) );
  NAND2_X1 U17741 ( .A1(n18847), .A2(n14724), .ZN(n14725) );
  OAI211_X1 U17742 ( .C1(n14738), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14728) );
  AOI21_X1 U17743 ( .B1(n15738), .B2(n18853), .A(n14728), .ZN(n14731) );
  NOR2_X1 U17744 ( .A1(n15741), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14729) );
  OR2_X1 U17745 ( .A1(n14496), .A2(n14729), .ZN(n15735) );
  OR2_X1 U17746 ( .A1(n15735), .A2(n18841), .ZN(n14730) );
  OAI211_X1 U17747 ( .C1(n15736), .C2(n15926), .A(n14731), .B(n14730), .ZN(
        P2_U3023) );
  NOR2_X1 U17748 ( .A1(n9708), .A2(n14732), .ZN(n14733) );
  XNOR2_X1 U17749 ( .A(n14734), .B(n14733), .ZN(n15746) );
  INV_X1 U17750 ( .A(n15746), .ZN(n14749) );
  NOR2_X1 U17751 ( .A1(n14735), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15742) );
  NOR3_X1 U17752 ( .A1(n15742), .A2(n15741), .A3(n18841), .ZN(n14747) );
  INV_X1 U17753 ( .A(n14736), .ZN(n14740) );
  NAND2_X1 U17754 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18815), .ZN(n14737) );
  OAI221_X1 U17755 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14740), 
        .C1(n14739), .C2(n14738), .A(n14737), .ZN(n14746) );
  OR2_X1 U17756 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  NAND2_X1 U17757 ( .A1(n14744), .A2(n14743), .ZN(n15714) );
  OAI22_X1 U17758 ( .A1(n15743), .A2(n15894), .B1(n18832), .B2(n15714), .ZN(
        n14745) );
  NOR3_X1 U17759 ( .A1(n14747), .A2(n14746), .A3(n14745), .ZN(n14748) );
  OAI21_X1 U17760 ( .B1(n14749), .B2(n15926), .A(n14748), .ZN(P2_U3024) );
  INV_X1 U17761 ( .A(n14750), .ZN(n14760) );
  OAI21_X1 U17762 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15839), .ZN(n14752) );
  NOR2_X1 U17763 ( .A1(n14752), .A2(n14751), .ZN(n14759) );
  AOI21_X1 U17764 ( .B1(n18847), .B2(n15721), .A(n14753), .ZN(n14756) );
  NAND2_X1 U17765 ( .A1(n14754), .A2(n18853), .ZN(n14755) );
  OAI211_X1 U17766 ( .C1(n15835), .C2(n14757), .A(n14756), .B(n14755), .ZN(
        n14758) );
  AOI211_X1 U17767 ( .C1(n14760), .C2(n18846), .A(n14759), .B(n14758), .ZN(
        n14761) );
  OAI21_X1 U17768 ( .B1(n14762), .B2(n15926), .A(n14761), .ZN(P2_U3026) );
  INV_X1 U17769 ( .A(n14763), .ZN(n14768) );
  AOI21_X1 U17770 ( .B1(n14767), .B2(n14765), .A(n14764), .ZN(n14766) );
  INV_X1 U17771 ( .A(n14769), .ZN(n14770) );
  AOI21_X1 U17772 ( .B1(n14773), .B2(n14771), .A(n14770), .ZN(n15751) );
  NAND2_X1 U17773 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n18815), .ZN(n14772) );
  OAI221_X1 U17774 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n14774), 
        .C1(n14773), .C2(n15835), .A(n14772), .ZN(n14781) );
  NAND2_X1 U17775 ( .A1(n14776), .A2(n14775), .ZN(n14779) );
  INV_X1 U17776 ( .A(n14777), .ZN(n14778) );
  NAND2_X1 U17777 ( .A1(n14779), .A2(n14778), .ZN(n18551) );
  OAI22_X1 U17778 ( .A1(n18552), .A2(n15894), .B1(n18832), .B2(n18551), .ZN(
        n14780) );
  AOI211_X1 U17779 ( .C1(n15751), .C2(n18846), .A(n14781), .B(n14780), .ZN(
        n14782) );
  OAI21_X1 U17780 ( .B1(n15750), .B2(n15926), .A(n14782), .ZN(P2_U3028) );
  NAND2_X1 U17781 ( .A1(n14783), .A2(n14850), .ZN(n15873) );
  NOR2_X1 U17782 ( .A1(n14784), .A2(n15873), .ZN(n15851) );
  AOI22_X1 U17783 ( .A1(n14785), .A2(n18846), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15851), .ZN(n14801) );
  INV_X1 U17784 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14790) );
  NOR2_X1 U17785 ( .A1(n14801), .A2(n14790), .ZN(n14791) );
  AOI21_X1 U17786 ( .B1(n14786), .B2(n18854), .A(n14848), .ZN(n15847) );
  OAI21_X1 U17787 ( .B1(n18846), .B2(n18836), .A(n14787), .ZN(n14788) );
  OAI211_X1 U17788 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n14789), .A(
        n15847), .B(n14788), .ZN(n14804) );
  OAI22_X1 U17789 ( .A1(n18832), .A2(n18564), .B1(n19510), .B2(n15908), .ZN(
        n14792) );
  AOI21_X1 U17790 ( .B1(n14793), .B2(n18853), .A(n14792), .ZN(n14794) );
  OAI211_X1 U17791 ( .C1(n14796), .C2(n15926), .A(n14795), .B(n14794), .ZN(
        P2_U3029) );
  INV_X1 U17792 ( .A(n18576), .ZN(n14800) );
  AOI21_X1 U17793 ( .B1(n14798), .B2(n15845), .A(n14797), .ZN(n18704) );
  AOI22_X1 U17794 ( .A1(n18847), .A2(n18704), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n18815), .ZN(n14799) );
  OAI21_X1 U17795 ( .B1(n14800), .B2(n15894), .A(n14799), .ZN(n14803) );
  NOR2_X1 U17796 ( .A1(n14801), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14802) );
  AOI211_X1 U17797 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n14804), .A(
        n14803), .B(n14802), .ZN(n14805) );
  OAI21_X1 U17798 ( .B1(n15926), .B2(n14806), .A(n14805), .ZN(P2_U3030) );
  AOI211_X1 U17799 ( .C1(n15770), .C2(n13315), .A(n14807), .B(n15873), .ZN(
        n14819) );
  AOI21_X1 U17800 ( .B1(n14808), .B2(n18854), .A(n14848), .ZN(n15872) );
  OR2_X1 U17801 ( .A1(n14810), .A2(n14809), .ZN(n14812) );
  NAND2_X1 U17802 ( .A1(n14812), .A2(n14811), .ZN(n18715) );
  INV_X1 U17803 ( .A(n18715), .ZN(n14816) );
  OAI21_X1 U17804 ( .B1(n15894), .B2(n14814), .A(n14813), .ZN(n14815) );
  AOI21_X1 U17805 ( .B1(n18847), .B2(n14816), .A(n14815), .ZN(n14817) );
  OAI21_X1 U17806 ( .B1(n15872), .B2(n13315), .A(n14817), .ZN(n14818) );
  AOI211_X1 U17807 ( .C1(n14820), .C2(n18846), .A(n14819), .B(n14818), .ZN(
        n14821) );
  OAI21_X1 U17808 ( .B1(n14822), .B2(n15926), .A(n14821), .ZN(P2_U3033) );
  NAND2_X1 U17809 ( .A1(n14824), .A2(n14823), .ZN(n14829) );
  INV_X1 U17810 ( .A(n14825), .ZN(n14826) );
  NOR2_X1 U17811 ( .A1(n14827), .A2(n14826), .ZN(n14828) );
  XNOR2_X1 U17812 ( .A(n14829), .B(n14828), .ZN(n15776) );
  NAND2_X1 U17813 ( .A1(n14551), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15788) );
  NOR2_X1 U17814 ( .A1(n15788), .A2(n15787), .ZN(n15790) );
  OAI21_X1 U17815 ( .B1(n15790), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15771), .ZN(n15777) );
  AOI21_X1 U17816 ( .B1(n14849), .B2(n18854), .A(n14848), .ZN(n14830) );
  INV_X1 U17817 ( .A(n14830), .ZN(n15886) );
  INV_X1 U17818 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19502) );
  NOR2_X1 U17819 ( .A1(n19502), .A2(n18662), .ZN(n14833) );
  NAND2_X1 U17820 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n14850), .ZN(
        n15883) );
  AOI221_X1 U17821 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n15787), .C2(n14831), .A(
        n15883), .ZN(n14832) );
  AOI211_X1 U17822 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15886), .A(
        n14833), .B(n14832), .ZN(n14840) );
  OR2_X1 U17823 ( .A1(n14835), .A2(n14834), .ZN(n14837) );
  NAND2_X1 U17824 ( .A1(n14837), .A2(n14836), .ZN(n18721) );
  INV_X1 U17825 ( .A(n18721), .ZN(n14838) );
  AOI22_X1 U17826 ( .A1(n18847), .A2(n14838), .B1(n18853), .B2(n18609), .ZN(
        n14839) );
  OAI211_X1 U17827 ( .C1(n15777), .C2(n18841), .A(n14840), .B(n14839), .ZN(
        n14841) );
  INV_X1 U17828 ( .A(n14841), .ZN(n14842) );
  OAI21_X1 U17829 ( .B1(n15776), .B2(n15926), .A(n14842), .ZN(P2_U3035) );
  INV_X1 U17830 ( .A(n14843), .ZN(n15781) );
  NOR2_X1 U17831 ( .A1(n14844), .A2(n15781), .ZN(n14846) );
  XOR2_X1 U17832 ( .A(n14846), .B(n14845), .Z(n15795) );
  OAI21_X1 U17833 ( .B1(n14551), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15788), .ZN(n15794) );
  INV_X1 U17834 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19499) );
  NOR2_X1 U17835 ( .A1(n19499), .A2(n18662), .ZN(n14847) );
  AOI221_X1 U17836 ( .B1(n14850), .B2(n14849), .C1(n14848), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n14847), .ZN(n14856) );
  OR2_X1 U17837 ( .A1(n14852), .A2(n14851), .ZN(n14853) );
  NAND2_X1 U17838 ( .A1(n14853), .A2(n15881), .ZN(n18726) );
  INV_X1 U17839 ( .A(n18726), .ZN(n14854) );
  AOI22_X1 U17840 ( .A1(n18847), .A2(n14854), .B1(n18853), .B2(n18632), .ZN(
        n14855) );
  OAI211_X1 U17841 ( .C1(n15794), .C2(n18841), .A(n14856), .B(n14855), .ZN(
        n14857) );
  INV_X1 U17842 ( .A(n14857), .ZN(n14858) );
  OAI21_X1 U17843 ( .B1(n15926), .B2(n15795), .A(n14858), .ZN(P2_U3037) );
  NOR2_X1 U17844 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15898), .ZN(
        n14866) );
  INV_X1 U17845 ( .A(n18657), .ZN(n14863) );
  NOR2_X1 U17846 ( .A1(n19495), .A2(n18662), .ZN(n14862) );
  XNOR2_X1 U17847 ( .A(n14860), .B(n14859), .ZN(n18731) );
  NOR2_X1 U17848 ( .A1(n18832), .A2(n18731), .ZN(n14861) );
  AOI211_X1 U17849 ( .C1(n14863), .C2(n18853), .A(n14862), .B(n14861), .ZN(
        n14864) );
  OAI21_X1 U17850 ( .B1(n15891), .B2(n15899), .A(n14864), .ZN(n14865) );
  AOI211_X1 U17851 ( .C1(n14867), .C2(n18844), .A(n14866), .B(n14865), .ZN(
        n14868) );
  OAI21_X1 U17852 ( .B1(n14869), .B2(n18841), .A(n14868), .ZN(P2_U3040) );
  CLKBUF_X1 U17853 ( .A(n14871), .Z(n14872) );
  INV_X1 U17854 ( .A(n14872), .ZN(n14873) );
  XOR2_X1 U17855 ( .A(n14870), .B(n14873), .Z(n15814) );
  AND2_X1 U17856 ( .A1(n14875), .A2(n14874), .ZN(n14877) );
  OAI22_X1 U17857 ( .A1(n14878), .A2(n13413), .B1(n14877), .B2(n14876), .ZN(
        n15815) );
  OAI211_X1 U17858 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n14892), .B(n14879), .ZN(n14885) );
  XNOR2_X1 U17859 ( .A(n14881), .B(n14880), .ZN(n18738) );
  AOI22_X1 U17860 ( .A1(n18815), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n14891), .ZN(n14882) );
  OAI21_X1 U17861 ( .B1(n18832), .B2(n18738), .A(n14882), .ZN(n14883) );
  AOI21_X1 U17862 ( .B1(n18853), .B2(n18672), .A(n14883), .ZN(n14884) );
  OAI211_X1 U17863 ( .C1(n15815), .C2(n18841), .A(n14885), .B(n14884), .ZN(
        n14886) );
  AOI21_X1 U17864 ( .B1(n15814), .B2(n18844), .A(n14886), .ZN(n14887) );
  INV_X1 U17865 ( .A(n14887), .ZN(P2_U3041) );
  XOR2_X1 U17866 ( .A(n14889), .B(n14888), .Z(n18802) );
  NAND2_X1 U17867 ( .A1(n18802), .A2(n18844), .ZN(n14901) );
  NOR2_X1 U17868 ( .A1(n19491), .A2(n18662), .ZN(n14890) );
  AOI221_X1 U17869 ( .B1(n14892), .B2(n14894), .C1(n14891), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n14890), .ZN(n14900) );
  AOI22_X1 U17870 ( .A1(n18801), .A2(n18853), .B1(n18847), .B2(n14893), .ZN(
        n14899) );
  XNOR2_X1 U17871 ( .A(n14895), .B(n14894), .ZN(n14897) );
  XNOR2_X1 U17872 ( .A(n14897), .B(n14896), .ZN(n18800) );
  NAND2_X1 U17873 ( .A1(n18800), .A2(n18846), .ZN(n14898) );
  NAND4_X1 U17874 ( .A1(n14901), .A2(n14900), .A3(n14899), .A4(n14898), .ZN(
        P2_U3042) );
  NOR3_X1 U17875 ( .A1(n14903), .A2(n14902), .A3(n14914), .ZN(n14906) );
  NOR2_X1 U17876 ( .A1(n12734), .A2(n14904), .ZN(n14905) );
  AOI211_X1 U17877 ( .C1(n10773), .C2(n14912), .A(n14906), .B(n14905), .ZN(
        n15929) );
  NOR2_X1 U17878 ( .A1(n14907), .A2(n20564), .ZN(n14925) );
  INV_X1 U17879 ( .A(n14925), .ZN(n14909) );
  OAI21_X1 U17880 ( .B1(n18669), .B2(n18850), .A(n14908), .ZN(n14926) );
  OAI222_X1 U17881 ( .A1(n19543), .A2(n15929), .B1(n14909), .B2(n14926), .C1(
        n15408), .C2(n19563), .ZN(n14910) );
  MUX2_X1 U17882 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14910), .S(
        n15175), .Z(P2_U3600) );
  INV_X1 U17883 ( .A(n14911), .ZN(n14935) );
  NAND2_X1 U17884 ( .A1(n14912), .A2(n14935), .ZN(n14930) );
  NAND2_X1 U17885 ( .A1(n14913), .A2(n15948), .ZN(n14933) );
  INV_X1 U17886 ( .A(n14914), .ZN(n14915) );
  NAND2_X1 U17887 ( .A1(n14915), .A2(n10776), .ZN(n14932) );
  NAND2_X1 U17888 ( .A1(n10578), .A2(n14932), .ZN(n14918) );
  NAND2_X1 U17889 ( .A1(n14933), .A2(n14918), .ZN(n14921) );
  OR2_X1 U17890 ( .A1(n14917), .A2(n14916), .ZN(n14929) );
  INV_X1 U17891 ( .A(n14918), .ZN(n14919) );
  NAND2_X1 U17892 ( .A1(n14929), .A2(n14919), .ZN(n14920) );
  OAI211_X1 U17893 ( .C1(n14922), .C2(n14930), .A(n14921), .B(n14920), .ZN(
        n14923) );
  AOI21_X1 U17894 ( .B1(n18830), .B2(n14940), .A(n14923), .ZN(n15933) );
  OAI22_X1 U17895 ( .A1(n19555), .A2(n15408), .B1(n15933), .B2(n19543), .ZN(
        n14924) );
  AOI21_X1 U17896 ( .B1(n14926), .B2(n14925), .A(n14924), .ZN(n14927) );
  MUX2_X1 U17897 ( .A(n10776), .B(n14927), .S(n15175), .Z(n14928) );
  INV_X1 U17898 ( .A(n14928), .ZN(P2_U3599) );
  INV_X1 U17899 ( .A(n14929), .ZN(n14931) );
  OAI211_X1 U17900 ( .C1(n14931), .C2(n10392), .A(n14930), .B(n14932), .ZN(
        n14938) );
  NAND2_X1 U17901 ( .A1(n14933), .A2(n14932), .ZN(n14934) );
  OAI211_X1 U17902 ( .C1(n14936), .C2(n14935), .A(n14934), .B(n10578), .ZN(
        n14937) );
  MUX2_X1 U17903 ( .A(n14938), .B(n14937), .S(n15934), .Z(n14939) );
  AOI21_X1 U17904 ( .B1(n12728), .B2(n14940), .A(n14939), .ZN(n15939) );
  OAI22_X1 U17905 ( .A1(n19160), .A2(n15408), .B1(n15939), .B2(n19543), .ZN(
        n14941) );
  MUX2_X1 U17906 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14941), .S(
        n15175), .Z(P2_U3596) );
  AOI22_X1 U17907 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14955) );
  INV_X2 U17908 ( .A(n9585), .ZN(n16764) );
  AOI22_X1 U17909 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14954) );
  NOR2_X2 U17910 ( .A1(n18277), .A2(n14943), .ZN(n14991) );
  CLKBUF_X3 U17911 ( .A(n14991), .Z(n16762) );
  AOI22_X1 U17912 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14942) );
  OAI21_X1 U17913 ( .B1(n9584), .B2(n20603), .A(n14942), .ZN(n14952) );
  AOI22_X1 U17914 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U17915 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14949) );
  INV_X2 U17916 ( .A(n15256), .ZN(n15273) );
  INV_X2 U17917 ( .A(n15273), .ZN(n16760) );
  AOI22_X1 U17918 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U17919 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9587), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14947) );
  NAND4_X1 U17920 ( .A1(n14950), .A2(n14949), .A3(n14948), .A4(n14947), .ZN(
        n14951) );
  NAND2_X1 U17921 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18326), .ZN(n18315) );
  AOI22_X1 U17922 ( .A1(n16802), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U17923 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14959) );
  AOI22_X1 U17924 ( .A1(n16778), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14958) );
  INV_X2 U17925 ( .A(n9584), .ZN(n16780) );
  AOI22_X1 U17926 ( .A1(n16780), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14957) );
  NAND4_X1 U17927 ( .A1(n14960), .A2(n14959), .A3(n14958), .A4(n14957), .ZN(
        n14966) );
  AOI22_X1 U17928 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16804), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U17929 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16619), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U17930 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9589), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14962) );
  AOI22_X1 U17931 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16779), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14961) );
  NAND4_X1 U17932 ( .A1(n14964), .A2(n14963), .A3(n14962), .A4(n14961), .ZN(
        n14965) );
  AOI22_X1 U17933 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14970) );
  AOI22_X1 U17934 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14969) );
  AOI22_X1 U17935 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14968) );
  AOI22_X1 U17936 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14967) );
  NAND4_X1 U17937 ( .A1(n14970), .A2(n14969), .A3(n14968), .A4(n14967), .ZN(
        n14976) );
  AOI22_X1 U17938 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14974) );
  AOI22_X1 U17939 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14973) );
  AOI22_X1 U17940 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9589), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U17941 ( .A1(n16786), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14971) );
  NAND4_X1 U17942 ( .A1(n14974), .A2(n14973), .A3(n14972), .A4(n14971), .ZN(
        n14975) );
  INV_X1 U17943 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17823) );
  INV_X1 U17944 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17818) );
  OAI22_X1 U17945 ( .A1(n18443), .A2(n18091), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15156) );
  OAI22_X1 U17946 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17823), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14979), .ZN(n14986) );
  NOR2_X1 U17947 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17823), .ZN(
        n14980) );
  NAND2_X1 U17948 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14979), .ZN(
        n14985) );
  AOI22_X1 U17949 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14986), .B1(
        n14980), .B2(n14985), .ZN(n14981) );
  AOI21_X1 U17950 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18450), .A(
        n15155), .ZN(n15182) );
  NAND3_X1 U17951 ( .A1(n14981), .A2(n15182), .A3(n15156), .ZN(n14989) );
  OAI21_X1 U17952 ( .B1(n14984), .B2(n14983), .A(n14981), .ZN(n14982) );
  INV_X1 U17953 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15170) );
  AND2_X1 U17954 ( .A1(n14985), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14987) );
  OAI22_X1 U17955 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15170), .B1(
        n14987), .B2(n14986), .ZN(n15157) );
  NOR2_X1 U17956 ( .A1(n15181), .A2(n15157), .ZN(n14988) );
  AOI22_X1 U17957 ( .A1(n16786), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15000) );
  AOI22_X1 U17958 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14999) );
  AOI22_X1 U17959 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14990) );
  OAI21_X1 U17960 ( .B1(n9647), .B2(n20605), .A(n14990), .ZN(n14997) );
  AOI22_X1 U17961 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U17962 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14994) );
  AOI22_X1 U17963 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U17964 ( .A1(n16780), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14992) );
  NAND4_X1 U17965 ( .A1(n14995), .A2(n14994), .A3(n14993), .A4(n14992), .ZN(
        n14996) );
  AOI211_X1 U17966 ( .C1(n16785), .C2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n14997), .B(n14996), .ZN(n14998) );
  NAND3_X1 U17967 ( .A1(n15000), .A2(n14999), .A3(n14998), .ZN(n15142) );
  AOI22_X1 U17968 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15010) );
  AOI22_X1 U17969 ( .A1(n16802), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U17970 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15001) );
  OAI21_X1 U17971 ( .B1(n15188), .B2(n20519), .A(n15001), .ZN(n15007) );
  AOI22_X1 U17972 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16786), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U17973 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9586), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15004) );
  AOI22_X1 U17974 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U17975 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15002) );
  NAND4_X1 U17976 ( .A1(n15005), .A2(n15004), .A3(n15003), .A4(n15002), .ZN(
        n15006) );
  AOI211_X1 U17977 ( .C1(n9590), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n15007), .B(n15006), .ZN(n15008) );
  NAND3_X1 U17978 ( .A1(n15010), .A2(n15009), .A3(n15008), .ZN(n16857) );
  NAND2_X1 U17979 ( .A1(n17848), .A2(n17857), .ZN(n15138) );
  AOI22_X1 U17980 ( .A1(n16778), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U17981 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15019) );
  INV_X1 U17982 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U17983 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15011) );
  OAI21_X1 U17984 ( .B1(n15188), .B2(n16829), .A(n15011), .ZN(n15017) );
  AOI22_X1 U17985 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15015) );
  AOI22_X1 U17986 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15014) );
  AOI22_X1 U17987 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U17988 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15012) );
  NAND4_X1 U17989 ( .A1(n15015), .A2(n15014), .A3(n15013), .A4(n15012), .ZN(
        n15016) );
  AOI211_X1 U17990 ( .C1(n16804), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15017), .B(n15016), .ZN(n15018) );
  NAND3_X1 U17991 ( .A1(n15020), .A2(n15019), .A3(n15018), .ZN(n15176) );
  AOI22_X1 U17992 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15030) );
  AOI22_X1 U17993 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15029) );
  AOI22_X1 U17994 ( .A1(n16780), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15021) );
  OAI21_X1 U17995 ( .B1(n15188), .B2(n16843), .A(n15021), .ZN(n15027) );
  AOI22_X1 U17996 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15025) );
  AOI22_X1 U17997 ( .A1(n16786), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U17998 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15023) );
  AOI22_X1 U17999 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15022) );
  NAND4_X1 U18000 ( .A1(n15025), .A2(n15024), .A3(n15023), .A4(n15022), .ZN(
        n15026) );
  AOI211_X1 U18001 ( .C1(n9591), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15027), .B(n15026), .ZN(n15028) );
  AOI22_X1 U18002 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16619), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15040) );
  AOI22_X1 U18003 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9587), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U18004 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15031) );
  OAI21_X1 U18005 ( .B1(n16612), .B2(n20624), .A(n15031), .ZN(n15037) );
  AOI22_X1 U18006 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15035) );
  AOI22_X1 U18007 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15034) );
  AOI22_X1 U18008 ( .A1(n16786), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U18009 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9592), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15032) );
  NAND4_X1 U18010 ( .A1(n15035), .A2(n15034), .A3(n15033), .A4(n15032), .ZN(
        n15036) );
  AOI211_X1 U18011 ( .C1(n16763), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n15037), .B(n15036), .ZN(n15038) );
  NAND3_X1 U18012 ( .A1(n15040), .A2(n15039), .A3(n15038), .ZN(n15148) );
  NAND2_X1 U18013 ( .A1(n15135), .A2(n15202), .ZN(n15162) );
  NOR2_X1 U18014 ( .A1(n17848), .A2(n16857), .ZN(n18280) );
  NAND3_X1 U18015 ( .A1(n17848), .A2(n17864), .A3(n15153), .ZN(n15041) );
  OAI21_X2 U18016 ( .B1(n18265), .B2(n15200), .A(n15041), .ZN(n15410) );
  NAND2_X1 U18017 ( .A1(n17864), .A2(n16841), .ZN(n16852) );
  INV_X1 U18018 ( .A(n16852), .ZN(n16845) );
  NAND2_X1 U18019 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16583) );
  INV_X1 U18020 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16550) );
  INV_X1 U18021 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16549) );
  INV_X1 U18022 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16637) );
  INV_X1 U18023 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16653) );
  INV_X1 U18024 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16321) );
  INV_X1 U18025 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16732) );
  INV_X1 U18026 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16777) );
  INV_X1 U18027 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16438) );
  INV_X1 U18028 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16820) );
  INV_X1 U18029 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16520) );
  NAND2_X1 U18030 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16523) );
  NOR2_X1 U18031 ( .A1(n16520), .A2(n16523), .ZN(n16838) );
  NAND2_X1 U18032 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16838), .ZN(n16830) );
  NOR2_X1 U18033 ( .A1(n16487), .A2(n16830), .ZN(n16818) );
  INV_X1 U18034 ( .A(n16795), .ZN(n16817) );
  NOR2_X2 U18035 ( .A1(n16438), .A2(n16817), .ZN(n16816) );
  NAND4_X1 U18036 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(P3_EBX_REG_15__SCAN_IN), .A4(P3_EBX_REG_14__SCAN_IN), .ZN(n15042)
         );
  NOR3_X2 U18037 ( .A1(n16321), .A2(n16705), .A3(n15042), .ZN(n16680) );
  NAND2_X1 U18038 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16680), .ZN(n16666) );
  NOR2_X2 U18039 ( .A1(n16653), .A2(n16666), .ZN(n16636) );
  NAND2_X1 U18040 ( .A1(n17864), .A2(n16636), .ZN(n16641) );
  NAND2_X1 U18041 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16600), .ZN(n16592) );
  INV_X1 U18042 ( .A(n16592), .ZN(n16597) );
  NOR2_X1 U18043 ( .A1(n16850), .A2(n16597), .ZN(n16590) );
  AOI21_X1 U18044 ( .B1(n16845), .B2(n16583), .A(n16590), .ZN(n16587) );
  INV_X1 U18045 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16220) );
  NOR2_X1 U18046 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16592), .ZN(n15115) );
  AOI22_X1 U18047 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15046) );
  AOI22_X1 U18048 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16786), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15045) );
  AOI22_X1 U18049 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15044) );
  AOI22_X1 U18050 ( .A1(n16780), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15043) );
  NAND4_X1 U18051 ( .A1(n15046), .A2(n15045), .A3(n15044), .A4(n15043), .ZN(
        n15052) );
  AOI22_X1 U18052 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15050) );
  AOI22_X1 U18053 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15049) );
  AOI22_X1 U18054 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15048) );
  AOI22_X1 U18055 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16779), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15047) );
  NAND4_X1 U18056 ( .A1(n15050), .A2(n15049), .A3(n15048), .A4(n15047), .ZN(
        n15051) );
  NOR2_X1 U18057 ( .A1(n15052), .A2(n15051), .ZN(n16589) );
  AOI22_X1 U18058 ( .A1(n16778), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U18059 ( .A1(n16802), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U18060 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15054) );
  AOI22_X1 U18061 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15053) );
  NAND4_X1 U18062 ( .A1(n15056), .A2(n15055), .A3(n15054), .A4(n15053), .ZN(
        n15062) );
  AOI22_X1 U18063 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15060) );
  AOI22_X1 U18064 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U18065 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U18066 ( .A1(n16786), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15057) );
  NAND4_X1 U18067 ( .A1(n15060), .A2(n15059), .A3(n15058), .A4(n15057), .ZN(
        n15061) );
  NOR2_X1 U18068 ( .A1(n15062), .A2(n15061), .ZN(n16598) );
  AOI22_X1 U18069 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U18070 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U18071 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15064) );
  AOI22_X1 U18072 ( .A1(n16780), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15063) );
  NAND4_X1 U18073 ( .A1(n15066), .A2(n15065), .A3(n15064), .A4(n15063), .ZN(
        n15073) );
  AOI22_X1 U18074 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15071) );
  AOI22_X1 U18075 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U18076 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U18077 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15068) );
  NAND4_X1 U18078 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        n15072) );
  NOR2_X1 U18079 ( .A1(n15073), .A2(n15072), .ZN(n16607) );
  AOI22_X1 U18080 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15077) );
  AOI22_X1 U18081 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U18082 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U18083 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15074) );
  NAND4_X1 U18084 ( .A1(n15077), .A2(n15076), .A3(n15075), .A4(n15074), .ZN(
        n15083) );
  AOI22_X1 U18085 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15081) );
  AOI22_X1 U18086 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U18087 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15079) );
  AOI22_X1 U18088 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15078) );
  NAND4_X1 U18089 ( .A1(n15081), .A2(n15080), .A3(n15079), .A4(n15078), .ZN(
        n15082) );
  NOR2_X1 U18090 ( .A1(n15083), .A2(n15082), .ZN(n16606) );
  NOR2_X1 U18091 ( .A1(n16607), .A2(n16606), .ZN(n16603) );
  AOI22_X1 U18092 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16763), .B1(
        n16779), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15093) );
  AOI22_X1 U18093 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n16802), .ZN(n15092) );
  INV_X1 U18094 ( .A(n15273), .ZN(n16796) );
  AOI22_X1 U18095 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n16796), .ZN(n15084) );
  OAI21_X1 U18096 ( .B1(n20625), .B2(n9585), .A(n15084), .ZN(n15090) );
  AOI22_X1 U18097 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9589), .ZN(n15088) );
  AOI22_X1 U18098 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9586), .B1(n9590), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15087) );
  AOI22_X1 U18099 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n16778), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15086) );
  AOI22_X1 U18100 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15085) );
  NAND4_X1 U18101 ( .A1(n15088), .A2(n15087), .A3(n15086), .A4(n15085), .ZN(
        n15089) );
  AOI211_X1 U18102 ( .C1(n16804), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n15090), .B(n15089), .ZN(n15091) );
  NAND3_X1 U18103 ( .A1(n15093), .A2(n15092), .A3(n15091), .ZN(n16602) );
  NAND2_X1 U18104 ( .A1(n16603), .A2(n16602), .ZN(n16601) );
  NOR2_X1 U18105 ( .A1(n16598), .A2(n16601), .ZN(n16595) );
  AOI22_X1 U18106 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15104) );
  AOI22_X1 U18107 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U18108 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15094) );
  OAI21_X1 U18109 ( .B1(n9646), .B2(n20624), .A(n15094), .ZN(n15101) );
  AOI22_X1 U18110 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U18111 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15098) );
  AOI22_X1 U18112 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U18113 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15096) );
  NAND4_X1 U18114 ( .A1(n15099), .A2(n15098), .A3(n15097), .A4(n15096), .ZN(
        n15100) );
  AOI211_X1 U18115 ( .C1(n9591), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n15101), .B(n15100), .ZN(n15102) );
  NAND3_X1 U18116 ( .A1(n15104), .A2(n15103), .A3(n15102), .ZN(n16594) );
  NAND2_X1 U18117 ( .A1(n16595), .A2(n16594), .ZN(n16593) );
  NOR2_X1 U18118 ( .A1(n16589), .A2(n16593), .ZN(n16588) );
  INV_X1 U18119 ( .A(n16588), .ZN(n16580) );
  AOI22_X1 U18120 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15108) );
  AOI22_X1 U18121 ( .A1(n16796), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15107) );
  AOI22_X1 U18122 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15106) );
  AOI22_X1 U18123 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15105) );
  NAND4_X1 U18124 ( .A1(n15108), .A2(n15107), .A3(n15106), .A4(n15105), .ZN(
        n15114) );
  AOI22_X1 U18125 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16786), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U18126 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15111) );
  AOI22_X1 U18127 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U18128 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15109) );
  NAND4_X1 U18129 ( .A1(n15112), .A2(n15111), .A3(n15110), .A4(n15109), .ZN(
        n15113) );
  NOR2_X1 U18130 ( .A1(n15114), .A2(n15113), .ZN(n16579) );
  XOR2_X1 U18131 ( .A(n16580), .B(n16579), .Z(n16870) );
  AOI22_X1 U18132 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n15115), .B1(n16850), 
        .B2(n16870), .ZN(n15116) );
  OAI21_X1 U18133 ( .B1(n16587), .B2(n16220), .A(n15116), .ZN(P3_U2675) );
  INV_X1 U18134 ( .A(n16705), .ZN(n15128) );
  AOI22_X1 U18135 ( .A1(n17864), .A2(n16746), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n16847), .ZN(n15127) );
  AOI22_X1 U18136 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U18137 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U18138 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15118) );
  AOI22_X1 U18139 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15117) );
  NAND4_X1 U18140 ( .A1(n15120), .A2(n15119), .A3(n15118), .A4(n15117), .ZN(
        n15126) );
  AOI22_X1 U18141 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U18142 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U18143 ( .A1(n15236), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15122) );
  AOI22_X1 U18144 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15121) );
  NAND4_X1 U18145 ( .A1(n15124), .A2(n15123), .A3(n15122), .A4(n15121), .ZN(
        n15125) );
  NOR2_X1 U18146 ( .A1(n15126), .A2(n15125), .ZN(n16948) );
  OAI22_X1 U18147 ( .A1(n15128), .A2(n15127), .B1(n16948), .B2(n16834), .ZN(
        P3_U2690) );
  INV_X1 U18148 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17826) );
  NAND2_X1 U18149 ( .A1(n17826), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17868) );
  INV_X1 U18150 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18419) );
  NOR2_X1 U18151 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18478) );
  AOI21_X1 U18152 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18478), .ZN(n18331) );
  NAND2_X1 U18153 ( .A1(n18475), .A2(n17830), .ZN(n18018) );
  INV_X1 U18154 ( .A(n18018), .ZN(n18171) );
  OAI21_X1 U18155 ( .B1(n18299), .B2(n18425), .A(n15170), .ZN(n15168) );
  NOR2_X1 U18156 ( .A1(n16778), .A2(n15168), .ZN(n17814) );
  INV_X1 U18157 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16153) );
  NAND3_X1 U18158 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n18418)
         );
  AOI21_X1 U18159 ( .B1(n17814), .B2(n16153), .A(n18418), .ZN(n15129) );
  NOR2_X1 U18160 ( .A1(n18171), .A2(n15129), .ZN(n17817) );
  INV_X1 U18161 ( .A(n17817), .ZN(n17822) );
  NAND2_X1 U18162 ( .A1(n17868), .A2(n17822), .ZN(n15132) );
  INV_X1 U18163 ( .A(n15132), .ZN(n15131) );
  INV_X1 U18164 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18485) );
  NAND3_X1 U18165 ( .A1(n18485), .A2(n18419), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18168) );
  INV_X1 U18166 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18429) );
  NAND2_X1 U18167 ( .A1(n18429), .A2(n18419), .ZN(n16542) );
  NAND2_X1 U18168 ( .A1(n18485), .A2(n18419), .ZN(n16147) );
  NAND2_X1 U18169 ( .A1(n16542), .A2(n16147), .ZN(n17815) );
  INV_X1 U18170 ( .A(n17815), .ZN(n18469) );
  INV_X1 U18171 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16170) );
  NOR2_X1 U18172 ( .A1(n18429), .A2(n16170), .ZN(n17318) );
  OAI22_X1 U18173 ( .A1(n18469), .A2(n17318), .B1(n17826), .B2(n18419), .ZN(
        n15134) );
  NAND3_X1 U18174 ( .A1(n18091), .A2(n17822), .A3(n15134), .ZN(n15130) );
  OAI221_X1 U18175 ( .B1(n18091), .B2(n15131), .C1(n18091), .C2(n18168), .A(
        n15130), .ZN(P3_U2864) );
  NAND2_X1 U18176 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18044) );
  NOR2_X1 U18177 ( .A1(n18469), .A2(n17318), .ZN(n15133) );
  AOI221_X1 U18178 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18044), .C1(n15133), 
        .C2(n18044), .A(n15132), .ZN(n17821) );
  INV_X1 U18179 ( .A(n18168), .ZN(n18117) );
  OAI221_X1 U18180 ( .B1(n18117), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18117), .C2(n15134), .A(n17822), .ZN(n17819) );
  AOI22_X1 U18181 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17821), .B1(
        n17819), .B2(n17818), .ZN(P3_U2865) );
  NOR2_X1 U18182 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18419), .ZN(n17829) );
  NOR2_X1 U18183 ( .A1(n15200), .A2(n18265), .ZN(n15165) );
  NAND2_X1 U18184 ( .A1(n15176), .A2(n16857), .ZN(n15141) );
  INV_X1 U18185 ( .A(n15141), .ZN(n15143) );
  INV_X1 U18186 ( .A(n15135), .ZN(n15147) );
  NAND2_X1 U18187 ( .A1(n15176), .A2(n17857), .ZN(n18269) );
  INV_X1 U18188 ( .A(n18269), .ZN(n15136) );
  NOR2_X1 U18189 ( .A1(n17864), .A2(n15136), .ZN(n15413) );
  NAND2_X1 U18190 ( .A1(n17834), .A2(n17001), .ZN(n15198) );
  NOR2_X1 U18191 ( .A1(n15413), .A2(n15198), .ZN(n15161) );
  INV_X1 U18192 ( .A(n15177), .ZN(n17838) );
  NAND2_X1 U18193 ( .A1(n17831), .A2(n18472), .ZN(n15199) );
  NAND2_X1 U18194 ( .A1(n17838), .A2(n15199), .ZN(n15140) );
  AOI21_X1 U18195 ( .B1(n17838), .B2(n17831), .A(n15136), .ZN(n15137) );
  AOI21_X1 U18196 ( .B1(n15138), .B2(n15141), .A(n15137), .ZN(n15139) );
  AOI21_X1 U18197 ( .B1(n15141), .B2(n15140), .A(n15139), .ZN(n15145) );
  OAI21_X1 U18198 ( .B1(n17864), .B2(n15143), .A(n15142), .ZN(n15144) );
  OAI211_X1 U18199 ( .C1(n15146), .C2(n15148), .A(n15145), .B(n15144), .ZN(
        n15160) );
  NAND2_X1 U18200 ( .A1(n15150), .A2(n15206), .ZN(n15201) );
  INV_X1 U18201 ( .A(n15201), .ZN(n15154) );
  NOR2_X1 U18202 ( .A1(n18472), .A2(n17001), .ZN(n15411) );
  INV_X1 U18203 ( .A(n15159), .ZN(n15151) );
  XOR2_X1 U18204 ( .A(n15156), .B(n15155), .Z(n15158) );
  NAND2_X1 U18205 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18466) );
  NAND2_X1 U18206 ( .A1(n18259), .A2(n18466), .ZN(n15163) );
  NOR2_X1 U18207 ( .A1(n18472), .A2(n17063), .ZN(n18317) );
  INV_X2 U18208 ( .A(n18483), .ZN(n18482) );
  NOR2_X1 U18209 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18336) );
  NOR3_X1 U18210 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18355), .A3(n18336), 
        .ZN(n18471) );
  OAI21_X1 U18211 ( .B1(n15159), .B2(n18317), .A(n18471), .ZN(n17000) );
  AOI211_X1 U18212 ( .C1(n16151), .C2(n15162), .A(n15161), .B(n15160), .ZN(
        n15183) );
  OAI21_X1 U18213 ( .B1(n15163), .B2(n17000), .A(n15183), .ZN(n15164) );
  NOR3_X1 U18214 ( .A1(n15165), .A2(n15412), .A3(n15164), .ZN(n18304) );
  OAI22_X1 U18215 ( .A1(n18304), .A2(n18315), .B1(n16153), .B2(n18418), .ZN(
        n15166) );
  INV_X1 U18216 ( .A(n18451), .ZN(n18448) );
  INV_X1 U18217 ( .A(n16542), .ZN(n18486) );
  INV_X1 U18218 ( .A(n15167), .ZN(n18276) );
  AND2_X1 U18219 ( .A1(n15168), .A2(n18276), .ZN(n18267) );
  NAND3_X1 U18220 ( .A1(n18448), .A2(n18486), .A3(n18267), .ZN(n15169) );
  OAI21_X1 U18221 ( .B1(n18448), .B2(n15170), .A(n15169), .ZN(P3_U3284) );
  AND4_X1 U18222 ( .A1(n15171), .A2(n13275), .A3(n18495), .A4(n15940), .ZN(
        n15172) );
  NAND2_X1 U18223 ( .A1(n15175), .A2(n15172), .ZN(n15173) );
  OAI21_X1 U18224 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(P2_U3595) );
  NAND2_X1 U18225 ( .A1(n17838), .A2(n15176), .ZN(n15180) );
  INV_X1 U18226 ( .A(n18259), .ZN(n16149) );
  INV_X1 U18227 ( .A(n18466), .ZN(n18473) );
  NOR2_X1 U18228 ( .A1(n17834), .A2(n15177), .ZN(n15207) );
  AOI211_X1 U18229 ( .C1(n17834), .C2(n15177), .A(n15207), .B(n18471), .ZN(
        n15178) );
  NOR2_X1 U18230 ( .A1(n18473), .A2(n15178), .ZN(n16150) );
  NAND2_X1 U18231 ( .A1(n15180), .A2(n16150), .ZN(n15179) );
  OAI22_X1 U18232 ( .A1(n15180), .A2(n18265), .B1(n16149), .B2(n15179), .ZN(
        n15185) );
  AOI21_X1 U18233 ( .B1(n15182), .B2(n15181), .A(n16149), .ZN(n18262) );
  NAND2_X1 U18234 ( .A1(n15207), .A2(n18262), .ZN(n15974) );
  OAI21_X1 U18235 ( .B1(n17857), .B2(n15974), .A(n15183), .ZN(n15184) );
  AOI22_X1 U18236 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15197) );
  AOI22_X1 U18237 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9586), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15196) );
  AOI22_X1 U18238 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15187) );
  OAI21_X1 U18239 ( .B1(n16612), .B2(n20603), .A(n15187), .ZN(n15194) );
  AOI22_X1 U18240 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15192) );
  AOI22_X1 U18241 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U18242 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U18243 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15189) );
  NAND4_X1 U18244 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15193) );
  AOI211_X1 U18245 ( .C1(n16619), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n15194), .B(n15193), .ZN(n15195) );
  NAND2_X1 U18246 ( .A1(n15199), .A2(n15198), .ZN(n18487) );
  INV_X1 U18247 ( .A(n15202), .ZN(n15204) );
  INV_X1 U18248 ( .A(n16169), .ZN(n15203) );
  NAND3_X1 U18249 ( .A1(n15204), .A2(n18472), .A3(n15203), .ZN(n15205) );
  NAND2_X1 U18250 ( .A1(n15206), .A2(n15205), .ZN(n18278) );
  NAND2_X1 U18251 ( .A1(n17722), .A2(n15207), .ZN(n18261) );
  INV_X1 U18252 ( .A(n18261), .ZN(n17784) );
  INV_X1 U18253 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17624) );
  INV_X1 U18254 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17607) );
  NOR2_X1 U18255 ( .A1(n17624), .A2(n17607), .ZN(n17599) );
  NAND2_X1 U18256 ( .A1(n17599), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17553) );
  INV_X1 U18257 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17249) );
  INV_X1 U18258 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17225) );
  NOR2_X1 U18259 ( .A1(n17249), .A2(n17225), .ZN(n17573) );
  NAND2_X1 U18260 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17573), .ZN(
        n17557) );
  NOR2_X1 U18261 ( .A1(n17553), .A2(n17557), .ZN(n17555) );
  INV_X1 U18262 ( .A(n17555), .ZN(n17507) );
  INV_X1 U18263 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17531) );
  INV_X1 U18264 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15208) );
  NOR2_X1 U18265 ( .A1(n17531), .A2(n15208), .ZN(n17496) );
  INV_X1 U18266 ( .A(n17496), .ZN(n15344) );
  INV_X1 U18267 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17537) );
  INV_X1 U18268 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17177) );
  NOR2_X1 U18269 ( .A1(n17537), .A2(n17177), .ZN(n17516) );
  NAND2_X1 U18270 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17516), .ZN(
        n17506) );
  NOR3_X1 U18271 ( .A1(n17507), .A2(n15344), .A3(n17506), .ZN(n16035) );
  INV_X1 U18272 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17616) );
  NAND2_X1 U18273 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17662) );
  INV_X1 U18274 ( .A(n17662), .ZN(n17694) );
  NAND2_X1 U18275 ( .A1(n17694), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17676) );
  NAND2_X1 U18276 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17293) );
  NOR2_X1 U18277 ( .A1(n17676), .A2(n17293), .ZN(n17298) );
  NAND2_X1 U18278 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17298), .ZN(
        n17615) );
  NOR2_X1 U18279 ( .A1(n17616), .A2(n17615), .ZN(n17594) );
  INV_X1 U18280 ( .A(n17594), .ZN(n17494) );
  INV_X1 U18281 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17737) );
  INV_X1 U18282 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17747) );
  INV_X1 U18283 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17733) );
  NOR3_X1 U18284 ( .A1(n17737), .A2(n17747), .A3(n17733), .ZN(n15210) );
  INV_X1 U18285 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18447) );
  INV_X1 U18286 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18430) );
  INV_X1 U18287 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20606) );
  OAI21_X1 U18288 ( .B1(n18447), .B2(n18430), .A(n20606), .ZN(n17779) );
  INV_X1 U18289 ( .A(n17779), .ZN(n15209) );
  NAND3_X1 U18290 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17592) );
  NOR2_X1 U18291 ( .A1(n15209), .A2(n17592), .ZN(n17718) );
  NAND2_X1 U18292 ( .A1(n15210), .A2(n17718), .ZN(n17614) );
  NOR2_X1 U18293 ( .A1(n17494), .A2(n17614), .ZN(n17595) );
  OAI21_X1 U18294 ( .B1(n18447), .B2(n18270), .A(n17806), .ZN(n17786) );
  NOR2_X1 U18295 ( .A1(n20606), .A2(n18430), .ZN(n17591) );
  INV_X1 U18296 ( .A(n17591), .ZN(n17759) );
  NOR2_X1 U18297 ( .A1(n17759), .A2(n17592), .ZN(n17719) );
  NAND2_X1 U18298 ( .A1(n17719), .A2(n15210), .ZN(n17661) );
  NOR2_X1 U18299 ( .A1(n17494), .A2(n17661), .ZN(n17596) );
  AOI22_X1 U18300 ( .A1(n18266), .A2(n17595), .B1(n17786), .B2(n17596), .ZN(
        n15211) );
  INV_X1 U18301 ( .A(n15211), .ZN(n16034) );
  NAND2_X1 U18302 ( .A1(n16035), .A2(n16034), .ZN(n16026) );
  INV_X1 U18303 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20633) );
  NOR2_X1 U18304 ( .A1(n20633), .A2(n17507), .ZN(n17544) );
  NAND2_X1 U18305 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17544), .ZN(
        n17173) );
  AOI22_X1 U18306 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15221) );
  AOI22_X1 U18307 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15220) );
  AOI22_X1 U18308 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15212) );
  OAI21_X1 U18309 ( .B1(n15273), .B2(n20519), .A(n15212), .ZN(n15218) );
  AOI22_X1 U18310 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16779), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U18311 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15215) );
  AOI22_X1 U18312 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15214) );
  AOI22_X1 U18313 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15213) );
  NAND4_X1 U18314 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15217) );
  AOI211_X1 U18315 ( .C1(n9592), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n15218), .B(n15217), .ZN(n15219) );
  NAND3_X1 U18316 ( .A1(n15221), .A2(n15220), .A3(n15219), .ZN(n15299) );
  AOI22_X1 U18317 ( .A1(n16796), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15225) );
  AOI22_X1 U18318 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15224) );
  AOI22_X1 U18319 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15223) );
  AOI22_X1 U18320 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15222) );
  NAND4_X1 U18321 ( .A1(n15225), .A2(n15224), .A3(n15223), .A4(n15222), .ZN(
        n15231) );
  AOI22_X1 U18322 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15229) );
  AOI22_X1 U18323 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U18324 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U18325 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15226) );
  NAND4_X1 U18326 ( .A1(n15229), .A2(n15228), .A3(n15227), .A4(n15226), .ZN(
        n15230) );
  AOI22_X1 U18327 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U18328 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15234) );
  INV_X2 U18329 ( .A(n9584), .ZN(n16734) );
  AOI22_X1 U18330 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15233) );
  AOI22_X1 U18331 ( .A1(n16796), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15232) );
  NAND4_X1 U18332 ( .A1(n15235), .A2(n15234), .A3(n15233), .A4(n15232), .ZN(
        n15242) );
  AOI22_X1 U18333 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U18334 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15236), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15239) );
  AOI22_X1 U18335 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15238) );
  AOI22_X1 U18336 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15237) );
  NAND4_X1 U18337 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        n15241) );
  AOI22_X1 U18338 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15250) );
  AOI22_X1 U18339 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16786), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15249) );
  AOI22_X1 U18340 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15243) );
  OAI21_X1 U18341 ( .B1(n15273), .B2(n16843), .A(n15243), .ZN(n15248) );
  AOI22_X1 U18342 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15247) );
  AOI22_X1 U18343 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15246) );
  AOI22_X1 U18344 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15245) );
  AOI22_X1 U18345 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15244) );
  AOI22_X1 U18346 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n16779), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n16778), .ZN(n15258) );
  AOI22_X1 U18347 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U18348 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15255) );
  AOI22_X1 U18349 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16800), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15254) );
  AOI22_X1 U18350 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16764), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U18351 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15259), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U18352 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U18353 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16619), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15268) );
  AOI22_X1 U18354 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15260) );
  OAI21_X1 U18355 ( .B1(n9585), .B2(n20605), .A(n15260), .ZN(n15266) );
  AOI22_X1 U18356 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9589), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15264) );
  AOI22_X1 U18357 ( .A1(n16778), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15263) );
  AOI22_X1 U18358 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15262) );
  AOI22_X1 U18359 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15261) );
  NAND4_X1 U18360 ( .A1(n15264), .A2(n15263), .A3(n15262), .A4(n15261), .ZN(
        n15265) );
  AOI211_X1 U18361 ( .C1(n16804), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15266), .B(n15265), .ZN(n15267) );
  NAND3_X1 U18362 ( .A1(n15269), .A2(n15268), .A3(n15267), .ZN(n15300) );
  XOR2_X1 U18363 ( .A(n15300), .B(n15270), .Z(n15289) );
  INV_X1 U18364 ( .A(n16984), .ZN(n15303) );
  XNOR2_X1 U18365 ( .A(n15303), .B(n15271), .ZN(n15287) );
  AND2_X1 U18366 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15287), .ZN(
        n15288) );
  NOR2_X1 U18367 ( .A1(n20606), .A2(n15285), .ZN(n15286) );
  AOI22_X1 U18368 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15283) );
  AOI22_X1 U18369 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15282) );
  INV_X1 U18370 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16799) );
  AOI22_X1 U18371 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15272) );
  OAI21_X1 U18372 ( .B1(n15273), .B2(n16799), .A(n15272), .ZN(n15281) );
  AOI22_X1 U18373 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15279) );
  AOI22_X1 U18374 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U18375 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15277) );
  AOI22_X1 U18376 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15276) );
  NAND4_X1 U18377 ( .A1(n15279), .A2(n15278), .A3(n15277), .A4(n15276), .ZN(
        n15280) );
  NAND2_X1 U18378 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17487), .ZN(
        n17486) );
  NOR2_X1 U18379 ( .A1(n15284), .A2(n17478), .ZN(n17467) );
  XOR2_X1 U18380 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15285), .Z(
        n17466) );
  INV_X1 U18381 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17778) );
  XOR2_X1 U18382 ( .A(n17778), .B(n15287), .Z(n17451) );
  INV_X1 U18383 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17769) );
  XOR2_X1 U18384 ( .A(n17769), .B(n15289), .Z(n17444) );
  XNOR2_X1 U18385 ( .A(n16977), .B(n15291), .ZN(n17429) );
  OAI21_X1 U18386 ( .B1(n15295), .B2(n17644), .A(n17359), .ZN(n15297) );
  NOR2_X1 U18387 ( .A1(n15296), .A2(n15297), .ZN(n15298) );
  NOR2_X2 U18388 ( .A1(n17733), .A2(n15337), .ZN(n17689) );
  NAND2_X1 U18389 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17536), .ZN(
        n17162) );
  NOR2_X1 U18390 ( .A1(n17531), .A2(n17162), .ZN(n17161) );
  NAND2_X1 U18391 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17161), .ZN(
        n17116) );
  NAND2_X1 U18392 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16039) );
  AOI221_X1 U18393 ( .B1(n17688), .B2(n16026), .C1(n17116), .C2(n16026), .A(
        n16039), .ZN(n15330) );
  NAND2_X1 U18394 ( .A1(n18264), .A2(n17793), .ZN(n17802) );
  INV_X1 U18395 ( .A(n15300), .ZN(n16981) );
  INV_X1 U18396 ( .A(n15306), .ZN(n16988) );
  NAND2_X1 U18397 ( .A1(n16988), .A2(n15305), .ZN(n15304) );
  NAND2_X1 U18398 ( .A1(n15304), .A2(n15303), .ZN(n15315) );
  INV_X1 U18399 ( .A(n16977), .ZN(n15301) );
  NAND2_X1 U18400 ( .A1(n15302), .A2(n15301), .ZN(n15321) );
  NOR2_X1 U18401 ( .A1(n9927), .A2(n15321), .ZN(n15324) );
  NAND2_X1 U18402 ( .A1(n15324), .A2(n17644), .ZN(n15325) );
  XOR2_X1 U18403 ( .A(n15302), .B(n15301), .Z(n15319) );
  AND2_X1 U18404 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15319), .ZN(
        n15320) );
  XNOR2_X1 U18405 ( .A(n15304), .B(n15303), .ZN(n15313) );
  NOR2_X1 U18406 ( .A1(n17778), .A2(n15313), .ZN(n15314) );
  NOR2_X1 U18407 ( .A1(n15307), .A2(n20606), .ZN(n15312) );
  XOR2_X1 U18408 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15307), .Z(
        n17469) );
  NOR2_X1 U18409 ( .A1(n15309), .A2(n18447), .ZN(n15310) );
  INV_X1 U18410 ( .A(n17487), .ZN(n15415) );
  NAND3_X1 U18411 ( .A1(n15415), .A2(n15309), .A3(n18447), .ZN(n15308) );
  OAI221_X1 U18412 ( .B1(n15310), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15415), .C2(n15309), .A(n15308), .ZN(n17468) );
  NOR2_X1 U18413 ( .A1(n17469), .A2(n17468), .ZN(n15311) );
  NOR2_X1 U18414 ( .A1(n15312), .A2(n15311), .ZN(n17455) );
  XOR2_X1 U18415 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15313), .Z(
        n17454) );
  NOR2_X1 U18416 ( .A1(n17455), .A2(n17454), .ZN(n17453) );
  XNOR2_X1 U18417 ( .A(n15315), .B(n16981), .ZN(n15317) );
  NOR2_X1 U18418 ( .A1(n15316), .A2(n15317), .ZN(n15318) );
  XOR2_X1 U18419 ( .A(n10030), .B(n15319), .Z(n17432) );
  NOR2_X1 U18420 ( .A1(n17433), .A2(n17432), .ZN(n17431) );
  XNOR2_X1 U18421 ( .A(n15321), .B(n9927), .ZN(n15323) );
  XNOR2_X1 U18422 ( .A(n15323), .B(n15322), .ZN(n17419) );
  XOR2_X1 U18423 ( .A(n15324), .B(n17646), .Z(n15326) );
  NOR2_X1 U18424 ( .A1(n15325), .A2(n15327), .ZN(n15329) );
  INV_X1 U18425 ( .A(n15325), .ZN(n15328) );
  INV_X1 U18426 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17685) );
  NOR2_X1 U18427 ( .A1(n17676), .A2(n17685), .ZN(n17647) );
  INV_X1 U18428 ( .A(n17647), .ZN(n17329) );
  INV_X1 U18429 ( .A(n17173), .ZN(n15340) );
  NOR2_X1 U18430 ( .A1(n15333), .A2(n16039), .ZN(n16042) );
  AOI22_X1 U18431 ( .A1(n17793), .A2(n15330), .B1(n17809), .B2(n16042), .ZN(
        n15399) );
  INV_X1 U18432 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16013) );
  OR3_X2 U18433 ( .A1(n16542), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_0__SCAN_IN), .ZN(n17712) );
  NOR2_X1 U18434 ( .A1(n18270), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17758) );
  NAND2_X1 U18435 ( .A1(n17555), .A2(n17596), .ZN(n17495) );
  NOR2_X1 U18436 ( .A1(n17506), .A2(n17495), .ZN(n17517) );
  NAND2_X1 U18437 ( .A1(n17806), .A2(n18270), .ZN(n17760) );
  INV_X1 U18438 ( .A(n17760), .ZN(n17720) );
  AOI21_X1 U18439 ( .B1(n17496), .B2(n17517), .A(n17720), .ZN(n15331) );
  AOI21_X1 U18440 ( .B1(n17595), .B2(n16035), .A(n18301), .ZN(n17500) );
  NOR4_X1 U18441 ( .A1(n17758), .A2(n15331), .A3(n17500), .A4(n17804), .ZN(
        n15332) );
  OAI21_X1 U18442 ( .B1(n18270), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15332), .ZN(n15393) );
  AOI21_X1 U18443 ( .B1(n17649), .B2(n9925), .A(n15393), .ZN(n16041) );
  OAI21_X1 U18444 ( .B1(n17722), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16041), .ZN(n15336) );
  NOR2_X1 U18445 ( .A1(n16039), .A2(n16013), .ZN(n15396) );
  INV_X1 U18446 ( .A(n15396), .ZN(n16028) );
  NOR2_X1 U18447 ( .A1(n16028), .A2(n17116), .ZN(n16002) );
  NOR2_X1 U18448 ( .A1(n16002), .A2(n17644), .ZN(n15334) );
  NAND2_X1 U18449 ( .A1(n17497), .A2(n15396), .ZN(n15993) );
  AOI22_X1 U18450 ( .A1(n15334), .A2(n17811), .B1(n17809), .B2(n15993), .ZN(
        n15400) );
  INV_X1 U18451 ( .A(n15400), .ZN(n15335) );
  AOI21_X1 U18452 ( .B1(n17712), .B2(n15336), .A(n15335), .ZN(n15347) );
  NAND2_X1 U18453 ( .A1(n17261), .A2(n17249), .ZN(n17235) );
  NOR2_X1 U18454 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17235), .ZN(
        n17220) );
  INV_X1 U18455 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17556) );
  NAND2_X1 U18456 ( .A1(n17220), .A2(n17556), .ZN(n17204) );
  NOR3_X1 U18457 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17204), .ZN(n15341) );
  NOR2_X1 U18458 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17313) );
  NOR2_X1 U18459 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17635) );
  NOR2_X1 U18460 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17349) );
  INV_X1 U18461 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17660) );
  NAND2_X1 U18462 ( .A1(n15338), .A2(n17631), .ZN(n17277) );
  INV_X1 U18463 ( .A(n15338), .ZN(n15339) );
  AOI221_X1 U18464 ( .B1(n17388), .B2(n17624), .C1(n17631), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15339), .ZN(n17273) );
  OAI221_X1 U18465 ( .B1(n15341), .B2(n15340), .C1(n15341), .C2(n17277), .A(
        n17205), .ZN(n17176) );
  INV_X1 U18466 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17254) );
  NAND2_X1 U18467 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17207), .ZN(
        n17182) );
  INV_X1 U18468 ( .A(n17175), .ZN(n17164) );
  NAND2_X1 U18469 ( .A1(n17359), .A2(n17164), .ZN(n15342) );
  OAI221_X1 U18470 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17359), 
        .C1(n17531), .C2(n15343), .A(n15342), .ZN(n17144) );
  NOR2_X1 U18471 ( .A1(n15343), .A2(n17359), .ZN(n17163) );
  INV_X1 U18472 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17118) );
  NOR2_X1 U18473 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17359), .ZN(
        n16036) );
  AOI21_X1 U18474 ( .B1(n15395), .B2(n15394), .A(n16036), .ZN(n15345) );
  XOR2_X1 U18475 ( .A(n15345), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16016) );
  AOI22_X1 U18476 ( .A1(n9597), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17681), 
        .B2(n16016), .ZN(n15346) );
  OAI221_X1 U18477 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15399), 
        .C1(n16013), .C2(n15347), .A(n15346), .ZN(P3_U2833) );
  AOI22_X1 U18478 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n18563), .ZN(n15355) );
  AOI22_X1 U18479 ( .A1(n15348), .A2(n18639), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18677), .ZN(n15354) );
  OAI22_X1 U18480 ( .A1(n15743), .A2(n18656), .B1(n18676), .B2(n15714), .ZN(
        n15349) );
  INV_X1 U18481 ( .A(n15349), .ZN(n15353) );
  OAI211_X1 U18482 ( .C1(n15351), .C2(n15749), .A(n18678), .B(n15350), .ZN(
        n15352) );
  NAND4_X1 U18483 ( .A1(n15355), .A2(n15354), .A3(n15353), .A4(n15352), .ZN(
        P2_U2833) );
  INV_X1 U18484 ( .A(n15364), .ZN(n15366) );
  NOR3_X1 U18485 ( .A1(n15357), .A2(n15356), .A3(n20259), .ZN(n15361) );
  INV_X1 U18486 ( .A(n15358), .ZN(n15359) );
  OAI22_X1 U18487 ( .A1(n15361), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n15360), .B2(n15359), .ZN(n15363) );
  NAND2_X1 U18488 ( .A1(n15361), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15362) );
  OAI211_X1 U18489 ( .C1(n15364), .C2(n20226), .A(n15363), .B(n15362), .ZN(
        n15365) );
  OAI21_X1 U18490 ( .B1(n15366), .B2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n15365), .ZN(n15367) );
  AOI222_X1 U18491 ( .A1(n20626), .A2(n15368), .B1(n20626), .B2(n15367), .C1(
        n15368), .C2(n15367), .ZN(n15378) );
  INV_X1 U18492 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15369) );
  NAND2_X1 U18493 ( .A1(n19617), .A2(n15369), .ZN(n15370) );
  NAND2_X1 U18494 ( .A1(n15371), .A2(n15370), .ZN(n15372) );
  AND4_X1 U18495 ( .A1(n15375), .A2(n15374), .A3(n15373), .A4(n15372), .ZN(
        n15376) );
  OAI211_X1 U18496 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15378), .A(
        n15377), .B(n15376), .ZN(n15383) );
  NOR3_X1 U18497 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11260), .A3(n20415), 
        .ZN(n15381) );
  NAND2_X1 U18498 ( .A1(n20291), .A2(n20415), .ZN(n15379) );
  OAI22_X1 U18499 ( .A1(n15384), .A2(n15381), .B1(n15380), .B2(n15379), .ZN(
        n15659) );
  AOI221_X1 U18500 ( .B1(n20401), .B2(n20400), .C1(n15383), .C2(n20400), .A(
        n15659), .ZN(n15663) );
  AOI21_X1 U18501 ( .B1(n15384), .B2(n15383), .A(n15382), .ZN(n15386) );
  OAI211_X1 U18502 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20415), .A(n15386), 
        .B(n15385), .ZN(n15387) );
  NOR2_X1 U18503 ( .A1(n15663), .A2(n15387), .ZN(n15392) );
  NAND2_X1 U18504 ( .A1(n15389), .A2(n15388), .ZN(n15390) );
  NAND2_X1 U18505 ( .A1(n20401), .A2(n15390), .ZN(n15391) );
  OAI22_X1 U18506 ( .A1(n15392), .A2(n20401), .B1(n15663), .B2(n15391), .ZN(
        P1_U3161) );
  INV_X1 U18507 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16027) );
  OAI221_X1 U18508 ( .B1(n15393), .B2(n17619), .C1(n15393), .C2(n16028), .A(
        n17712), .ZN(n16022) );
  NAND2_X1 U18509 ( .A1(n15396), .A2(n16027), .ZN(n16004) );
  NOR2_X1 U18510 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15394), .ZN(
        n15975) );
  INV_X1 U18511 ( .A(n15975), .ZN(n15397) );
  INV_X1 U18512 ( .A(n15395), .ZN(n16038) );
  NAND2_X1 U18513 ( .A1(n15396), .A2(n16038), .ZN(n15977) );
  OAI21_X1 U18514 ( .B1(n17388), .B2(n15397), .A(n15977), .ZN(n15398) );
  NAND2_X1 U18515 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15398), .ZN(
        n15976) );
  INV_X1 U18516 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20422) );
  INV_X1 U18517 ( .A(HOLD), .ZN(n20407) );
  NOR2_X1 U18518 ( .A1(n20422), .A2(n20407), .ZN(n15403) );
  AOI22_X1 U18519 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15402) );
  NAND2_X1 U18520 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20491), .ZN(n20406) );
  OAI211_X1 U18521 ( .C1(n15403), .C2(n15402), .A(n15401), .B(n20406), .ZN(
        P1_U3195) );
  AND2_X1 U18522 ( .A1(n19758), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U18523 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15404) );
  NOR2_X1 U18524 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19596) );
  NAND2_X1 U18525 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18921), .ZN(n19461) );
  NOR2_X1 U18526 ( .A1(n19602), .A2(n19461), .ZN(n15960) );
  NOR4_X1 U18527 ( .A1(n15404), .A2(n19596), .A3(n15960), .A4(n15962), .ZN(
        P2_U3178) );
  INV_X1 U18528 ( .A(n15961), .ZN(n19583) );
  INV_X1 U18529 ( .A(n19596), .ZN(n15406) );
  NAND2_X1 U18530 ( .A1(n15406), .A2(n15405), .ZN(n15407) );
  AOI221_X1 U18531 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15962), .C1(n19583), .C2(
        n15962), .A(n19405), .ZN(n19579) );
  INV_X1 U18532 ( .A(n19579), .ZN(n19576) );
  NOR2_X1 U18533 ( .A1(n15409), .A2(n19576), .ZN(P2_U3047) );
  INV_X1 U18534 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n17824) );
  NAND2_X1 U18535 ( .A1(n15413), .A2(n16856), .ZN(n16992) );
  INV_X1 U18536 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17060) );
  AOI21_X1 U18537 ( .B1(n16856), .B2(n17864), .A(P3_EAX_REG_0__SCAN_IN), .ZN(
        n15416) );
  OAI222_X1 U18538 ( .A1(n17824), .A2(n16992), .B1(n16940), .B2(n15416), .C1(
        n16989), .C2(n15415), .ZN(P3_U2735) );
  OAI22_X1 U18539 ( .A1(n15417), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n18531), .B2(n18832), .ZN(n15418) );
  AOI211_X1 U18540 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15420), .A(
        n15419), .B(n15418), .ZN(n15424) );
  INV_X1 U18541 ( .A(n15421), .ZN(n18519) );
  AOI22_X1 U18542 ( .A1(n15422), .A2(n18846), .B1(n18853), .B2(n18519), .ZN(
        n15423) );
  OAI211_X1 U18543 ( .C1(n15425), .C2(n15926), .A(n15424), .B(n15423), .ZN(
        P2_U3025) );
  OR2_X1 U18544 ( .A1(n19695), .A2(n15426), .ZN(n15430) );
  INV_X1 U18545 ( .A(n15427), .ZN(n15428) );
  AOI22_X1 U18546 ( .A1(n15428), .A2(n19641), .B1(n19710), .B2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15429) );
  AND2_X1 U18547 ( .A1(n15430), .A2(n15429), .ZN(n15437) );
  INV_X1 U18548 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15431) );
  OAI21_X1 U18549 ( .B1(n13855), .B2(n15432), .A(n15431), .ZN(n15433) );
  AOI22_X1 U18550 ( .A1(n15435), .A2(n19667), .B1(n15434), .B2(n15433), .ZN(
        n15436) );
  OAI211_X1 U18551 ( .C1(n19673), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        P1_U2817) );
  OAI22_X1 U18552 ( .A1(n19695), .A2(n15440), .B1(n19686), .B2(n15439), .ZN(
        n15448) );
  OAI22_X1 U18553 ( .A1(n15443), .A2(n20451), .B1(n15442), .B2(n15441), .ZN(
        n15447) );
  OAI22_X1 U18554 ( .A1(n15445), .A2(n15480), .B1(n15444), .B2(n19673), .ZN(
        n15446) );
  NOR3_X1 U18555 ( .A1(n15448), .A2(n15447), .A3(n15446), .ZN(n15449) );
  OAI21_X1 U18556 ( .B1(n15450), .B2(n19713), .A(n15449), .ZN(P1_U2819) );
  INV_X1 U18557 ( .A(n15451), .ZN(n15510) );
  INV_X1 U18558 ( .A(n15452), .ZN(n15453) );
  INV_X1 U18559 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20449) );
  NAND3_X1 U18560 ( .A1(n15454), .A2(n15453), .A3(n20449), .ZN(n15458) );
  INV_X1 U18561 ( .A(n15514), .ZN(n15456) );
  NOR2_X1 U18562 ( .A1(n19686), .A2(n11590), .ZN(n15455) );
  AOI211_X1 U18563 ( .C1(n19641), .C2(n15456), .A(n19650), .B(n15455), .ZN(
        n15457) );
  OAI211_X1 U18564 ( .C1(n15459), .C2(n19695), .A(n15458), .B(n15457), .ZN(
        n15460) );
  AOI21_X1 U18565 ( .B1(n15510), .B2(n19667), .A(n15460), .ZN(n15464) );
  OAI21_X1 U18566 ( .B1(n15462), .B2(n15461), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15463) );
  OAI211_X1 U18567 ( .C1(n15465), .C2(n19673), .A(n15464), .B(n15463), .ZN(
        P1_U2821) );
  OAI21_X1 U18568 ( .B1(n19686), .B2(n15466), .A(n19693), .ZN(n15467) );
  AOI21_X1 U18569 ( .B1(n19708), .B2(P1_EBX_REG_15__SCAN_IN), .A(n15467), .ZN(
        n15468) );
  OAI21_X1 U18570 ( .B1(n15486), .B2(n20443), .A(n15468), .ZN(n15469) );
  AOI211_X1 U18571 ( .C1(n15528), .C2(n19667), .A(n15470), .B(n15469), .ZN(
        n15474) );
  XNOR2_X1 U18572 ( .A(n15472), .B(n15471), .ZN(n15585) );
  AOI22_X1 U18573 ( .A1(n15527), .A2(n19641), .B1(n19707), .B2(n15585), .ZN(
        n15473) );
  NAND2_X1 U18574 ( .A1(n15474), .A2(n15473), .ZN(P1_U2825) );
  AOI21_X1 U18575 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15475), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15485) );
  INV_X1 U18576 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15477) );
  OAI22_X1 U18577 ( .A1(n19695), .A2(n15477), .B1(n19686), .B2(n15476), .ZN(
        n15478) );
  AOI211_X1 U18578 ( .C1(n15592), .C2(n19707), .A(n19650), .B(n15478), .ZN(
        n15484) );
  OAI22_X1 U18579 ( .A1(n15481), .A2(n15480), .B1(n15479), .B2(n19713), .ZN(
        n15482) );
  INV_X1 U18580 ( .A(n15482), .ZN(n15483) );
  OAI211_X1 U18581 ( .C1(n15486), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        P1_U2826) );
  AOI22_X1 U18582 ( .A1(n19708), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19710), .ZN(n15496) );
  AND2_X1 U18583 ( .A1(n15488), .A2(n15487), .ZN(n15489) );
  NOR2_X1 U18584 ( .A1(n15490), .A2(n15489), .ZN(n15599) );
  AOI21_X1 U18585 ( .B1(n15599), .B2(n19707), .A(n19650), .ZN(n15495) );
  AOI22_X1 U18586 ( .A1(n15535), .A2(n19641), .B1(n19667), .B2(n15534), .ZN(
        n15494) );
  AND2_X1 U18587 ( .A1(n15491), .A2(n19634), .ZN(n15502) );
  OAI221_X1 U18588 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n15502), .A(n15492), .ZN(n15493) );
  NAND4_X1 U18589 ( .A1(n15496), .A2(n15495), .A3(n15494), .A4(n15493), .ZN(
        P1_U2828) );
  AOI21_X1 U18590 ( .B1(n19710), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19650), .ZN(n15497) );
  INV_X1 U18591 ( .A(n15497), .ZN(n15501) );
  OAI22_X1 U18592 ( .A1(n15499), .A2(n19673), .B1(n15498), .B2(n19695), .ZN(
        n15500) );
  AOI211_X1 U18593 ( .C1(n15502), .C2(n14106), .A(n15501), .B(n15500), .ZN(
        n15505) );
  AOI22_X1 U18594 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15503), .B1(n19667), 
        .B2(n15539), .ZN(n15504) );
  OAI211_X1 U18595 ( .C1(n15543), .C2(n19713), .A(n15505), .B(n15504), .ZN(
        P1_U2829) );
  AOI22_X1 U18596 ( .A1(n15528), .A2(n11912), .B1(n19725), .B2(n15585), .ZN(
        n15506) );
  OAI21_X1 U18597 ( .B1(n19728), .B2(n15507), .A(n15506), .ZN(P1_U2857) );
  INV_X1 U18598 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U18599 ( .A1(n15534), .A2(n11912), .B1(n19725), .B2(n15599), .ZN(
        n15508) );
  OAI21_X1 U18600 ( .B1(n19728), .B2(n15509), .A(n15508), .ZN(P1_U2860) );
  AOI22_X1 U18601 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U18602 ( .A1(n15511), .A2(n19795), .B1(n19794), .B2(n15510), .ZN(
        n15512) );
  OAI211_X1 U18603 ( .C1(n19810), .C2(n15514), .A(n15513), .B(n15512), .ZN(
        P1_U2980) );
  AOI21_X1 U18604 ( .B1(n13910), .B2(n15515), .A(n9827), .ZN(n15517) );
  NOR2_X1 U18605 ( .A1(n15517), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15516) );
  MUX2_X1 U18606 ( .A(n15517), .B(n15516), .S(n10117), .Z(n15518) );
  XNOR2_X1 U18607 ( .A(n15518), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15581) );
  AOI22_X1 U18608 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U18609 ( .A1(n15520), .A2(n19794), .B1(n15536), .B2(n15519), .ZN(
        n15521) );
  OAI211_X1 U18610 ( .C1(n19804), .C2(n15581), .A(n15522), .B(n15521), .ZN(
        P1_U2982) );
  MUX2_X1 U18611 ( .A(n13192), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .S(
        n9615), .Z(n15526) );
  NOR2_X1 U18612 ( .A1(n15524), .A2(n15523), .ZN(n15525) );
  XOR2_X1 U18613 ( .A(n15526), .B(n15525), .Z(n15588) );
  AOI22_X1 U18614 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15530) );
  AOI22_X1 U18615 ( .A1(n15528), .A2(n19794), .B1(n15527), .B2(n15536), .ZN(
        n15529) );
  OAI211_X1 U18616 ( .C1(n15588), .C2(n19804), .A(n15530), .B(n15529), .ZN(
        P1_U2984) );
  AOI21_X1 U18617 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n15610) );
  AOI22_X1 U18618 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U18619 ( .A1(n15536), .A2(n15535), .B1(n19794), .B2(n15534), .ZN(
        n15537) );
  OAI211_X1 U18620 ( .C1(n15610), .C2(n19804), .A(n15538), .B(n15537), .ZN(
        P1_U2987) );
  AOI22_X1 U18621 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U18622 ( .A1(n19795), .A2(n15540), .B1(n19794), .B2(n15539), .ZN(
        n15541) );
  OAI211_X1 U18623 ( .C1(n19810), .C2(n15543), .A(n15542), .B(n15541), .ZN(
        P1_U2988) );
  AOI22_X1 U18624 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15549) );
  NAND2_X1 U18625 ( .A1(n15545), .A2(n15544), .ZN(n15546) );
  XNOR2_X1 U18626 ( .A(n15547), .B(n15546), .ZN(n15635) );
  AOI22_X1 U18627 ( .A1(n15635), .A2(n19795), .B1(n19794), .B2(n19647), .ZN(
        n15548) );
  OAI211_X1 U18628 ( .C1(n19810), .C2(n19651), .A(n15549), .B(n15548), .ZN(
        P1_U2992) );
  AOI22_X1 U18629 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15554) );
  XNOR2_X1 U18630 ( .A(n15550), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15551) );
  XNOR2_X1 U18631 ( .A(n15552), .B(n15551), .ZN(n15645) );
  AOI22_X1 U18632 ( .A1(n15645), .A2(n19795), .B1(n19794), .B2(n19722), .ZN(
        n15553) );
  OAI211_X1 U18633 ( .C1(n19810), .C2(n19669), .A(n15554), .B(n15553), .ZN(
        P1_U2993) );
  AOI22_X1 U18634 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15561) );
  OAI21_X1 U18635 ( .B1(n15557), .B2(n15556), .A(n15555), .ZN(n15558) );
  INV_X1 U18636 ( .A(n15558), .ZN(n15653) );
  INV_X1 U18637 ( .A(n15559), .ZN(n19676) );
  AOI22_X1 U18638 ( .A1(n15653), .A2(n19795), .B1(n19794), .B2(n19676), .ZN(
        n15560) );
  OAI211_X1 U18639 ( .C1(n19810), .C2(n19683), .A(n15561), .B(n15560), .ZN(
        P1_U2994) );
  AOI21_X1 U18640 ( .B1(n15563), .B2(n15562), .A(n15591), .ZN(n15573) );
  NOR2_X1 U18641 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15583), .ZN(
        n15564) );
  AOI22_X1 U18642 ( .A1(n12502), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n15565), 
        .B2(n15564), .ZN(n15571) );
  INV_X1 U18643 ( .A(n15566), .ZN(n15569) );
  INV_X1 U18644 ( .A(n15567), .ZN(n15568) );
  AOI22_X1 U18645 ( .A1(n15569), .A2(n19823), .B1(n19825), .B2(n15568), .ZN(
        n15570) );
  OAI211_X1 U18646 ( .C1(n15573), .C2(n15572), .A(n15571), .B(n15570), .ZN(
        P1_U3013) );
  AOI221_X1 U18647 ( .B1(n15575), .B2(n15574), .C1(n15583), .C2(n15574), .A(
        n15573), .ZN(n15578) );
  NOR2_X1 U18648 ( .A1(n15576), .A2(n19834), .ZN(n15577) );
  NOR2_X1 U18649 ( .A1(n15578), .A2(n15577), .ZN(n15580) );
  NAND2_X1 U18650 ( .A1(n12502), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15579) );
  OAI211_X1 U18651 ( .C1(n15581), .C2(n19838), .A(n15580), .B(n15579), .ZN(
        P1_U3014) );
  AOI22_X1 U18652 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15582), .B1(
        n12502), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15587) );
  NOR2_X1 U18653 ( .A1(n15589), .A2(n15583), .ZN(n15584) );
  AOI22_X1 U18654 ( .A1(n15585), .A2(n19825), .B1(n13192), .B2(n15584), .ZN(
        n15586) );
  OAI211_X1 U18655 ( .C1(n15588), .C2(n19838), .A(n15587), .B(n15586), .ZN(
        P1_U3016) );
  NAND2_X1 U18656 ( .A1(n15590), .A2(n15589), .ZN(n15596) );
  AOI22_X1 U18657 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15591), .B1(
        n12502), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15595) );
  AOI22_X1 U18658 ( .A1(n15593), .A2(n19823), .B1(n19825), .B2(n15592), .ZN(
        n15594) );
  OAI211_X1 U18659 ( .C1(n15606), .C2(n15596), .A(n15595), .B(n15594), .ZN(
        P1_U3017) );
  AOI221_X1 U18660 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15598), 
        .C1(n15597), .C2(n15598), .A(n13196), .ZN(n15604) );
  INV_X1 U18661 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15602) );
  NAND2_X1 U18662 ( .A1(n15599), .A2(n19825), .ZN(n15600) );
  OAI21_X1 U18663 ( .B1(n15602), .B2(n15601), .A(n15600), .ZN(n15603) );
  NOR2_X1 U18664 ( .A1(n15604), .A2(n15603), .ZN(n15609) );
  NOR2_X1 U18665 ( .A1(n15606), .A2(n15605), .ZN(n15644) );
  NAND3_X1 U18666 ( .A1(n15607), .A2(n15644), .A3(n13196), .ZN(n15608) );
  OAI211_X1 U18667 ( .C1(n15610), .C2(n19838), .A(n15609), .B(n15608), .ZN(
        P1_U3019) );
  OAI211_X1 U18668 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15611), .B(n15650), .ZN(n15618) );
  AOI21_X1 U18669 ( .B1(n15613), .B2(n19825), .A(n15612), .ZN(n15617) );
  AOI22_X1 U18670 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15615), .B1(
        n19823), .B2(n15614), .ZN(n15616) );
  OAI211_X1 U18671 ( .C1(n15619), .C2(n15618), .A(n15617), .B(n15616), .ZN(
        P1_U3021) );
  NAND2_X1 U18672 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15644), .ZN(
        n15638) );
  INV_X1 U18673 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15621) );
  INV_X1 U18674 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U18675 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15621), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15620), .ZN(n15633) );
  AOI21_X1 U18676 ( .B1(n15623), .B2(n19825), .A(n15622), .ZN(n15632) );
  NAND2_X1 U18677 ( .A1(n15624), .A2(n19815), .ZN(n15656) );
  INV_X1 U18678 ( .A(n15656), .ZN(n15627) );
  OAI21_X1 U18679 ( .B1(n15626), .B2(n19815), .A(n15625), .ZN(n15652) );
  AOI21_X1 U18680 ( .B1(n15628), .B2(n15627), .A(n15652), .ZN(n15649) );
  OAI21_X1 U18681 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15629), .A(
        n15649), .ZN(n15634) );
  AOI22_X1 U18682 ( .A1(n15630), .A2(n19823), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n15634), .ZN(n15631) );
  OAI211_X1 U18683 ( .C1(n15638), .C2(n15633), .A(n15632), .B(n15631), .ZN(
        P1_U3023) );
  AOI22_X1 U18684 ( .A1(n19654), .A2(n19825), .B1(n12502), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U18685 ( .A1(n15635), .A2(n19823), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15634), .ZN(n15636) );
  OAI211_X1 U18686 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n15638), .A(
        n15637), .B(n15636), .ZN(P1_U3024) );
  INV_X1 U18687 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15648) );
  AOI21_X1 U18688 ( .B1(n15641), .B2(n15640), .A(n15639), .ZN(n15643) );
  OR2_X1 U18689 ( .A1(n15643), .A2(n15642), .ZN(n19662) );
  INV_X1 U18690 ( .A(n19662), .ZN(n19721) );
  AOI22_X1 U18691 ( .A1(n19721), .A2(n19825), .B1(n12502), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15647) );
  AOI22_X1 U18692 ( .A1(n15645), .A2(n19823), .B1(n15648), .B2(n15644), .ZN(
        n15646) );
  OAI211_X1 U18693 ( .C1(n15649), .C2(n15648), .A(n15647), .B(n15646), .ZN(
        P1_U3025) );
  NAND2_X1 U18694 ( .A1(n19811), .A2(n15650), .ZN(n19829) );
  INV_X1 U18695 ( .A(n19674), .ZN(n15651) );
  AOI22_X1 U18696 ( .A1(n15651), .A2(n19825), .B1(n12502), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U18697 ( .A1(n15653), .A2(n19823), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15652), .ZN(n15654) );
  OAI211_X1 U18698 ( .C1(n15656), .C2(n19829), .A(n15655), .B(n15654), .ZN(
        P1_U3026) );
  NAND4_X1 U18699 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n11260), .A4(n20415), .ZN(n15657) );
  NAND2_X1 U18700 ( .A1(n15658), .A2(n15657), .ZN(n20402) );
  OAI21_X1 U18701 ( .B1(n15660), .B2(n20402), .A(n15659), .ZN(n15661) );
  OAI221_X1 U18702 ( .B1(n20494), .B2(n20232), .C1(n20494), .C2(n20415), .A(
        n15661), .ZN(n15662) );
  AOI221_X1 U18703 ( .B1(n15663), .B2(n20400), .C1(n20401), .C2(n20400), .A(
        n15662), .ZN(P1_U3162) );
  NOR2_X1 U18704 ( .A1(n15663), .A2(n20401), .ZN(n15665) );
  OAI22_X1 U18705 ( .A1(n20232), .A2(n15665), .B1(n15664), .B2(n20401), .ZN(
        P1_U3466) );
  AOI22_X1 U18706 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n18563), .ZN(n15678) );
  INV_X1 U18707 ( .A(n15666), .ZN(n15667) );
  AOI22_X1 U18708 ( .A1(n15667), .A2(n18639), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18677), .ZN(n15677) );
  INV_X1 U18709 ( .A(n15668), .ZN(n15669) );
  OAI22_X1 U18710 ( .A1(n15670), .A2(n18656), .B1(n15669), .B2(n18676), .ZN(
        n15671) );
  INV_X1 U18711 ( .A(n15671), .ZN(n15676) );
  OAI211_X1 U18712 ( .C1(n15674), .C2(n15673), .A(n18678), .B(n15672), .ZN(
        n15675) );
  NAND4_X1 U18713 ( .A1(n15678), .A2(n15677), .A3(n15676), .A4(n15675), .ZN(
        P2_U2829) );
  NAND2_X1 U18714 ( .A1(n15695), .A2(n18669), .ZN(n15679) );
  XOR2_X1 U18715 ( .A(n15680), .B(n15679), .Z(n15689) );
  AOI22_X1 U18716 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n18563), .ZN(n15682) );
  NAND2_X1 U18717 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18677), .ZN(
        n15681) );
  OAI211_X1 U18718 ( .C1(n15683), .C2(n18676), .A(n15682), .B(n15681), .ZN(
        n15686) );
  NOR2_X1 U18719 ( .A1(n15684), .A2(n18656), .ZN(n15685) );
  AOI211_X1 U18720 ( .C1(n18639), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        n15688) );
  OAI21_X1 U18721 ( .B1(n19465), .B2(n15689), .A(n15688), .ZN(P2_U2830) );
  AOI22_X1 U18722 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n18667), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n18563), .ZN(n15701) );
  OAI22_X1 U18723 ( .A1(n15690), .A2(n18687), .B1(n18663), .B2(n10014), .ZN(
        n15691) );
  INV_X1 U18724 ( .A(n15691), .ZN(n15700) );
  OAI22_X1 U18725 ( .A1(n15693), .A2(n18656), .B1(n15692), .B2(n18676), .ZN(
        n15694) );
  INV_X1 U18726 ( .A(n15694), .ZN(n15699) );
  OAI211_X1 U18727 ( .C1(n15697), .C2(n15696), .A(n18678), .B(n15695), .ZN(
        n15698) );
  NAND4_X1 U18728 ( .A1(n15701), .A2(n15700), .A3(n15699), .A4(n15698), .ZN(
        P2_U2831) );
  OAI22_X1 U18729 ( .A1(n18679), .A2(n12101), .B1(n12104), .B2(n18681), .ZN(
        n15702) );
  AOI21_X1 U18730 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18677), .A(
        n15702), .ZN(n15704) );
  NAND2_X1 U18731 ( .A1(n15738), .A2(n18689), .ZN(n15703) );
  OAI211_X1 U18732 ( .C1(n15705), .C2(n18687), .A(n15704), .B(n15703), .ZN(
        n15706) );
  INV_X1 U18733 ( .A(n15706), .ZN(n15711) );
  OAI211_X1 U18734 ( .C1(n15709), .C2(n15708), .A(n18678), .B(n15707), .ZN(
        n15710) );
  OAI211_X1 U18735 ( .C1(n18676), .C2(n15712), .A(n15711), .B(n15710), .ZN(
        P2_U2832) );
  AOI22_X1 U18736 ( .A1(n18701), .A2(n15713), .B1(n18756), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U18737 ( .A1(n18703), .A2(BUF1_REG_22__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15718) );
  INV_X1 U18738 ( .A(n15714), .ZN(n15715) );
  AOI22_X1 U18739 ( .A1(n15716), .A2(n18761), .B1(n18757), .B2(n15715), .ZN(
        n15717) );
  NAND3_X1 U18740 ( .A1(n15719), .A2(n15718), .A3(n15717), .ZN(P2_U2897) );
  AOI22_X1 U18741 ( .A1(n18701), .A2(n15720), .B1(n18756), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U18742 ( .A1(n18703), .A2(BUF1_REG_20__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15727) );
  INV_X1 U18743 ( .A(n15721), .ZN(n15722) );
  OAI22_X1 U18744 ( .A1(n15724), .A2(n18733), .B1(n15723), .B2(n15722), .ZN(
        n15725) );
  INV_X1 U18745 ( .A(n15725), .ZN(n15726) );
  NAND3_X1 U18746 ( .A1(n15728), .A2(n15727), .A3(n15726), .ZN(P2_U2899) );
  AOI22_X1 U18747 ( .A1(n18701), .A2(n18748), .B1(n18756), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15733) );
  AOI22_X1 U18748 ( .A1(n18703), .A2(BUF1_REG_18__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n15732) );
  INV_X1 U18749 ( .A(n18551), .ZN(n15729) );
  AOI22_X1 U18750 ( .A1(n15730), .A2(n18761), .B1(n18757), .B2(n15729), .ZN(
        n15731) );
  NAND3_X1 U18751 ( .A1(n15733), .A2(n15732), .A3(n15731), .ZN(P2_U2901) );
  AOI22_X1 U18752 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n18815), .B1(n15824), 
        .B2(n15734), .ZN(n15740) );
  OAI22_X1 U18753 ( .A1(n15736), .A2(n15817), .B1(n15816), .B2(n15735), .ZN(
        n15737) );
  AOI21_X1 U18754 ( .B1(n18819), .B2(n15738), .A(n15737), .ZN(n15739) );
  OAI211_X1 U18755 ( .C1(n15833), .C2(n20563), .A(n15740), .B(n15739), .ZN(
        P2_U2991) );
  AOI22_X1 U18756 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18815), .ZN(n15748) );
  NOR3_X1 U18757 ( .A1(n15742), .A2(n15741), .A3(n15816), .ZN(n15745) );
  NOR2_X1 U18758 ( .A1(n15743), .A2(n15828), .ZN(n15744) );
  AOI211_X1 U18759 ( .C1(n15746), .C2(n18811), .A(n15745), .B(n15744), .ZN(
        n15747) );
  OAI211_X1 U18760 ( .C1(n18817), .C2(n15749), .A(n15748), .B(n15747), .ZN(
        P2_U2992) );
  AOI22_X1 U18761 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18815), .ZN(n15753) );
  AOI22_X1 U18762 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18815), .ZN(n15765) );
  INV_X1 U18763 ( .A(n15754), .ZN(n15759) );
  OAI21_X1 U18764 ( .B1(n15758), .B2(n15756), .A(n15755), .ZN(n15757) );
  OAI21_X1 U18765 ( .B1(n15759), .B2(n15758), .A(n15757), .ZN(n15867) );
  INV_X1 U18766 ( .A(n15760), .ZN(n15761) );
  AOI21_X1 U18767 ( .B1(n15870), .B2(n15762), .A(n15761), .ZN(n15863) );
  AOI222_X1 U18768 ( .A1(n15867), .A2(n18811), .B1(n18819), .B2(n15763), .C1(
        n18814), .C2(n15863), .ZN(n15764) );
  OAI211_X1 U18769 ( .C1(n18817), .C2(n15766), .A(n15765), .B(n15764), .ZN(
        P2_U3000) );
  AOI22_X1 U18770 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18815), .ZN(n15774) );
  NAND2_X1 U18771 ( .A1(n9637), .A2(n15767), .ZN(n15769) );
  XOR2_X1 U18772 ( .A(n15769), .B(n15768), .Z(n15877) );
  XNOR2_X1 U18773 ( .A(n15771), .B(n15770), .ZN(n15880) );
  OAI22_X1 U18774 ( .A1(n15880), .A2(n15816), .B1(n15828), .B2(n15875), .ZN(
        n15772) );
  AOI21_X1 U18775 ( .B1(n15877), .B2(n18811), .A(n15772), .ZN(n15773) );
  OAI211_X1 U18776 ( .C1(n18817), .C2(n15775), .A(n15774), .B(n15773), .ZN(
        P2_U3002) );
  AOI22_X1 U18777 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18815), .B1(n15824), 
        .B2(n18608), .ZN(n15780) );
  OAI22_X1 U18778 ( .A1(n15777), .A2(n15816), .B1(n15776), .B2(n15817), .ZN(
        n15778) );
  AOI21_X1 U18779 ( .B1(n18819), .B2(n18609), .A(n15778), .ZN(n15779) );
  OAI211_X1 U18780 ( .C1(n15833), .C2(n18602), .A(n15780), .B(n15779), .ZN(
        P2_U3003) );
  AOI22_X1 U18781 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18815), .ZN(n15793) );
  NOR2_X1 U18782 ( .A1(n15782), .A2(n15781), .ZN(n15786) );
  NAND2_X1 U18783 ( .A1(n15784), .A2(n15783), .ZN(n15785) );
  XNOR2_X1 U18784 ( .A(n15786), .B(n15785), .ZN(n15890) );
  INV_X1 U18785 ( .A(n15890), .ZN(n15791) );
  AND2_X1 U18786 ( .A1(n15788), .A2(n15787), .ZN(n15789) );
  NOR2_X1 U18787 ( .A1(n15790), .A2(n15789), .ZN(n15887) );
  AOI222_X1 U18788 ( .A1(n15791), .A2(n18811), .B1(n18819), .B2(n18618), .C1(
        n18814), .C2(n15887), .ZN(n15792) );
  OAI211_X1 U18789 ( .C1(n18817), .C2(n18615), .A(n15793), .B(n15792), .ZN(
        P2_U3004) );
  AOI22_X1 U18790 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18815), .B1(n15824), 
        .B2(n18631), .ZN(n15798) );
  OAI22_X1 U18791 ( .A1(n15795), .A2(n15817), .B1(n15794), .B2(n15816), .ZN(
        n15796) );
  AOI21_X1 U18792 ( .B1(n18819), .B2(n18632), .A(n15796), .ZN(n15797) );
  OAI211_X1 U18793 ( .C1(n15833), .C2(n18625), .A(n15798), .B(n15797), .ZN(
        P2_U3005) );
  AOI22_X1 U18794 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18815), .ZN(n15812) );
  INV_X1 U18795 ( .A(n15799), .ZN(n15800) );
  XNOR2_X1 U18796 ( .A(n15801), .B(n15800), .ZN(n15892) );
  NAND2_X1 U18797 ( .A1(n15892), .A2(n18814), .ZN(n15809) );
  NAND2_X1 U18798 ( .A1(n14589), .A2(n15802), .ZN(n15807) );
  INV_X1 U18799 ( .A(n15803), .ZN(n15804) );
  NOR2_X1 U18800 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  XNOR2_X1 U18801 ( .A(n15807), .B(n15806), .ZN(n15897) );
  NAND2_X1 U18802 ( .A1(n15897), .A2(n18811), .ZN(n15808) );
  OAI211_X1 U18803 ( .C1(n15828), .C2(n15893), .A(n15809), .B(n15808), .ZN(
        n15810) );
  INV_X1 U18804 ( .A(n15810), .ZN(n15811) );
  OAI211_X1 U18805 ( .C1(n18817), .C2(n15813), .A(n15812), .B(n15811), .ZN(
        P2_U3006) );
  AOI22_X1 U18806 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18815), .B1(n15824), 
        .B2(n18671), .ZN(n15821) );
  INV_X1 U18807 ( .A(n15814), .ZN(n15818) );
  OAI22_X1 U18808 ( .A1(n15818), .A2(n15817), .B1(n15816), .B2(n15815), .ZN(
        n15819) );
  AOI21_X1 U18809 ( .B1(n18819), .B2(n18672), .A(n15819), .ZN(n15820) );
  OAI211_X1 U18810 ( .C1(n15833), .C2(n15822), .A(n15821), .B(n15820), .ZN(
        P2_U3009) );
  AOI22_X1 U18811 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n18815), .B1(n15824), 
        .B2(n15823), .ZN(n15832) );
  NAND3_X1 U18812 ( .A1(n15826), .A2(n18814), .A3(n15825), .ZN(n15827) );
  OAI21_X1 U18813 ( .B1(n15828), .B2(n9935), .A(n15827), .ZN(n15829) );
  AOI21_X1 U18814 ( .B1(n15830), .B2(n18811), .A(n15829), .ZN(n15831) );
  OAI211_X1 U18815 ( .C1(n15834), .C2(n15833), .A(n15832), .B(n15831), .ZN(
        P2_U3011) );
  NOR2_X1 U18816 ( .A1(n12088), .A2(n18662), .ZN(n15837) );
  OAI22_X1 U18817 ( .A1(n15835), .A2(n15838), .B1(n18832), .B2(n18538), .ZN(
        n15836) );
  AOI211_X1 U18818 ( .C1(n15839), .C2(n15838), .A(n15837), .B(n15836), .ZN(
        n15843) );
  INV_X1 U18819 ( .A(n18539), .ZN(n15840) );
  AOI22_X1 U18820 ( .A1(n15841), .A2(n18846), .B1(n18853), .B2(n15840), .ZN(
        n15842) );
  OAI211_X1 U18821 ( .C1(n15926), .C2(n15844), .A(n15843), .B(n15842), .ZN(
        P2_U3027) );
  NOR2_X1 U18822 ( .A1(n12074), .A2(n18662), .ZN(n15849) );
  OAI21_X1 U18823 ( .B1(n15846), .B2(n9677), .A(n15845), .ZN(n18710) );
  OAI22_X1 U18824 ( .A1(n15847), .A2(n15850), .B1(n18832), .B2(n18710), .ZN(
        n15848) );
  AOI211_X1 U18825 ( .C1(n15851), .C2(n15850), .A(n15849), .B(n15848), .ZN(
        n15856) );
  INV_X1 U18826 ( .A(n15852), .ZN(n18585) );
  OAI22_X1 U18827 ( .A1(n15853), .A2(n18841), .B1(n15894), .B2(n18585), .ZN(
        n15854) );
  INV_X1 U18828 ( .A(n15854), .ZN(n15855) );
  OAI211_X1 U18829 ( .C1(n15926), .C2(n15857), .A(n15856), .B(n15855), .ZN(
        P2_U3031) );
  AOI211_X1 U18830 ( .C1(n15870), .C2(n15859), .A(n15858), .B(n15873), .ZN(
        n15862) );
  INV_X1 U18831 ( .A(n15860), .ZN(n18713) );
  OAI22_X1 U18832 ( .A1(n18832), .A2(n18713), .B1(n19506), .B2(n15908), .ZN(
        n15861) );
  NOR2_X1 U18833 ( .A1(n15862), .A2(n15861), .ZN(n15869) );
  INV_X1 U18834 ( .A(n15863), .ZN(n15865) );
  OAI22_X1 U18835 ( .A1(n15865), .A2(n18841), .B1(n15894), .B2(n15864), .ZN(
        n15866) );
  AOI21_X1 U18836 ( .B1(n18844), .B2(n15867), .A(n15866), .ZN(n15868) );
  OAI211_X1 U18837 ( .C1(n15872), .C2(n15870), .A(n15869), .B(n15868), .ZN(
        P2_U3032) );
  NAND2_X1 U18838 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18815), .ZN(n15871) );
  OAI221_X1 U18839 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15873), 
        .C1(n15770), .C2(n15872), .A(n15871), .ZN(n15874) );
  AOI21_X1 U18840 ( .B1(n18716), .B2(n18847), .A(n15874), .ZN(n15879) );
  INV_X1 U18841 ( .A(n15875), .ZN(n15876) );
  AOI22_X1 U18842 ( .A1(n15877), .A2(n18844), .B1(n18853), .B2(n15876), .ZN(
        n15878) );
  OAI211_X1 U18843 ( .C1(n18841), .C2(n15880), .A(n15879), .B(n15878), .ZN(
        P2_U3034) );
  NOR2_X1 U18844 ( .A1(n12029), .A2(n18662), .ZN(n15885) );
  XNOR2_X1 U18845 ( .A(n15882), .B(n15881), .ZN(n18724) );
  OAI22_X1 U18846 ( .A1(n15883), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18724), .B2(n18832), .ZN(n15884) );
  AOI211_X1 U18847 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n15886), .A(
        n15885), .B(n15884), .ZN(n15889) );
  AOI22_X1 U18848 ( .A1(n15887), .A2(n18846), .B1(n18853), .B2(n18618), .ZN(
        n15888) );
  OAI211_X1 U18849 ( .C1(n15890), .C2(n15926), .A(n15889), .B(n15888), .ZN(
        P2_U3036) );
  OAI21_X1 U18850 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15898), .A(
        n15891), .ZN(n15910) );
  AOI22_X1 U18851 ( .A1(n15910), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n18847), .B2(n18727), .ZN(n15904) );
  INV_X1 U18852 ( .A(n15892), .ZN(n15895) );
  OAI22_X1 U18853 ( .A1(n15895), .A2(n18841), .B1(n15894), .B2(n15893), .ZN(
        n15896) );
  AOI21_X1 U18854 ( .B1(n18844), .B2(n15897), .A(n15896), .ZN(n15903) );
  NAND2_X1 U18855 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18815), .ZN(n15902) );
  INV_X1 U18856 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15900) );
  NOR2_X1 U18857 ( .A1(n15899), .A2(n15898), .ZN(n15912) );
  OAI221_X1 U18858 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15900), .C2(n15911), .A(
        n15912), .ZN(n15901) );
  NAND4_X1 U18859 ( .A1(n15904), .A2(n15903), .A3(n15902), .A4(n15901), .ZN(
        P2_U3038) );
  OAI21_X1 U18860 ( .B1(n15907), .B2(n15906), .A(n15905), .ZN(n18730) );
  OAI22_X1 U18861 ( .A1(n18832), .A2(n18730), .B1(n19497), .B2(n15908), .ZN(
        n15909) );
  AOI221_X1 U18862 ( .B1(n15912), .B2(n15911), .C1(n15910), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15909), .ZN(n15916) );
  INV_X1 U18863 ( .A(n18642), .ZN(n15913) );
  AOI22_X1 U18864 ( .A1(n15914), .A2(n18844), .B1(n18853), .B2(n15913), .ZN(
        n15915) );
  OAI211_X1 U18865 ( .C1(n18841), .C2(n15917), .A(n15916), .B(n15915), .ZN(
        P2_U3039) );
  NAND2_X1 U18866 ( .A1(n18853), .A2(n18690), .ZN(n15918) );
  OAI21_X1 U18867 ( .B1(n18851), .B2(n12207), .A(n15918), .ZN(n15922) );
  INV_X1 U18868 ( .A(n18683), .ZN(n15919) );
  OAI22_X1 U18869 ( .A1(n18841), .A2(n15920), .B1(n18832), .B2(n15919), .ZN(
        n15921) );
  AOI211_X1 U18870 ( .C1(n12207), .C2(n18854), .A(n15922), .B(n15921), .ZN(
        n15924) );
  OAI211_X1 U18871 ( .C1(n15926), .C2(n15925), .A(n15924), .B(n15923), .ZN(
        P2_U3046) );
  INV_X1 U18872 ( .A(n15927), .ZN(n15928) );
  OAI211_X1 U18873 ( .C1(n15929), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15928), .ZN(n15931) );
  NAND2_X1 U18874 ( .A1(n15929), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15930) );
  NAND2_X1 U18875 ( .A1(n15931), .A2(n15930), .ZN(n15932) );
  NOR2_X1 U18876 ( .A1(n15958), .A2(n15932), .ZN(n15937) );
  MUX2_X1 U18877 ( .A(n15933), .B(n10776), .S(n15958), .Z(n15954) );
  INV_X1 U18878 ( .A(n15937), .ZN(n15935) );
  MUX2_X1 U18879 ( .A(n15939), .B(n15934), .S(n15958), .Z(n15955) );
  OAI221_X1 U18880 ( .B1(n15954), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .C1(n15954), .C2(n15935), .A(n15955), .ZN(n15936) );
  AOI22_X1 U18881 ( .A1(n15937), .A2(n19560), .B1(n19554), .B2(n15936), .ZN(
        n15938) );
  AOI211_X1 U18882 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n15939), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n15938), .ZN(n15957) );
  OR2_X1 U18883 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n15951) );
  NAND2_X1 U18884 ( .A1(n13275), .A2(n15940), .ZN(n15942) );
  OAI22_X1 U18885 ( .A1(n10815), .A2(n15942), .B1(n18868), .B2(n15941), .ZN(
        n15950) );
  INV_X1 U18886 ( .A(n15943), .ZN(n15949) );
  AOI22_X1 U18887 ( .A1(n15949), .A2(n15946), .B1(n15945), .B2(n15944), .ZN(
        n15947) );
  OAI21_X1 U18888 ( .B1(n15949), .B2(n15948), .A(n15947), .ZN(n19586) );
  AOI211_X1 U18889 ( .C1(n15952), .C2(n15951), .A(n15950), .B(n19586), .ZN(
        n15953) );
  OAI21_X1 U18890 ( .B1(n15955), .B2(n15954), .A(n15953), .ZN(n15956) );
  AOI211_X1 U18891 ( .C1(n15958), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n15957), .B(n15956), .ZN(n15972) );
  AOI211_X1 U18892 ( .C1(n15962), .C2(n15961), .A(n15960), .B(n15959), .ZN(
        n15971) );
  INV_X1 U18893 ( .A(n19599), .ZN(n15963) );
  NOR3_X1 U18894 ( .A1(n15964), .A2(n15963), .A3(n18921), .ZN(n15966) );
  OAI221_X1 U18895 ( .B1(n15967), .B2(n15972), .C1(n15967), .C2(n20564), .A(
        n15966), .ZN(n19464) );
  INV_X1 U18896 ( .A(n19464), .ZN(n15969) );
  INV_X1 U18897 ( .A(n19602), .ZN(n19595) );
  AOI22_X1 U18898 ( .A1(n19595), .A2(n15966), .B1(n19596), .B2(n15965), .ZN(
        n15968) );
  AOI22_X1 U18899 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15969), .B1(n15968), 
        .B2(n15967), .ZN(n15970) );
  OAI211_X1 U18900 ( .C1(n15972), .C2(n19458), .A(n15971), .B(n15970), .ZN(
        P2_U3176) );
  OAI21_X1 U18901 ( .B1(n19571), .B2(n19464), .A(n15973), .ZN(P2_U3593) );
  NOR2_X2 U18902 ( .A1(n17834), .A2(n16152), .ZN(n17481) );
  NOR2_X1 U18903 ( .A1(n17388), .A2(n15975), .ZN(n15983) );
  NAND2_X1 U18904 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17388), .ZN(
        n15978) );
  OAI211_X1 U18905 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17388), .A(
        n15976), .B(n15978), .ZN(n15982) );
  OAI21_X1 U18906 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16027), .A(
        n15977), .ZN(n15980) );
  OAI22_X1 U18907 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17388), .B1(
        n15978), .B2(n16027), .ZN(n15979) );
  OAI21_X1 U18908 ( .B1(n15983), .B2(n15980), .A(n15979), .ZN(n15981) );
  OAI21_X1 U18909 ( .B1(n15983), .B2(n15982), .A(n15981), .ZN(n16033) );
  INV_X1 U18910 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16174) );
  NAND2_X1 U18911 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17394) );
  NAND3_X1 U18912 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16365) );
  NOR2_X1 U18913 ( .A1(n17394), .A2(n16365), .ZN(n17306) );
  NAND2_X1 U18914 ( .A1(n17391), .A2(n17306), .ZN(n17321) );
  NAND2_X1 U18915 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17323) );
  NAND2_X1 U18916 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17200) );
  NAND2_X1 U18917 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17195), .ZN(
        n17156) );
  NAND2_X1 U18918 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17157) );
  NAND2_X1 U18919 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17126) );
  NAND2_X1 U18920 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16008), .ZN(
        n15984) );
  NAND2_X1 U18921 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16010), .ZN(
        n15998) );
  INV_X1 U18922 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18406) );
  NOR2_X1 U18923 ( .A1(n18406), .A2(n17712), .ZN(n16024) );
  INV_X1 U18924 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16198) );
  INV_X1 U18925 ( .A(n15984), .ZN(n15987) );
  NAND2_X1 U18926 ( .A1(n18475), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18334) );
  AOI21_X1 U18927 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n15985), .A(
        n18205), .ZN(n17322) );
  INV_X1 U18928 ( .A(n17322), .ZN(n17279) );
  NAND2_X1 U18929 ( .A1(n15987), .A2(n17279), .ZN(n16000) );
  NOR2_X1 U18930 ( .A1(n16198), .A2(n16000), .ZN(n15991) );
  NOR2_X1 U18931 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17267), .ZN(
        n16012) );
  NOR2_X1 U18932 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16000), .ZN(
        n15989) );
  NOR2_X1 U18933 ( .A1(n17484), .A2(n17125), .ZN(n16181) );
  INV_X1 U18934 ( .A(n16181), .ZN(n16190) );
  OR2_X1 U18935 ( .A1(n16190), .A2(n17126), .ZN(n16191) );
  INV_X1 U18936 ( .A(n18334), .ZN(n17240) );
  INV_X1 U18937 ( .A(n15986), .ZN(n18019) );
  NOR2_X1 U18938 ( .A1(n18019), .A2(n15987), .ZN(n16007) );
  AOI211_X1 U18939 ( .C1(n16191), .C2(n17240), .A(n17457), .B(n16007), .ZN(
        n15988) );
  INV_X1 U18940 ( .A(n15988), .ZN(n16009) );
  NOR3_X1 U18941 ( .A1(n16012), .A2(n15989), .A3(n16009), .ZN(n15999) );
  INV_X1 U18942 ( .A(n15999), .ZN(n15990) );
  MUX2_X1 U18943 ( .A(n15991), .B(n15990), .S(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n15992) );
  AOI211_X1 U18944 ( .C1(n17285), .C2(n9609), .A(n16024), .B(n15992), .ZN(
        n15997) );
  INV_X1 U18945 ( .A(n15993), .ZN(n16003) );
  NAND2_X1 U18946 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16003), .ZN(
        n15994) );
  INV_X1 U18947 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18431) );
  XOR2_X1 U18948 ( .A(n15994), .B(n18431), .Z(n16025) );
  NAND2_X1 U18949 ( .A1(n17646), .A2(n17481), .ZN(n17117) );
  NAND2_X1 U18950 ( .A1(n16002), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15995) );
  XOR2_X1 U18951 ( .A(n15995), .B(n18431), .Z(n16029) );
  AOI22_X1 U18952 ( .A1(n9601), .A2(n16025), .B1(n17399), .B2(n16029), .ZN(
        n15996) );
  OAI211_X1 U18953 ( .C1(n17402), .C2(n16033), .A(n15997), .B(n15996), .ZN(
        P3_U2799) );
  OAI21_X1 U18954 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16010), .A(
        n15998), .ZN(n16196) );
  AOI21_X1 U18955 ( .B1(n16198), .B2(n16000), .A(n15999), .ZN(n16001) );
  AOI21_X1 U18956 ( .B1(P3_REIP_REG_30__SCAN_IN), .B2(n9597), .A(n16001), .ZN(
        n16006) );
  NOR2_X1 U18957 ( .A1(n16002), .A2(n17117), .ZN(n16015) );
  NOR2_X1 U18958 ( .A1(n16003), .A2(n17492), .ZN(n16017) );
  NAND2_X1 U18959 ( .A1(n16035), .A2(n17212), .ZN(n17141) );
  AOI22_X1 U18960 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16009), .B1(
        n16008), .B2(n16007), .ZN(n16021) );
  INV_X1 U18961 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16215) );
  AOI21_X1 U18962 ( .B1(n16215), .B2(n16191), .A(n16010), .ZN(n16209) );
  INV_X1 U18963 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18404) );
  NOR2_X1 U18964 ( .A1(n17712), .A2(n18404), .ZN(n16011) );
  AOI221_X1 U18965 ( .B1(n16012), .B2(n16209), .C1(n17285), .C2(n16209), .A(
        n16011), .ZN(n16020) );
  OAI21_X1 U18966 ( .B1(n16039), .B2(n17116), .A(n16013), .ZN(n16014) );
  AOI22_X1 U18967 ( .A1(n17342), .A2(n16016), .B1(n16015), .B2(n16014), .ZN(
        n16019) );
  OAI21_X1 U18968 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16042), .A(
        n16017), .ZN(n16018) );
  NAND4_X1 U18969 ( .A1(n16021), .A2(n16020), .A3(n16019), .A4(n16018), .ZN(
        P3_U2801) );
  NOR2_X1 U18970 ( .A1(n17804), .A2(n17722), .ZN(n17762) );
  INV_X1 U18971 ( .A(n17762), .ZN(n17796) );
  AOI221_X1 U18972 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16022), 
        .C1(n17796), .C2(n16022), .A(n18431), .ZN(n16023) );
  AOI211_X1 U18973 ( .C1(n16025), .C2(n17809), .A(n16024), .B(n16023), .ZN(
        n16032) );
  NOR4_X1 U18974 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16028), .A3(
        n16027), .A4(n16026), .ZN(n16030) );
  OAI221_X1 U18975 ( .B1(n16030), .B2(n16029), .C1(n16030), .C2(n17725), .A(
        n17793), .ZN(n16031) );
  OAI211_X1 U18976 ( .C1(n16033), .C2(n17727), .A(n16032), .B(n16031), .ZN(
        P3_U2831) );
  INV_X1 U18977 ( .A(n18264), .ZN(n17789) );
  OAI22_X1 U18978 ( .A1(n17691), .A2(n17789), .B1(n17688), .B2(n17356), .ZN(
        n17593) );
  AOI21_X1 U18979 ( .B1(n17594), .B2(n17593), .A(n16034), .ZN(n17546) );
  NOR2_X1 U18980 ( .A1(n17546), .A2(n17804), .ZN(n17567) );
  INV_X1 U18981 ( .A(n16035), .ZN(n17493) );
  NOR3_X1 U18982 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n9925), .A3(
        n17493), .ZN(n17124) );
  AOI22_X1 U18983 ( .A1(n9597), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17567), 
        .B2(n17124), .ZN(n16048) );
  NAND3_X1 U18984 ( .A1(n17132), .A2(n17811), .A3(n16036), .ZN(n16047) );
  AOI22_X1 U18985 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17359), .B1(
        n17388), .B2(n17118), .ZN(n17121) );
  NAND3_X1 U18986 ( .A1(n17131), .A2(n17681), .A3(n17121), .ZN(n16046) );
  AOI21_X1 U18987 ( .B1(n17388), .B2(n16037), .A(n17131), .ZN(n17120) );
  NOR2_X1 U18988 ( .A1(n17121), .A2(n17120), .ZN(n17119) );
  NOR4_X1 U18989 ( .A1(n17646), .A2(n16038), .A3(n17119), .A4(n18261), .ZN(
        n16044) );
  OAI21_X1 U18990 ( .B1(n16039), .B2(n17116), .A(n17725), .ZN(n16040) );
  OAI211_X1 U18991 ( .C1(n16042), .C2(n17789), .A(n16041), .B(n16040), .ZN(
        n16043) );
  OAI211_X1 U18992 ( .C1(n16044), .C2(n16043), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17712), .ZN(n16045) );
  NOR3_X1 U18993 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16050) );
  NOR4_X1 U18994 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16049) );
  NAND4_X1 U18995 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16050), .A3(n16049), .A4(
        U215), .ZN(U213) );
  INV_X1 U18996 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16140) );
  INV_X2 U18997 ( .A(U214), .ZN(n16103) );
  NOR2_X1 U18998 ( .A1(n16103), .A2(n16051), .ZN(n16087) );
  INV_X1 U18999 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20599) );
  OAI222_X1 U19000 ( .A1(U212), .A2(n16140), .B1(n16105), .B2(n18910), .C1(
        U214), .C2(n20599), .ZN(U216) );
  INV_X1 U19001 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16053) );
  INV_X2 U19002 ( .A(U212), .ZN(n16102) );
  AOI22_X1 U19003 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16102), .ZN(n16052) );
  OAI21_X1 U19004 ( .B1(n16053), .B2(n16105), .A(n16052), .ZN(U217) );
  AOI222_X1 U19005 ( .A1(n16102), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n16087), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n16103), .C2(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n16054) );
  INV_X1 U19006 ( .A(n16054), .ZN(U218) );
  INV_X1 U19007 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20584) );
  AOI22_X1 U19008 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16102), .ZN(n16055) );
  OAI21_X1 U19009 ( .B1(n20584), .B2(n16105), .A(n16055), .ZN(U219) );
  INV_X1 U19010 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16057) );
  AOI22_X1 U19011 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16102), .ZN(n16056) );
  OAI21_X1 U19012 ( .B1(n16057), .B2(n16105), .A(n16056), .ZN(U220) );
  INV_X1 U19013 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16059) );
  AOI22_X1 U19014 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16102), .ZN(n16058) );
  OAI21_X1 U19015 ( .B1(n16059), .B2(n16105), .A(n16058), .ZN(U221) );
  INV_X1 U19016 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16061) );
  AOI22_X1 U19017 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16102), .ZN(n16060) );
  OAI21_X1 U19018 ( .B1(n16061), .B2(n16105), .A(n16060), .ZN(U222) );
  AOI222_X1 U19019 ( .A1(n16102), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(n16087), 
        .B2(BUF1_REG_24__SCAN_IN), .C1(n16103), .C2(P1_DATAO_REG_24__SCAN_IN), 
        .ZN(n16062) );
  INV_X1 U19020 ( .A(n16062), .ZN(U223) );
  AOI22_X1 U19021 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16102), .ZN(n16063) );
  OAI21_X1 U19022 ( .B1(n16064), .B2(n16105), .A(n16063), .ZN(U224) );
  INV_X1 U19023 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16066) );
  AOI22_X1 U19024 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16102), .ZN(n16065) );
  OAI21_X1 U19025 ( .B1(n16066), .B2(n16105), .A(n16065), .ZN(U225) );
  INV_X1 U19026 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16068) );
  AOI22_X1 U19027 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16102), .ZN(n16067) );
  OAI21_X1 U19028 ( .B1(n16068), .B2(n16105), .A(n16067), .ZN(U226) );
  AOI22_X1 U19029 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16102), .ZN(n16069) );
  OAI21_X1 U19030 ( .B1(n13737), .B2(n16105), .A(n16069), .ZN(U227) );
  INV_X1 U19031 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16071) );
  AOI22_X1 U19032 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16102), .ZN(n16070) );
  OAI21_X1 U19033 ( .B1(n16071), .B2(n16105), .A(n16070), .ZN(U228) );
  AOI22_X1 U19034 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16102), .ZN(n16072) );
  OAI21_X1 U19035 ( .B1(n13745), .B2(n16105), .A(n16072), .ZN(U229) );
  INV_X1 U19036 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U19037 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16102), .ZN(n16073) );
  OAI21_X1 U19038 ( .B1(n16074), .B2(n16105), .A(n16073), .ZN(U230) );
  INV_X1 U19039 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16076) );
  AOI22_X1 U19040 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16102), .ZN(n16075) );
  OAI21_X1 U19041 ( .B1(n16076), .B2(n16105), .A(n16075), .ZN(U231) );
  AOI22_X1 U19042 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16102), .ZN(n16077) );
  OAI21_X1 U19043 ( .B1(n12372), .B2(n16105), .A(n16077), .ZN(U232) );
  INV_X1 U19044 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16079) );
  AOI22_X1 U19045 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16102), .ZN(n16078) );
  OAI21_X1 U19046 ( .B1(n16079), .B2(n16105), .A(n16078), .ZN(U233) );
  AOI22_X1 U19047 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16102), .ZN(n16080) );
  OAI21_X1 U19048 ( .B1(n12180), .B2(n16105), .A(n16080), .ZN(U234) );
  INV_X1 U19049 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16082) );
  AOI22_X1 U19050 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16102), .ZN(n16081) );
  OAI21_X1 U19051 ( .B1(n16082), .B2(n16105), .A(n16081), .ZN(U235) );
  AOI22_X1 U19052 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16102), .ZN(n16083) );
  OAI21_X1 U19053 ( .B1(n12176), .B2(n16105), .A(n16083), .ZN(U236) );
  AOI22_X1 U19054 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16102), .ZN(n16084) );
  OAI21_X1 U19055 ( .B1(n16085), .B2(n16105), .A(n16084), .ZN(U237) );
  AOI22_X1 U19056 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16102), .ZN(n16086) );
  OAI21_X1 U19057 ( .B1(n12185), .B2(n16105), .A(n16086), .ZN(U238) );
  AOI222_X1 U19058 ( .A1(n16102), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n16087), 
        .B2(BUF1_REG_8__SCAN_IN), .C1(n16103), .C2(P1_DATAO_REG_8__SCAN_IN), 
        .ZN(n16088) );
  INV_X1 U19059 ( .A(n16088), .ZN(U239) );
  INV_X1 U19060 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U19061 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16102), .ZN(n16089) );
  OAI21_X1 U19062 ( .B1(n16090), .B2(n16105), .A(n16089), .ZN(U240) );
  INV_X1 U19063 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16092) );
  AOI22_X1 U19064 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16102), .ZN(n16091) );
  OAI21_X1 U19065 ( .B1(n16092), .B2(n16105), .A(n16091), .ZN(U241) );
  INV_X1 U19066 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20637) );
  AOI22_X1 U19067 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16102), .ZN(n16093) );
  OAI21_X1 U19068 ( .B1(n20637), .B2(n16105), .A(n16093), .ZN(U242) );
  INV_X1 U19069 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16095) );
  AOI22_X1 U19070 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16102), .ZN(n16094) );
  OAI21_X1 U19071 ( .B1(n16095), .B2(n16105), .A(n16094), .ZN(U243) );
  INV_X1 U19072 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16097) );
  AOI22_X1 U19073 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16102), .ZN(n16096) );
  OAI21_X1 U19074 ( .B1(n16097), .B2(n16105), .A(n16096), .ZN(U244) );
  INV_X1 U19075 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16099) );
  AOI22_X1 U19076 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16102), .ZN(n16098) );
  OAI21_X1 U19077 ( .B1(n16099), .B2(n16105), .A(n16098), .ZN(U245) );
  INV_X1 U19078 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19079 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16102), .ZN(n16100) );
  OAI21_X1 U19080 ( .B1(n16101), .B2(n16105), .A(n16100), .ZN(U246) );
  INV_X1 U19081 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U19082 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16103), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16102), .ZN(n16104) );
  OAI21_X1 U19083 ( .B1(n16106), .B2(n16105), .A(n16104), .ZN(U247) );
  OAI22_X1 U19084 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16138), .ZN(n16107) );
  INV_X1 U19085 ( .A(n16107), .ZN(U251) );
  OAI22_X1 U19086 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16138), .ZN(n16108) );
  INV_X1 U19087 ( .A(n16108), .ZN(U252) );
  OAI22_X1 U19088 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16138), .ZN(n16109) );
  INV_X1 U19089 ( .A(n16109), .ZN(U253) );
  OAI22_X1 U19090 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16138), .ZN(n16110) );
  INV_X1 U19091 ( .A(n16110), .ZN(U254) );
  OAI22_X1 U19092 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16138), .ZN(n16111) );
  INV_X1 U19093 ( .A(n16111), .ZN(U255) );
  OAI22_X1 U19094 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16138), .ZN(n16112) );
  INV_X1 U19095 ( .A(n16112), .ZN(U256) );
  OAI22_X1 U19096 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16138), .ZN(n16113) );
  INV_X1 U19097 ( .A(n16113), .ZN(U257) );
  OAI22_X1 U19098 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16138), .ZN(n16114) );
  INV_X1 U19099 ( .A(n16114), .ZN(U258) );
  OAI22_X1 U19100 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16138), .ZN(n16115) );
  INV_X1 U19101 ( .A(n16115), .ZN(U259) );
  OAI22_X1 U19102 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16130), .ZN(n16116) );
  INV_X1 U19103 ( .A(n16116), .ZN(U260) );
  OAI22_X1 U19104 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16130), .ZN(n16117) );
  INV_X1 U19105 ( .A(n16117), .ZN(U261) );
  OAI22_X1 U19106 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16138), .ZN(n16118) );
  INV_X1 U19107 ( .A(n16118), .ZN(U262) );
  OAI22_X1 U19108 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16130), .ZN(n16119) );
  INV_X1 U19109 ( .A(n16119), .ZN(U263) );
  OAI22_X1 U19110 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16138), .ZN(n16120) );
  INV_X1 U19111 ( .A(n16120), .ZN(U264) );
  OAI22_X1 U19112 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16138), .ZN(n16121) );
  INV_X1 U19113 ( .A(n16121), .ZN(U265) );
  OAI22_X1 U19114 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16130), .ZN(n16122) );
  INV_X1 U19115 ( .A(n16122), .ZN(U266) );
  OAI22_X1 U19116 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16130), .ZN(n16123) );
  INV_X1 U19117 ( .A(n16123), .ZN(U267) );
  OAI22_X1 U19118 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16130), .ZN(n16124) );
  INV_X1 U19119 ( .A(n16124), .ZN(U268) );
  OAI22_X1 U19120 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16130), .ZN(n16125) );
  INV_X1 U19121 ( .A(n16125), .ZN(U269) );
  OAI22_X1 U19122 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16130), .ZN(n16126) );
  INV_X1 U19123 ( .A(n16126), .ZN(U270) );
  OAI22_X1 U19124 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16130), .ZN(n16127) );
  INV_X1 U19125 ( .A(n16127), .ZN(U271) );
  OAI22_X1 U19126 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16138), .ZN(n16128) );
  INV_X1 U19127 ( .A(n16128), .ZN(U272) );
  OAI22_X1 U19128 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16138), .ZN(n16129) );
  INV_X1 U19129 ( .A(n16129), .ZN(U273) );
  OAI22_X1 U19130 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16130), .ZN(n16131) );
  INV_X1 U19131 ( .A(n16131), .ZN(U274) );
  OAI22_X1 U19132 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16138), .ZN(n16132) );
  INV_X1 U19133 ( .A(n16132), .ZN(U275) );
  OAI22_X1 U19134 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16138), .ZN(n16133) );
  INV_X1 U19135 ( .A(n16133), .ZN(U276) );
  OAI22_X1 U19136 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16138), .ZN(n16134) );
  INV_X1 U19137 ( .A(n16134), .ZN(U277) );
  OAI22_X1 U19138 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16138), .ZN(n16135) );
  INV_X1 U19139 ( .A(n16135), .ZN(U278) );
  OAI22_X1 U19140 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16138), .ZN(n16136) );
  INV_X1 U19141 ( .A(n16136), .ZN(U279) );
  INV_X1 U19142 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n20591) );
  INV_X1 U19143 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18895) );
  AOI22_X1 U19144 ( .A1(n16138), .A2(n20591), .B1(n18895), .B2(U215), .ZN(U280) );
  OAI22_X1 U19145 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16138), .ZN(n16137) );
  INV_X1 U19146 ( .A(n16137), .ZN(U281) );
  INV_X1 U19147 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18908) );
  AOI22_X1 U19148 ( .A1(n16138), .A2(n16140), .B1(n18908), .B2(U215), .ZN(U282) );
  INV_X1 U19149 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16139) );
  AOI222_X1 U19150 ( .A1(n20599), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16140), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16139), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16141) );
  INV_X2 U19151 ( .A(n16143), .ZN(n16142) );
  INV_X1 U19152 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18368) );
  INV_X1 U19153 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19501) );
  AOI22_X1 U19154 ( .A1(n16142), .A2(n18368), .B1(n19501), .B2(n16143), .ZN(
        U347) );
  INV_X1 U19155 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18366) );
  INV_X1 U19156 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19500) );
  AOI22_X1 U19157 ( .A1(n16142), .A2(n18366), .B1(n19500), .B2(n16143), .ZN(
        U348) );
  INV_X1 U19158 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18364) );
  INV_X1 U19159 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U19160 ( .A1(n16142), .A2(n18364), .B1(n20555), .B2(n16143), .ZN(
        U349) );
  INV_X1 U19161 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18363) );
  AOI22_X1 U19162 ( .A1(n16142), .A2(n18363), .B1(n20544), .B2(n16143), .ZN(
        U350) );
  INV_X1 U19163 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18361) );
  INV_X1 U19164 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19496) );
  AOI22_X1 U19165 ( .A1(n16142), .A2(n18361), .B1(n19496), .B2(n16143), .ZN(
        U351) );
  INV_X1 U19166 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18358) );
  INV_X1 U19167 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19494) );
  AOI22_X1 U19168 ( .A1(n16142), .A2(n18358), .B1(n19494), .B2(n16143), .ZN(
        U352) );
  INV_X1 U19169 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18357) );
  INV_X1 U19170 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19492) );
  AOI22_X1 U19171 ( .A1(n16142), .A2(n18357), .B1(n19492), .B2(n16143), .ZN(
        U353) );
  INV_X1 U19172 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18354) );
  INV_X1 U19173 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19490) );
  AOI22_X1 U19174 ( .A1(n16142), .A2(n18354), .B1(n19490), .B2(n16143), .ZN(
        U354) );
  INV_X1 U19175 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18407) );
  INV_X1 U19176 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19532) );
  AOI22_X1 U19177 ( .A1(n16142), .A2(n18407), .B1(n19532), .B2(n16143), .ZN(
        U355) );
  INV_X1 U19178 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18405) );
  INV_X1 U19179 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19530) );
  AOI22_X1 U19180 ( .A1(n16142), .A2(n18405), .B1(n19530), .B2(n16143), .ZN(
        U356) );
  INV_X1 U19181 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18402) );
  INV_X1 U19182 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U19183 ( .A1(n16142), .A2(n18402), .B1(n19528), .B2(n16143), .ZN(
        U357) );
  INV_X1 U19184 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18401) );
  INV_X1 U19185 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19526) );
  AOI22_X1 U19186 ( .A1(n16142), .A2(n18401), .B1(n19526), .B2(n16143), .ZN(
        U358) );
  INV_X1 U19187 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18399) );
  INV_X1 U19188 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19525) );
  AOI22_X1 U19189 ( .A1(n16142), .A2(n18399), .B1(n19525), .B2(n16143), .ZN(
        U359) );
  INV_X1 U19190 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18397) );
  INV_X1 U19191 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19523) );
  AOI22_X1 U19192 ( .A1(n16142), .A2(n18397), .B1(n19523), .B2(n16143), .ZN(
        U360) );
  INV_X1 U19193 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18394) );
  INV_X1 U19194 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19521) );
  AOI22_X1 U19195 ( .A1(n16142), .A2(n18394), .B1(n19521), .B2(n16143), .ZN(
        U361) );
  INV_X1 U19196 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18392) );
  INV_X1 U19197 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19520) );
  AOI22_X1 U19198 ( .A1(n16142), .A2(n18392), .B1(n19520), .B2(n16143), .ZN(
        U362) );
  INV_X1 U19199 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18391) );
  INV_X1 U19200 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19519) );
  AOI22_X1 U19201 ( .A1(n16142), .A2(n18391), .B1(n19519), .B2(n16143), .ZN(
        U363) );
  INV_X1 U19202 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18389) );
  INV_X1 U19203 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19518) );
  AOI22_X1 U19204 ( .A1(n16142), .A2(n18389), .B1(n19518), .B2(n16143), .ZN(
        U364) );
  INV_X1 U19205 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18352) );
  AOI22_X1 U19206 ( .A1(n16142), .A2(n18352), .B1(n20527), .B2(n16143), .ZN(
        U365) );
  INV_X1 U19207 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18386) );
  INV_X1 U19208 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19516) );
  AOI22_X1 U19209 ( .A1(n16142), .A2(n18386), .B1(n19516), .B2(n16143), .ZN(
        U366) );
  INV_X1 U19210 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18385) );
  INV_X1 U19211 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19514) );
  AOI22_X1 U19212 ( .A1(n16142), .A2(n18385), .B1(n19514), .B2(n16143), .ZN(
        U367) );
  INV_X1 U19213 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20576) );
  INV_X1 U19214 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19513) );
  AOI22_X1 U19215 ( .A1(n16142), .A2(n20576), .B1(n19513), .B2(n16143), .ZN(
        U368) );
  INV_X1 U19216 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18382) );
  INV_X1 U19217 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19511) );
  AOI22_X1 U19218 ( .A1(n16142), .A2(n18382), .B1(n19511), .B2(n16143), .ZN(
        U369) );
  INV_X1 U19219 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18380) );
  INV_X1 U19220 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19509) );
  AOI22_X1 U19221 ( .A1(n16142), .A2(n18380), .B1(n19509), .B2(n16143), .ZN(
        U370) );
  INV_X1 U19222 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18378) );
  INV_X1 U19223 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19508) );
  AOI22_X1 U19224 ( .A1(n16142), .A2(n18378), .B1(n19508), .B2(n16143), .ZN(
        U371) );
  INV_X1 U19225 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18375) );
  INV_X1 U19226 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19507) );
  AOI22_X1 U19227 ( .A1(n16142), .A2(n18375), .B1(n19507), .B2(n16143), .ZN(
        U372) );
  INV_X1 U19228 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18374) );
  INV_X1 U19229 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19505) );
  AOI22_X1 U19230 ( .A1(n16142), .A2(n18374), .B1(n19505), .B2(n16143), .ZN(
        U373) );
  INV_X1 U19231 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18372) );
  INV_X1 U19232 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19504) );
  AOI22_X1 U19233 ( .A1(n16142), .A2(n18372), .B1(n19504), .B2(n16143), .ZN(
        U374) );
  INV_X1 U19234 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18370) );
  INV_X1 U19235 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19503) );
  AOI22_X1 U19236 ( .A1(n16142), .A2(n18370), .B1(n19503), .B2(n16143), .ZN(
        U375) );
  INV_X1 U19237 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18350) );
  INV_X1 U19238 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19487) );
  AOI22_X1 U19239 ( .A1(n16142), .A2(n18350), .B1(n19487), .B2(n16143), .ZN(
        U376) );
  INV_X1 U19240 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18349) );
  NAND2_X1 U19241 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18349), .ZN(n18339) );
  AOI22_X1 U19242 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18339), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18347), .ZN(n18416) );
  AOI21_X1 U19243 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18416), .ZN(n16144) );
  INV_X1 U19244 ( .A(n16144), .ZN(P3_U2633) );
  INV_X1 U19245 ( .A(n18326), .ZN(n16171) );
  AND2_X1 U19246 ( .A1(n17063), .A2(n16151), .ZN(n16145) );
  OAI21_X1 U19247 ( .B1(n16145), .B2(n17062), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16146) );
  OAI21_X1 U19248 ( .B1(n16147), .B2(n16171), .A(n16146), .ZN(P3_U2634) );
  AOI21_X1 U19249 ( .B1(n18347), .B2(n18349), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16148) );
  AOI22_X1 U19250 ( .A1(n18482), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16148), 
        .B2(n18483), .ZN(P3_U2635) );
  OAI21_X1 U19251 ( .B1(n18336), .B2(BS16), .A(n18416), .ZN(n18414) );
  OAI21_X1 U19252 ( .B1(n18416), .B2(n16170), .A(n18414), .ZN(P3_U2636) );
  AOI211_X1 U19253 ( .C1(n17063), .C2(n16151), .A(n16150), .B(n16149), .ZN(
        n18311) );
  NOR2_X1 U19254 ( .A1(n18311), .A2(n18315), .ZN(n18462) );
  OAI21_X1 U19255 ( .B1(n18462), .B2(n16153), .A(n16152), .ZN(P3_U2637) );
  NOR4_X1 U19256 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16157) );
  NOR4_X1 U19257 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16156) );
  NOR4_X1 U19258 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16155) );
  NOR4_X1 U19259 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16154) );
  NAND4_X1 U19260 ( .A1(n16157), .A2(n16156), .A3(n16155), .A4(n16154), .ZN(
        n16163) );
  NOR4_X1 U19261 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16161) );
  AOI211_X1 U19262 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16160) );
  NOR4_X1 U19263 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16159) );
  NOR4_X1 U19264 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16158) );
  NAND4_X1 U19265 ( .A1(n16161), .A2(n16160), .A3(n16159), .A4(n16158), .ZN(
        n16162) );
  NOR2_X1 U19266 ( .A1(n16163), .A2(n16162), .ZN(n18456) );
  INV_X1 U19267 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16165) );
  NOR3_X1 U19268 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16166) );
  OAI21_X1 U19269 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16166), .A(n18456), .ZN(
        n16164) );
  OAI21_X1 U19270 ( .B1(n18456), .B2(n16165), .A(n16164), .ZN(P3_U2638) );
  INV_X1 U19271 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18452) );
  INV_X1 U19272 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18415) );
  AOI21_X1 U19273 ( .B1(n18452), .B2(n18415), .A(n16166), .ZN(n16168) );
  INV_X1 U19274 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16167) );
  INV_X1 U19275 ( .A(n18456), .ZN(n18459) );
  AOI22_X1 U19276 ( .A1(n18456), .A2(n16168), .B1(n16167), .B2(n18459), .ZN(
        P3_U2639) );
  INV_X1 U19277 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16551) );
  NOR3_X1 U19278 ( .A1(n16551), .A2(n17834), .A3(n17831), .ZN(n16173) );
  OAI211_X2 U19279 ( .C1(P3_STATEBS16_REG_SCAN_IN), .C2(n18473), .A(n18488), 
        .B(n16173), .ZN(n16539) );
  NOR2_X1 U19280 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16539), .ZN(n16177) );
  NOR2_X1 U19281 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16524) );
  NAND2_X1 U19282 ( .A1(n16524), .A2(n16520), .ZN(n16519) );
  NOR2_X1 U19283 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16519), .ZN(n16498) );
  NAND2_X1 U19284 ( .A1(n16498), .A2(n16487), .ZN(n16486) );
  NAND2_X1 U19285 ( .A1(n16470), .A2(n20629), .ZN(n16456) );
  NAND2_X1 U19286 ( .A1(n16445), .A2(n16438), .ZN(n16437) );
  NAND2_X1 U19287 ( .A1(n16417), .A2(n16777), .ZN(n16413) );
  NAND2_X1 U19288 ( .A1(n16402), .A2(n16732), .ZN(n16392) );
  INV_X1 U19289 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16730) );
  NAND2_X1 U19290 ( .A1(n16374), .A2(n16730), .ZN(n16370) );
  INV_X1 U19291 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16345) );
  NAND2_X1 U19292 ( .A1(n16354), .A2(n16345), .ZN(n16344) );
  NAND2_X1 U19293 ( .A1(n16329), .A2(n16321), .ZN(n16320) );
  NAND2_X1 U19294 ( .A1(n16311), .A2(n16653), .ZN(n16303) );
  INV_X1 U19295 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16546) );
  NAND2_X1 U19296 ( .A1(n16292), .A2(n16546), .ZN(n16283) );
  NAND2_X1 U19297 ( .A1(n16268), .A2(n16549), .ZN(n16262) );
  NOR2_X1 U19298 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16262), .ZN(n16246) );
  INV_X1 U19299 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16241) );
  NAND2_X1 U19300 ( .A1(n16246), .A2(n16241), .ZN(n16240) );
  NOR2_X1 U19301 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16240), .ZN(n16229) );
  NAND2_X1 U19302 ( .A1(n16229), .A2(n16220), .ZN(n16219) );
  NOR2_X1 U19303 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16219), .ZN(n16206) );
  INV_X1 U19304 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18408) );
  NAND2_X1 U19305 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16221) );
  NOR2_X1 U19306 ( .A1(n18404), .A2(n16221), .ZN(n16180) );
  INV_X1 U19307 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18398) );
  OAI211_X1 U19308 ( .C1(n18471), .C2(n18472), .A(n18466), .B(n16170), .ZN(
        n16172) );
  INV_X1 U19309 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20587) );
  INV_X1 U19310 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18376) );
  INV_X1 U19311 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18373) );
  INV_X1 U19312 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18369) );
  INV_X1 U19313 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20608) );
  INV_X1 U19314 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18356) );
  NAND3_X1 U19315 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16480) );
  NOR2_X1 U19316 ( .A1(n18356), .A2(n16480), .ZN(n16475) );
  NAND2_X1 U19317 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16475), .ZN(n16432) );
  INV_X1 U19318 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18362) );
  INV_X1 U19319 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18360) );
  NOR2_X1 U19320 ( .A1(n18362), .A2(n18360), .ZN(n16447) );
  INV_X1 U19321 ( .A(n16447), .ZN(n16433) );
  NOR3_X1 U19322 ( .A1(n20608), .A2(n16432), .A3(n16433), .ZN(n16408) );
  NAND3_X1 U19323 ( .A1(n16408), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_9__SCAN_IN), .ZN(n16401) );
  NOR2_X1 U19324 ( .A1(n18369), .A2(n16401), .ZN(n16391) );
  NAND2_X1 U19325 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16391), .ZN(n16366) );
  NOR3_X1 U19326 ( .A1(n18376), .A2(n18373), .A3(n16366), .ZN(n16277) );
  INV_X1 U19327 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18390) );
  INV_X1 U19328 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18387) );
  INV_X1 U19329 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18381) );
  NAND2_X1 U19330 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16341) );
  NOR2_X1 U19331 ( .A1(n18381), .A2(n16341), .ZN(n16310) );
  NAND3_X1 U19332 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16310), .ZN(n16297) );
  NOR2_X1 U19333 ( .A1(n18387), .A2(n16297), .ZN(n16278) );
  NAND2_X1 U19334 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16278), .ZN(n16284) );
  NOR2_X1 U19335 ( .A1(n18390), .A2(n16284), .ZN(n16266) );
  NAND3_X1 U19336 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16277), .A3(n16266), 
        .ZN(n16259) );
  NOR2_X1 U19337 ( .A1(n20587), .A2(n16259), .ZN(n16245) );
  AND2_X1 U19338 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16245), .ZN(n16179) );
  NAND2_X1 U19339 ( .A1(n16530), .A2(n16179), .ZN(n16237) );
  NOR2_X1 U19340 ( .A1(n18398), .A2(n16237), .ZN(n16232) );
  NAND2_X1 U19341 ( .A1(n16180), .A2(n16232), .ZN(n16178) );
  NOR3_X1 U19342 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18408), .A3(n16178), 
        .ZN(n16176) );
  INV_X1 U19343 ( .A(n18166), .ZN(n18324) );
  NOR2_X1 U19344 ( .A1(n16171), .A2(n18324), .ZN(n18320) );
  INV_X1 U19345 ( .A(n16172), .ZN(n18316) );
  INV_X1 U19346 ( .A(n16276), .ZN(n16538) );
  OAI22_X1 U19347 ( .A1(n16174), .A2(n16450), .B1(n16551), .B2(n16538), .ZN(
        n16175) );
  AOI211_X1 U19348 ( .C1(n16177), .C2(n16206), .A(n16176), .B(n16175), .ZN(
        n16195) );
  NOR2_X1 U19349 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16178), .ZN(n16199) );
  NOR2_X1 U19350 ( .A1(n16529), .A2(n16530), .ZN(n16545) );
  INV_X1 U19351 ( .A(n16529), .ZN(n16541) );
  OAI221_X1 U19352 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n16510), .C1(n16179), 
        .C2(n16510), .A(n16541), .ZN(n16226) );
  INV_X1 U19353 ( .A(n16226), .ZN(n16244) );
  OAI21_X1 U19354 ( .B1(n16545), .B2(n16180), .A(n16244), .ZN(n16212) );
  OAI21_X1 U19355 ( .B1(n16199), .B2(n16212), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16194) );
  INV_X1 U19356 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U19357 ( .A1(n16181), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n17138), .B2(n16190), .ZN(n17134) );
  INV_X1 U19358 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16182) );
  NAND2_X1 U19359 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17145), .ZN(
        n17114) );
  AOI21_X1 U19360 ( .B1(n16182), .B2(n17114), .A(n16181), .ZN(n17146) );
  INV_X1 U19361 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17171) );
  INV_X1 U19362 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17187) );
  NOR2_X1 U19363 ( .A1(n17484), .A2(n17199), .ZN(n16187) );
  INV_X1 U19364 ( .A(n16187), .ZN(n16188) );
  NOR2_X1 U19365 ( .A1(n17187), .A2(n17155), .ZN(n16185) );
  INV_X1 U19366 ( .A(n16185), .ZN(n16184) );
  NOR2_X1 U19367 ( .A1(n17171), .A2(n16184), .ZN(n16183) );
  OAI21_X1 U19368 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16183), .A(
        n17114), .ZN(n17159) );
  INV_X1 U19369 ( .A(n17159), .ZN(n16249) );
  OAI22_X1 U19370 ( .A1(n17171), .A2(n16185), .B1(n16184), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17168) );
  AOI21_X1 U19371 ( .B1(n17187), .B2(n17155), .A(n16185), .ZN(n17185) );
  INV_X1 U19372 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17217) );
  NOR2_X1 U19373 ( .A1(n17217), .A2(n16188), .ZN(n16186) );
  OAI21_X1 U19374 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16186), .A(
        n17155), .ZN(n17202) );
  INV_X1 U19375 ( .A(n17202), .ZN(n16281) );
  OAI22_X1 U19376 ( .A1(n17217), .A2(n16187), .B1(n16188), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17213) );
  INV_X1 U19377 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17244) );
  NAND2_X1 U19378 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17241), .ZN(
        n17239) );
  INV_X1 U19379 ( .A(n17239), .ZN(n16323) );
  NAND2_X1 U19380 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16323), .ZN(
        n16322) );
  NOR2_X1 U19381 ( .A1(n17244), .A2(n16322), .ZN(n17197) );
  OAI21_X1 U19382 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17197), .A(
        n16188), .ZN(n16189) );
  INV_X1 U19383 ( .A(n16189), .ZN(n17231) );
  NAND2_X1 U19384 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17281), .ZN(
        n16331) );
  INV_X1 U19385 ( .A(n16331), .ZN(n17283) );
  NAND2_X1 U19386 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17283), .ZN(
        n16353) );
  NOR2_X1 U19387 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16353), .ZN(
        n16307) );
  INV_X4 U19388 ( .A(n16496), .ZN(n16467) );
  AOI21_X1 U19389 ( .B1(n17197), .B2(n16307), .A(n16467), .ZN(n16299) );
  NOR2_X1 U19390 ( .A1(n16298), .A2(n16467), .ZN(n16291) );
  NOR2_X1 U19391 ( .A1(n17213), .A2(n16291), .ZN(n16290) );
  NOR2_X1 U19392 ( .A1(n16290), .A2(n16467), .ZN(n16280) );
  NOR2_X1 U19393 ( .A1(n16279), .A2(n16467), .ZN(n16270) );
  NOR2_X1 U19394 ( .A1(n16269), .A2(n16467), .ZN(n16257) );
  NOR2_X1 U19395 ( .A1(n16256), .A2(n16467), .ZN(n16248) );
  NOR2_X1 U19396 ( .A1(n16247), .A2(n16467), .ZN(n16236) );
  NOR2_X1 U19397 ( .A1(n16235), .A2(n16467), .ZN(n16228) );
  NOR2_X1 U19398 ( .A1(n17134), .A2(n16228), .ZN(n16227) );
  NOR2_X1 U19399 ( .A1(n16190), .A2(n17138), .ZN(n16192) );
  OAI21_X1 U19400 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16192), .A(
        n16191), .ZN(n16216) );
  AOI21_X1 U19401 ( .B1(n16227), .B2(n16216), .A(n16467), .ZN(n16208) );
  NAND4_X1 U19402 ( .A1(n9609), .A2(n9720), .A3(n16207), .A4(n16196), .ZN(
        n16193) );
  NAND3_X1 U19403 ( .A1(n16195), .A2(n16194), .A3(n16193), .ZN(P3_U2640) );
  NOR2_X1 U19404 ( .A1(n16207), .A2(n16467), .ZN(n16197) );
  XOR2_X1 U19405 ( .A(n16197), .B(n16196), .Z(n16204) );
  NOR2_X1 U19406 ( .A1(n16198), .A2(n16450), .ZN(n16200) );
  AOI211_X1 U19407 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n16212), .A(n16200), 
        .B(n16199), .ZN(n16203) );
  XNOR2_X1 U19408 ( .A(P3_EBX_REG_30__SCAN_IN), .B(n16206), .ZN(n16201) );
  AOI22_X1 U19409 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16276), .B1(n16525), 
        .B2(n16201), .ZN(n16202) );
  OAI211_X1 U19410 ( .C1(n18330), .C2(n16204), .A(n16203), .B(n16202), .ZN(
        P3_U2641) );
  NOR2_X1 U19411 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16221), .ZN(n16205) );
  AOI22_X1 U19412 ( .A1(n16531), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16232), 
        .B2(n16205), .ZN(n16214) );
  AOI211_X1 U19413 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16219), .A(n16206), .B(
        n16539), .ZN(n16211) );
  AOI211_X1 U19414 ( .C1(n16209), .C2(n16208), .A(n16207), .B(n18330), .ZN(
        n16210) );
  AOI211_X1 U19415 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16212), .A(n16211), 
        .B(n16210), .ZN(n16213) );
  OAI211_X1 U19416 ( .C1(n16215), .C2(n16450), .A(n16214), .B(n16213), .ZN(
        P3_U2642) );
  AOI22_X1 U19417 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16225) );
  NOR2_X1 U19418 ( .A1(n16467), .A2(n16227), .ZN(n16217) );
  INV_X1 U19419 ( .A(n16216), .ZN(n17115) );
  XOR2_X1 U19420 ( .A(n16217), .B(n17115), .Z(n16218) );
  AOI22_X1 U19421 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16226), .B1(n9720), 
        .B2(n16218), .ZN(n16224) );
  OAI211_X1 U19422 ( .C1(n16229), .C2(n16220), .A(n16525), .B(n16219), .ZN(
        n16223) );
  OAI211_X1 U19423 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16232), .B(n16221), .ZN(n16222) );
  NAND4_X1 U19424 ( .A1(n16225), .A2(n16224), .A3(n16223), .A4(n16222), .ZN(
        P3_U2643) );
  AOI22_X1 U19425 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16226), .B1(n16531), 
        .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16234) );
  INV_X1 U19426 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18400) );
  AOI211_X1 U19427 ( .C1(n17134), .C2(n16228), .A(n16227), .B(n18330), .ZN(
        n16231) );
  AOI211_X1 U19428 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16240), .A(n16229), .B(
        n16539), .ZN(n16230) );
  AOI211_X1 U19429 ( .C1(n16232), .C2(n18400), .A(n16231), .B(n16230), .ZN(
        n16233) );
  OAI211_X1 U19430 ( .C1(n17138), .C2(n16450), .A(n16234), .B(n16233), .ZN(
        P3_U2644) );
  AOI211_X1 U19431 ( .C1(n17146), .C2(n16236), .A(n16235), .B(n18330), .ZN(
        n16239) );
  OAI22_X1 U19432 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16237), .B1(n16241), 
        .B2(n16538), .ZN(n16238) );
  AOI211_X1 U19433 ( .C1(n16533), .C2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16239), .B(n16238), .ZN(n16243) );
  OAI211_X1 U19434 ( .C1(n16246), .C2(n16241), .A(n16525), .B(n16240), .ZN(
        n16242) );
  OAI211_X1 U19435 ( .C1(n16244), .C2(n18398), .A(n16243), .B(n16242), .ZN(
        P3_U2645) );
  NAND2_X1 U19436 ( .A1(n16530), .A2(n16245), .ZN(n16255) );
  AOI22_X1 U19437 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16254) );
  AOI21_X1 U19438 ( .B1(n16530), .B2(n16259), .A(n16529), .ZN(n16267) );
  OAI21_X1 U19439 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16510), .A(n16267), 
        .ZN(n16252) );
  AOI211_X1 U19440 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16262), .A(n16246), .B(
        n16539), .ZN(n16251) );
  AOI211_X1 U19441 ( .C1(n16249), .C2(n16248), .A(n16247), .B(n18330), .ZN(
        n16250) );
  AOI211_X1 U19442 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16252), .A(n16251), 
        .B(n16250), .ZN(n16253) );
  OAI211_X1 U19443 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16255), .A(n16254), 
        .B(n16253), .ZN(P3_U2646) );
  AOI211_X1 U19444 ( .C1(n17168), .C2(n16257), .A(n16256), .B(n18330), .ZN(
        n16261) );
  NAND2_X1 U19445 ( .A1(n16530), .A2(n20587), .ZN(n16258) );
  OAI22_X1 U19446 ( .A1(n16538), .A2(n16549), .B1(n16259), .B2(n16258), .ZN(
        n16260) );
  AOI211_X1 U19447 ( .C1(n16533), .C2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16261), .B(n16260), .ZN(n16264) );
  OAI211_X1 U19448 ( .C1(n16268), .C2(n16549), .A(n16525), .B(n16262), .ZN(
        n16263) );
  OAI211_X1 U19449 ( .C1(n16267), .C2(n20587), .A(n16264), .B(n16263), .ZN(
        P3_U2647) );
  NAND2_X1 U19450 ( .A1(n16530), .A2(n16277), .ZN(n16352) );
  NOR2_X1 U19451 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16352), .ZN(n16265) );
  AOI22_X1 U19452 ( .A1(n16531), .A2(P3_EBX_REG_23__SCAN_IN), .B1(n16266), 
        .B2(n16265), .ZN(n16275) );
  INV_X1 U19453 ( .A(n16267), .ZN(n16273) );
  AOI211_X1 U19454 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16283), .A(n16268), .B(
        n16539), .ZN(n16272) );
  AOI211_X1 U19455 ( .C1(n17185), .C2(n16270), .A(n16269), .B(n18330), .ZN(
        n16271) );
  AOI211_X1 U19456 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16273), .A(n16272), 
        .B(n16271), .ZN(n16274) );
  OAI211_X1 U19457 ( .C1(n17187), .C2(n16450), .A(n16275), .B(n16274), .ZN(
        P3_U2648) );
  AOI22_X1 U19458 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16533), .B1(
        n16276), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16288) );
  NAND2_X1 U19459 ( .A1(n16541), .A2(n16277), .ZN(n16368) );
  INV_X1 U19460 ( .A(n16368), .ZN(n16342) );
  AOI21_X1 U19461 ( .B1(n16278), .B2(n16342), .A(n16545), .ZN(n16302) );
  INV_X1 U19462 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18388) );
  INV_X1 U19463 ( .A(n16352), .ZN(n16360) );
  AND3_X1 U19464 ( .A1(n18388), .A2(n16278), .A3(n16360), .ZN(n16289) );
  AOI211_X1 U19465 ( .C1(n16281), .C2(n16280), .A(n16279), .B(n18330), .ZN(
        n16282) );
  AOI221_X1 U19466 ( .B1(n16302), .B2(P3_REIP_REG_22__SCAN_IN), .C1(n16289), 
        .C2(P3_REIP_REG_22__SCAN_IN), .A(n16282), .ZN(n16287) );
  OAI211_X1 U19467 ( .C1(n16292), .C2(n16546), .A(n16525), .B(n16283), .ZN(
        n16286) );
  OR3_X1 U19468 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16284), .A3(n16352), .ZN(
        n16285) );
  NAND4_X1 U19469 ( .A1(n16288), .A2(n16287), .A3(n16286), .A4(n16285), .ZN(
        P3_U2649) );
  AOI21_X1 U19470 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16531), .A(n16289), .ZN(
        n16296) );
  AOI211_X1 U19471 ( .C1(n17213), .C2(n16291), .A(n16290), .B(n18330), .ZN(
        n16294) );
  AOI211_X1 U19472 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16303), .A(n16292), .B(
        n16539), .ZN(n16293) );
  AOI211_X1 U19473 ( .C1(n16302), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16294), 
        .B(n16293), .ZN(n16295) );
  OAI211_X1 U19474 ( .C1(n17217), .C2(n16450), .A(n16296), .B(n16295), .ZN(
        P3_U2650) );
  AOI22_X1 U19475 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16306) );
  NOR2_X1 U19476 ( .A1(n16297), .A2(n16352), .ZN(n16301) );
  AOI211_X1 U19477 ( .C1(n17231), .C2(n16299), .A(n16298), .B(n18330), .ZN(
        n16300) );
  AOI221_X1 U19478 ( .B1(n16302), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16301), 
        .C2(n18387), .A(n16300), .ZN(n16305) );
  OAI211_X1 U19479 ( .C1(n16311), .C2(n16653), .A(n16525), .B(n16303), .ZN(
        n16304) );
  NAND3_X1 U19480 ( .A1(n16306), .A2(n16305), .A3(n16304), .ZN(P3_U2651) );
  AOI21_X1 U19481 ( .B1(n17244), .B2(n16322), .A(n17197), .ZN(n17246) );
  INV_X1 U19482 ( .A(n16307), .ZN(n16356) );
  OAI21_X1 U19483 ( .B1(n16322), .B2(n16356), .A(n9609), .ZN(n16308) );
  XNOR2_X1 U19484 ( .A(n17246), .B(n16308), .ZN(n16309) );
  AOI22_X1 U19485 ( .A1(n16531), .A2(P3_EBX_REG_19__SCAN_IN), .B1(n9720), .B2(
        n16309), .ZN(n16317) );
  AOI21_X1 U19486 ( .B1(n16310), .B2(n16342), .A(n16545), .ZN(n16338) );
  NOR2_X1 U19487 ( .A1(n17244), .A2(n16450), .ZN(n16313) );
  AOI211_X1 U19488 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16320), .A(n16311), .B(
        n16539), .ZN(n16312) );
  AOI211_X1 U19489 ( .C1(n16338), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16313), 
        .B(n16312), .ZN(n16316) );
  NOR3_X1 U19490 ( .A1(n18381), .A2(n16341), .A3(n16352), .ZN(n16319) );
  NAND2_X1 U19491 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16314) );
  OAI211_X1 U19492 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16319), .B(n16314), .ZN(n16315) );
  NAND4_X1 U19493 ( .A1(n16317), .A2(n16316), .A3(n17712), .A4(n16315), .ZN(
        P3_U2652) );
  INV_X1 U19494 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18383) );
  INV_X1 U19495 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17259) );
  OAI22_X1 U19496 ( .A1(n17259), .A2(n16450), .B1(n16538), .B2(n16321), .ZN(
        n16318) );
  AOI221_X1 U19497 ( .B1(n16338), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16319), 
        .C2(n18383), .A(n16318), .ZN(n16328) );
  OAI211_X1 U19498 ( .C1(n16329), .C2(n16321), .A(n16525), .B(n16320), .ZN(
        n16327) );
  OAI21_X1 U19499 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16323), .A(
        n16322), .ZN(n17256) );
  OAI21_X1 U19500 ( .B1(n17239), .B2(n16356), .A(n9609), .ZN(n16325) );
  AOI21_X1 U19501 ( .B1(n17256), .B2(n16325), .A(n18330), .ZN(n16324) );
  OAI21_X1 U19502 ( .B1(n17256), .B2(n16325), .A(n16324), .ZN(n16326) );
  NAND4_X1 U19503 ( .A1(n16328), .A2(n17712), .A3(n16327), .A4(n16326), .ZN(
        P3_U2653) );
  AOI211_X1 U19504 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16344), .A(n16329), .B(
        n16539), .ZN(n16330) );
  AOI211_X1 U19505 ( .C1(n16531), .C2(P3_EBX_REG_17__SCAN_IN), .A(n9597), .B(
        n16330), .ZN(n16340) );
  NOR2_X1 U19506 ( .A1(n16341), .A2(n16352), .ZN(n16337) );
  NAND2_X1 U19507 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17280) );
  NOR2_X1 U19508 ( .A1(n17280), .A2(n16331), .ZN(n16332) );
  OAI21_X1 U19509 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16332), .A(
        n17239), .ZN(n17268) );
  INV_X1 U19510 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16333) );
  AOI21_X1 U19511 ( .B1(n16333), .B2(n16353), .A(n16332), .ZN(n17284) );
  OAI21_X1 U19512 ( .B1(n17284), .B2(n16356), .A(n9609), .ZN(n16335) );
  OAI21_X1 U19513 ( .B1(n17268), .B2(n16335), .A(n9720), .ZN(n16334) );
  AOI21_X1 U19514 ( .B1(n17268), .B2(n16335), .A(n16334), .ZN(n16336) );
  AOI221_X1 U19515 ( .B1(n16338), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16337), 
        .C2(n18381), .A(n16336), .ZN(n16339) );
  OAI211_X1 U19516 ( .C1(n17226), .C2(n16450), .A(n16340), .B(n16339), .ZN(
        P3_U2654) );
  OAI21_X1 U19517 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), 
        .A(n16341), .ZN(n16351) );
  AOI22_X1 U19518 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16350) );
  NOR2_X1 U19519 ( .A1(n16545), .A2(n16342), .ZN(n16361) );
  NAND2_X1 U19520 ( .A1(n9609), .A2(n16356), .ZN(n16343) );
  XOR2_X1 U19521 ( .A(n16343), .B(n17284), .Z(n16347) );
  OAI211_X1 U19522 ( .C1(n16354), .C2(n16345), .A(n16525), .B(n16344), .ZN(
        n16346) );
  OAI21_X1 U19523 ( .B1(n16347), .B2(n18330), .A(n16346), .ZN(n16348) );
  AOI211_X1 U19524 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n16361), .A(n9597), .B(
        n16348), .ZN(n16349) );
  OAI211_X1 U19525 ( .C1(n16352), .C2(n16351), .A(n16350), .B(n16349), .ZN(
        P3_U2655) );
  NOR2_X1 U19526 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18330), .ZN(
        n16526) );
  INV_X1 U19527 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16358) );
  NAND2_X1 U19528 ( .A1(n16467), .A2(n9720), .ZN(n16483) );
  INV_X1 U19529 ( .A(n16483), .ZN(n16527) );
  AOI21_X1 U19530 ( .B1(n16526), .B2(n16358), .A(n16527), .ZN(n16364) );
  OAI21_X1 U19531 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17283), .A(
        n16353), .ZN(n17294) );
  AOI211_X1 U19532 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16370), .A(n16354), .B(
        n16539), .ZN(n16355) );
  AOI21_X1 U19533 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16531), .A(n16355), .ZN(
        n16363) );
  INV_X1 U19534 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18377) );
  NOR2_X1 U19535 ( .A1(n16467), .A2(n18330), .ZN(n16532) );
  NAND3_X1 U19536 ( .A1(n16532), .A2(n16356), .A3(n17294), .ZN(n16357) );
  OAI211_X1 U19537 ( .C1(n16358), .C2(n16450), .A(n17712), .B(n16357), .ZN(
        n16359) );
  AOI221_X1 U19538 ( .B1(n16361), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n16360), 
        .C2(n18377), .A(n16359), .ZN(n16362) );
  OAI211_X1 U19539 ( .C1(n16364), .C2(n17294), .A(n16363), .B(n16362), .ZN(
        P3_U2656) );
  AOI22_X1 U19540 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16373) );
  NAND2_X1 U19541 ( .A1(n17391), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17392) );
  NOR2_X1 U19542 ( .A1(n17484), .A2(n17392), .ZN(n16443) );
  NAND2_X1 U19543 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16443), .ZN(
        n16430) );
  NOR2_X1 U19544 ( .A1(n16365), .A2(n16430), .ZN(n17320) );
  INV_X1 U19545 ( .A(n17320), .ZN(n16397) );
  OR2_X1 U19546 ( .A1(n17323), .A2(n16397), .ZN(n16375) );
  AOI21_X1 U19547 ( .B1(n17308), .B2(n16375), .A(n17283), .ZN(n17310) );
  INV_X1 U19548 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16469) );
  NAND3_X1 U19549 ( .A1(n16469), .A2(n17391), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16444) );
  INV_X1 U19550 ( .A(n16444), .ZN(n16448) );
  NAND2_X1 U19551 ( .A1(n17306), .A2(n16448), .ZN(n16388) );
  OAI21_X1 U19552 ( .B1(n17323), .B2(n16388), .A(n9609), .ZN(n16378) );
  XNOR2_X1 U19553 ( .A(n17310), .B(n16378), .ZN(n16369) );
  OR2_X1 U19554 ( .A1(n16510), .A2(n16366), .ZN(n16387) );
  OAI22_X1 U19555 ( .A1(n16545), .A2(n18376), .B1(n16387), .B2(n18373), .ZN(
        n16367) );
  AOI22_X1 U19556 ( .A1(n9720), .A2(n16369), .B1(n16368), .B2(n16367), .ZN(
        n16372) );
  OAI211_X1 U19557 ( .C1(n16374), .C2(n16730), .A(n16525), .B(n16370), .ZN(
        n16371) );
  NAND4_X1 U19558 ( .A1(n16373), .A2(n16372), .A3(n17712), .A4(n16371), .ZN(
        P3_U2657) );
  INV_X1 U19559 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18371) );
  OAI21_X1 U19560 ( .B1(n16391), .B2(n16510), .A(n16541), .ZN(n16405) );
  AOI21_X1 U19561 ( .B1(n16530), .B2(n18371), .A(n16405), .ZN(n16386) );
  AOI211_X1 U19562 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16392), .A(n16374), .B(
        n16539), .ZN(n16384) );
  INV_X1 U19563 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16379) );
  INV_X1 U19564 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17333) );
  NOR2_X1 U19565 ( .A1(n17333), .A2(n16397), .ZN(n16376) );
  OAI21_X1 U19566 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16376), .A(
        n16375), .ZN(n17326) );
  NAND2_X1 U19567 ( .A1(n9720), .A2(n17326), .ZN(n16377) );
  OAI22_X1 U19568 ( .A1(n16538), .A2(n16379), .B1(n16378), .B2(n16377), .ZN(
        n16383) );
  INV_X1 U19569 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16380) );
  AOI21_X1 U19570 ( .B1(n16526), .B2(n16380), .A(n16527), .ZN(n16381) );
  OAI22_X1 U19571 ( .A1(n16381), .A2(n17326), .B1(n16380), .B2(n16450), .ZN(
        n16382) );
  NOR4_X1 U19572 ( .A1(n9597), .A2(n16384), .A3(n16383), .A4(n16382), .ZN(
        n16385) );
  OAI221_X1 U19573 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n16387), .C1(n18373), 
        .C2(n16386), .A(n16385), .ZN(P3_U2658) );
  AOI22_X1 U19574 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16396) );
  AOI22_X1 U19575 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16397), .B1(
        n17320), .B2(n17333), .ZN(n17345) );
  NAND2_X1 U19576 ( .A1(n9609), .A2(n16388), .ZN(n16398) );
  XOR2_X1 U19577 ( .A(n17345), .B(n16398), .Z(n16389) );
  AOI21_X1 U19578 ( .B1(n9720), .B2(n16389), .A(n9597), .ZN(n16395) );
  NOR2_X1 U19579 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16510), .ZN(n16390) );
  AOI22_X1 U19580 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16405), .B1(n16391), 
        .B2(n16390), .ZN(n16394) );
  OAI211_X1 U19581 ( .C1(n16402), .C2(n16732), .A(n16525), .B(n16392), .ZN(
        n16393) );
  NAND4_X1 U19582 ( .A1(n16396), .A2(n16395), .A3(n16394), .A4(n16393), .ZN(
        P3_U2659) );
  INV_X1 U19583 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17351) );
  INV_X1 U19584 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17367) );
  INV_X1 U19585 ( .A(n16430), .ZN(n16419) );
  NAND2_X1 U19586 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16419), .ZN(
        n16418) );
  NOR2_X1 U19587 ( .A1(n17367), .A2(n16418), .ZN(n16411) );
  OAI21_X1 U19588 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16411), .A(
        n16397), .ZN(n17352) );
  AOI22_X1 U19589 ( .A1(n9720), .A2(n17352), .B1(n16411), .B2(n16526), .ZN(
        n16399) );
  AOI22_X1 U19590 ( .A1(n16399), .A2(n16483), .B1(n17352), .B2(n16398), .ZN(
        n16400) );
  AOI21_X1 U19591 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16531), .A(n16400), .ZN(
        n16407) );
  OAI21_X1 U19592 ( .B1(n16510), .B2(n16401), .A(n18369), .ZN(n16404) );
  AOI211_X1 U19593 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16413), .A(n16402), .B(
        n16539), .ZN(n16403) );
  AOI211_X1 U19594 ( .C1(n16405), .C2(n16404), .A(n9597), .B(n16403), .ZN(
        n16406) );
  OAI211_X1 U19595 ( .C1(n17351), .C2(n16450), .A(n16407), .B(n16406), .ZN(
        P3_U2660) );
  OAI21_X1 U19596 ( .B1(n16408), .B2(n16510), .A(n16541), .ZN(n16435) );
  INV_X1 U19597 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18367) );
  INV_X1 U19598 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18365) );
  NAND2_X1 U19599 ( .A1(n16530), .A2(n16408), .ZN(n16429) );
  AOI221_X1 U19600 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n18367), .C2(n18365), .A(n16429), .ZN(n16410) );
  OAI22_X1 U19601 ( .A1(n17367), .A2(n16450), .B1(n16538), .B2(n16777), .ZN(
        n16409) );
  AOI211_X1 U19602 ( .C1(n16435), .C2(P3_REIP_REG_10__SCAN_IN), .A(n16410), 
        .B(n16409), .ZN(n16416) );
  AOI21_X1 U19603 ( .B1(n17367), .B2(n16418), .A(n16411), .ZN(n17363) );
  NOR2_X1 U19604 ( .A1(n17394), .A2(n16444), .ZN(n16422) );
  AOI21_X1 U19605 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16422), .A(
        n16467), .ZN(n16421) );
  AOI21_X1 U19606 ( .B1(n17363), .B2(n16421), .A(n18330), .ZN(n16412) );
  OAI21_X1 U19607 ( .B1(n17363), .B2(n16421), .A(n16412), .ZN(n16415) );
  OAI211_X1 U19608 ( .C1(n16417), .C2(n16777), .A(n16525), .B(n16413), .ZN(
        n16414) );
  NAND4_X1 U19609 ( .A1(n16416), .A2(n17712), .A3(n16415), .A4(n16414), .ZN(
        P3_U2661) );
  INV_X1 U19610 ( .A(n16435), .ZN(n16428) );
  AOI211_X1 U19611 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16437), .A(n16417), .B(
        n16539), .ZN(n16426) );
  INV_X1 U19612 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16420) );
  OAI21_X1 U19613 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16419), .A(
        n16418), .ZN(n17386) );
  OAI22_X1 U19614 ( .A1(n16538), .A2(n16420), .B1(n17386), .B2(n16483), .ZN(
        n16425) );
  INV_X1 U19615 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17375) );
  OAI211_X1 U19616 ( .C1(n16422), .C2(n17386), .A(n9720), .B(n16421), .ZN(
        n16423) );
  OAI21_X1 U19617 ( .B1(n16450), .B2(n17375), .A(n16423), .ZN(n16424) );
  NOR4_X1 U19618 ( .A1(n9597), .A2(n16426), .A3(n16425), .A4(n16424), .ZN(
        n16427) );
  OAI221_X1 U19619 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16429), .C1(n18365), 
        .C2(n16428), .A(n16427), .ZN(P3_U2662) );
  AOI22_X1 U19620 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n16441) );
  AOI21_X1 U19621 ( .B1(n16443), .B2(n16469), .A(n16467), .ZN(n16431) );
  OAI21_X1 U19622 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16443), .A(
        n16430), .ZN(n17397) );
  XNOR2_X1 U19623 ( .A(n16431), .B(n17397), .ZN(n16436) );
  INV_X1 U19624 ( .A(n16432), .ZN(n16473) );
  NAND2_X1 U19625 ( .A1(n16530), .A2(n16473), .ZN(n16464) );
  OAI21_X1 U19626 ( .B1(n16433), .B2(n16464), .A(n20608), .ZN(n16434) );
  AOI22_X1 U19627 ( .A1(n9720), .A2(n16436), .B1(n16435), .B2(n16434), .ZN(
        n16440) );
  OAI211_X1 U19628 ( .C1(n16445), .C2(n16438), .A(n16525), .B(n16437), .ZN(
        n16439) );
  NAND4_X1 U19629 ( .A1(n16441), .A2(n16440), .A3(n17712), .A4(n16439), .ZN(
        P3_U2663) );
  INV_X1 U19630 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17406) );
  INV_X1 U19631 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16466) );
  NAND3_X1 U19632 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16442), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16482) );
  NOR2_X1 U19633 ( .A1(n16466), .A2(n16482), .ZN(n16465) );
  NAND2_X1 U19634 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16465), .ZN(
        n16455) );
  AOI21_X1 U19635 ( .B1(n17406), .B2(n16455), .A(n16443), .ZN(n17411) );
  NAND3_X1 U19636 ( .A1(n9720), .A2(n9609), .A3(n16444), .ZN(n16459) );
  AOI211_X1 U19637 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16456), .A(n16445), .B(
        n16539), .ZN(n16446) );
  AOI21_X1 U19638 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n16531), .A(n16446), .ZN(
        n16454) );
  OAI21_X1 U19639 ( .B1(n16473), .B2(n16510), .A(n16541), .ZN(n16476) );
  AOI211_X1 U19640 ( .C1(n18362), .C2(n18360), .A(n16447), .B(n16464), .ZN(
        n16452) );
  OAI211_X1 U19641 ( .C1(n16448), .C2(n16467), .A(n9720), .B(n17411), .ZN(
        n16449) );
  OAI211_X1 U19642 ( .C1(n17406), .C2(n16450), .A(n17712), .B(n16449), .ZN(
        n16451) );
  AOI211_X1 U19643 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n16476), .A(n16452), .B(
        n16451), .ZN(n16453) );
  OAI211_X1 U19644 ( .C1(n17411), .C2(n16459), .A(n16454), .B(n16453), .ZN(
        P3_U2664) );
  AOI22_X1 U19645 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16463) );
  OAI21_X1 U19646 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16465), .A(
        n16455), .ZN(n17423) );
  INV_X1 U19647 ( .A(n17423), .ZN(n16460) );
  OAI22_X1 U19648 ( .A1(n16527), .A2(n16526), .B1(n17422), .B2(n16467), .ZN(
        n16458) );
  OAI211_X1 U19649 ( .C1(n16470), .C2(n20629), .A(n16525), .B(n16456), .ZN(
        n16457) );
  OAI221_X1 U19650 ( .B1(n16460), .B2(n16459), .C1(n17423), .C2(n16458), .A(
        n16457), .ZN(n16461) );
  AOI211_X1 U19651 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n16476), .A(n9597), .B(
        n16461), .ZN(n16462) );
  OAI211_X1 U19652 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n16464), .A(n16463), .B(
        n16462), .ZN(P3_U2665) );
  AOI22_X1 U19653 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16533), .B1(
        n16531), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n16479) );
  AOI21_X1 U19654 ( .B1(n16466), .B2(n16482), .A(n16465), .ZN(n17434) );
  INV_X1 U19655 ( .A(n16482), .ZN(n16468) );
  AOI21_X1 U19656 ( .B1(n16469), .B2(n16468), .A(n16467), .ZN(n16484) );
  XOR2_X1 U19657 ( .A(n17434), .B(n16484), .Z(n16472) );
  AOI211_X1 U19658 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16486), .A(n16470), .B(
        n16539), .ZN(n16471) );
  NOR2_X1 U19659 ( .A1(n16473), .A2(n16510), .ZN(n16474) );
  AOI22_X1 U19660 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16476), .B1(n16475), 
        .B2(n16474), .ZN(n16477) );
  NAND3_X1 U19661 ( .A1(n16479), .A2(n16478), .A3(n16477), .ZN(P3_U2666) );
  AOI21_X1 U19662 ( .B1(n16530), .B2(n16480), .A(n16529), .ZN(n16504) );
  NOR3_X1 U19663 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16510), .A3(n16480), .ZN(
        n16481) );
  AOI21_X1 U19664 ( .B1(n16533), .B2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16481), .ZN(n16495) );
  NOR2_X1 U19665 ( .A1(n17484), .A2(n17441), .ZN(n16497) );
  OAI21_X1 U19666 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16497), .A(
        n16482), .ZN(n17449) );
  OAI22_X1 U19667 ( .A1(n16538), .A2(n16487), .B1(n17449), .B2(n16483), .ZN(
        n16493) );
  NOR2_X1 U19668 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17484), .ZN(
        n16514) );
  NOR2_X1 U19669 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17441), .ZN(
        n16485) );
  AOI22_X1 U19670 ( .A1(n16514), .A2(n16485), .B1(n16484), .B2(n17449), .ZN(
        n16491) );
  OAI211_X1 U19671 ( .C1(n16498), .C2(n16487), .A(n16525), .B(n16486), .ZN(
        n16490) );
  NOR2_X1 U19672 ( .A1(n17001), .A2(n16488), .ZN(n18490) );
  OAI21_X1 U19673 ( .B1(n16796), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18490), .ZN(n16489) );
  OAI211_X1 U19674 ( .C1(n16491), .C2(n18330), .A(n16490), .B(n16489), .ZN(
        n16492) );
  NOR3_X1 U19675 ( .A1(n9597), .A2(n16493), .A3(n16492), .ZN(n16494) );
  OAI211_X1 U19676 ( .C1(n18356), .C2(n16504), .A(n16495), .B(n16494), .ZN(
        P3_U2667) );
  INV_X1 U19677 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16509) );
  NAND2_X1 U19678 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16511) );
  OAI21_X1 U19679 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16511), .A(
        n9609), .ZN(n16499) );
  NOR2_X1 U19680 ( .A1(n18330), .A2(n16499), .ZN(n16513) );
  INV_X1 U19681 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17458) );
  AOI21_X1 U19682 ( .B1(n17458), .B2(n16511), .A(n16497), .ZN(n16501) );
  INV_X1 U19683 ( .A(n16501), .ZN(n17464) );
  AOI211_X1 U19684 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16519), .A(n16498), .B(
        n16539), .ZN(n16506) );
  INV_X1 U19685 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18353) );
  NOR2_X1 U19686 ( .A1(n18450), .A2(n18299), .ZN(n18298) );
  OAI21_X1 U19687 ( .B1(n18298), .B2(n18425), .A(n9648), .ZN(n18422) );
  AOI22_X1 U19688 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16533), .B1(
        n18490), .B2(n18422), .ZN(n16503) );
  NAND3_X1 U19689 ( .A1(n16501), .A2(n9720), .A3(n16499), .ZN(n16502) );
  OAI211_X1 U19690 ( .C1(n16504), .C2(n18353), .A(n16503), .B(n16502), .ZN(
        n16505) );
  AOI211_X1 U19691 ( .C1(n16513), .C2(n17464), .A(n16506), .B(n16505), .ZN(
        n16508) );
  NAND4_X1 U19692 ( .A1(n16530), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .A4(n18353), .ZN(n16507) );
  OAI211_X1 U19693 ( .C1(n16509), .C2(n16538), .A(n16508), .B(n16507), .ZN(
        P3_U2668) );
  INV_X1 U19694 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18351) );
  AOI221_X1 U19695 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_2__SCAN_IN), 
        .C1(n18452), .C2(n18351), .A(n16510), .ZN(n16518) );
  NOR2_X1 U19696 ( .A1(n18450), .A2(n18443), .ZN(n18281) );
  NOR2_X1 U19697 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18281), .ZN(
        n18302) );
  NOR2_X1 U19698 ( .A1(n18302), .A2(n18298), .ZN(n18432) );
  OAI21_X1 U19699 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16511), .ZN(n17470) );
  INV_X1 U19700 ( .A(n17470), .ZN(n16512) );
  AOI22_X1 U19701 ( .A1(n18432), .A2(n18490), .B1(n16512), .B2(n16527), .ZN(
        n16516) );
  OAI21_X1 U19702 ( .B1(n16514), .B2(n17470), .A(n16513), .ZN(n16515) );
  OAI211_X1 U19703 ( .C1(n16520), .C2(n16538), .A(n16516), .B(n16515), .ZN(
        n16517) );
  AOI211_X1 U19704 ( .C1(n16533), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16518), .B(n16517), .ZN(n16522) );
  OAI211_X1 U19705 ( .C1(n16524), .C2(n16520), .A(n16525), .B(n16519), .ZN(
        n16521) );
  OAI211_X1 U19706 ( .C1(n18351), .C2(n16541), .A(n16522), .B(n16521), .ZN(
        P3_U2669) );
  INV_X1 U19707 ( .A(n16523), .ZN(n16840) );
  NOR2_X1 U19708 ( .A1(n16524), .A2(n16840), .ZN(n16844) );
  AOI22_X1 U19709 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n18443), .B2(n18450), .ZN(
        n18440) );
  AOI22_X1 U19710 ( .A1(n16525), .A2(n16844), .B1(n18440), .B2(n18490), .ZN(
        n16537) );
  OR2_X1 U19711 ( .A1(n16527), .A2(n16526), .ZN(n16528) );
  AOI22_X1 U19712 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16529), .B1(n17484), 
        .B2(n16528), .ZN(n16536) );
  AOI22_X1 U19713 ( .A1(n16531), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n16530), .B2(
        n18452), .ZN(n16535) );
  OAI221_X1 U19714 ( .B1(n16533), .B2(n16532), .C1(n16533), .C2(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16534) );
  NAND4_X1 U19715 ( .A1(n16537), .A2(n16536), .A3(n16535), .A4(n16534), .ZN(
        P3_U2670) );
  INV_X1 U19716 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18458) );
  NAND2_X1 U19717 ( .A1(n16539), .A2(n16538), .ZN(n16540) );
  AOI22_X1 U19718 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16540), .B1(n18490), .B2(
        n18450), .ZN(n16544) );
  NAND3_X1 U19719 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16542), .A3(
        n16541), .ZN(n16543) );
  OAI211_X1 U19720 ( .C1(n16545), .C2(n18458), .A(n16544), .B(n16543), .ZN(
        P3_U2671) );
  INV_X1 U19721 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16586) );
  NOR3_X1 U19722 ( .A1(n16546), .A2(n16637), .A3(n16583), .ZN(n16547) );
  NAND4_X1 U19723 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n16636), .A4(n16547), .ZN(n16548) );
  NOR4_X1 U19724 ( .A1(n16586), .A2(n16550), .A3(n16549), .A4(n16548), .ZN(
        n16577) );
  NAND2_X1 U19725 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16577), .ZN(n16576) );
  NAND2_X1 U19726 ( .A1(n16576), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16553) );
  NAND2_X1 U19727 ( .A1(n17864), .A2(n16551), .ZN(n16552) );
  OAI22_X1 U19728 ( .A1(n16850), .A2(n16553), .B1(n16576), .B2(n16552), .ZN(
        P3_U2672) );
  AOI22_X1 U19729 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16557) );
  AOI22_X1 U19730 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16556) );
  AOI22_X1 U19731 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16555) );
  AOI22_X1 U19732 ( .A1(n16786), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16554) );
  NAND4_X1 U19733 ( .A1(n16557), .A2(n16556), .A3(n16555), .A4(n16554), .ZN(
        n16563) );
  AOI22_X1 U19734 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16561) );
  AOI22_X1 U19735 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16560) );
  AOI22_X1 U19736 ( .A1(n16778), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16559) );
  AOI22_X1 U19737 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16558) );
  NAND4_X1 U19738 ( .A1(n16561), .A2(n16560), .A3(n16559), .A4(n16558), .ZN(
        n16562) );
  NOR2_X1 U19739 ( .A1(n16563), .A2(n16562), .ZN(n16575) );
  AOI22_X1 U19740 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16567) );
  AOI22_X1 U19741 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16566) );
  AOI22_X1 U19742 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16565) );
  AOI22_X1 U19743 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16564) );
  NAND4_X1 U19744 ( .A1(n16567), .A2(n16566), .A3(n16565), .A4(n16564), .ZN(
        n16573) );
  AOI22_X1 U19745 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16571) );
  AOI22_X1 U19746 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16570) );
  AOI22_X1 U19747 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U19748 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16568) );
  NAND4_X1 U19749 ( .A1(n16571), .A2(n16570), .A3(n16569), .A4(n16568), .ZN(
        n16572) );
  NOR2_X1 U19750 ( .A1(n16573), .A2(n16572), .ZN(n16581) );
  NOR3_X1 U19751 ( .A1(n16581), .A2(n16580), .A3(n16579), .ZN(n16574) );
  XOR2_X1 U19752 ( .A(n16575), .B(n16574), .Z(n16863) );
  OAI211_X1 U19753 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16577), .A(n16576), .B(
        n16847), .ZN(n16578) );
  OAI21_X1 U19754 ( .B1(n16863), .B2(n16847), .A(n16578), .ZN(P3_U2673) );
  NOR2_X1 U19755 ( .A1(n16580), .A2(n16579), .ZN(n16582) );
  XNOR2_X1 U19756 ( .A(n16582), .B(n16581), .ZN(n16867) );
  NOR3_X1 U19757 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16592), .A3(n16583), .ZN(
        n16584) );
  AOI21_X1 U19758 ( .B1(n16850), .B2(n16867), .A(n16584), .ZN(n16585) );
  OAI21_X1 U19759 ( .B1(n16587), .B2(n16586), .A(n16585), .ZN(P3_U2674) );
  AOI21_X1 U19760 ( .B1(n16589), .B2(n16593), .A(n16588), .ZN(n16875) );
  AOI22_X1 U19761 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16590), .B1(n16850), 
        .B2(n16875), .ZN(n16591) );
  OAI21_X1 U19762 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16592), .A(n16591), .ZN(
        P3_U2676) );
  AOI21_X1 U19763 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16847), .A(n16600), .ZN(
        n16596) );
  OAI21_X1 U19764 ( .B1(n16595), .B2(n16594), .A(n16593), .ZN(n16884) );
  OAI22_X1 U19765 ( .A1(n16597), .A2(n16596), .B1(n16847), .B2(n16884), .ZN(
        P3_U2677) );
  INV_X1 U19766 ( .A(n16605), .ZN(n16609) );
  AOI22_X1 U19767 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16847), .B1(
        P3_EBX_REG_24__SCAN_IN), .B2(n16609), .ZN(n16599) );
  XNOR2_X1 U19768 ( .A(n16598), .B(n16601), .ZN(n16889) );
  OAI22_X1 U19769 ( .A1(n16600), .A2(n16599), .B1(n16847), .B2(n16889), .ZN(
        P3_U2678) );
  OAI21_X1 U19770 ( .B1(n16603), .B2(n16602), .A(n16601), .ZN(n16894) );
  NAND3_X1 U19771 ( .A1(n16605), .A2(P3_EBX_REG_24__SCAN_IN), .A3(n16847), 
        .ZN(n16604) );
  OAI221_X1 U19772 ( .B1(n16605), .B2(P3_EBX_REG_24__SCAN_IN), .C1(n16847), 
        .C2(n16894), .A(n16604), .ZN(P3_U2679) );
  AOI21_X1 U19773 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16847), .A(n16625), .ZN(
        n16608) );
  XNOR2_X1 U19774 ( .A(n16607), .B(n16606), .ZN(n16899) );
  OAI22_X1 U19775 ( .A1(n16609), .A2(n16608), .B1(n16847), .B2(n16899), .ZN(
        P3_U2680) );
  AOI21_X1 U19776 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16847), .A(n16610), .ZN(
        n16624) );
  AOI22_X1 U19777 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16622) );
  AOI22_X1 U19778 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16621) );
  AOI22_X1 U19779 ( .A1(n16796), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16611) );
  OAI21_X1 U19780 ( .B1(n16612), .B2(n20519), .A(n16611), .ZN(n16618) );
  AOI22_X1 U19781 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16616) );
  AOI22_X1 U19782 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16615) );
  AOI22_X1 U19783 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16779), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16614) );
  AOI22_X1 U19784 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16613) );
  NAND4_X1 U19785 ( .A1(n16616), .A2(n16615), .A3(n16614), .A4(n16613), .ZN(
        n16617) );
  AOI211_X1 U19786 ( .C1(n16619), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n16618), .B(n16617), .ZN(n16620) );
  NAND3_X1 U19787 ( .A1(n16622), .A2(n16621), .A3(n16620), .ZN(n16900) );
  INV_X1 U19788 ( .A(n16900), .ZN(n16623) );
  OAI22_X1 U19789 ( .A1(n16625), .A2(n16624), .B1(n16623), .B2(n16834), .ZN(
        P3_U2681) );
  AOI22_X1 U19790 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16629) );
  AOI22_X1 U19791 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16628) );
  AOI22_X1 U19792 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16627) );
  AOI22_X1 U19793 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16626) );
  NAND4_X1 U19794 ( .A1(n16629), .A2(n16628), .A3(n16627), .A4(n16626), .ZN(
        n16635) );
  AOI22_X1 U19795 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16633) );
  AOI22_X1 U19796 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16632) );
  AOI22_X1 U19797 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16631) );
  AOI22_X1 U19798 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16630) );
  NAND4_X1 U19799 ( .A1(n16633), .A2(n16632), .A3(n16631), .A4(n16630), .ZN(
        n16634) );
  NOR2_X1 U19800 ( .A1(n16635), .A2(n16634), .ZN(n16910) );
  INV_X1 U19801 ( .A(n16910), .ZN(n16639) );
  OAI21_X1 U19802 ( .B1(n16637), .B2(n16636), .A(n16834), .ZN(n16638) );
  OAI21_X1 U19803 ( .B1(n16847), .B2(n16639), .A(n16638), .ZN(n16640) );
  OAI21_X1 U19804 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16641), .A(n16640), .ZN(
        P3_U2682) );
  AOI22_X1 U19805 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16645) );
  AOI22_X1 U19806 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16644) );
  AOI22_X1 U19807 ( .A1(n15275), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16643) );
  AOI22_X1 U19808 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16642) );
  NAND4_X1 U19809 ( .A1(n16645), .A2(n16644), .A3(n16643), .A4(n16642), .ZN(
        n16651) );
  AOI22_X1 U19810 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16779), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16649) );
  AOI22_X1 U19811 ( .A1(n16796), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16648) );
  AOI22_X1 U19812 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16647) );
  AOI22_X1 U19813 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14991), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16646) );
  NAND4_X1 U19814 ( .A1(n16649), .A2(n16648), .A3(n16647), .A4(n16646), .ZN(
        n16650) );
  NOR2_X1 U19815 ( .A1(n16651), .A2(n16650), .ZN(n16914) );
  INV_X1 U19816 ( .A(n16666), .ZN(n16652) );
  OAI33_X1 U19817 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16901), .A3(n16666), 
        .B1(n16653), .B2(n16850), .B3(n16652), .ZN(n16654) );
  INV_X1 U19818 ( .A(n16654), .ZN(n16655) );
  OAI21_X1 U19819 ( .B1(n16914), .B2(n16847), .A(n16655), .ZN(P3_U2683) );
  AOI22_X1 U19820 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16659) );
  AOI22_X1 U19821 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16658) );
  AOI22_X1 U19822 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16786), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16657) );
  AOI22_X1 U19823 ( .A1(n15236), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16656) );
  NAND4_X1 U19824 ( .A1(n16659), .A2(n16658), .A3(n16657), .A4(n16656), .ZN(
        n16665) );
  AOI22_X1 U19825 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16663) );
  AOI22_X1 U19826 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16662) );
  AOI22_X1 U19827 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16661) );
  AOI22_X1 U19828 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9586), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16660) );
  NAND4_X1 U19829 ( .A1(n16663), .A2(n16662), .A3(n16661), .A4(n16660), .ZN(
        n16664) );
  NOR2_X1 U19830 ( .A1(n16665), .A2(n16664), .ZN(n16919) );
  OAI211_X1 U19831 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16680), .A(n16666), .B(
        n16847), .ZN(n16667) );
  OAI21_X1 U19832 ( .B1(n16919), .B2(n16847), .A(n16667), .ZN(P3_U2684) );
  INV_X1 U19833 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16668) );
  NAND3_X1 U19834 ( .A1(n17864), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n16746), 
        .ZN(n16729) );
  NOR3_X1 U19835 ( .A1(n16668), .A2(n16730), .A3(n16729), .ZN(n16717) );
  AND2_X1 U19836 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16717), .ZN(n16704) );
  AND2_X1 U19837 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16704), .ZN(n16692) );
  AOI21_X1 U19838 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16847), .A(n16692), .ZN(
        n16679) );
  AOI22_X1 U19839 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14991), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16672) );
  AOI22_X1 U19840 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16671) );
  AOI22_X1 U19841 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16670) );
  AOI22_X1 U19842 ( .A1(n16780), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16669) );
  NAND4_X1 U19843 ( .A1(n16672), .A2(n16671), .A3(n16670), .A4(n16669), .ZN(
        n16678) );
  AOI22_X1 U19844 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16676) );
  AOI22_X1 U19845 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16675) );
  AOI22_X1 U19846 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16674) );
  AOI22_X1 U19847 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16673) );
  NAND4_X1 U19848 ( .A1(n16676), .A2(n16675), .A3(n16674), .A4(n16673), .ZN(
        n16677) );
  NOR2_X1 U19849 ( .A1(n16678), .A2(n16677), .ZN(n16924) );
  OAI22_X1 U19850 ( .A1(n16680), .A2(n16679), .B1(n16924), .B2(n16834), .ZN(
        P3_U2685) );
  AOI21_X1 U19851 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16847), .A(n16704), .ZN(
        n16691) );
  AOI22_X1 U19852 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16778), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16684) );
  AOI22_X1 U19853 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14991), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16683) );
  AOI22_X1 U19854 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16786), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16682) );
  AOI22_X1 U19855 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n16800), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n16780), .ZN(n16681) );
  NAND4_X1 U19856 ( .A1(n16684), .A2(n16683), .A3(n16682), .A4(n16681), .ZN(
        n16690) );
  AOI22_X1 U19857 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9592), .ZN(n16688) );
  AOI22_X1 U19858 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9589), .B1(n9591), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16687) );
  AOI22_X1 U19859 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9586), .ZN(n16686) );
  AOI22_X1 U19860 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15236), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16685) );
  NAND4_X1 U19861 ( .A1(n16688), .A2(n16687), .A3(n16686), .A4(n16685), .ZN(
        n16689) );
  NOR2_X1 U19862 ( .A1(n16690), .A2(n16689), .ZN(n16929) );
  OAI22_X1 U19863 ( .A1(n16692), .A2(n16691), .B1(n16929), .B2(n16834), .ZN(
        P3_U2686) );
  AOI21_X1 U19864 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n16847), .A(n16717), .ZN(
        n16703) );
  AOI22_X1 U19865 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16696) );
  AOI22_X1 U19866 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16695) );
  AOI22_X1 U19867 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16694) );
  AOI22_X1 U19868 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16693) );
  NAND4_X1 U19869 ( .A1(n16696), .A2(n16695), .A3(n16694), .A4(n16693), .ZN(
        n16702) );
  AOI22_X1 U19870 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16700) );
  AOI22_X1 U19871 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16699) );
  AOI22_X1 U19872 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16698) );
  AOI22_X1 U19873 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16697) );
  NAND4_X1 U19874 ( .A1(n16700), .A2(n16699), .A3(n16698), .A4(n16697), .ZN(
        n16701) );
  NOR2_X1 U19875 ( .A1(n16702), .A2(n16701), .ZN(n16935) );
  OAI22_X1 U19876 ( .A1(n16704), .A2(n16703), .B1(n16935), .B2(n16834), .ZN(
        P3_U2687) );
  NOR2_X1 U19877 ( .A1(n16730), .A2(n16705), .ZN(n16728) );
  OAI21_X1 U19878 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16728), .A(n16834), .ZN(
        n16716) );
  AOI22_X1 U19879 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9592), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16709) );
  AOI22_X1 U19880 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16708) );
  AOI22_X1 U19881 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16707) );
  AOI22_X1 U19882 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16706) );
  NAND4_X1 U19883 ( .A1(n16709), .A2(n16708), .A3(n16707), .A4(n16706), .ZN(
        n16715) );
  AOI22_X1 U19884 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16713) );
  AOI22_X1 U19885 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16796), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16712) );
  AOI22_X1 U19886 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16711) );
  AOI22_X1 U19887 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16710) );
  NAND4_X1 U19888 ( .A1(n16713), .A2(n16712), .A3(n16711), .A4(n16710), .ZN(
        n16714) );
  NOR2_X1 U19889 ( .A1(n16715), .A2(n16714), .ZN(n16939) );
  OAI22_X1 U19890 ( .A1(n16717), .A2(n16716), .B1(n16939), .B2(n16834), .ZN(
        P3_U2688) );
  AOI22_X1 U19891 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16727) );
  AOI22_X1 U19892 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16726) );
  AOI22_X1 U19893 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16796), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16718) );
  OAI21_X1 U19894 ( .B1(n9584), .B2(n20519), .A(n16718), .ZN(n16724) );
  AOI22_X1 U19895 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16722) );
  AOI22_X1 U19896 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16721) );
  AOI22_X1 U19897 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16720) );
  AOI22_X1 U19898 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16719) );
  NAND4_X1 U19899 ( .A1(n16722), .A2(n16721), .A3(n16720), .A4(n16719), .ZN(
        n16723) );
  AOI211_X1 U19900 ( .C1(n16800), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n16724), .B(n16723), .ZN(n16725) );
  NAND3_X1 U19901 ( .A1(n16727), .A2(n16726), .A3(n16725), .ZN(n16943) );
  AOI21_X1 U19902 ( .B1(n16730), .B2(n16729), .A(n16728), .ZN(n16731) );
  MUX2_X1 U19903 ( .A(n16943), .B(n16731), .S(n16834), .Z(P3_U2689) );
  AOI21_X1 U19904 ( .B1(n16732), .B2(n16757), .A(n16850), .ZN(n16733) );
  INV_X1 U19905 ( .A(n16733), .ZN(n16745) );
  AOI22_X1 U19906 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16738) );
  AOI22_X1 U19907 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16737) );
  AOI22_X1 U19908 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16736) );
  AOI22_X1 U19909 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16735) );
  NAND4_X1 U19910 ( .A1(n16738), .A2(n16737), .A3(n16736), .A4(n16735), .ZN(
        n16744) );
  AOI22_X1 U19911 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16742) );
  AOI22_X1 U19912 ( .A1(n16800), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16741) );
  AOI22_X1 U19913 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9592), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16740) );
  AOI22_X1 U19914 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16739) );
  NAND4_X1 U19915 ( .A1(n16742), .A2(n16741), .A3(n16740), .A4(n16739), .ZN(
        n16743) );
  NOR2_X1 U19916 ( .A1(n16744), .A2(n16743), .ZN(n16952) );
  OAI22_X1 U19917 ( .A1(n16746), .A2(n16745), .B1(n16952), .B2(n16834), .ZN(
        P3_U2691) );
  AOI22_X1 U19918 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16750) );
  AOI22_X1 U19919 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16796), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16749) );
  AOI22_X1 U19920 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16780), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16748) );
  AOI22_X1 U19921 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16747) );
  NAND4_X1 U19922 ( .A1(n16750), .A2(n16749), .A3(n16748), .A4(n16747), .ZN(
        n16756) );
  AOI22_X1 U19923 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16754) );
  AOI22_X1 U19924 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16753) );
  AOI22_X1 U19925 ( .A1(n16762), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16752) );
  AOI22_X1 U19926 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16751) );
  NAND4_X1 U19927 ( .A1(n16754), .A2(n16753), .A3(n16752), .A4(n16751), .ZN(
        n16755) );
  NOR2_X1 U19928 ( .A1(n16756), .A2(n16755), .ZN(n16955) );
  OAI21_X1 U19929 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16758), .A(n16757), .ZN(
        n16759) );
  AOI22_X1 U19930 ( .A1(n16850), .A2(n16955), .B1(n16759), .B2(n16847), .ZN(
        P3_U2692) );
  NAND2_X1 U19931 ( .A1(n16847), .A2(n16774), .ZN(n16793) );
  AOI22_X1 U19932 ( .A1(n16779), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16760), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16773) );
  AOI22_X1 U19933 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16772) );
  AOI22_X1 U19934 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16761) );
  OAI21_X1 U19935 ( .B1(n9584), .B2(n16843), .A(n16761), .ZN(n16770) );
  AOI22_X1 U19936 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16762), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16768) );
  AOI22_X1 U19937 ( .A1(n16763), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16767) );
  AOI22_X1 U19938 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16766) );
  AOI22_X1 U19939 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16764), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16765) );
  NAND4_X1 U19940 ( .A1(n16768), .A2(n16767), .A3(n16766), .A4(n16765), .ZN(
        n16769) );
  AOI211_X1 U19941 ( .C1(n16785), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n16770), .B(n16769), .ZN(n16771) );
  NAND3_X1 U19942 ( .A1(n16773), .A2(n16772), .A3(n16771), .ZN(n16958) );
  NOR3_X1 U19943 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16901), .A3(n16774), .ZN(
        n16775) );
  AOI21_X1 U19944 ( .B1(n16850), .B2(n16958), .A(n16775), .ZN(n16776) );
  OAI21_X1 U19945 ( .B1(n16777), .B2(n16793), .A(n16776), .ZN(P3_U2693) );
  AOI22_X1 U19946 ( .A1(n16619), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16784) );
  AOI22_X1 U19947 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n16764), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n16778), .ZN(n16783) );
  AOI22_X1 U19948 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9592), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n16796), .ZN(n16782) );
  AOI22_X1 U19949 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16780), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n16779), .ZN(n16781) );
  NAND4_X1 U19950 ( .A1(n16784), .A2(n16783), .A3(n16782), .A4(n16781), .ZN(
        n16792) );
  AOI22_X1 U19951 ( .A1(n16785), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n16800), .ZN(n16790) );
  AOI22_X1 U19952 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9588), .ZN(n16789) );
  AOI22_X1 U19953 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16786), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16788) );
  AOI22_X1 U19954 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9589), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n16802), .ZN(n16787) );
  NAND4_X1 U19955 ( .A1(n16790), .A2(n16789), .A3(n16788), .A4(n16787), .ZN(
        n16791) );
  NOR2_X1 U19956 ( .A1(n16792), .A2(n16791), .ZN(n16963) );
  NOR2_X1 U19957 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16816), .ZN(n16794) );
  OAI22_X1 U19958 ( .A1(n16963), .A2(n16834), .B1(n16794), .B2(n16793), .ZN(
        P3_U2694) );
  OAI21_X1 U19959 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16795), .A(n16834), .ZN(
        n16815) );
  AOI22_X1 U19960 ( .A1(n16796), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16813) );
  AOI22_X1 U19961 ( .A1(n16797), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16812) );
  AOI22_X1 U19962 ( .A1(n16764), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16778), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16798) );
  OAI21_X1 U19963 ( .B1(n9584), .B2(n16799), .A(n16798), .ZN(n16810) );
  AOI22_X1 U19964 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U19965 ( .A1(n16801), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16800), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16807) );
  AOI22_X1 U19966 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16806) );
  AOI22_X1 U19967 ( .A1(n16804), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16763), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16805) );
  NAND4_X1 U19968 ( .A1(n16808), .A2(n16807), .A3(n16806), .A4(n16805), .ZN(
        n16809) );
  AOI211_X1 U19969 ( .C1(n16779), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n16810), .B(n16809), .ZN(n16811) );
  NAND3_X1 U19970 ( .A1(n16813), .A2(n16812), .A3(n16811), .ZN(n16966) );
  INV_X1 U19971 ( .A(n16966), .ZN(n16814) );
  OAI22_X1 U19972 ( .A1(n16816), .A2(n16815), .B1(n16814), .B2(n16834), .ZN(
        P3_U2695) );
  NAND2_X1 U19973 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16817), .ZN(n16823) );
  INV_X1 U19974 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16822) );
  INV_X1 U19975 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16819) );
  NAND2_X1 U19976 ( .A1(n16818), .A2(n16845), .ZN(n16831) );
  NOR2_X1 U19977 ( .A1(n16819), .A2(n16831), .ZN(n16824) );
  NAND3_X1 U19978 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16824), .A3(n16820), .ZN(
        n16821) );
  OAI221_X1 U19979 ( .B1(n16850), .B2(n16823), .C1(n16847), .C2(n16822), .A(
        n16821), .ZN(P3_U2696) );
  AOI22_X1 U19980 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16826), .B1(n16824), .B2(
        n20629), .ZN(n16825) );
  AOI22_X1 U19981 ( .A1(n16850), .A2(n20519), .B1(n16825), .B2(n16847), .ZN(
        P3_U2697) );
  OAI21_X1 U19982 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16827), .A(n16826), .ZN(
        n16828) );
  AOI22_X1 U19983 ( .A1(n16850), .A2(n16829), .B1(n16828), .B2(n16847), .ZN(
        P3_U2698) );
  INV_X1 U19984 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16833) );
  NOR2_X1 U19985 ( .A1(n16830), .A2(n16852), .ZN(n16837) );
  OAI211_X1 U19986 ( .C1(n16837), .C2(P3_EBX_REG_4__SCAN_IN), .A(n16847), .B(
        n16831), .ZN(n16832) );
  OAI21_X1 U19987 ( .B1(n16847), .B2(n16833), .A(n16832), .ZN(P3_U2699) );
  AOI22_X1 U19988 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16847), .B1(n16838), .B2(
        n16845), .ZN(n16836) );
  INV_X1 U19989 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16835) );
  OAI22_X1 U19990 ( .A1(n16837), .A2(n16836), .B1(n16835), .B2(n16834), .ZN(
        P3_U2700) );
  NAND2_X1 U19991 ( .A1(n16838), .A2(n16845), .ZN(n16839) );
  OAI221_X1 U19992 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n16841), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n16840), .A(n16839), .ZN(n16842) );
  AOI22_X1 U19993 ( .A1(n16850), .A2(n16843), .B1(n16842), .B2(n16847), .ZN(
        P3_U2701) );
  INV_X1 U19994 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U19995 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n16849), .B1(n16845), .B2(
        n16844), .ZN(n16846) );
  OAI21_X1 U19996 ( .B1(n16848), .B2(n16847), .A(n16846), .ZN(P3_U2702) );
  AOI22_X1 U19997 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16850), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n16849), .ZN(n16851) );
  OAI21_X1 U19998 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n16852), .A(n16851), .ZN(
        P3_U2703) );
  INV_X1 U19999 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17004) );
  INV_X1 U20000 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17009) );
  INV_X1 U20001 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17111) );
  INV_X1 U20002 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17043) );
  INV_X1 U20003 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17046) );
  INV_X1 U20004 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17049) );
  INV_X1 U20005 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17051) );
  NOR4_X1 U20006 ( .A1(n17043), .A2(n17046), .A3(n17049), .A4(n17051), .ZN(
        n16853) );
  NAND4_X1 U20007 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(n16853), .ZN(n16941) );
  INV_X1 U20008 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17034) );
  INV_X1 U20009 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17036) );
  INV_X1 U20010 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17092) );
  NAND2_X1 U20011 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n16942) );
  NOR4_X1 U20012 ( .A1(n17034), .A2(n17036), .A3(n17092), .A4(n16942), .ZN(
        n16854) );
  NOR2_X2 U20013 ( .A1(n17111), .A2(n16944), .ZN(n16936) );
  INV_X1 U20014 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17015) );
  INV_X1 U20015 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17017) );
  NAND4_X1 U20016 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n16855)
         );
  NAND2_X1 U20017 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n16896), .ZN(n16895) );
  NAND2_X1 U20018 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n16891), .ZN(n16890) );
  NOR2_X2 U20019 ( .A1(n17009), .A2(n16885), .ZN(n16880) );
  NAND2_X1 U20020 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n16880), .ZN(n16876) );
  NAND2_X1 U20021 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n16864), .ZN(n16860) );
  NAND2_X1 U20022 ( .A1(n16860), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n16859) );
  NAND2_X1 U20023 ( .A1(n16857), .A2(n16996), .ZN(n16879) );
  NAND2_X1 U20024 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n16930), .ZN(n16858) );
  OAI221_X1 U20025 ( .B1(n16860), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n16859), 
        .C2(n16996), .A(n16858), .ZN(P3_U2704) );
  NAND2_X1 U20026 ( .A1(n17853), .A2(n16996), .ZN(n16905) );
  AOI22_X1 U20027 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16930), .ZN(n16862) );
  OAI211_X1 U20028 ( .C1(n16864), .C2(P3_EAX_REG_30__SCAN_IN), .A(n9610), .B(
        n16860), .ZN(n16861) );
  OAI211_X1 U20029 ( .C1(n16863), .C2(n16989), .A(n16862), .B(n16861), .ZN(
        P3_U2705) );
  INV_X1 U20030 ( .A(n16864), .ZN(n16866) );
  OAI21_X1 U20031 ( .B1(n16996), .B2(n17004), .A(n16871), .ZN(n16865) );
  AOI22_X1 U20032 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n16930), .B1(n16866), .B2(
        n16865), .ZN(n16869) );
  AOI22_X1 U20033 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n16931), .B1(n16867), .B2(
        n16993), .ZN(n16868) );
  NAND2_X1 U20034 ( .A1(n16869), .A2(n16868), .ZN(P3_U2706) );
  INV_X1 U20035 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20036 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n16930), .B1(n16870), .B2(
        n16993), .ZN(n16874) );
  OAI211_X1 U20037 ( .C1(n16872), .C2(P3_EAX_REG_28__SCAN_IN), .A(n9610), .B(
        n16871), .ZN(n16873) );
  OAI211_X1 U20038 ( .C1(n16905), .C2(n17100), .A(n16874), .B(n16873), .ZN(
        P3_U2707) );
  INV_X1 U20039 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U20040 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n16931), .B1(n16875), .B2(
        n16993), .ZN(n16878) );
  OAI211_X1 U20041 ( .C1(n16880), .C2(P3_EAX_REG_27__SCAN_IN), .A(n9610), .B(
        n16876), .ZN(n16877) );
  OAI211_X1 U20042 ( .C1(n16879), .C2(n17841), .A(n16878), .B(n16877), .ZN(
        P3_U2708) );
  AOI22_X1 U20043 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16930), .ZN(n16883) );
  AOI211_X1 U20044 ( .C1(n17009), .C2(n16885), .A(n16880), .B(n16996), .ZN(
        n16881) );
  INV_X1 U20045 ( .A(n16881), .ZN(n16882) );
  OAI211_X1 U20046 ( .C1(n16884), .C2(n16989), .A(n16883), .B(n16882), .ZN(
        P3_U2709) );
  AOI22_X1 U20047 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16930), .ZN(n16888) );
  OAI211_X1 U20048 ( .C1(n16886), .C2(P3_EAX_REG_25__SCAN_IN), .A(n9610), .B(
        n16885), .ZN(n16887) );
  OAI211_X1 U20049 ( .C1(n16889), .C2(n16989), .A(n16888), .B(n16887), .ZN(
        P3_U2710) );
  AOI22_X1 U20050 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16930), .ZN(n16893) );
  OAI211_X1 U20051 ( .C1(n16891), .C2(P3_EAX_REG_24__SCAN_IN), .A(n9610), .B(
        n16890), .ZN(n16892) );
  OAI211_X1 U20052 ( .C1(n16894), .C2(n16989), .A(n16893), .B(n16892), .ZN(
        P3_U2711) );
  AOI22_X1 U20053 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16930), .ZN(n16898) );
  OAI211_X1 U20054 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n16896), .A(n9610), .B(
        n16895), .ZN(n16897) );
  OAI211_X1 U20055 ( .C1(n16899), .C2(n16989), .A(n16898), .B(n16897), .ZN(
        P3_U2712) );
  INV_X1 U20056 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n17856) );
  AOI22_X1 U20057 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n16930), .B1(n16993), .B2(
        n16900), .ZN(n16904) );
  INV_X1 U20058 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17021) );
  NOR2_X1 U20059 ( .A1(n16901), .A2(n16932), .ZN(n16926) );
  NAND2_X1 U20060 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n16926), .ZN(n16925) );
  NAND2_X1 U20061 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n16915), .ZN(n16911) );
  NAND2_X1 U20062 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n16907), .ZN(n16906) );
  OAI21_X1 U20063 ( .B1(n17015), .B2(n16996), .A(n16906), .ZN(n16902) );
  OAI21_X1 U20064 ( .B1(n17015), .B2(n16906), .A(n16902), .ZN(n16903) );
  OAI211_X1 U20065 ( .C1(n17856), .C2(n16905), .A(n16904), .B(n16903), .ZN(
        P3_U2713) );
  AOI22_X1 U20066 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16930), .ZN(n16909) );
  OAI211_X1 U20067 ( .C1(n16907), .C2(P3_EAX_REG_21__SCAN_IN), .A(n9610), .B(
        n16906), .ZN(n16908) );
  OAI211_X1 U20068 ( .C1(n16910), .C2(n16989), .A(n16909), .B(n16908), .ZN(
        P3_U2714) );
  AOI22_X1 U20069 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16930), .ZN(n16913) );
  OAI211_X1 U20070 ( .C1(n16915), .C2(P3_EAX_REG_20__SCAN_IN), .A(n9610), .B(
        n16911), .ZN(n16912) );
  OAI211_X1 U20071 ( .C1(n16914), .C2(n16989), .A(n16913), .B(n16912), .ZN(
        P3_U2715) );
  AOI22_X1 U20072 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16930), .ZN(n16918) );
  AOI211_X1 U20073 ( .C1(n17021), .C2(n16920), .A(n16915), .B(n16996), .ZN(
        n16916) );
  INV_X1 U20074 ( .A(n16916), .ZN(n16917) );
  OAI211_X1 U20075 ( .C1(n16919), .C2(n16989), .A(n16918), .B(n16917), .ZN(
        P3_U2716) );
  AOI22_X1 U20076 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16930), .ZN(n16923) );
  OAI211_X1 U20077 ( .C1(n16921), .C2(P3_EAX_REG_18__SCAN_IN), .A(n9610), .B(
        n16920), .ZN(n16922) );
  OAI211_X1 U20078 ( .C1(n16924), .C2(n16989), .A(n16923), .B(n16922), .ZN(
        P3_U2717) );
  AOI22_X1 U20079 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16930), .ZN(n16928) );
  OAI211_X1 U20080 ( .C1(n16926), .C2(P3_EAX_REG_17__SCAN_IN), .A(n9610), .B(
        n16925), .ZN(n16927) );
  OAI211_X1 U20081 ( .C1(n16929), .C2(n16989), .A(n16928), .B(n16927), .ZN(
        P3_U2718) );
  AOI22_X1 U20082 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n16931), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16930), .ZN(n16934) );
  OAI211_X1 U20083 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n16936), .A(n9610), .B(
        n16932), .ZN(n16933) );
  OAI211_X1 U20084 ( .C1(n16935), .C2(n16989), .A(n16934), .B(n16933), .ZN(
        P3_U2719) );
  INV_X1 U20085 ( .A(n16992), .ZN(n16994) );
  AOI211_X1 U20086 ( .C1(n17111), .C2(n16944), .A(n16996), .B(n16936), .ZN(
        n16937) );
  AOI21_X1 U20087 ( .B1(n16994), .B2(BUF2_REG_15__SCAN_IN), .A(n16937), .ZN(
        n16938) );
  OAI21_X1 U20088 ( .B1(n16939), .B2(n16989), .A(n16938), .ZN(P3_U2720) );
  NAND2_X1 U20089 ( .A1(n17864), .A2(n16940), .ZN(n16999) );
  NOR2_X1 U20090 ( .A1(n16941), .A2(n16999), .ZN(n16973) );
  NAND2_X1 U20091 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n16973), .ZN(n16967) );
  NAND2_X1 U20092 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n16961), .ZN(n16951) );
  NOR2_X1 U20093 ( .A1(n17034), .A2(n16951), .ZN(n16954) );
  NAND2_X1 U20094 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n16954), .ZN(n16947) );
  AOI22_X1 U20095 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n16994), .B1(n16993), .B2(
        n16943), .ZN(n16946) );
  NAND3_X1 U20096 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n9610), .A3(n16944), .ZN(
        n16945) );
  OAI211_X1 U20097 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n16947), .A(n16946), .B(
        n16945), .ZN(P3_U2721) );
  INV_X1 U20098 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17104) );
  INV_X1 U20099 ( .A(n16947), .ZN(n16950) );
  AOI21_X1 U20100 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n9610), .A(n16954), .ZN(
        n16949) );
  OAI222_X1 U20101 ( .A1(n16992), .A2(n17104), .B1(n16950), .B2(n16949), .C1(
        n16989), .C2(n16948), .ZN(P3_U2722) );
  INV_X1 U20102 ( .A(n16951), .ZN(n16957) );
  AOI21_X1 U20103 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n9610), .A(n16957), .ZN(
        n16953) );
  OAI222_X1 U20104 ( .A1(n16992), .A2(n17100), .B1(n16954), .B2(n16953), .C1(
        n16989), .C2(n16952), .ZN(P3_U2723) );
  INV_X1 U20105 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17098) );
  AOI21_X1 U20106 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n9610), .A(n16961), .ZN(
        n16956) );
  OAI222_X1 U20107 ( .A1(n16992), .A2(n17098), .B1(n16957), .B2(n16956), .C1(
        n16989), .C2(n16955), .ZN(P3_U2724) );
  INV_X1 U20108 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17040) );
  NOR2_X1 U20109 ( .A1(n17040), .A2(n16967), .ZN(n16965) );
  OAI21_X1 U20110 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n16965), .A(n9610), .ZN(
        n16960) );
  AOI22_X1 U20111 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n16994), .B1(n16993), .B2(
        n16958), .ZN(n16959) );
  OAI21_X1 U20112 ( .B1(n16961), .B2(n16960), .A(n16959), .ZN(P3_U2725) );
  INV_X1 U20113 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17094) );
  OAI21_X1 U20114 ( .B1(n17040), .B2(n16996), .A(n16967), .ZN(n16962) );
  INV_X1 U20115 ( .A(n16962), .ZN(n16964) );
  OAI222_X1 U20116 ( .A1(n16992), .A2(n17094), .B1(n16965), .B2(n16964), .C1(
        n16989), .C2(n16963), .ZN(P3_U2726) );
  AOI22_X1 U20117 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n16994), .B1(n16993), .B2(
        n16966), .ZN(n16970) );
  OAI211_X1 U20118 ( .C1(n16968), .C2(P3_EAX_REG_8__SCAN_IN), .A(n9610), .B(
        n16967), .ZN(n16969) );
  NAND2_X1 U20119 ( .A1(n16970), .A2(n16969), .ZN(P3_U2727) );
  INV_X1 U20120 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n17861) );
  NAND2_X1 U20121 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n16971) );
  NOR2_X1 U20122 ( .A1(n16971), .A2(n16999), .ZN(n16991) );
  NAND2_X1 U20123 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n16991), .ZN(n16980) );
  NOR2_X1 U20124 ( .A1(n17051), .A2(n16980), .ZN(n16983) );
  NAND2_X1 U20125 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n16983), .ZN(n16974) );
  NOR2_X1 U20126 ( .A1(n17046), .A2(n16974), .ZN(n16975) );
  AOI21_X1 U20127 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n9610), .A(n16975), .ZN(
        n16972) );
  OAI222_X1 U20128 ( .A1(n16992), .A2(n17861), .B1(n16973), .B2(n16972), .C1(
        n16989), .C2(n17646), .ZN(P3_U2728) );
  INV_X1 U20129 ( .A(n16974), .ZN(n16978) );
  AOI21_X1 U20130 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n9610), .A(n16978), .ZN(
        n16976) );
  OAI222_X1 U20131 ( .A1(n16992), .A2(n17856), .B1(n16976), .B2(n16975), .C1(
        n16989), .C2(n9927), .ZN(P3_U2729) );
  INV_X1 U20132 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n17852) );
  AOI21_X1 U20133 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n9610), .A(n16983), .ZN(
        n16979) );
  OAI222_X1 U20134 ( .A1(n16992), .A2(n17852), .B1(n16979), .B2(n16978), .C1(
        n16989), .C2(n16977), .ZN(P3_U2730) );
  INV_X1 U20135 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n17847) );
  INV_X1 U20136 ( .A(n16980), .ZN(n16986) );
  AOI21_X1 U20137 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n9610), .A(n16986), .ZN(
        n16982) );
  OAI222_X1 U20138 ( .A1(n17847), .A2(n16992), .B1(n16983), .B2(n16982), .C1(
        n16989), .C2(n16981), .ZN(P3_U2731) );
  INV_X1 U20139 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17842) );
  AOI21_X1 U20140 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n9610), .A(n16991), .ZN(
        n16985) );
  OAI222_X1 U20141 ( .A1(n17842), .A2(n16992), .B1(n16986), .B2(n16985), .C1(
        n16989), .C2(n16984), .ZN(P3_U2732) );
  INV_X1 U20142 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n17837) );
  INV_X1 U20143 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17084) );
  INV_X1 U20144 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17055) );
  OAI22_X1 U20145 ( .A1(n16999), .A2(n17084), .B1(n17055), .B2(n16996), .ZN(
        n16987) );
  INV_X1 U20146 ( .A(n16987), .ZN(n16990) );
  OAI222_X1 U20147 ( .A1(n17837), .A2(n16992), .B1(n16991), .B2(n16990), .C1(
        n16989), .C2(n16988), .ZN(P3_U2733) );
  NAND3_X1 U20148 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n9610), .A3(n16995), .ZN(
        n16997) );
  OAI211_X1 U20149 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n16999), .A(n16998), .B(
        n16997), .ZN(P3_U2734) );
  NOR2_X1 U20150 ( .A1(n18429), .A2(n18334), .ZN(n17044) );
  CLKBUF_X1 U20151 ( .A(n17044), .Z(n18467) );
  AND2_X1 U20152 ( .A1(n17047), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20153 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17081) );
  NAND2_X1 U20154 ( .A1(n17028), .A2(n17001), .ZN(n17026) );
  AOI22_X1 U20155 ( .A1(n18467), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17002) );
  OAI21_X1 U20156 ( .B1(n17081), .B2(n17026), .A(n17002), .ZN(P3_U2737) );
  AOI22_X1 U20157 ( .A1(n18467), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17003) );
  OAI21_X1 U20158 ( .B1(n17004), .B2(n17026), .A(n17003), .ZN(P3_U2738) );
  INV_X1 U20159 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20600) );
  AOI22_X1 U20160 ( .A1(n18467), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17005) );
  OAI21_X1 U20161 ( .B1(n20600), .B2(n17026), .A(n17005), .ZN(P3_U2739) );
  INV_X1 U20162 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20163 ( .A1(n18467), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17006) );
  OAI21_X1 U20164 ( .B1(n17007), .B2(n17026), .A(n17006), .ZN(P3_U2740) );
  AOI22_X1 U20165 ( .A1(n18467), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17008) );
  OAI21_X1 U20166 ( .B1(n17009), .B2(n17026), .A(n17008), .ZN(P3_U2741) );
  INV_X1 U20167 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20168 ( .A1(n18467), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17010) );
  OAI21_X1 U20169 ( .B1(n17011), .B2(n17026), .A(n17010), .ZN(P3_U2742) );
  INV_X1 U20170 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20171 ( .A1(n18467), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17012) );
  OAI21_X1 U20172 ( .B1(n17074), .B2(n17026), .A(n17012), .ZN(P3_U2743) );
  INV_X1 U20173 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20628) );
  AOI22_X1 U20174 ( .A1(n18467), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17013) );
  OAI21_X1 U20175 ( .B1(n20628), .B2(n17026), .A(n17013), .ZN(P3_U2744) );
  AOI22_X1 U20176 ( .A1(n18467), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17014) );
  OAI21_X1 U20177 ( .B1(n17015), .B2(n17026), .A(n17014), .ZN(P3_U2745) );
  AOI22_X1 U20178 ( .A1(n17044), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17016) );
  OAI21_X1 U20179 ( .B1(n17017), .B2(n17026), .A(n17016), .ZN(P3_U2746) );
  INV_X1 U20180 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20181 ( .A1(n17044), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17018) );
  OAI21_X1 U20182 ( .B1(n17019), .B2(n17026), .A(n17018), .ZN(P3_U2747) );
  AOI22_X1 U20183 ( .A1(n17044), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17020) );
  OAI21_X1 U20184 ( .B1(n17021), .B2(n17026), .A(n17020), .ZN(P3_U2748) );
  INV_X1 U20185 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20186 ( .A1(n17044), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17022) );
  OAI21_X1 U20187 ( .B1(n17023), .B2(n17026), .A(n17022), .ZN(P3_U2749) );
  INV_X1 U20188 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20189 ( .A1(n17044), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17024) );
  OAI21_X1 U20190 ( .B1(n17066), .B2(n17026), .A(n17024), .ZN(P3_U2750) );
  INV_X1 U20191 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20192 ( .A1(n17044), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17025) );
  OAI21_X1 U20193 ( .B1(n17027), .B2(n17026), .A(n17025), .ZN(P3_U2751) );
  AOI22_X1 U20194 ( .A1(n17044), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17029) );
  OAI21_X1 U20195 ( .B1(n17111), .B2(n17059), .A(n17029), .ZN(P3_U2752) );
  INV_X1 U20196 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20197 ( .A1(n17044), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17030) );
  OAI21_X1 U20198 ( .B1(n17106), .B2(n17059), .A(n17030), .ZN(P3_U2753) );
  INV_X1 U20199 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20200 ( .A1(n17044), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17031) );
  OAI21_X1 U20201 ( .B1(n17032), .B2(n17059), .A(n17031), .ZN(P3_U2754) );
  AOI22_X1 U20202 ( .A1(n17044), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17033) );
  OAI21_X1 U20203 ( .B1(n17034), .B2(n17059), .A(n17033), .ZN(P3_U2755) );
  AOI22_X1 U20204 ( .A1(n18467), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17035) );
  OAI21_X1 U20205 ( .B1(n17036), .B2(n17059), .A(n17035), .ZN(P3_U2756) );
  INV_X1 U20206 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20207 ( .A1(n18467), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17037) );
  OAI21_X1 U20208 ( .B1(n17038), .B2(n17059), .A(n17037), .ZN(P3_U2757) );
  AOI22_X1 U20209 ( .A1(n18467), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17039) );
  OAI21_X1 U20210 ( .B1(n17040), .B2(n17059), .A(n17039), .ZN(P3_U2758) );
  AOI22_X1 U20211 ( .A1(n18467), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17041) );
  OAI21_X1 U20212 ( .B1(n17092), .B2(n17059), .A(n17041), .ZN(P3_U2759) );
  AOI22_X1 U20213 ( .A1(n18467), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17042) );
  OAI21_X1 U20214 ( .B1(n17043), .B2(n17059), .A(n17042), .ZN(P3_U2760) );
  AOI22_X1 U20215 ( .A1(n17044), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17045) );
  OAI21_X1 U20216 ( .B1(n17046), .B2(n17059), .A(n17045), .ZN(P3_U2761) );
  AOI22_X1 U20217 ( .A1(n18467), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17047), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17048) );
  OAI21_X1 U20218 ( .B1(n17049), .B2(n17059), .A(n17048), .ZN(P3_U2762) );
  AOI22_X1 U20219 ( .A1(n18467), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17050) );
  OAI21_X1 U20220 ( .B1(n17051), .B2(n17059), .A(n17050), .ZN(P3_U2763) );
  INV_X1 U20221 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20222 ( .A1(n18467), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17052) );
  OAI21_X1 U20223 ( .B1(n17053), .B2(n17059), .A(n17052), .ZN(P3_U2764) );
  AOI22_X1 U20224 ( .A1(n18467), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17054) );
  OAI21_X1 U20225 ( .B1(n17055), .B2(n17059), .A(n17054), .ZN(P3_U2765) );
  AOI22_X1 U20226 ( .A1(n18467), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17056) );
  OAI21_X1 U20227 ( .B1(n17084), .B2(n17059), .A(n17056), .ZN(P3_U2766) );
  AOI22_X1 U20228 ( .A1(n18467), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17057), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17058) );
  OAI21_X1 U20229 ( .B1(n17060), .B2(n17059), .A(n17058), .ZN(P3_U2767) );
  AOI211_X1 U20230 ( .C1(n18473), .C2(n18472), .A(n17063), .B(n17062), .ZN(
        n17061) );
  INV_X2 U20231 ( .A(n17061), .ZN(n17107) );
  OR3_X1 U20232 ( .A1(n18472), .A2(n17063), .A3(n17062), .ZN(n17110) );
  AOI22_X1 U20233 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17107), .ZN(n17064) );
  OAI21_X1 U20234 ( .B1(n17824), .B2(n17103), .A(n17064), .ZN(P3_U2768) );
  AOI22_X1 U20235 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17108), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17107), .ZN(n17065) );
  OAI21_X1 U20236 ( .B1(n17066), .B2(n17110), .A(n17065), .ZN(P3_U2769) );
  AOI22_X1 U20237 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17107), .ZN(n17067) );
  OAI21_X1 U20238 ( .B1(n17837), .B2(n17103), .A(n17067), .ZN(P3_U2770) );
  AOI22_X1 U20239 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17107), .ZN(n17068) );
  OAI21_X1 U20240 ( .B1(n17842), .B2(n17103), .A(n17068), .ZN(P3_U2771) );
  AOI22_X1 U20241 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17107), .ZN(n17069) );
  OAI21_X1 U20242 ( .B1(n17847), .B2(n17103), .A(n17069), .ZN(P3_U2772) );
  AOI22_X1 U20243 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17107), .ZN(n17070) );
  OAI21_X1 U20244 ( .B1(n17852), .B2(n17103), .A(n17070), .ZN(P3_U2773) );
  AOI22_X1 U20245 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17107), .ZN(n17071) );
  OAI21_X1 U20246 ( .B1(n17856), .B2(n17103), .A(n17071), .ZN(P3_U2774) );
  AOI22_X1 U20247 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17107), .ZN(n17072) );
  OAI21_X1 U20248 ( .B1(n17861), .B2(n17103), .A(n17072), .ZN(P3_U2775) );
  AOI22_X1 U20249 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17108), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17107), .ZN(n17073) );
  OAI21_X1 U20250 ( .B1(n17074), .B2(n17110), .A(n17073), .ZN(P3_U2776) );
  AOI22_X1 U20251 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17107), .ZN(n17075) );
  OAI21_X1 U20252 ( .B1(n17094), .B2(n17103), .A(n17075), .ZN(P3_U2777) );
  INV_X1 U20253 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20254 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17107), .ZN(n17076) );
  OAI21_X1 U20255 ( .B1(n17096), .B2(n17103), .A(n17076), .ZN(P3_U2778) );
  AOI22_X1 U20256 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17107), .ZN(n17077) );
  OAI21_X1 U20257 ( .B1(n17098), .B2(n17103), .A(n17077), .ZN(P3_U2779) );
  AOI22_X1 U20258 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17107), .ZN(n17078) );
  OAI21_X1 U20259 ( .B1(n17100), .B2(n17103), .A(n17078), .ZN(P3_U2780) );
  AOI22_X1 U20260 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17101), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17107), .ZN(n17079) );
  OAI21_X1 U20261 ( .B1(n17104), .B2(n17103), .A(n17079), .ZN(P3_U2781) );
  AOI22_X1 U20262 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17108), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17107), .ZN(n17080) );
  OAI21_X1 U20263 ( .B1(n17081), .B2(n17110), .A(n17080), .ZN(P3_U2782) );
  AOI22_X1 U20264 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17107), .ZN(n17082) );
  OAI21_X1 U20265 ( .B1(n17824), .B2(n17103), .A(n17082), .ZN(P3_U2783) );
  AOI22_X1 U20266 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17108), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17107), .ZN(n17083) );
  OAI21_X1 U20267 ( .B1(n17084), .B2(n17110), .A(n17083), .ZN(P3_U2784) );
  AOI22_X1 U20268 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17107), .ZN(n17085) );
  OAI21_X1 U20269 ( .B1(n17837), .B2(n17103), .A(n17085), .ZN(P3_U2785) );
  AOI22_X1 U20270 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17107), .ZN(n17086) );
  OAI21_X1 U20271 ( .B1(n17842), .B2(n17103), .A(n17086), .ZN(P3_U2786) );
  AOI22_X1 U20272 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17107), .ZN(n17087) );
  OAI21_X1 U20273 ( .B1(n17847), .B2(n17103), .A(n17087), .ZN(P3_U2787) );
  AOI22_X1 U20274 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17107), .ZN(n17088) );
  OAI21_X1 U20275 ( .B1(n17852), .B2(n17103), .A(n17088), .ZN(P3_U2788) );
  AOI22_X1 U20276 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17107), .ZN(n17089) );
  OAI21_X1 U20277 ( .B1(n17856), .B2(n17103), .A(n17089), .ZN(P3_U2789) );
  AOI22_X1 U20278 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17107), .ZN(n17090) );
  OAI21_X1 U20279 ( .B1(n17861), .B2(n17103), .A(n17090), .ZN(P3_U2790) );
  AOI22_X1 U20280 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17108), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17107), .ZN(n17091) );
  OAI21_X1 U20281 ( .B1(n17092), .B2(n17110), .A(n17091), .ZN(P3_U2791) );
  AOI22_X1 U20282 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17107), .ZN(n17093) );
  OAI21_X1 U20283 ( .B1(n17094), .B2(n17103), .A(n17093), .ZN(P3_U2792) );
  AOI22_X1 U20284 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17107), .ZN(n17095) );
  OAI21_X1 U20285 ( .B1(n17096), .B2(n17103), .A(n17095), .ZN(P3_U2793) );
  AOI22_X1 U20286 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17107), .ZN(n17097) );
  OAI21_X1 U20287 ( .B1(n17098), .B2(n17103), .A(n17097), .ZN(P3_U2794) );
  AOI22_X1 U20288 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17107), .ZN(n17099) );
  OAI21_X1 U20289 ( .B1(n17100), .B2(n17103), .A(n17099), .ZN(P3_U2795) );
  AOI22_X1 U20290 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17101), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17107), .ZN(n17102) );
  OAI21_X1 U20291 ( .B1(n17104), .B2(n17103), .A(n17102), .ZN(P3_U2796) );
  AOI22_X1 U20292 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17108), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17107), .ZN(n17105) );
  OAI21_X1 U20293 ( .B1(n17106), .B2(n17110), .A(n17105), .ZN(P3_U2797) );
  AOI22_X1 U20294 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17108), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17107), .ZN(n17109) );
  OAI21_X1 U20295 ( .B1(n17111), .B2(n17110), .A(n17109), .ZN(P3_U2798) );
  AOI21_X1 U20296 ( .B1(n17125), .B2(n17318), .A(n17457), .ZN(n17112) );
  INV_X1 U20297 ( .A(n17112), .ZN(n17113) );
  AOI21_X1 U20298 ( .B1(n17240), .B2(n17114), .A(n17113), .ZN(n17149) );
  OAI21_X1 U20299 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17267), .A(
        n17149), .ZN(n17135) );
  AOI22_X1 U20300 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17135), .B1(
        n17285), .B2(n17115), .ZN(n17130) );
  NOR2_X1 U20301 ( .A1(n9601), .A2(n17399), .ZN(n17232) );
  INV_X1 U20302 ( .A(n17116), .ZN(n17498) );
  OAI22_X1 U20303 ( .A1(n17497), .A2(n17492), .B1(n17498), .B2(n17117), .ZN(
        n17152) );
  NOR2_X1 U20304 ( .A1(n9925), .A2(n17152), .ZN(n17142) );
  NOR3_X1 U20305 ( .A1(n17232), .A2(n17142), .A3(n17118), .ZN(n17123) );
  AOI211_X1 U20306 ( .C1(n17121), .C2(n17120), .A(n17119), .B(n17402), .ZN(
        n17122) );
  AOI211_X1 U20307 ( .C1(n17124), .C2(n17212), .A(n17123), .B(n17122), .ZN(
        n17129) );
  NAND2_X1 U20308 ( .A1(n9597), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17128) );
  NOR2_X1 U20309 ( .A1(n17322), .A2(n17125), .ZN(n17139) );
  OAI211_X1 U20310 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17139), .B(n17126), .ZN(n17127) );
  NAND4_X1 U20311 ( .A1(n17130), .A2(n17129), .A3(n17128), .A4(n17127), .ZN(
        P3_U2802) );
  NOR2_X1 U20312 ( .A1(n17132), .A2(n17131), .ZN(n17133) );
  XOR2_X1 U20313 ( .A(n17133), .B(n17388), .Z(n17505) );
  AOI22_X1 U20314 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17135), .B1(
        n17285), .B2(n17134), .ZN(n17136) );
  NAND2_X1 U20315 ( .A1(n9597), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17503) );
  OAI211_X1 U20316 ( .C1(n17505), .C2(n17402), .A(n17136), .B(n17503), .ZN(
        n17137) );
  AOI21_X1 U20317 ( .B1(n17139), .B2(n17138), .A(n17137), .ZN(n17140) );
  OAI221_X1 U20318 ( .B1(n17142), .B2(n9925), .C1(n17142), .C2(n17141), .A(
        n17140), .ZN(P3_U2803) );
  AOI21_X1 U20319 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17144), .A(
        n17143), .ZN(n17515) );
  NAND2_X1 U20320 ( .A1(n17555), .A2(n17212), .ZN(n17211) );
  NOR4_X1 U20321 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17531), .A3(
        n17506), .A4(n17211), .ZN(n17151) );
  AOI21_X1 U20322 ( .B1(n17145), .B2(n18205), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17148) );
  OAI21_X1 U20323 ( .B1(n17285), .B2(n15985), .A(n17146), .ZN(n17147) );
  NAND2_X1 U20324 ( .A1(n9597), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17513) );
  OAI211_X1 U20325 ( .C1(n17149), .C2(n17148), .A(n17147), .B(n17513), .ZN(
        n17150) );
  AOI211_X1 U20326 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17152), .A(
        n17151), .B(n17150), .ZN(n17153) );
  OAI21_X1 U20327 ( .B1(n17515), .B2(n17402), .A(n17153), .ZN(P3_U2804) );
  XOR2_X1 U20328 ( .A(n17154), .B(n17531), .Z(n17521) );
  AND2_X1 U20329 ( .A1(n17156), .A2(n18205), .ZN(n17194) );
  AOI211_X1 U20330 ( .C1(n17240), .C2(n17155), .A(n17457), .B(n17194), .ZN(
        n17188) );
  OAI21_X1 U20331 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17267), .A(
        n17188), .ZN(n17170) );
  NOR2_X1 U20332 ( .A1(n17322), .A2(n17156), .ZN(n17172) );
  OAI211_X1 U20333 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17172), .B(n17157), .ZN(n17158) );
  NAND2_X1 U20334 ( .A1(n9597), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17529) );
  OAI211_X1 U20335 ( .C1(n17346), .C2(n17159), .A(n17158), .B(n17529), .ZN(
        n17160) );
  AOI21_X1 U20336 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17170), .A(
        n17160), .ZN(n17167) );
  AOI21_X1 U20337 ( .B1(n17531), .B2(n17162), .A(n17161), .ZN(n17522) );
  AOI21_X1 U20338 ( .B1(n17164), .B2(n17359), .A(n17163), .ZN(n17165) );
  XOR2_X1 U20339 ( .A(n17165), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17527) );
  AOI22_X1 U20340 ( .A1(n17399), .A2(n17522), .B1(n17342), .B2(n17527), .ZN(
        n17166) );
  OAI211_X1 U20341 ( .C1(n17492), .C2(n17521), .A(n17167), .B(n17166), .ZN(
        P3_U2805) );
  INV_X1 U20342 ( .A(n17168), .ZN(n17181) );
  NOR2_X1 U20343 ( .A1(n17712), .A2(n20587), .ZN(n17169) );
  AOI221_X1 U20344 ( .B1(n17172), .B2(n17171), .C1(n17170), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17169), .ZN(n17180) );
  NOR2_X1 U20345 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17173), .ZN(
        n17532) );
  INV_X1 U20346 ( .A(n17536), .ZN(n17174) );
  AOI22_X1 U20347 ( .A1(n9601), .A2(n17533), .B1(n17399), .B2(n17174), .ZN(
        n17189) );
  AOI21_X1 U20348 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17176), .A(
        n17175), .ZN(n17543) );
  OAI22_X1 U20349 ( .A1(n17189), .A2(n17177), .B1(n17543), .B2(n17402), .ZN(
        n17178) );
  AOI21_X1 U20350 ( .B1(n17212), .B2(n17532), .A(n17178), .ZN(n17179) );
  OAI211_X1 U20351 ( .C1(n17346), .C2(n17181), .A(n17180), .B(n17179), .ZN(
        P3_U2806) );
  AOI22_X1 U20352 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17359), .B1(
        n17182), .B2(n17204), .ZN(n17183) );
  NAND2_X1 U20353 ( .A1(n17205), .A2(n17183), .ZN(n17184) );
  XOR2_X1 U20354 ( .A(n17184), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17551) );
  NAND2_X1 U20355 ( .A1(n9597), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17550) );
  OAI21_X1 U20356 ( .B1(n17285), .B2(n15985), .A(n17185), .ZN(n17186) );
  OAI211_X1 U20357 ( .C1(n17188), .C2(n17187), .A(n17550), .B(n17186), .ZN(
        n17193) );
  NOR2_X1 U20358 ( .A1(n20633), .A2(n17211), .ZN(n17191) );
  INV_X1 U20359 ( .A(n17189), .ZN(n17190) );
  MUX2_X1 U20360 ( .A(n17191), .B(n17190), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17192) );
  AOI211_X1 U20361 ( .C1(n17195), .C2(n17194), .A(n17193), .B(n17192), .ZN(
        n17196) );
  OAI21_X1 U20362 ( .B1(n17402), .B2(n17551), .A(n17196), .ZN(P3_U2807) );
  OAI21_X1 U20363 ( .B1(n17197), .B2(n18334), .A(n17488), .ZN(n17198) );
  AOI21_X1 U20364 ( .B1(n17318), .B2(n17199), .A(n17198), .ZN(n17229) );
  OAI21_X1 U20365 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17267), .A(
        n17229), .ZN(n17216) );
  NOR2_X1 U20366 ( .A1(n17322), .A2(n17199), .ZN(n17218) );
  OAI211_X1 U20367 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17218), .B(n17200), .ZN(n17201) );
  NAND2_X1 U20368 ( .A1(n9597), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17565) );
  OAI211_X1 U20369 ( .C1(n17346), .C2(n17202), .A(n17201), .B(n17565), .ZN(
        n17203) );
  AOI21_X1 U20370 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17216), .A(
        n17203), .ZN(n17210) );
  INV_X1 U20371 ( .A(n9650), .ZN(n17639) );
  AOI22_X1 U20372 ( .A1(n9601), .A2(n17639), .B1(n17399), .B2(n17631), .ZN(
        n17291) );
  OAI21_X1 U20373 ( .B1(n17555), .B2(n17232), .A(n17291), .ZN(n17222) );
  INV_X1 U20374 ( .A(n17204), .ZN(n17206) );
  OAI21_X1 U20375 ( .B1(n17207), .B2(n17206), .A(n17205), .ZN(n17208) );
  XOR2_X1 U20376 ( .A(n17208), .B(n20633), .Z(n17564) );
  AOI22_X1 U20377 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17222), .B1(
        n17342), .B2(n17564), .ZN(n17209) );
  OAI211_X1 U20378 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17211), .A(
        n17210), .B(n17209), .ZN(P3_U2808) );
  NAND2_X1 U20379 ( .A1(n17573), .A2(n17556), .ZN(n17578) );
  INV_X1 U20380 ( .A(n17553), .ZN(n17569) );
  NAND2_X1 U20381 ( .A1(n17569), .A2(n17212), .ZN(n17253) );
  INV_X1 U20382 ( .A(n17213), .ZN(n17214) );
  OAI22_X1 U20383 ( .A1(n17712), .A2(n18388), .B1(n17346), .B2(n17214), .ZN(
        n17215) );
  AOI221_X1 U20384 ( .B1(n17218), .B2(n17217), .C1(n17216), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17215), .ZN(n17224) );
  NAND3_X1 U20385 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17388), .A3(
        n17219), .ZN(n17234) );
  INV_X1 U20386 ( .A(n17234), .ZN(n17247) );
  AOI22_X1 U20387 ( .A1(n17573), .A2(n17247), .B1(n17263), .B2(n17220), .ZN(
        n17221) );
  XOR2_X1 U20388 ( .A(n17556), .B(n17221), .Z(n17568) );
  AOI22_X1 U20389 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17222), .B1(
        n17342), .B2(n17568), .ZN(n17223) );
  OAI211_X1 U20390 ( .C1(n17578), .C2(n17253), .A(n17224), .B(n17223), .ZN(
        P3_U2809) );
  NAND2_X1 U20391 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17225), .ZN(
        n17585) );
  NAND2_X1 U20392 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17242) );
  NOR4_X1 U20393 ( .A1(n17226), .A2(n17266), .A3(n17242), .A4(n18019), .ZN(
        n17227) );
  NOR2_X1 U20394 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17227), .ZN(
        n17228) );
  OAI22_X1 U20395 ( .A1(n17229), .A2(n17228), .B1(n17712), .B2(n18387), .ZN(
        n17230) );
  AOI221_X1 U20396 ( .B1(n17285), .B2(n17231), .C1(n15985), .C2(n17231), .A(
        n17230), .ZN(n17238) );
  NOR2_X1 U20397 ( .A1(n17553), .A2(n17249), .ZN(n17580) );
  OAI21_X1 U20398 ( .B1(n17232), .B2(n17580), .A(n17291), .ZN(n17250) );
  AOI221_X1 U20399 ( .B1(n17249), .B2(n17235), .C1(n17234), .C2(n17235), .A(
        n17233), .ZN(n17236) );
  XOR2_X1 U20400 ( .A(n17236), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n17579) );
  AOI22_X1 U20401 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17250), .B1(
        n17342), .B2(n17579), .ZN(n17237) );
  OAI211_X1 U20402 ( .C1(n17585), .C2(n17253), .A(n17238), .B(n17237), .ZN(
        P3_U2810) );
  INV_X1 U20403 ( .A(n17318), .ZN(n17456) );
  OAI21_X1 U20404 ( .B1(n17241), .B2(n17456), .A(n17488), .ZN(n17271) );
  AOI21_X1 U20405 ( .B1(n17240), .B2(n17239), .A(n17271), .ZN(n17255) );
  AND2_X1 U20406 ( .A1(n17279), .A2(n17241), .ZN(n17260) );
  OAI211_X1 U20407 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17260), .B(n17242), .ZN(n17243) );
  NAND2_X1 U20408 ( .A1(n9597), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17588) );
  OAI211_X1 U20409 ( .C1(n17255), .C2(n17244), .A(n17243), .B(n17588), .ZN(
        n17245) );
  AOI21_X1 U20410 ( .B1(n17285), .B2(n17246), .A(n17245), .ZN(n17252) );
  AOI21_X1 U20411 ( .B1(n17261), .B2(n17263), .A(n17247), .ZN(n17248) );
  XOR2_X1 U20412 ( .A(n17249), .B(n17248), .Z(n17586) );
  AOI22_X1 U20413 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17250), .B1(
        n17342), .B2(n17586), .ZN(n17251) );
  OAI211_X1 U20414 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17253), .A(
        n17252), .B(n17251), .ZN(P3_U2811) );
  NAND2_X1 U20415 ( .A1(n17599), .A2(n17254), .ZN(n17606) );
  INV_X1 U20416 ( .A(n17255), .ZN(n17258) );
  NAND2_X1 U20417 ( .A1(n9597), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17604) );
  OAI21_X1 U20418 ( .B1(n17346), .B2(n17256), .A(n17604), .ZN(n17257) );
  AOI221_X1 U20419 ( .B1(n17260), .B2(n17259), .C1(n17258), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17257), .ZN(n17265) );
  OAI21_X1 U20420 ( .B1(n17599), .B2(n17292), .A(n17291), .ZN(n17274) );
  AOI21_X1 U20421 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17388), .A(
        n17261), .ZN(n17262) );
  XOR2_X1 U20422 ( .A(n17263), .B(n17262), .Z(n17602) );
  AOI22_X1 U20423 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17274), .B1(
        n17342), .B2(n17602), .ZN(n17264) );
  OAI211_X1 U20424 ( .C1(n17292), .C2(n17606), .A(n17265), .B(n17264), .ZN(
        P3_U2812) );
  NAND2_X1 U20425 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17607), .ZN(
        n17613) );
  NOR2_X1 U20426 ( .A1(n17266), .A2(n18019), .ZN(n17270) );
  NAND2_X1 U20427 ( .A1(n9597), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17611) );
  OAI21_X1 U20428 ( .B1(n17471), .B2(n17268), .A(n17611), .ZN(n17269) );
  AOI221_X1 U20429 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17271), .C1(
        n17270), .C2(n17271), .A(n17269), .ZN(n17276) );
  OAI21_X1 U20430 ( .B1(n17273), .B2(n17607), .A(n17272), .ZN(n17610) );
  AOI22_X1 U20431 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17274), .B1(
        n17342), .B2(n17610), .ZN(n17275) );
  OAI211_X1 U20432 ( .C1(n17292), .C2(n17613), .A(n17276), .B(n17275), .ZN(
        P3_U2813) );
  NAND2_X1 U20433 ( .A1(n17388), .A2(n17689), .ZN(n17378) );
  OAI22_X1 U20434 ( .A1(n17378), .A2(n17494), .B1(n17277), .B2(n17388), .ZN(
        n17278) );
  XOR2_X1 U20435 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17278), .Z(
        n17621) );
  NAND2_X1 U20436 ( .A1(n17281), .A2(n17279), .ZN(n17295) );
  OAI21_X1 U20437 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17280), .ZN(n17288) );
  OAI21_X1 U20438 ( .B1(n17456), .B2(n17281), .A(n17488), .ZN(n17282) );
  INV_X1 U20439 ( .A(n17282), .ZN(n17307) );
  OAI21_X1 U20440 ( .B1(n17283), .B2(n18334), .A(n17307), .ZN(n17297) );
  AOI22_X1 U20441 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17297), .B1(
        n17285), .B2(n17284), .ZN(n17287) );
  NAND2_X1 U20442 ( .A1(n9597), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17286) );
  OAI211_X1 U20443 ( .C1(n17295), .C2(n17288), .A(n17287), .B(n17286), .ZN(
        n17289) );
  AOI21_X1 U20444 ( .B1(n17342), .B2(n17621), .A(n17289), .ZN(n17290) );
  OAI221_X1 U20445 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17292), 
        .C1(n17624), .C2(n17291), .A(n17290), .ZN(P3_U2814) );
  NAND2_X1 U20446 ( .A1(n17647), .A2(n17689), .ZN(n17668) );
  NOR2_X1 U20447 ( .A1(n17293), .A2(n17668), .ZN(n17311) );
  NOR2_X1 U20448 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17311), .ZN(
        n17633) );
  NAND2_X1 U20449 ( .A1(n17399), .A2(n17631), .ZN(n17304) );
  NOR2_X1 U20450 ( .A1(n17712), .A2(n18377), .ZN(n17626) );
  OAI22_X1 U20451 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17295), .B1(
        n17294), .B2(n17346), .ZN(n17296) );
  AOI211_X1 U20452 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17297), .A(
        n17626), .B(n17296), .ZN(n17303) );
  NAND2_X1 U20453 ( .A1(n17359), .A2(n17387), .ZN(n17379) );
  INV_X1 U20454 ( .A(n17379), .ZN(n17348) );
  NAND3_X1 U20455 ( .A1(n17349), .A2(n17348), .A3(n17660), .ZN(n17336) );
  INV_X1 U20456 ( .A(n17336), .ZN(n17312) );
  INV_X1 U20457 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U20458 ( .A1(n17689), .A2(n17298), .B1(n17312), .B2(n17332), .ZN(
        n17299) );
  AOI221_X1 U20459 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17685), 
        .C1(n17359), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17299), .ZN(
        n17300) );
  XOR2_X1 U20460 ( .A(n17300), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n17636) );
  NOR2_X1 U20461 ( .A1(n9650), .A2(n17492), .ZN(n17301) );
  NAND2_X1 U20462 ( .A1(n17305), .A2(n17616), .ZN(n17638) );
  AOI22_X1 U20463 ( .A1(n17342), .A2(n17636), .B1(n17301), .B2(n17638), .ZN(
        n17302) );
  OAI211_X1 U20464 ( .C1(n17633), .C2(n17304), .A(n17303), .B(n17302), .ZN(
        P3_U2815) );
  OAI221_X1 U20465 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17665), .A(n17305), .ZN(
        n17659) );
  NOR3_X1 U20466 ( .A1(n17421), .A2(n17422), .A3(n18019), .ZN(n17407) );
  NAND2_X1 U20467 ( .A1(n17306), .A2(n17407), .ZN(n17355) );
  AOI221_X1 U20468 ( .B1(n17323), .B2(n17308), .C1(n17355), .C2(n17308), .A(
        n17307), .ZN(n17309) );
  NOR2_X1 U20469 ( .A1(n17712), .A2(n18376), .ZN(n17657) );
  AOI211_X1 U20470 ( .C1(n17310), .C2(n17480), .A(n17309), .B(n17657), .ZN(
        n17317) );
  INV_X1 U20471 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17648) );
  NAND2_X1 U20472 ( .A1(n17647), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17628) );
  AOI221_X1 U20473 ( .B1(n17356), .B2(n17648), .C1(n17628), .C2(n17648), .A(
        n17311), .ZN(n17643) );
  NOR2_X1 U20474 ( .A1(n17329), .A2(n17378), .ZN(n17314) );
  AOI22_X1 U20475 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17314), .B1(
        n17313), .B2(n17312), .ZN(n17315) );
  XOR2_X1 U20476 ( .A(n17648), .B(n17315), .Z(n17645) );
  AOI22_X1 U20477 ( .A1(n17399), .A2(n17643), .B1(n17342), .B2(n17645), .ZN(
        n17316) );
  OAI211_X1 U20478 ( .C1(n17492), .C2(n17659), .A(n17317), .B(n17316), .ZN(
        P3_U2816) );
  AOI22_X1 U20479 ( .A1(n9601), .A2(n9761), .B1(n17399), .B2(n17668), .ZN(
        n17338) );
  NAND2_X1 U20480 ( .A1(n17318), .A2(n17321), .ZN(n17319) );
  OAI211_X1 U20481 ( .C1(n17320), .C2(n18334), .A(n17319), .B(n17488), .ZN(
        n17335) );
  NOR2_X1 U20482 ( .A1(n17322), .A2(n17321), .ZN(n17334) );
  OAI211_X1 U20483 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17334), .B(n17323), .ZN(n17325) );
  NAND2_X1 U20484 ( .A1(n9597), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17324) );
  OAI211_X1 U20485 ( .C1(n17346), .C2(n17326), .A(n17325), .B(n17324), .ZN(
        n17327) );
  AOI21_X1 U20486 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17335), .A(
        n17327), .ZN(n17331) );
  OAI22_X1 U20487 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17336), .B1(
        n17378), .B2(n17329), .ZN(n17328) );
  XNOR2_X1 U20488 ( .A(n17332), .B(n17328), .ZN(n17671) );
  NOR2_X1 U20489 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17329), .ZN(
        n17670) );
  AOI22_X1 U20490 ( .A1(n17342), .A2(n17671), .B1(n17670), .B2(n17383), .ZN(
        n17330) );
  OAI211_X1 U20491 ( .C1(n17338), .C2(n17332), .A(n17331), .B(n17330), .ZN(
        P3_U2817) );
  NOR2_X1 U20492 ( .A1(n17712), .A2(n18371), .ZN(n17682) );
  AOI221_X1 U20493 ( .B1(n17335), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C1(
        n17334), .C2(n17333), .A(n17682), .ZN(n17344) );
  NOR2_X1 U20494 ( .A1(n17662), .A2(n17378), .ZN(n17347) );
  INV_X1 U20495 ( .A(n17347), .ZN(n17361) );
  OAI21_X1 U20496 ( .B1(n17660), .B2(n17361), .A(n17336), .ZN(n17337) );
  XOR2_X1 U20497 ( .A(n17337), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17680) );
  INV_X1 U20498 ( .A(n17383), .ZN(n17365) );
  NOR2_X1 U20499 ( .A1(n17365), .A2(n17676), .ZN(n17340) );
  INV_X1 U20500 ( .A(n17338), .ZN(n17339) );
  MUX2_X1 U20501 ( .A(n17340), .B(n17339), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17341) );
  AOI21_X1 U20502 ( .B1(n17342), .B2(n17680), .A(n17341), .ZN(n17343) );
  OAI211_X1 U20503 ( .C1(n17346), .C2(n17345), .A(n17344), .B(n17343), .ZN(
        P3_U2818) );
  AOI21_X1 U20504 ( .B1(n17349), .B2(n17348), .A(n17347), .ZN(n17350) );
  XOR2_X1 U20505 ( .A(n17350), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n17700) );
  INV_X1 U20506 ( .A(n17407), .ZN(n17374) );
  NOR3_X1 U20507 ( .A1(n17394), .A2(n17375), .A3(n17374), .ZN(n17366) );
  NAND2_X1 U20508 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17366), .ZN(
        n17369) );
  OAI21_X1 U20509 ( .B1(n17485), .B2(n17351), .A(n17369), .ZN(n17354) );
  OAI22_X1 U20510 ( .A1(n17471), .A2(n17352), .B1(n17712), .B2(n18369), .ZN(
        n17353) );
  AOI21_X1 U20511 ( .B1(n17355), .B2(n17354), .A(n17353), .ZN(n17358) );
  AOI22_X1 U20512 ( .A1(n9601), .A2(n17691), .B1(n17399), .B2(n17356), .ZN(
        n17381) );
  OAI21_X1 U20513 ( .B1(n17694), .B2(n17365), .A(n17381), .ZN(n17371) );
  NOR2_X1 U20514 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17662), .ZN(
        n17686) );
  AOI22_X1 U20515 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17371), .B1(
        n17686), .B2(n17383), .ZN(n17357) );
  OAI211_X1 U20516 ( .C1(n17700), .C2(n17402), .A(n17358), .B(n17357), .ZN(
        P3_U2819) );
  INV_X1 U20517 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17709) );
  INV_X1 U20518 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17364) );
  OAI221_X1 U20519 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17379), .C1(
        n17709), .C2(n17378), .A(n17364), .ZN(n17362) );
  NAND4_X1 U20520 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17387), .A3(
        n17709), .A4(n17359), .ZN(n17360) );
  NAND3_X1 U20521 ( .A1(n17362), .A2(n17361), .A3(n17360), .ZN(n17708) );
  AOI22_X1 U20522 ( .A1(n9597), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17363), 
        .B2(n17480), .ZN(n17373) );
  OAI21_X1 U20523 ( .B1(n17365), .B2(n17709), .A(n17364), .ZN(n17370) );
  INV_X1 U20524 ( .A(n17366), .ZN(n17377) );
  OAI21_X1 U20525 ( .B1(n17485), .B2(n17367), .A(n17377), .ZN(n17368) );
  AOI22_X1 U20526 ( .A1(n17371), .A2(n17370), .B1(n17369), .B2(n17368), .ZN(
        n17372) );
  OAI211_X1 U20527 ( .C1(n17402), .C2(n17708), .A(n17373), .B(n17372), .ZN(
        P3_U2820) );
  OAI22_X1 U20528 ( .A1(n17485), .A2(n17375), .B1(n17394), .B2(n17374), .ZN(
        n17376) );
  AOI22_X1 U20529 ( .A1(n9597), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17377), .B2(
        n17376), .ZN(n17385) );
  NAND2_X1 U20530 ( .A1(n17379), .A2(n17378), .ZN(n17380) );
  XOR2_X1 U20531 ( .A(n17380), .B(n17709), .Z(n17717) );
  OAI22_X1 U20532 ( .A1(n17381), .A2(n17709), .B1(n17717), .B2(n17402), .ZN(
        n17382) );
  AOI21_X1 U20533 ( .B1(n17709), .B2(n17383), .A(n17382), .ZN(n17384) );
  OAI211_X1 U20534 ( .C1(n17471), .C2(n17386), .A(n17385), .B(n17384), .ZN(
        P3_U2821) );
  NOR2_X1 U20535 ( .A1(n17689), .A2(n17387), .ZN(n17724) );
  XOR2_X1 U20536 ( .A(n17724), .B(n17388), .Z(n17728) );
  AOI21_X1 U20537 ( .B1(n17390), .B2(n17733), .A(n17389), .ZN(n17730) );
  OAI21_X1 U20538 ( .B1(n17391), .B2(n17456), .A(n17488), .ZN(n17408) );
  INV_X1 U20539 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17393) );
  AOI21_X1 U20540 ( .B1(n17393), .B2(n17392), .A(n18019), .ZN(n17395) );
  AOI22_X1 U20541 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17408), .B1(
        n17395), .B2(n17394), .ZN(n17396) );
  NAND2_X1 U20542 ( .A1(n9597), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17731) );
  OAI211_X1 U20543 ( .C1(n17471), .C2(n17397), .A(n17396), .B(n17731), .ZN(
        n17398) );
  AOI21_X1 U20544 ( .B1(n9601), .B2(n17730), .A(n17398), .ZN(n17401) );
  NAND2_X1 U20545 ( .A1(n17728), .A2(n17399), .ZN(n17400) );
  OAI211_X1 U20546 ( .C1(n17728), .C2(n17402), .A(n17401), .B(n17400), .ZN(
        P3_U2822) );
  NAND2_X1 U20547 ( .A1(n17404), .A2(n17403), .ZN(n17405) );
  XOR2_X1 U20548 ( .A(n17405), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n17743) );
  NOR2_X1 U20549 ( .A1(n17712), .A2(n18362), .ZN(n17735) );
  AOI221_X1 U20550 ( .B1(n17408), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17407), .C2(n17406), .A(n17735), .ZN(n17413) );
  AOI21_X1 U20551 ( .B1(n17737), .B2(n17410), .A(n17409), .ZN(n17740) );
  AOI22_X1 U20552 ( .A1(n17481), .A2(n17740), .B1(n17411), .B2(n17480), .ZN(
        n17412) );
  OAI211_X1 U20553 ( .C1(n17492), .C2(n17743), .A(n17413), .B(n17412), .ZN(
        P3_U2823) );
  AOI21_X1 U20554 ( .B1(n17416), .B2(n17415), .A(n17414), .ZN(n17745) );
  NOR2_X1 U20555 ( .A1(n17421), .A2(n18019), .ZN(n17417) );
  AOI22_X1 U20556 ( .A1(n17481), .A2(n17745), .B1(n17417), .B2(n17422), .ZN(
        n17426) );
  AOI21_X1 U20557 ( .B1(n17419), .B2(n17747), .A(n17418), .ZN(n17746) );
  INV_X1 U20558 ( .A(n17485), .ZN(n17420) );
  OAI21_X1 U20559 ( .B1(n18019), .B2(n17421), .A(n17420), .ZN(n17437) );
  OAI22_X1 U20560 ( .A1(n17471), .A2(n17423), .B1(n17422), .B2(n17437), .ZN(
        n17424) );
  AOI21_X1 U20561 ( .B1(n9601), .B2(n17746), .A(n17424), .ZN(n17425) );
  OAI211_X1 U20562 ( .C1(n17712), .C2(n18360), .A(n17426), .B(n17425), .ZN(
        P3_U2824) );
  NOR2_X1 U20563 ( .A1(n17457), .A2(n17441), .ZN(n17459) );
  AOI21_X1 U20564 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17459), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17438) );
  OAI21_X1 U20565 ( .B1(n17429), .B2(n17428), .A(n17427), .ZN(n17430) );
  XOR2_X1 U20566 ( .A(n17430), .B(n10030), .Z(n17752) );
  AOI22_X1 U20567 ( .A1(n17481), .A2(n17752), .B1(n9597), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17436) );
  AOI21_X1 U20568 ( .B1(n17433), .B2(n17432), .A(n17431), .ZN(n17753) );
  AOI22_X1 U20569 ( .A1(n9601), .A2(n17753), .B1(n17434), .B2(n17480), .ZN(
        n17435) );
  OAI211_X1 U20570 ( .C1(n17438), .C2(n17437), .A(n17436), .B(n17435), .ZN(
        P3_U2825) );
  AOI21_X1 U20571 ( .B1(n17769), .B2(n17440), .A(n17439), .ZN(n17766) );
  NOR2_X1 U20572 ( .A1(n17712), .A2(n18356), .ZN(n17763) );
  NOR3_X1 U20573 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17441), .A3(
        n18019), .ZN(n17442) );
  AOI211_X1 U20574 ( .C1(n9601), .C2(n17766), .A(n17763), .B(n17442), .ZN(
        n17448) );
  AOI21_X1 U20575 ( .B1(n17445), .B2(n17444), .A(n17443), .ZN(n17764) );
  NOR2_X1 U20576 ( .A1(n17485), .A2(n17459), .ZN(n17446) );
  AOI22_X1 U20577 ( .A1(n17481), .A2(n17764), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17446), .ZN(n17447) );
  OAI211_X1 U20578 ( .C1(n17471), .C2(n17449), .A(n17448), .B(n17447), .ZN(
        P3_U2826) );
  AOI21_X1 U20579 ( .B1(n17452), .B2(n17451), .A(n17450), .ZN(n17771) );
  AOI22_X1 U20580 ( .A1(n17481), .A2(n17771), .B1(n9597), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17463) );
  AOI21_X1 U20581 ( .B1(n17455), .B2(n17454), .A(n17453), .ZN(n17775) );
  INV_X1 U20582 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17474) );
  NOR4_X1 U20583 ( .A1(n17457), .A2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17474), .A4(n17456), .ZN(n17461) );
  NOR3_X1 U20584 ( .A1(n17485), .A2(n17459), .A3(n17458), .ZN(n17460) );
  AOI211_X1 U20585 ( .C1(n9601), .C2(n17775), .A(n17461), .B(n17460), .ZN(
        n17462) );
  OAI211_X1 U20586 ( .C1(n17471), .C2(n17464), .A(n17463), .B(n17462), .ZN(
        P3_U2827) );
  AOI21_X1 U20587 ( .B1(n17467), .B2(n17466), .A(n17465), .ZN(n17785) );
  NOR2_X1 U20588 ( .A1(n17712), .A2(n18351), .ZN(n17791) );
  XNOR2_X1 U20589 ( .A(n17469), .B(n17468), .ZN(n17790) );
  OAI22_X1 U20590 ( .A1(n17471), .A2(n17470), .B1(n17492), .B2(n17790), .ZN(
        n17472) );
  AOI211_X1 U20591 ( .C1(n17481), .C2(n17785), .A(n17791), .B(n17472), .ZN(
        n17473) );
  OAI221_X1 U20592 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18019), .C1(
        n17474), .C2(n17488), .A(n17473), .ZN(P3_U2828) );
  NOR2_X1 U20593 ( .A1(n17487), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17475) );
  XOR2_X1 U20594 ( .A(n17475), .B(n17479), .Z(n17803) );
  INV_X1 U20595 ( .A(n17803), .ZN(n17476) );
  AOI22_X1 U20596 ( .A1(n9601), .A2(n17476), .B1(n9597), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17483) );
  AOI21_X1 U20597 ( .B1(n17479), .B2(n17486), .A(n17478), .ZN(n17799) );
  AOI22_X1 U20598 ( .A1(n17481), .A2(n17799), .B1(n17484), .B2(n17480), .ZN(
        n17482) );
  OAI211_X1 U20599 ( .C1(n17485), .C2(n17484), .A(n17483), .B(n17482), .ZN(
        P3_U2829) );
  OAI21_X1 U20600 ( .B1(n17487), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17486), .ZN(n17808) );
  INV_X1 U20601 ( .A(n17808), .ZN(n17810) );
  NAND3_X1 U20602 ( .A1(n18429), .A2(n18334), .A3(n17488), .ZN(n17489) );
  AOI22_X1 U20603 ( .A1(n9597), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17489), .ZN(n17490) );
  OAI221_X1 U20604 ( .B1(n17810), .B2(n17492), .C1(n17808), .C2(n17491), .A(
        n17490), .ZN(P3_U2830) );
  AOI221_X1 U20605 ( .B1(n17546), .B2(n9925), .C1(n17493), .C2(n9925), .A(
        n17804), .ZN(n17502) );
  NOR3_X1 U20606 ( .A1(n18447), .A2(n17494), .A3(n17661), .ZN(n17618) );
  AOI21_X1 U20607 ( .B1(n17555), .B2(n17618), .A(n18270), .ZN(n17560) );
  AOI221_X1 U20608 ( .B1(n20633), .B2(n17760), .C1(n17495), .C2(n17760), .A(
        n17560), .ZN(n17535) );
  OAI21_X1 U20609 ( .B1(n17720), .B2(n17516), .A(n17535), .ZN(n17519) );
  OAI22_X1 U20610 ( .A1(n17806), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18270), .B2(n17496), .ZN(n17499) );
  OAI211_X1 U20611 ( .C1(n17806), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17509), .ZN(n17501) );
  AOI22_X1 U20612 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17761), .B1(
        n17502), .B2(n17501), .ZN(n17504) );
  OAI211_X1 U20613 ( .C1(n17505), .C2(n17727), .A(n17504), .B(n17503), .ZN(
        P3_U2835) );
  OR2_X1 U20614 ( .A1(n17531), .A2(n17506), .ZN(n17508) );
  OR2_X1 U20615 ( .A1(n17507), .A2(n17546), .ZN(n17562) );
  NOR2_X1 U20616 ( .A1(n17508), .A2(n17562), .ZN(n17511) );
  INV_X1 U20617 ( .A(n17509), .ZN(n17510) );
  MUX2_X1 U20618 ( .A(n17511), .B(n17510), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17512) );
  AOI22_X1 U20619 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17761), .B1(
        n17793), .B2(n17512), .ZN(n17514) );
  OAI211_X1 U20620 ( .C1(n17515), .C2(n17727), .A(n17514), .B(n17513), .ZN(
        P3_U2836) );
  NAND3_X1 U20621 ( .A1(n17544), .A2(n17595), .A3(n17516), .ZN(n17520) );
  INV_X1 U20622 ( .A(n17520), .ZN(n17518) );
  AOI22_X1 U20623 ( .A1(n18266), .A2(n17518), .B1(n17786), .B2(n17517), .ZN(
        n17526) );
  AOI21_X1 U20624 ( .B1(n18266), .B2(n17520), .A(n17519), .ZN(n17525) );
  INV_X1 U20625 ( .A(n17521), .ZN(n17523) );
  AOI22_X1 U20626 ( .A1(n18264), .A2(n17523), .B1(n17725), .B2(n17522), .ZN(
        n17524) );
  OAI221_X1 U20627 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17526), 
        .C1(n17531), .C2(n17525), .A(n17524), .ZN(n17528) );
  AOI22_X1 U20628 ( .A1(n17793), .A2(n17528), .B1(n17681), .B2(n17527), .ZN(
        n17530) );
  OAI211_X1 U20629 ( .C1(n17805), .C2(n17531), .A(n17530), .B(n17529), .ZN(
        P3_U2837) );
  AOI22_X1 U20630 ( .A1(n9597), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17567), 
        .B2(n17532), .ZN(n17542) );
  AOI21_X1 U20631 ( .B1(n18264), .B2(n17533), .A(n17761), .ZN(n17534) );
  OAI211_X1 U20632 ( .C1(n17536), .C2(n17688), .A(n17535), .B(n17534), .ZN(
        n17540) );
  NAND2_X1 U20633 ( .A1(n17544), .A2(n17595), .ZN(n17538) );
  AOI211_X1 U20634 ( .C1(n18266), .C2(n17538), .A(n17537), .B(n17540), .ZN(
        n17539) );
  NOR2_X1 U20635 ( .A1(n9597), .A2(n17539), .ZN(n17547) );
  OAI211_X1 U20636 ( .C1(n17619), .C2(n17540), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17547), .ZN(n17541) );
  OAI211_X1 U20637 ( .C1(n17543), .C2(n17727), .A(n17542), .B(n17541), .ZN(
        P3_U2838) );
  INV_X1 U20638 ( .A(n17544), .ZN(n17545) );
  NOR3_X1 U20639 ( .A1(n17546), .A2(n17761), .A3(n17545), .ZN(n17548) );
  OAI21_X1 U20640 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17548), .A(
        n17547), .ZN(n17549) );
  OAI211_X1 U20641 ( .C1(n17551), .C2(n17727), .A(n17550), .B(n17549), .ZN(
        P3_U2839) );
  INV_X1 U20642 ( .A(n17595), .ZN(n17552) );
  OAI21_X1 U20643 ( .B1(n17553), .B2(n17552), .A(n18266), .ZN(n17554) );
  OAI221_X1 U20644 ( .B1(n17806), .B2(n17596), .C1(n17806), .C2(n17580), .A(
        n17554), .ZN(n17571) );
  NOR2_X1 U20645 ( .A1(n18264), .A2(n17725), .ZN(n17693) );
  OAI22_X1 U20646 ( .A1(n17806), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17555), .B2(n17693), .ZN(n17575) );
  AOI22_X1 U20647 ( .A1(n17725), .A2(n17631), .B1(n18264), .B2(n17639), .ZN(
        n17570) );
  AOI22_X1 U20648 ( .A1(n18266), .A2(n17557), .B1(n18294), .B2(n17556), .ZN(
        n17558) );
  NAND3_X1 U20649 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17570), .A3(
        n17558), .ZN(n17559) );
  NOR4_X1 U20650 ( .A1(n17560), .A2(n17571), .A3(n17575), .A4(n17559), .ZN(
        n17561) );
  AOI211_X1 U20651 ( .C1(n20633), .C2(n17562), .A(n17561), .B(n17804), .ZN(
        n17563) );
  AOI21_X1 U20652 ( .B1(n17681), .B2(n17564), .A(n17563), .ZN(n17566) );
  OAI211_X1 U20653 ( .C1(n17805), .C2(n20633), .A(n17566), .B(n17565), .ZN(
        P3_U2840) );
  NAND2_X1 U20654 ( .A1(n17569), .A2(n17567), .ZN(n17590) );
  AOI22_X1 U20655 ( .A1(n9597), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17681), 
        .B2(n17568), .ZN(n17577) );
  NOR2_X1 U20656 ( .A1(n18266), .A2(n18282), .ZN(n17795) );
  AOI21_X1 U20657 ( .B1(n17569), .B2(n17618), .A(n18270), .ZN(n17572) );
  NAND2_X1 U20658 ( .A1(n17793), .A2(n17570), .ZN(n17620) );
  NOR3_X1 U20659 ( .A1(n17572), .A2(n17620), .A3(n17571), .ZN(n17581) );
  OAI21_X1 U20660 ( .B1(n17573), .B2(n17795), .A(n17581), .ZN(n17574) );
  OAI211_X1 U20661 ( .C1(n17575), .C2(n17574), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17712), .ZN(n17576) );
  OAI211_X1 U20662 ( .C1(n17578), .C2(n17590), .A(n17577), .B(n17576), .ZN(
        P3_U2841) );
  AOI22_X1 U20663 ( .A1(n9597), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17681), 
        .B2(n17579), .ZN(n17584) );
  AOI221_X1 U20664 ( .B1(n17693), .B2(n17581), .C1(n17580), .C2(n17581), .A(
        n9597), .ZN(n17587) );
  NOR3_X1 U20665 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17795), .A3(
        n18485), .ZN(n17582) );
  OAI21_X1 U20666 ( .B1(n17587), .B2(n17582), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17583) );
  OAI211_X1 U20667 ( .C1(n17585), .C2(n17590), .A(n17584), .B(n17583), .ZN(
        P3_U2842) );
  AOI22_X1 U20668 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17587), .B1(
        n17681), .B2(n17586), .ZN(n17589) );
  OAI211_X1 U20669 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17590), .A(
        n17589), .B(n17588), .ZN(P3_U2843) );
  AOI22_X1 U20670 ( .A1(n18266), .A2(n17779), .B1(n17786), .B2(n17591), .ZN(
        n17772) );
  NOR2_X1 U20671 ( .A1(n17772), .A2(n17592), .ZN(n17748) );
  NAND2_X1 U20672 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17748), .ZN(
        n17736) );
  NOR3_X1 U20673 ( .A1(n17737), .A2(n17733), .A3(n17736), .ZN(n17627) );
  NOR2_X1 U20674 ( .A1(n17627), .A2(n17593), .ZN(n17677) );
  NAND2_X1 U20675 ( .A1(n17594), .A2(n17710), .ZN(n17625) );
  AOI21_X1 U20676 ( .B1(n17599), .B2(n17595), .A(n18301), .ZN(n17601) );
  INV_X1 U20677 ( .A(n17596), .ZN(n17597) );
  NOR3_X1 U20678 ( .A1(n17758), .A2(n17597), .A3(n17624), .ZN(n17598) );
  OAI22_X1 U20679 ( .A1(n17599), .A2(n17693), .B1(n17720), .B2(n17598), .ZN(
        n17600) );
  NOR3_X1 U20680 ( .A1(n17601), .A2(n17620), .A3(n17600), .ZN(n17608) );
  AOI221_X1 U20681 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17608), 
        .C1(n17720), .C2(n17608), .A(n9597), .ZN(n17603) );
  AOI22_X1 U20682 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17603), .B1(
        n17681), .B2(n17602), .ZN(n17605) );
  OAI211_X1 U20683 ( .C1(n17625), .C2(n17606), .A(n17605), .B(n17604), .ZN(
        P3_U2844) );
  NOR3_X1 U20684 ( .A1(n9597), .A2(n17608), .A3(n17607), .ZN(n17609) );
  AOI21_X1 U20685 ( .B1(n17681), .B2(n17610), .A(n17609), .ZN(n17612) );
  OAI211_X1 U20686 ( .C1(n17625), .C2(n17613), .A(n17612), .B(n17611), .ZN(
        P3_U2845) );
  INV_X1 U20687 ( .A(n17649), .ZN(n17704) );
  NAND2_X1 U20688 ( .A1(n18294), .A2(n17661), .ZN(n17702) );
  NAND2_X1 U20689 ( .A1(n18266), .A2(n17614), .ZN(n17692) );
  NAND2_X1 U20690 ( .A1(n17702), .A2(n17692), .ZN(n17714) );
  NOR2_X1 U20691 ( .A1(n17615), .A2(n17714), .ZN(n17651) );
  NOR2_X1 U20692 ( .A1(n18282), .A2(n17616), .ZN(n17617) );
  OAI22_X1 U20693 ( .A1(n17704), .A2(n17651), .B1(n17618), .B2(n17617), .ZN(
        n17630) );
  OAI221_X1 U20694 ( .B1(n17620), .B2(n17619), .C1(n17620), .C2(n17630), .A(
        n17712), .ZN(n17623) );
  AOI22_X1 U20695 ( .A1(n9597), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17681), 
        .B2(n17621), .ZN(n17622) );
  OAI221_X1 U20696 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17625), 
        .C1(n17624), .C2(n17623), .A(n17622), .ZN(P3_U2846) );
  AOI21_X1 U20697 ( .B1(n17761), .B2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17626), .ZN(n17642) );
  INV_X1 U20698 ( .A(n17627), .ZN(n17629) );
  NOR2_X1 U20699 ( .A1(n17629), .A2(n17628), .ZN(n17652) );
  OAI21_X1 U20700 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17652), .A(
        n17630), .ZN(n17634) );
  NAND2_X1 U20701 ( .A1(n17725), .A2(n17631), .ZN(n17632) );
  OAI22_X1 U20702 ( .A1(n17635), .A2(n17634), .B1(n17633), .B2(n17632), .ZN(
        n17637) );
  AOI22_X1 U20703 ( .A1(n17793), .A2(n17637), .B1(n17681), .B2(n17636), .ZN(
        n17641) );
  NAND3_X1 U20704 ( .A1(n17809), .A2(n17639), .A3(n17638), .ZN(n17640) );
  NAND3_X1 U20705 ( .A1(n17642), .A2(n17641), .A3(n17640), .ZN(P3_U2847) );
  OAI221_X1 U20706 ( .B1(n17646), .B2(n17645), .C1(n17644), .C2(n17643), .A(
        n17784), .ZN(n17655) );
  NOR2_X1 U20707 ( .A1(n18447), .A2(n17661), .ZN(n17687) );
  AOI21_X1 U20708 ( .B1(n17647), .B2(n17687), .A(n18270), .ZN(n17667) );
  NOR2_X1 U20709 ( .A1(n17649), .A2(n17648), .ZN(n17650) );
  OAI22_X1 U20710 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17795), .B1(
        n17651), .B2(n17650), .ZN(n17653) );
  OAI22_X1 U20711 ( .A1(n17667), .A2(n17653), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17652), .ZN(n17654) );
  AOI21_X1 U20712 ( .B1(n17655), .B2(n17654), .A(n17804), .ZN(n17656) );
  AOI211_X1 U20713 ( .C1(n17761), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17657), .B(n17656), .ZN(n17658) );
  OAI21_X1 U20714 ( .B1(n17802), .B2(n17659), .A(n17658), .ZN(P3_U2848) );
  AOI21_X1 U20715 ( .B1(n18294), .B2(n17660), .A(n17685), .ZN(n17674) );
  OAI21_X1 U20716 ( .B1(n17662), .B2(n17661), .A(n18294), .ZN(n17663) );
  INV_X1 U20717 ( .A(n17663), .ZN(n17664) );
  AOI21_X1 U20718 ( .B1(n18266), .B2(n17676), .A(n17664), .ZN(n17696) );
  OAI211_X1 U20719 ( .C1(n17665), .C2(n17789), .A(n17696), .B(n17692), .ZN(
        n17666) );
  AOI211_X1 U20720 ( .C1(n17725), .C2(n17668), .A(n17667), .B(n17666), .ZN(
        n17675) );
  OAI211_X1 U20721 ( .C1(n17704), .C2(n17674), .A(n17793), .B(n17675), .ZN(
        n17669) );
  NAND2_X1 U20722 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17669), .ZN(
        n17673) );
  AOI22_X1 U20723 ( .A1(n17681), .A2(n17671), .B1(n17710), .B2(n17670), .ZN(
        n17672) );
  OAI221_X1 U20724 ( .B1(n9597), .B2(n17673), .C1(n17712), .C2(n18373), .A(
        n17672), .ZN(P3_U2849) );
  AOI21_X1 U20725 ( .B1(n17675), .B2(n17674), .A(n17804), .ZN(n17679) );
  OAI21_X1 U20726 ( .B1(n17677), .B2(n17676), .A(n17685), .ZN(n17678) );
  AOI22_X1 U20727 ( .A1(n17681), .A2(n17680), .B1(n17679), .B2(n17678), .ZN(
        n17684) );
  INV_X1 U20728 ( .A(n17682), .ZN(n17683) );
  OAI211_X1 U20729 ( .C1(n17805), .C2(n17685), .A(n17684), .B(n17683), .ZN(
        P3_U2850) );
  AOI22_X1 U20730 ( .A1(n9597), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17710), 
        .B2(n17686), .ZN(n17699) );
  OAI22_X1 U20731 ( .A1(n17689), .A2(n17688), .B1(n18270), .B2(n17687), .ZN(
        n17690) );
  AOI211_X1 U20732 ( .C1(n17691), .C2(n18264), .A(n17804), .B(n17690), .ZN(
        n17711) );
  OAI211_X1 U20733 ( .C1(n17694), .C2(n17693), .A(n17711), .B(n17692), .ZN(
        n17695) );
  AOI21_X1 U20734 ( .B1(n18282), .B2(n17709), .A(n17695), .ZN(n17703) );
  OAI211_X1 U20735 ( .C1(n18270), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17696), .B(n17703), .ZN(n17697) );
  NAND3_X1 U20736 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17712), .A3(
        n17697), .ZN(n17698) );
  OAI211_X1 U20737 ( .C1(n17700), .C2(n17727), .A(n17699), .B(n17698), .ZN(
        P3_U2851) );
  NOR2_X1 U20738 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17709), .ZN(
        n17701) );
  AOI22_X1 U20739 ( .A1(n9597), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17710), 
        .B2(n17701), .ZN(n17707) );
  OAI211_X1 U20740 ( .C1(n17704), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17703), .B(n17702), .ZN(n17705) );
  NAND3_X1 U20741 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17712), .A3(
        n17705), .ZN(n17706) );
  OAI211_X1 U20742 ( .C1(n17708), .C2(n17727), .A(n17707), .B(n17706), .ZN(
        P3_U2852) );
  AOI22_X1 U20743 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n9597), .B1(n17710), .B2(
        n17709), .ZN(n17716) );
  INV_X1 U20744 ( .A(n17711), .ZN(n17713) );
  OAI211_X1 U20745 ( .C1(n17714), .C2(n17713), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n17712), .ZN(n17715) );
  OAI211_X1 U20746 ( .C1(n17717), .C2(n17727), .A(n17716), .B(n17715), .ZN(
        P3_U2853) );
  OAI22_X1 U20747 ( .A1(n17720), .A2(n17719), .B1(n17718), .B2(n18301), .ZN(
        n17721) );
  NOR2_X1 U20748 ( .A1(n17758), .A2(n17721), .ZN(n17744) );
  OAI211_X1 U20749 ( .C1(n17722), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n17744), .ZN(n17738) );
  AOI21_X1 U20750 ( .B1(n17762), .B2(n17738), .A(n17761), .ZN(n17734) );
  NOR3_X1 U20751 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17737), .A3(
        n17736), .ZN(n17723) );
  AOI21_X1 U20752 ( .B1(n17725), .B2(n17724), .A(n17723), .ZN(n17726) );
  OAI22_X1 U20753 ( .A1(n17728), .A2(n17727), .B1(n17726), .B2(n17804), .ZN(
        n17729) );
  AOI21_X1 U20754 ( .B1(n17809), .B2(n17730), .A(n17729), .ZN(n17732) );
  OAI211_X1 U20755 ( .C1(n17734), .C2(n17733), .A(n17732), .B(n17731), .ZN(
        P3_U2854) );
  AOI21_X1 U20756 ( .B1(n17761), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17735), .ZN(n17742) );
  AOI21_X1 U20757 ( .B1(n17737), .B2(n17736), .A(n17804), .ZN(n17739) );
  AOI22_X1 U20758 ( .A1(n17811), .A2(n17740), .B1(n17739), .B2(n17738), .ZN(
        n17741) );
  OAI211_X1 U20759 ( .C1(n17802), .C2(n17743), .A(n17742), .B(n17741), .ZN(
        P3_U2855) );
  OAI21_X1 U20760 ( .B1(n17744), .B2(n17804), .A(n17805), .ZN(n17754) );
  AOI22_X1 U20761 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17754), .B1(
        n9597), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U20762 ( .A1(n17809), .A2(n17746), .B1(n17811), .B2(n17745), .ZN(
        n17750) );
  NAND3_X1 U20763 ( .A1(n17793), .A2(n17748), .A3(n17747), .ZN(n17749) );
  NAND3_X1 U20764 ( .A1(n17751), .A2(n17750), .A3(n17749), .ZN(P3_U2856) );
  AOI22_X1 U20765 ( .A1(n9597), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17811), .B2(
        n17752), .ZN(n17757) );
  AOI22_X1 U20766 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17754), .B1(
        n17809), .B2(n17753), .ZN(n17756) );
  NOR3_X1 U20767 ( .A1(n17772), .A2(n17804), .A3(n17778), .ZN(n17765) );
  NAND3_X1 U20768 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17765), .A3(
        n10030), .ZN(n17755) );
  NAND3_X1 U20769 ( .A1(n17757), .A2(n17756), .A3(n17755), .ZN(P3_U2857) );
  AOI21_X1 U20770 ( .B1(n17760), .B2(n17759), .A(n17758), .ZN(n17781) );
  OAI211_X1 U20771 ( .C1(n18301), .C2(n17779), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n17781), .ZN(n17773) );
  AOI21_X1 U20772 ( .B1(n17762), .B2(n17773), .A(n17761), .ZN(n17770) );
  AOI21_X1 U20773 ( .B1(n17764), .B2(n17811), .A(n17763), .ZN(n17768) );
  AOI22_X1 U20774 ( .A1(n17766), .A2(n17809), .B1(n17765), .B2(n17769), .ZN(
        n17767) );
  OAI211_X1 U20775 ( .C1(n17770), .C2(n17769), .A(n17768), .B(n17767), .ZN(
        P3_U2858) );
  AOI22_X1 U20776 ( .A1(n9597), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n17811), .B2(
        n17771), .ZN(n17777) );
  AOI21_X1 U20777 ( .B1(n17772), .B2(n17778), .A(n17804), .ZN(n17774) );
  AOI22_X1 U20778 ( .A1(n17809), .A2(n17775), .B1(n17774), .B2(n17773), .ZN(
        n17776) );
  OAI211_X1 U20779 ( .C1(n17778), .C2(n17805), .A(n17777), .B(n17776), .ZN(
        P3_U2859) );
  NOR2_X1 U20780 ( .A1(n18301), .A2(n17779), .ZN(n17783) );
  NAND2_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17780) );
  AOI221_X1 U20782 ( .B1(n18301), .B2(n17781), .C1(n17780), .C2(n17781), .A(
        n20606), .ZN(n17782) );
  AOI211_X1 U20783 ( .C1(n17785), .C2(n17784), .A(n17783), .B(n17782), .ZN(
        n17788) );
  NAND3_X1 U20784 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17786), .A3(
        n20606), .ZN(n17787) );
  OAI211_X1 U20785 ( .C1(n17790), .C2(n17789), .A(n17788), .B(n17787), .ZN(
        n17792) );
  AOI21_X1 U20786 ( .B1(n17793), .B2(n17792), .A(n17791), .ZN(n17794) );
  OAI21_X1 U20787 ( .B1(n20606), .B2(n17805), .A(n17794), .ZN(P3_U2860) );
  OR3_X1 U20788 ( .A1(n17804), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n17795), .ZN(n17812) );
  AOI21_X1 U20789 ( .B1(n17805), .B2(n17812), .A(n18430), .ZN(n17798) );
  AOI211_X1 U20790 ( .C1(n17806), .C2(n18447), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17796), .ZN(n17797) );
  AOI211_X1 U20791 ( .C1(n17799), .C2(n17811), .A(n17798), .B(n17797), .ZN(
        n17801) );
  NAND2_X1 U20792 ( .A1(n9597), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n17800) );
  OAI211_X1 U20793 ( .C1(n17803), .C2(n17802), .A(n17801), .B(n17800), .ZN(
        P3_U2861) );
  AOI221_X1 U20794 ( .B1(n17806), .B2(n17805), .C1(n17804), .C2(n17805), .A(
        n18447), .ZN(n17807) );
  AOI221_X1 U20795 ( .B1(n17811), .B2(n17810), .C1(n17809), .C2(n17808), .A(
        n17807), .ZN(n17813) );
  OAI211_X1 U20796 ( .C1(n18458), .C2(n17712), .A(n17813), .B(n17812), .ZN(
        P3_U2862) );
  OAI211_X1 U20797 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n17814), .A(
        P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .ZN(n18323)
         );
  OAI21_X1 U20798 ( .B1(n17817), .B2(n17815), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17816) );
  OAI221_X1 U20799 ( .B1(n17817), .B2(n18323), .C1(n17817), .C2(n17868), .A(
        n17816), .ZN(P3_U2863) );
  INV_X1 U20800 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18308) );
  NAND2_X1 U20801 ( .A1(n17818), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18090) );
  INV_X1 U20802 ( .A(n18090), .ZN(n18116) );
  NOR2_X1 U20803 ( .A1(n17818), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17997) );
  NOR2_X1 U20804 ( .A1(n18116), .A2(n17997), .ZN(n17820) );
  OAI22_X1 U20805 ( .A1(n17821), .A2(n18308), .B1(n17820), .B2(n17819), .ZN(
        P3_U2866) );
  NOR2_X1 U20806 ( .A1(n17823), .A2(n17822), .ZN(P3_U2867) );
  NAND2_X1 U20807 ( .A1(n18205), .A2(BUF2_REG_16__SCAN_IN), .ZN(n20665) );
  NOR2_X1 U20808 ( .A1(n18091), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18067) );
  INV_X1 U20809 ( .A(n18067), .ZN(n17973) );
  NAND2_X1 U20810 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17827) );
  NOR2_X2 U20811 ( .A1(n17973), .A2(n17827), .ZN(n18196) );
  INV_X1 U20812 ( .A(n18196), .ZN(n17884) );
  NOR2_X2 U20813 ( .A1(n18018), .A2(n17824), .ZN(n20659) );
  NOR2_X1 U20814 ( .A1(n18091), .A2(n17826), .ZN(n18273) );
  INV_X1 U20815 ( .A(n17827), .ZN(n17825) );
  NAND2_X1 U20816 ( .A1(n18273), .A2(n17825), .ZN(n17903) );
  INV_X1 U20817 ( .A(n17903), .ZN(n18253) );
  NAND2_X1 U20818 ( .A1(n18091), .A2(n17826), .ZN(n18017) );
  INV_X1 U20819 ( .A(n18017), .ZN(n18274) );
  NOR2_X1 U20820 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17911) );
  NAND2_X1 U20821 ( .A1(n18274), .A2(n17911), .ZN(n17924) );
  NOR2_X1 U20822 ( .A1(n18253), .A2(n17928), .ZN(n17889) );
  NOR2_X1 U20823 ( .A1(n18166), .A2(n17889), .ZN(n17862) );
  NAND2_X1 U20824 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18205), .ZN(n18209) );
  INV_X1 U20825 ( .A(n18209), .ZN(n20658) );
  NOR2_X1 U20826 ( .A1(n17827), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18204) );
  NAND2_X1 U20827 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18204), .ZN(
        n18241) );
  INV_X1 U20828 ( .A(n18241), .ZN(n18251) );
  AOI22_X1 U20829 ( .A1(n20659), .A2(n17862), .B1(n20658), .B2(n18251), .ZN(
        n17833) );
  NOR2_X1 U20830 ( .A1(n17826), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n17952) );
  NOR2_X1 U20831 ( .A1(n18067), .A2(n17952), .ZN(n18119) );
  NOR2_X1 U20832 ( .A1(n18119), .A2(n17827), .ZN(n18165) );
  AOI211_X1 U20833 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n17889), .B(n18018), .ZN(
        n17828) );
  AOI21_X1 U20834 ( .B1(n18165), .B2(n18205), .A(n17828), .ZN(n17865) );
  NAND2_X1 U20835 ( .A1(n17830), .A2(n17829), .ZN(n17863) );
  NOR2_X1 U20836 ( .A1(n17863), .A2(n17831), .ZN(n18206) );
  AOI22_X1 U20837 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17865), .B1(
        n18206), .B2(n17928), .ZN(n17832) );
  OAI211_X1 U20838 ( .C1(n20665), .C2(n17884), .A(n17833), .B(n17832), .ZN(
        P3_U2868) );
  NAND2_X1 U20839 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18205), .ZN(n18177) );
  NAND2_X1 U20840 ( .A1(n18205), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18215) );
  INV_X1 U20841 ( .A(n18215), .ZN(n18174) );
  AOI22_X1 U20842 ( .A1(n18196), .A2(n18174), .B1(n17862), .B2(n18210), .ZN(
        n17836) );
  NOR2_X2 U20843 ( .A1(n17834), .A2(n17863), .ZN(n18212) );
  AOI22_X1 U20844 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17865), .B1(
        n17928), .B2(n18212), .ZN(n17835) );
  OAI211_X1 U20845 ( .C1(n18241), .C2(n18177), .A(n17836), .B(n17835), .ZN(
        P3_U2869) );
  NAND2_X1 U20846 ( .A1(n18205), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18221) );
  NAND2_X1 U20847 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18205), .ZN(n18181) );
  INV_X1 U20848 ( .A(n18181), .ZN(n18217) );
  NOR2_X2 U20849 ( .A1(n18018), .A2(n17837), .ZN(n18216) );
  AOI22_X1 U20850 ( .A1(n18251), .A2(n18217), .B1(n17862), .B2(n18216), .ZN(
        n17840) );
  NOR2_X2 U20851 ( .A1(n17838), .A2(n17863), .ZN(n18218) );
  AOI22_X1 U20852 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n17865), .B1(
        n17928), .B2(n18218), .ZN(n17839) );
  OAI211_X1 U20853 ( .C1(n17884), .C2(n18221), .A(n17840), .B(n17839), .ZN(
        P3_U2870) );
  NOR2_X1 U20854 ( .A1(n17841), .A2(n18019), .ZN(n18223) );
  INV_X1 U20855 ( .A(n18223), .ZN(n18185) );
  NAND2_X1 U20856 ( .A1(n18205), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18227) );
  INV_X1 U20857 ( .A(n18227), .ZN(n18182) );
  NOR2_X2 U20858 ( .A1(n18018), .A2(n17842), .ZN(n18222) );
  AOI22_X1 U20859 ( .A1(n18196), .A2(n18182), .B1(n17862), .B2(n18222), .ZN(
        n17845) );
  NOR2_X2 U20860 ( .A1(n17843), .A2(n17863), .ZN(n18224) );
  AOI22_X1 U20861 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n17865), .B1(
        n17928), .B2(n18224), .ZN(n17844) );
  OAI211_X1 U20862 ( .C1(n18241), .C2(n18185), .A(n17845), .B(n17844), .ZN(
        P3_U2871) );
  INV_X1 U20863 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n17846) );
  NOR2_X1 U20864 ( .A1(n18019), .A2(n17846), .ZN(n18229) );
  INV_X1 U20865 ( .A(n18229), .ZN(n18103) );
  NAND2_X1 U20866 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18205), .ZN(n18233) );
  INV_X1 U20867 ( .A(n18233), .ZN(n18100) );
  NOR2_X2 U20868 ( .A1(n18018), .A2(n17847), .ZN(n18228) );
  AOI22_X1 U20869 ( .A1(n18251), .A2(n18100), .B1(n17862), .B2(n18228), .ZN(
        n17850) );
  NOR2_X2 U20870 ( .A1(n17848), .A2(n17863), .ZN(n18230) );
  AOI22_X1 U20871 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n17865), .B1(
        n17928), .B2(n18230), .ZN(n17849) );
  OAI211_X1 U20872 ( .C1(n17884), .C2(n18103), .A(n17850), .B(n17849), .ZN(
        P3_U2872) );
  INV_X1 U20873 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n17851) );
  NOR2_X1 U20874 ( .A1(n17851), .A2(n18019), .ZN(n18104) );
  INV_X1 U20875 ( .A(n18104), .ZN(n18240) );
  NAND2_X1 U20876 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18205), .ZN(n18107) );
  INV_X1 U20877 ( .A(n18107), .ZN(n18236) );
  NOR2_X2 U20878 ( .A1(n17852), .A2(n18018), .ZN(n18234) );
  AOI22_X1 U20879 ( .A1(n18251), .A2(n18236), .B1(n17862), .B2(n18234), .ZN(
        n17855) );
  NOR2_X2 U20880 ( .A1(n17853), .A2(n17863), .ZN(n18237) );
  AOI22_X1 U20881 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n17865), .B1(
        n17928), .B2(n18237), .ZN(n17854) );
  OAI211_X1 U20882 ( .C1(n17884), .C2(n18240), .A(n17855), .B(n17854), .ZN(
        P3_U2873) );
  NAND2_X1 U20883 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18205), .ZN(n18159) );
  NAND2_X1 U20884 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18205), .ZN(n18247) );
  INV_X1 U20885 ( .A(n18247), .ZN(n18156) );
  NOR2_X2 U20886 ( .A1(n17856), .A2(n18018), .ZN(n18242) );
  AOI22_X1 U20887 ( .A1(n18251), .A2(n18156), .B1(n17862), .B2(n18242), .ZN(
        n17859) );
  NOR2_X2 U20888 ( .A1(n17857), .A2(n17863), .ZN(n18244) );
  AOI22_X1 U20889 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17865), .B1(
        n17928), .B2(n18244), .ZN(n17858) );
  OAI211_X1 U20890 ( .C1(n17884), .C2(n18159), .A(n17859), .B(n17858), .ZN(
        P3_U2874) );
  INV_X1 U20891 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n17860) );
  NOR2_X1 U20892 ( .A1(n17860), .A2(n18019), .ZN(n18250) );
  NAND2_X1 U20893 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18205), .ZN(n18258) );
  INV_X1 U20894 ( .A(n18258), .ZN(n18195) );
  NOR2_X2 U20895 ( .A1(n17861), .A2(n18018), .ZN(n18249) );
  AOI22_X1 U20896 ( .A1(n18251), .A2(n18195), .B1(n17862), .B2(n18249), .ZN(
        n17867) );
  NOR2_X2 U20897 ( .A1(n17864), .A2(n17863), .ZN(n18252) );
  AOI22_X1 U20898 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17865), .B1(
        n17928), .B2(n18252), .ZN(n17866) );
  OAI211_X1 U20899 ( .C1(n17884), .C2(n18200), .A(n17867), .B(n17866), .ZN(
        P3_U2875) );
  INV_X1 U20900 ( .A(n18206), .ZN(n20662) );
  INV_X1 U20901 ( .A(n17911), .ZN(n17949) );
  INV_X1 U20902 ( .A(n17952), .ZN(n18042) );
  NOR2_X2 U20903 ( .A1(n17949), .A2(n18042), .ZN(n20657) );
  INV_X1 U20904 ( .A(n20657), .ZN(n17948) );
  INV_X1 U20905 ( .A(n20665), .ZN(n18201) );
  NAND2_X1 U20906 ( .A1(n18091), .A2(n18324), .ZN(n18043) );
  NOR2_X1 U20907 ( .A1(n17949), .A2(n18043), .ZN(n17885) );
  AOI22_X1 U20908 ( .A1(n18201), .A2(n18253), .B1(n20659), .B2(n17885), .ZN(
        n17871) );
  NOR2_X1 U20909 ( .A1(n18308), .A2(n18044), .ZN(n18202) );
  INV_X1 U20910 ( .A(n17868), .ZN(n17869) );
  NOR2_X1 U20911 ( .A1(n18018), .A2(n17869), .ZN(n18203) );
  INV_X1 U20912 ( .A(n18203), .ZN(n17910) );
  NOR2_X1 U20913 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17910), .ZN(
        n17950) );
  AOI22_X1 U20914 ( .A1(n18205), .A2(n18202), .B1(n17911), .B2(n17950), .ZN(
        n17886) );
  AOI22_X1 U20915 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n17886), .B1(
        n20658), .B2(n18196), .ZN(n17870) );
  OAI211_X1 U20916 ( .C1(n20662), .C2(n17948), .A(n17871), .B(n17870), .ZN(
        P3_U2876) );
  AOI22_X1 U20917 ( .A1(n18253), .A2(n18174), .B1(n18210), .B2(n17885), .ZN(
        n17873) );
  AOI22_X1 U20918 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17886), .B1(
        n20657), .B2(n18212), .ZN(n17872) );
  OAI211_X1 U20919 ( .C1(n17884), .C2(n18177), .A(n17873), .B(n17872), .ZN(
        P3_U2877) );
  AOI22_X1 U20920 ( .A1(n18196), .A2(n18217), .B1(n18216), .B2(n17885), .ZN(
        n17875) );
  AOI22_X1 U20921 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n17886), .B1(
        n20657), .B2(n18218), .ZN(n17874) );
  OAI211_X1 U20922 ( .C1(n17903), .C2(n18221), .A(n17875), .B(n17874), .ZN(
        P3_U2878) );
  AOI22_X1 U20923 ( .A1(n18253), .A2(n18182), .B1(n18222), .B2(n17885), .ZN(
        n17877) );
  AOI22_X1 U20924 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n17886), .B1(
        n20657), .B2(n18224), .ZN(n17876) );
  OAI211_X1 U20925 ( .C1(n17884), .C2(n18185), .A(n17877), .B(n17876), .ZN(
        P3_U2879) );
  AOI22_X1 U20926 ( .A1(n18196), .A2(n18100), .B1(n18228), .B2(n17885), .ZN(
        n17879) );
  AOI22_X1 U20927 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n17886), .B1(
        n20657), .B2(n18230), .ZN(n17878) );
  OAI211_X1 U20928 ( .C1(n17903), .C2(n18103), .A(n17879), .B(n17878), .ZN(
        P3_U2880) );
  AOI22_X1 U20929 ( .A1(n18253), .A2(n18104), .B1(n18234), .B2(n17885), .ZN(
        n17881) );
  AOI22_X1 U20930 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n17886), .B1(
        n20657), .B2(n18237), .ZN(n17880) );
  OAI211_X1 U20931 ( .C1(n17884), .C2(n18107), .A(n17881), .B(n17880), .ZN(
        P3_U2881) );
  INV_X1 U20932 ( .A(n18159), .ZN(n18243) );
  AOI22_X1 U20933 ( .A1(n18253), .A2(n18243), .B1(n18242), .B2(n17885), .ZN(
        n17883) );
  AOI22_X1 U20934 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n17886), .B1(
        n20657), .B2(n18244), .ZN(n17882) );
  OAI211_X1 U20935 ( .C1(n17884), .C2(n18247), .A(n17883), .B(n17882), .ZN(
        P3_U2882) );
  AOI22_X1 U20936 ( .A1(n18196), .A2(n18195), .B1(n18249), .B2(n17885), .ZN(
        n17888) );
  AOI22_X1 U20937 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17886), .B1(
        n20657), .B2(n18252), .ZN(n17887) );
  OAI211_X1 U20938 ( .C1(n17903), .C2(n18200), .A(n17888), .B(n17887), .ZN(
        P3_U2883) );
  NOR2_X2 U20939 ( .A1(n17949), .A2(n17973), .ZN(n17968) );
  INV_X1 U20940 ( .A(n17968), .ZN(n20664) );
  OR2_X1 U20941 ( .A1(n17949), .A2(n18119), .ZN(n17932) );
  NOR2_X1 U20942 ( .A1(n18166), .A2(n17932), .ZN(n17906) );
  AOI22_X1 U20943 ( .A1(n18201), .A2(n17928), .B1(n20659), .B2(n17906), .ZN(
        n17892) );
  OAI21_X1 U20944 ( .B1(n17889), .B2(n18168), .A(n17932), .ZN(n17890) );
  OAI211_X1 U20945 ( .C1(n17968), .C2(n18419), .A(n18171), .B(n17890), .ZN(
        n17907) );
  AOI22_X1 U20946 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n17907), .B1(
        n20658), .B2(n18253), .ZN(n17891) );
  OAI211_X1 U20947 ( .C1(n20664), .C2(n20662), .A(n17892), .B(n17891), .ZN(
        P3_U2884) );
  AOI22_X1 U20948 ( .A1(n17928), .A2(n18174), .B1(n18210), .B2(n17906), .ZN(
        n17894) );
  AOI22_X1 U20949 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17907), .B1(
        n17968), .B2(n18212), .ZN(n17893) );
  OAI211_X1 U20950 ( .C1(n17903), .C2(n18177), .A(n17894), .B(n17893), .ZN(
        P3_U2885) );
  INV_X1 U20951 ( .A(n18221), .ZN(n18178) );
  AOI22_X1 U20952 ( .A1(n17928), .A2(n18178), .B1(n18216), .B2(n17906), .ZN(
        n17896) );
  AOI22_X1 U20953 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n17907), .B1(
        n17968), .B2(n18218), .ZN(n17895) );
  OAI211_X1 U20954 ( .C1(n17903), .C2(n18181), .A(n17896), .B(n17895), .ZN(
        P3_U2886) );
  AOI22_X1 U20955 ( .A1(n17928), .A2(n18182), .B1(n18222), .B2(n17906), .ZN(
        n17898) );
  AOI22_X1 U20956 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n17907), .B1(
        n17968), .B2(n18224), .ZN(n17897) );
  OAI211_X1 U20957 ( .C1(n17903), .C2(n18185), .A(n17898), .B(n17897), .ZN(
        P3_U2887) );
  AOI22_X1 U20958 ( .A1(n17928), .A2(n18229), .B1(n18228), .B2(n17906), .ZN(
        n17900) );
  AOI22_X1 U20959 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n17907), .B1(
        n17968), .B2(n18230), .ZN(n17899) );
  OAI211_X1 U20960 ( .C1(n17903), .C2(n18233), .A(n17900), .B(n17899), .ZN(
        P3_U2888) );
  AOI22_X1 U20961 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n17907), .B1(
        n18234), .B2(n17906), .ZN(n17902) );
  AOI22_X1 U20962 ( .A1(n17968), .A2(n18237), .B1(n17928), .B2(n18104), .ZN(
        n17901) );
  OAI211_X1 U20963 ( .C1(n17903), .C2(n18107), .A(n17902), .B(n17901), .ZN(
        P3_U2889) );
  AOI22_X1 U20964 ( .A1(n18253), .A2(n18156), .B1(n18242), .B2(n17906), .ZN(
        n17905) );
  AOI22_X1 U20965 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n17907), .B1(
        n17968), .B2(n18244), .ZN(n17904) );
  OAI211_X1 U20966 ( .C1(n17924), .C2(n18159), .A(n17905), .B(n17904), .ZN(
        P3_U2890) );
  AOI22_X1 U20967 ( .A1(n18253), .A2(n18195), .B1(n18249), .B2(n17906), .ZN(
        n17909) );
  AOI22_X1 U20968 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17907), .B1(
        n17968), .B2(n18252), .ZN(n17908) );
  OAI211_X1 U20969 ( .C1(n17924), .C2(n18200), .A(n17909), .B(n17908), .ZN(
        P3_U2891) );
  AOI22_X1 U20970 ( .A1(n20659), .A2(n17927), .B1(n20658), .B2(n17928), .ZN(
        n17913) );
  AOI21_X1 U20971 ( .B1(n18091), .B2(n18168), .A(n17910), .ZN(n17996) );
  NAND2_X1 U20972 ( .A1(n17911), .A2(n17996), .ZN(n17929) );
  NAND2_X1 U20973 ( .A1(n18273), .A2(n17911), .ZN(n17988) );
  INV_X1 U20974 ( .A(n17988), .ZN(n17992) );
  AOI22_X1 U20975 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18206), .ZN(n17912) );
  OAI211_X1 U20976 ( .C1(n20665), .C2(n17948), .A(n17913), .B(n17912), .ZN(
        P3_U2892) );
  INV_X1 U20977 ( .A(n18177), .ZN(n18211) );
  AOI22_X1 U20978 ( .A1(n17928), .A2(n18211), .B1(n18210), .B2(n17927), .ZN(
        n17915) );
  AOI22_X1 U20979 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18212), .ZN(n17914) );
  OAI211_X1 U20980 ( .C1(n17948), .C2(n18215), .A(n17915), .B(n17914), .ZN(
        P3_U2893) );
  AOI22_X1 U20981 ( .A1(n20657), .A2(n18178), .B1(n18216), .B2(n17927), .ZN(
        n17917) );
  AOI22_X1 U20982 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18218), .ZN(n17916) );
  OAI211_X1 U20983 ( .C1(n17924), .C2(n18181), .A(n17917), .B(n17916), .ZN(
        P3_U2894) );
  AOI22_X1 U20984 ( .A1(n17928), .A2(n18223), .B1(n18222), .B2(n17927), .ZN(
        n17919) );
  AOI22_X1 U20985 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18224), .ZN(n17918) );
  OAI211_X1 U20986 ( .C1(n17948), .C2(n18227), .A(n17919), .B(n17918), .ZN(
        P3_U2895) );
  AOI22_X1 U20987 ( .A1(n20657), .A2(n18229), .B1(n18228), .B2(n17927), .ZN(
        n17921) );
  AOI22_X1 U20988 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18230), .ZN(n17920) );
  OAI211_X1 U20989 ( .C1(n17924), .C2(n18233), .A(n17921), .B(n17920), .ZN(
        P3_U2896) );
  AOI22_X1 U20990 ( .A1(n20657), .A2(n18104), .B1(n18234), .B2(n17927), .ZN(
        n17923) );
  AOI22_X1 U20991 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18237), .ZN(n17922) );
  OAI211_X1 U20992 ( .C1(n17924), .C2(n18107), .A(n17923), .B(n17922), .ZN(
        P3_U2897) );
  AOI22_X1 U20993 ( .A1(n17928), .A2(n18156), .B1(n18242), .B2(n17927), .ZN(
        n17926) );
  AOI22_X1 U20994 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18244), .ZN(n17925) );
  OAI211_X1 U20995 ( .C1(n17948), .C2(n18159), .A(n17926), .B(n17925), .ZN(
        P3_U2898) );
  AOI22_X1 U20996 ( .A1(n17928), .A2(n18195), .B1(n18249), .B2(n17927), .ZN(
        n17931) );
  AOI22_X1 U20997 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17929), .B1(
        n17992), .B2(n18252), .ZN(n17930) );
  OAI211_X1 U20998 ( .C1(n17948), .C2(n18200), .A(n17931), .B(n17930), .ZN(
        P3_U2899) );
  NAND2_X1 U20999 ( .A1(n18274), .A2(n17997), .ZN(n20663) );
  NOR2_X1 U21000 ( .A1(n18013), .A2(n17992), .ZN(n17974) );
  NOR2_X1 U21001 ( .A1(n18166), .A2(n17974), .ZN(n20660) );
  AOI22_X1 U21002 ( .A1(n20660), .A2(n18210), .B1(n20657), .B2(n18211), .ZN(
        n17935) );
  OAI22_X1 U21003 ( .A1(n17974), .A2(n18018), .B1(n18019), .B2(n17932), .ZN(
        n17933) );
  OAI21_X1 U21004 ( .B1(n18013), .B2(n18419), .A(n17933), .ZN(n20668) );
  AOI22_X1 U21005 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20668), .B1(
        n18013), .B2(n18212), .ZN(n17934) );
  OAI211_X1 U21006 ( .C1(n20664), .C2(n18215), .A(n17935), .B(n17934), .ZN(
        P3_U2901) );
  AOI22_X1 U21007 ( .A1(n17968), .A2(n18178), .B1(n20660), .B2(n18216), .ZN(
        n17937) );
  AOI22_X1 U21008 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20668), .B1(
        n18013), .B2(n18218), .ZN(n17936) );
  OAI211_X1 U21009 ( .C1(n17948), .C2(n18181), .A(n17937), .B(n17936), .ZN(
        P3_U2902) );
  AOI22_X1 U21010 ( .A1(n20660), .A2(n18222), .B1(n20657), .B2(n18223), .ZN(
        n17939) );
  AOI22_X1 U21011 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20668), .B1(
        n18013), .B2(n18224), .ZN(n17938) );
  OAI211_X1 U21012 ( .C1(n20664), .C2(n18227), .A(n17939), .B(n17938), .ZN(
        P3_U2903) );
  AOI22_X1 U21013 ( .A1(n20660), .A2(n18228), .B1(n20657), .B2(n18100), .ZN(
        n17941) );
  AOI22_X1 U21014 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20668), .B1(
        n18013), .B2(n18230), .ZN(n17940) );
  OAI211_X1 U21015 ( .C1(n20664), .C2(n18103), .A(n17941), .B(n17940), .ZN(
        P3_U2904) );
  AOI22_X1 U21016 ( .A1(n20660), .A2(n18234), .B1(n20657), .B2(n18236), .ZN(
        n17943) );
  AOI22_X1 U21017 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20668), .B1(
        n18013), .B2(n18237), .ZN(n17942) );
  OAI211_X1 U21018 ( .C1(n20664), .C2(n18240), .A(n17943), .B(n17942), .ZN(
        P3_U2905) );
  AOI22_X1 U21019 ( .A1(n17968), .A2(n18243), .B1(n20660), .B2(n18242), .ZN(
        n17945) );
  AOI22_X1 U21020 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20668), .B1(
        n18013), .B2(n18244), .ZN(n17944) );
  OAI211_X1 U21021 ( .C1(n17948), .C2(n18247), .A(n17945), .B(n17944), .ZN(
        P3_U2906) );
  AOI22_X1 U21022 ( .A1(n17968), .A2(n18250), .B1(n20660), .B2(n18249), .ZN(
        n17947) );
  AOI22_X1 U21023 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20668), .B1(
        n18013), .B2(n18252), .ZN(n17946) );
  OAI211_X1 U21024 ( .C1(n17948), .C2(n18258), .A(n17947), .B(n17946), .ZN(
        P3_U2907) );
  INV_X1 U21025 ( .A(n17997), .ZN(n17972) );
  NOR2_X1 U21026 ( .A1(n17972), .A2(n18043), .ZN(n17967) );
  AOI22_X1 U21027 ( .A1(n18201), .A2(n17992), .B1(n20659), .B2(n17967), .ZN(
        n17954) );
  NOR2_X1 U21028 ( .A1(n18091), .A2(n17949), .ZN(n17951) );
  AOI22_X1 U21029 ( .A1(n18205), .A2(n17951), .B1(n17997), .B2(n17950), .ZN(
        n17969) );
  NAND2_X1 U21030 ( .A1(n17997), .A2(n17952), .ZN(n18034) );
  AOI22_X1 U21031 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n17969), .B1(
        n18206), .B2(n18038), .ZN(n17953) );
  OAI211_X1 U21032 ( .C1(n20664), .C2(n18209), .A(n17954), .B(n17953), .ZN(
        P3_U2908) );
  AOI22_X1 U21033 ( .A1(n17992), .A2(n18174), .B1(n18210), .B2(n17967), .ZN(
        n17956) );
  AOI22_X1 U21034 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17969), .B1(
        n18212), .B2(n18038), .ZN(n17955) );
  OAI211_X1 U21035 ( .C1(n20664), .C2(n18177), .A(n17956), .B(n17955), .ZN(
        P3_U2909) );
  AOI22_X1 U21036 ( .A1(n17992), .A2(n18178), .B1(n18216), .B2(n17967), .ZN(
        n17958) );
  AOI22_X1 U21037 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n17969), .B1(
        n18218), .B2(n18038), .ZN(n17957) );
  OAI211_X1 U21038 ( .C1(n20664), .C2(n18181), .A(n17958), .B(n17957), .ZN(
        P3_U2910) );
  AOI22_X1 U21039 ( .A1(n17992), .A2(n18182), .B1(n18222), .B2(n17967), .ZN(
        n17960) );
  AOI22_X1 U21040 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n17969), .B1(
        n18224), .B2(n18038), .ZN(n17959) );
  OAI211_X1 U21041 ( .C1(n20664), .C2(n18185), .A(n17960), .B(n17959), .ZN(
        P3_U2911) );
  AOI22_X1 U21042 ( .A1(n17968), .A2(n18100), .B1(n18228), .B2(n17967), .ZN(
        n17962) );
  AOI22_X1 U21043 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n17969), .B1(
        n18230), .B2(n18038), .ZN(n17961) );
  OAI211_X1 U21044 ( .C1(n17988), .C2(n18103), .A(n17962), .B(n17961), .ZN(
        P3_U2912) );
  AOI22_X1 U21045 ( .A1(n17968), .A2(n18236), .B1(n18234), .B2(n17967), .ZN(
        n17964) );
  AOI22_X1 U21046 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n17969), .B1(
        n18237), .B2(n18038), .ZN(n17963) );
  OAI211_X1 U21047 ( .C1(n17988), .C2(n18240), .A(n17964), .B(n17963), .ZN(
        P3_U2913) );
  AOI22_X1 U21048 ( .A1(n17968), .A2(n18156), .B1(n18242), .B2(n17967), .ZN(
        n17966) );
  AOI22_X1 U21049 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n17969), .B1(
        n18244), .B2(n18038), .ZN(n17965) );
  OAI211_X1 U21050 ( .C1(n17988), .C2(n18159), .A(n17966), .B(n17965), .ZN(
        P3_U2914) );
  AOI22_X1 U21051 ( .A1(n17968), .A2(n18195), .B1(n18249), .B2(n17967), .ZN(
        n17971) );
  AOI22_X1 U21052 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17969), .B1(
        n18252), .B2(n18038), .ZN(n17970) );
  OAI211_X1 U21053 ( .C1(n17988), .C2(n18200), .A(n17971), .B(n17970), .ZN(
        P3_U2915) );
  NOR2_X2 U21054 ( .A1(n17973), .A2(n17972), .ZN(n18059) );
  INV_X1 U21055 ( .A(n18059), .ZN(n18066) );
  AOI21_X1 U21056 ( .B1(n18034), .B2(n18066), .A(n18166), .ZN(n17991) );
  AOI22_X1 U21057 ( .A1(n17992), .A2(n20658), .B1(n20659), .B2(n17991), .ZN(
        n17977) );
  AOI221_X1 U21058 ( .B1(n17974), .B2(n18034), .C1(n18168), .C2(n18034), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n17975) );
  OAI21_X1 U21059 ( .B1(n18059), .B2(n17975), .A(n18171), .ZN(n17993) );
  AOI22_X1 U21060 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n17993), .B1(
        n18206), .B2(n18059), .ZN(n17976) );
  OAI211_X1 U21061 ( .C1(n20665), .C2(n20663), .A(n17977), .B(n17976), .ZN(
        P3_U2916) );
  AOI22_X1 U21062 ( .A1(n17992), .A2(n18211), .B1(n18210), .B2(n17991), .ZN(
        n17979) );
  AOI22_X1 U21063 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17993), .B1(
        n18212), .B2(n18059), .ZN(n17978) );
  OAI211_X1 U21064 ( .C1(n20663), .C2(n18215), .A(n17979), .B(n17978), .ZN(
        P3_U2917) );
  AOI22_X1 U21065 ( .A1(n18013), .A2(n18178), .B1(n18216), .B2(n17991), .ZN(
        n17981) );
  AOI22_X1 U21066 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n17993), .B1(
        n18218), .B2(n18059), .ZN(n17980) );
  OAI211_X1 U21067 ( .C1(n17988), .C2(n18181), .A(n17981), .B(n17980), .ZN(
        P3_U2918) );
  AOI22_X1 U21068 ( .A1(n17992), .A2(n18223), .B1(n18222), .B2(n17991), .ZN(
        n17983) );
  AOI22_X1 U21069 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n17993), .B1(
        n18224), .B2(n18059), .ZN(n17982) );
  OAI211_X1 U21070 ( .C1(n20663), .C2(n18227), .A(n17983), .B(n17982), .ZN(
        P3_U2919) );
  AOI22_X1 U21071 ( .A1(n18013), .A2(n18229), .B1(n18228), .B2(n17991), .ZN(
        n17985) );
  AOI22_X1 U21072 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n17993), .B1(
        n18230), .B2(n18059), .ZN(n17984) );
  OAI211_X1 U21073 ( .C1(n17988), .C2(n18233), .A(n17985), .B(n17984), .ZN(
        P3_U2920) );
  AOI22_X1 U21074 ( .A1(n18013), .A2(n18104), .B1(n18234), .B2(n17991), .ZN(
        n17987) );
  AOI22_X1 U21075 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n17993), .B1(
        n18237), .B2(n18059), .ZN(n17986) );
  OAI211_X1 U21076 ( .C1(n17988), .C2(n18107), .A(n17987), .B(n17986), .ZN(
        P3_U2921) );
  AOI22_X1 U21077 ( .A1(n17992), .A2(n18156), .B1(n18242), .B2(n17991), .ZN(
        n17990) );
  AOI22_X1 U21078 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n17993), .B1(
        n18244), .B2(n18059), .ZN(n17989) );
  OAI211_X1 U21079 ( .C1(n20663), .C2(n18159), .A(n17990), .B(n17989), .ZN(
        P3_U2922) );
  AOI22_X1 U21080 ( .A1(n17992), .A2(n18195), .B1(n18249), .B2(n17991), .ZN(
        n17995) );
  AOI22_X1 U21081 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17993), .B1(
        n18252), .B2(n18059), .ZN(n17994) );
  OAI211_X1 U21082 ( .C1(n20663), .C2(n18200), .A(n17995), .B(n17994), .ZN(
        P3_U2923) );
  AOI22_X1 U21083 ( .A1(n18201), .A2(n18038), .B1(n20659), .B2(n18012), .ZN(
        n17999) );
  NAND2_X1 U21084 ( .A1(n17997), .A2(n17996), .ZN(n18014) );
  NAND2_X1 U21085 ( .A1(n18273), .A2(n17997), .ZN(n18089) );
  INV_X1 U21086 ( .A(n18089), .ZN(n18076) );
  AOI22_X1 U21087 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18014), .B1(
        n18206), .B2(n18076), .ZN(n17998) );
  OAI211_X1 U21088 ( .C1(n20663), .C2(n18209), .A(n17999), .B(n17998), .ZN(
        P3_U2924) );
  AOI22_X1 U21089 ( .A1(n18013), .A2(n18211), .B1(n18210), .B2(n18012), .ZN(
        n18001) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18014), .B1(
        n18212), .B2(n18076), .ZN(n18000) );
  OAI211_X1 U21091 ( .C1(n18215), .C2(n18034), .A(n18001), .B(n18000), .ZN(
        P3_U2925) );
  AOI22_X1 U21092 ( .A1(n18178), .A2(n18038), .B1(n18216), .B2(n18012), .ZN(
        n18003) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18014), .B1(
        n18218), .B2(n18076), .ZN(n18002) );
  OAI211_X1 U21094 ( .C1(n20663), .C2(n18181), .A(n18003), .B(n18002), .ZN(
        P3_U2926) );
  AOI22_X1 U21095 ( .A1(n18222), .A2(n18012), .B1(n18182), .B2(n18038), .ZN(
        n18005) );
  AOI22_X1 U21096 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18014), .B1(
        n18224), .B2(n18076), .ZN(n18004) );
  OAI211_X1 U21097 ( .C1(n20663), .C2(n18185), .A(n18005), .B(n18004), .ZN(
        P3_U2927) );
  AOI22_X1 U21098 ( .A1(n18229), .A2(n18038), .B1(n18228), .B2(n18012), .ZN(
        n18007) );
  AOI22_X1 U21099 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18014), .B1(
        n18230), .B2(n18076), .ZN(n18006) );
  OAI211_X1 U21100 ( .C1(n20663), .C2(n18233), .A(n18007), .B(n18006), .ZN(
        P3_U2928) );
  AOI22_X1 U21101 ( .A1(n18013), .A2(n18236), .B1(n18234), .B2(n18012), .ZN(
        n18009) );
  AOI22_X1 U21102 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18014), .B1(
        n18237), .B2(n18076), .ZN(n18008) );
  OAI211_X1 U21103 ( .C1(n18240), .C2(n18034), .A(n18009), .B(n18008), .ZN(
        P3_U2929) );
  AOI22_X1 U21104 ( .A1(n18013), .A2(n18156), .B1(n18242), .B2(n18012), .ZN(
        n18011) );
  AOI22_X1 U21105 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18014), .B1(
        n18244), .B2(n18076), .ZN(n18010) );
  OAI211_X1 U21106 ( .C1(n18159), .C2(n18034), .A(n18011), .B(n18010), .ZN(
        P3_U2930) );
  AOI22_X1 U21107 ( .A1(n18013), .A2(n18195), .B1(n18249), .B2(n18012), .ZN(
        n18016) );
  AOI22_X1 U21108 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18014), .B1(
        n18252), .B2(n18076), .ZN(n18015) );
  OAI211_X1 U21109 ( .C1(n18200), .C2(n18034), .A(n18016), .B(n18015), .ZN(
        P3_U2931) );
  NOR2_X2 U21110 ( .A1(n18017), .A2(n18090), .ZN(n18112) );
  INV_X1 U21111 ( .A(n18112), .ZN(n18110) );
  NOR2_X1 U21112 ( .A1(n18076), .A2(n18112), .ZN(n18068) );
  NOR2_X1 U21113 ( .A1(n18166), .A2(n18068), .ZN(n18037) );
  AOI22_X1 U21114 ( .A1(n20659), .A2(n18037), .B1(n20658), .B2(n18038), .ZN(
        n18023) );
  NOR2_X1 U21115 ( .A1(n18038), .A2(n18059), .ZN(n18020) );
  OAI22_X1 U21116 ( .A1(n18020), .A2(n18019), .B1(n18068), .B2(n18018), .ZN(
        n18021) );
  OAI21_X1 U21117 ( .B1(n18112), .B2(n18419), .A(n18021), .ZN(n18039) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18039), .B1(
        n18201), .B2(n18059), .ZN(n18022) );
  OAI211_X1 U21119 ( .C1(n20662), .C2(n18110), .A(n18023), .B(n18022), .ZN(
        P3_U2932) );
  AOI22_X1 U21120 ( .A1(n18210), .A2(n18037), .B1(n18174), .B2(n18059), .ZN(
        n18025) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18039), .B1(
        n18212), .B2(n18112), .ZN(n18024) );
  OAI211_X1 U21122 ( .C1(n18177), .C2(n18034), .A(n18025), .B(n18024), .ZN(
        P3_U2933) );
  AOI22_X1 U21123 ( .A1(n18217), .A2(n18038), .B1(n18216), .B2(n18037), .ZN(
        n18027) );
  AOI22_X1 U21124 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18039), .B1(
        n18218), .B2(n18112), .ZN(n18026) );
  OAI211_X1 U21125 ( .C1(n18221), .C2(n18066), .A(n18027), .B(n18026), .ZN(
        P3_U2934) );
  AOI22_X1 U21126 ( .A1(n18223), .A2(n18038), .B1(n18222), .B2(n18037), .ZN(
        n18029) );
  AOI22_X1 U21127 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18039), .B1(
        n18224), .B2(n18112), .ZN(n18028) );
  OAI211_X1 U21128 ( .C1(n18227), .C2(n18066), .A(n18029), .B(n18028), .ZN(
        P3_U2935) );
  AOI22_X1 U21129 ( .A1(n18100), .A2(n18038), .B1(n18228), .B2(n18037), .ZN(
        n18031) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18039), .B1(
        n18230), .B2(n18112), .ZN(n18030) );
  OAI211_X1 U21131 ( .C1(n18103), .C2(n18066), .A(n18031), .B(n18030), .ZN(
        P3_U2936) );
  AOI22_X1 U21132 ( .A1(n18104), .A2(n18059), .B1(n18234), .B2(n18037), .ZN(
        n18033) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18039), .B1(
        n18237), .B2(n18112), .ZN(n18032) );
  OAI211_X1 U21134 ( .C1(n18107), .C2(n18034), .A(n18033), .B(n18032), .ZN(
        P3_U2937) );
  AOI22_X1 U21135 ( .A1(n18156), .A2(n18038), .B1(n18242), .B2(n18037), .ZN(
        n18036) );
  AOI22_X1 U21136 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18039), .B1(
        n18244), .B2(n18112), .ZN(n18035) );
  OAI211_X1 U21137 ( .C1(n18159), .C2(n18066), .A(n18036), .B(n18035), .ZN(
        P3_U2938) );
  AOI22_X1 U21138 ( .A1(n18195), .A2(n18038), .B1(n18249), .B2(n18037), .ZN(
        n18041) );
  AOI22_X1 U21139 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18039), .B1(
        n18252), .B2(n18112), .ZN(n18040) );
  OAI211_X1 U21140 ( .C1(n18200), .C2(n18066), .A(n18041), .B(n18040), .ZN(
        P3_U2939) );
  NOR2_X2 U21141 ( .A1(n18042), .A2(n18090), .ZN(n18137) );
  NOR2_X1 U21142 ( .A1(n18090), .A2(n18043), .ZN(n18062) );
  AOI22_X1 U21143 ( .A1(n20659), .A2(n18062), .B1(n20658), .B2(n18059), .ZN(
        n18048) );
  NOR2_X1 U21144 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18044), .ZN(
        n18046) );
  NOR2_X1 U21145 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18090), .ZN(
        n18045) );
  AOI22_X1 U21146 ( .A1(n18205), .A2(n18046), .B1(n18203), .B2(n18045), .ZN(
        n18063) );
  AOI22_X1 U21147 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18063), .B1(
        n18201), .B2(n18076), .ZN(n18047) );
  OAI211_X1 U21148 ( .C1(n20662), .C2(n18135), .A(n18048), .B(n18047), .ZN(
        P3_U2940) );
  AOI22_X1 U21149 ( .A1(n18210), .A2(n18062), .B1(n18174), .B2(n18076), .ZN(
        n18050) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18063), .B1(
        n18212), .B2(n18137), .ZN(n18049) );
  OAI211_X1 U21151 ( .C1(n18177), .C2(n18066), .A(n18050), .B(n18049), .ZN(
        P3_U2941) );
  AOI22_X1 U21152 ( .A1(n18178), .A2(n18076), .B1(n18216), .B2(n18062), .ZN(
        n18052) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18063), .B1(
        n18218), .B2(n18137), .ZN(n18051) );
  OAI211_X1 U21154 ( .C1(n18181), .C2(n18066), .A(n18052), .B(n18051), .ZN(
        P3_U2942) );
  AOI22_X1 U21155 ( .A1(n18223), .A2(n18059), .B1(n18222), .B2(n18062), .ZN(
        n18054) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18063), .B1(
        n18224), .B2(n18137), .ZN(n18053) );
  OAI211_X1 U21157 ( .C1(n18227), .C2(n18089), .A(n18054), .B(n18053), .ZN(
        P3_U2943) );
  AOI22_X1 U21158 ( .A1(n18229), .A2(n18076), .B1(n18228), .B2(n18062), .ZN(
        n18056) );
  AOI22_X1 U21159 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18063), .B1(
        n18230), .B2(n18137), .ZN(n18055) );
  OAI211_X1 U21160 ( .C1(n18233), .C2(n18066), .A(n18056), .B(n18055), .ZN(
        P3_U2944) );
  AOI22_X1 U21161 ( .A1(n18104), .A2(n18076), .B1(n18234), .B2(n18062), .ZN(
        n18058) );
  AOI22_X1 U21162 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18063), .B1(
        n18237), .B2(n18137), .ZN(n18057) );
  OAI211_X1 U21163 ( .C1(n18107), .C2(n18066), .A(n18058), .B(n18057), .ZN(
        P3_U2945) );
  AOI22_X1 U21164 ( .A1(n18156), .A2(n18059), .B1(n18242), .B2(n18062), .ZN(
        n18061) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18063), .B1(
        n18244), .B2(n18137), .ZN(n18060) );
  OAI211_X1 U21166 ( .C1(n18159), .C2(n18089), .A(n18061), .B(n18060), .ZN(
        P3_U2946) );
  AOI22_X1 U21167 ( .A1(n18250), .A2(n18076), .B1(n18249), .B2(n18062), .ZN(
        n18065) );
  AOI22_X1 U21168 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18063), .B1(
        n18252), .B2(n18137), .ZN(n18064) );
  OAI211_X1 U21169 ( .C1(n18258), .C2(n18066), .A(n18065), .B(n18064), .ZN(
        P3_U2947) );
  AOI22_X1 U21170 ( .A1(n18201), .A2(n18112), .B1(n20659), .B2(n18085), .ZN(
        n18071) );
  NAND2_X1 U21171 ( .A1(n18067), .A2(n18116), .ZN(n18153) );
  AOI221_X1 U21172 ( .B1(n18068), .B2(n18135), .C1(n18168), .C2(n18135), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18069) );
  OAI21_X1 U21173 ( .B1(n18161), .B2(n18069), .A(n18171), .ZN(n18086) );
  AOI22_X1 U21174 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18086), .B1(
        n18206), .B2(n18161), .ZN(n18070) );
  OAI211_X1 U21175 ( .C1(n18209), .C2(n18089), .A(n18071), .B(n18070), .ZN(
        P3_U2948) );
  AOI22_X1 U21176 ( .A1(n18211), .A2(n18076), .B1(n18210), .B2(n18085), .ZN(
        n18073) );
  AOI22_X1 U21177 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18086), .B1(
        n18212), .B2(n18161), .ZN(n18072) );
  OAI211_X1 U21178 ( .C1(n18215), .C2(n18110), .A(n18073), .B(n18072), .ZN(
        P3_U2949) );
  AOI22_X1 U21179 ( .A1(n18178), .A2(n18112), .B1(n18216), .B2(n18085), .ZN(
        n18075) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18086), .B1(
        n18218), .B2(n18161), .ZN(n18074) );
  OAI211_X1 U21181 ( .C1(n18181), .C2(n18089), .A(n18075), .B(n18074), .ZN(
        P3_U2950) );
  AOI22_X1 U21182 ( .A1(n18223), .A2(n18076), .B1(n18222), .B2(n18085), .ZN(
        n18078) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18086), .B1(
        n18224), .B2(n18161), .ZN(n18077) );
  OAI211_X1 U21184 ( .C1(n18227), .C2(n18110), .A(n18078), .B(n18077), .ZN(
        P3_U2951) );
  AOI22_X1 U21185 ( .A1(n18229), .A2(n18112), .B1(n18228), .B2(n18085), .ZN(
        n18080) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18086), .B1(
        n18230), .B2(n18161), .ZN(n18079) );
  OAI211_X1 U21187 ( .C1(n18233), .C2(n18089), .A(n18080), .B(n18079), .ZN(
        P3_U2952) );
  AOI22_X1 U21188 ( .A1(n18104), .A2(n18112), .B1(n18234), .B2(n18085), .ZN(
        n18082) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18086), .B1(
        n18237), .B2(n18161), .ZN(n18081) );
  OAI211_X1 U21190 ( .C1(n18107), .C2(n18089), .A(n18082), .B(n18081), .ZN(
        P3_U2953) );
  AOI22_X1 U21191 ( .A1(n18243), .A2(n18112), .B1(n18242), .B2(n18085), .ZN(
        n18084) );
  AOI22_X1 U21192 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18086), .B1(
        n18244), .B2(n18161), .ZN(n18083) );
  OAI211_X1 U21193 ( .C1(n18247), .C2(n18089), .A(n18084), .B(n18083), .ZN(
        P3_U2954) );
  AOI22_X1 U21194 ( .A1(n18250), .A2(n18112), .B1(n18249), .B2(n18085), .ZN(
        n18088) );
  AOI22_X1 U21195 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18086), .B1(
        n18252), .B2(n18161), .ZN(n18087) );
  OAI211_X1 U21196 ( .C1(n18258), .C2(n18089), .A(n18088), .B(n18087), .ZN(
        P3_U2955) );
  NOR2_X1 U21197 ( .A1(n18091), .A2(n18090), .ZN(n18142) );
  AND2_X1 U21198 ( .A1(n18324), .A2(n18142), .ZN(n18111) );
  AOI22_X1 U21199 ( .A1(n20659), .A2(n18111), .B1(n20658), .B2(n18112), .ZN(
        n18093) );
  OAI211_X1 U21200 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18205), .A(
        n18203), .B(n18116), .ZN(n18113) );
  NAND2_X1 U21201 ( .A1(n18273), .A2(n18116), .ZN(n18192) );
  INV_X1 U21202 ( .A(n18192), .ZN(n18194) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18113), .B1(
        n18206), .B2(n18194), .ZN(n18092) );
  OAI211_X1 U21204 ( .C1(n20665), .C2(n18135), .A(n18093), .B(n18092), .ZN(
        P3_U2956) );
  AOI22_X1 U21205 ( .A1(n18210), .A2(n18111), .B1(n18174), .B2(n18137), .ZN(
        n18095) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18113), .B1(
        n18212), .B2(n18194), .ZN(n18094) );
  OAI211_X1 U21207 ( .C1(n18177), .C2(n18110), .A(n18095), .B(n18094), .ZN(
        P3_U2957) );
  AOI22_X1 U21208 ( .A1(n18217), .A2(n18112), .B1(n18216), .B2(n18111), .ZN(
        n18097) );
  AOI22_X1 U21209 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18113), .B1(
        n18218), .B2(n18194), .ZN(n18096) );
  OAI211_X1 U21210 ( .C1(n18221), .C2(n18135), .A(n18097), .B(n18096), .ZN(
        P3_U2958) );
  AOI22_X1 U21211 ( .A1(n18223), .A2(n18112), .B1(n18222), .B2(n18111), .ZN(
        n18099) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18113), .B1(
        n18224), .B2(n18194), .ZN(n18098) );
  OAI211_X1 U21213 ( .C1(n18227), .C2(n18135), .A(n18099), .B(n18098), .ZN(
        P3_U2959) );
  AOI22_X1 U21214 ( .A1(n18100), .A2(n18112), .B1(n18228), .B2(n18111), .ZN(
        n18102) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18113), .B1(
        n18230), .B2(n18194), .ZN(n18101) );
  OAI211_X1 U21216 ( .C1(n18103), .C2(n18135), .A(n18102), .B(n18101), .ZN(
        P3_U2960) );
  AOI22_X1 U21217 ( .A1(n18104), .A2(n18137), .B1(n18234), .B2(n18111), .ZN(
        n18106) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18113), .B1(
        n18237), .B2(n18194), .ZN(n18105) );
  OAI211_X1 U21219 ( .C1(n18107), .C2(n18110), .A(n18106), .B(n18105), .ZN(
        P3_U2961) );
  AOI22_X1 U21220 ( .A1(n18243), .A2(n18137), .B1(n18242), .B2(n18111), .ZN(
        n18109) );
  AOI22_X1 U21221 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18113), .B1(
        n18244), .B2(n18194), .ZN(n18108) );
  OAI211_X1 U21222 ( .C1(n18247), .C2(n18110), .A(n18109), .B(n18108), .ZN(
        P3_U2962) );
  AOI22_X1 U21223 ( .A1(n18195), .A2(n18112), .B1(n18249), .B2(n18111), .ZN(
        n18115) );
  AOI22_X1 U21224 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18113), .B1(
        n18252), .B2(n18194), .ZN(n18114) );
  OAI211_X1 U21225 ( .C1(n18200), .C2(n18135), .A(n18115), .B(n18114), .ZN(
        P3_U2963) );
  INV_X1 U21226 ( .A(n18204), .ZN(n18141) );
  NOR2_X2 U21227 ( .A1(n18141), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18235) );
  INV_X1 U21228 ( .A(n18235), .ZN(n18257) );
  AOI21_X1 U21229 ( .B1(n18192), .B2(n18257), .A(n18166), .ZN(n18136) );
  AOI22_X1 U21230 ( .A1(n18201), .A2(n18161), .B1(n20659), .B2(n18136), .ZN(
        n18122) );
  NAND2_X1 U21231 ( .A1(n18117), .A2(n18116), .ZN(n18118) );
  AOI221_X1 U21232 ( .B1(n18119), .B2(n18192), .C1(n18118), .C2(n18192), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18120) );
  OAI21_X1 U21233 ( .B1(n18235), .B2(n18120), .A(n18171), .ZN(n18138) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18138), .B1(
        n18206), .B2(n18235), .ZN(n18121) );
  OAI211_X1 U21235 ( .C1(n18209), .C2(n18135), .A(n18122), .B(n18121), .ZN(
        P3_U2964) );
  AOI22_X1 U21236 ( .A1(n18211), .A2(n18137), .B1(n18210), .B2(n18136), .ZN(
        n18124) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18138), .B1(
        n18212), .B2(n18235), .ZN(n18123) );
  OAI211_X1 U21238 ( .C1(n18215), .C2(n18153), .A(n18124), .B(n18123), .ZN(
        P3_U2965) );
  AOI22_X1 U21239 ( .A1(n18217), .A2(n18137), .B1(n18216), .B2(n18136), .ZN(
        n18126) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18138), .B1(
        n18218), .B2(n18235), .ZN(n18125) );
  OAI211_X1 U21241 ( .C1(n18221), .C2(n18153), .A(n18126), .B(n18125), .ZN(
        P3_U2966) );
  AOI22_X1 U21242 ( .A1(n18222), .A2(n18136), .B1(n18182), .B2(n18161), .ZN(
        n18128) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18138), .B1(
        n18224), .B2(n18235), .ZN(n18127) );
  OAI211_X1 U21244 ( .C1(n18185), .C2(n18135), .A(n18128), .B(n18127), .ZN(
        P3_U2967) );
  AOI22_X1 U21245 ( .A1(n18229), .A2(n18161), .B1(n18228), .B2(n18136), .ZN(
        n18130) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18138), .B1(
        n18230), .B2(n18235), .ZN(n18129) );
  OAI211_X1 U21247 ( .C1(n18233), .C2(n18135), .A(n18130), .B(n18129), .ZN(
        P3_U2968) );
  AOI22_X1 U21248 ( .A1(n18236), .A2(n18137), .B1(n18234), .B2(n18136), .ZN(
        n18132) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18138), .B1(
        n18237), .B2(n18235), .ZN(n18131) );
  OAI211_X1 U21250 ( .C1(n18240), .C2(n18153), .A(n18132), .B(n18131), .ZN(
        P3_U2969) );
  AOI22_X1 U21251 ( .A1(n18243), .A2(n18161), .B1(n18242), .B2(n18136), .ZN(
        n18134) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18138), .B1(
        n18244), .B2(n18235), .ZN(n18133) );
  OAI211_X1 U21253 ( .C1(n18247), .C2(n18135), .A(n18134), .B(n18133), .ZN(
        P3_U2970) );
  AOI22_X1 U21254 ( .A1(n18195), .A2(n18137), .B1(n18249), .B2(n18136), .ZN(
        n18140) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18138), .B1(
        n18252), .B2(n18235), .ZN(n18139) );
  OAI211_X1 U21256 ( .C1(n18200), .C2(n18153), .A(n18140), .B(n18139), .ZN(
        P3_U2971) );
  NOR2_X1 U21257 ( .A1(n18166), .A2(n18141), .ZN(n18160) );
  AOI22_X1 U21258 ( .A1(n18201), .A2(n18194), .B1(n20659), .B2(n18160), .ZN(
        n18144) );
  AOI22_X1 U21259 ( .A1(n18205), .A2(n18142), .B1(n18204), .B2(n18203), .ZN(
        n18162) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18162), .B1(
        n18206), .B2(n18251), .ZN(n18143) );
  OAI211_X1 U21261 ( .C1(n18209), .C2(n18153), .A(n18144), .B(n18143), .ZN(
        P3_U2972) );
  AOI22_X1 U21262 ( .A1(n18211), .A2(n18161), .B1(n18210), .B2(n18160), .ZN(
        n18146) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18162), .B1(
        n18251), .B2(n18212), .ZN(n18145) );
  OAI211_X1 U21264 ( .C1(n18215), .C2(n18192), .A(n18146), .B(n18145), .ZN(
        P3_U2973) );
  AOI22_X1 U21265 ( .A1(n18178), .A2(n18194), .B1(n18216), .B2(n18160), .ZN(
        n18148) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18162), .B1(
        n18251), .B2(n18218), .ZN(n18147) );
  OAI211_X1 U21267 ( .C1(n18181), .C2(n18153), .A(n18148), .B(n18147), .ZN(
        P3_U2974) );
  AOI22_X1 U21268 ( .A1(n18223), .A2(n18161), .B1(n18222), .B2(n18160), .ZN(
        n18150) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18162), .B1(
        n18251), .B2(n18224), .ZN(n18149) );
  OAI211_X1 U21270 ( .C1(n18227), .C2(n18192), .A(n18150), .B(n18149), .ZN(
        P3_U2975) );
  AOI22_X1 U21271 ( .A1(n18229), .A2(n18194), .B1(n18228), .B2(n18160), .ZN(
        n18152) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18162), .B1(
        n18251), .B2(n18230), .ZN(n18151) );
  OAI211_X1 U21273 ( .C1(n18233), .C2(n18153), .A(n18152), .B(n18151), .ZN(
        P3_U2976) );
  AOI22_X1 U21274 ( .A1(n18236), .A2(n18161), .B1(n18234), .B2(n18160), .ZN(
        n18155) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18162), .B1(
        n18251), .B2(n18237), .ZN(n18154) );
  OAI211_X1 U21276 ( .C1(n18240), .C2(n18192), .A(n18155), .B(n18154), .ZN(
        P3_U2977) );
  AOI22_X1 U21277 ( .A1(n18156), .A2(n18161), .B1(n18242), .B2(n18160), .ZN(
        n18158) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18162), .B1(
        n18251), .B2(n18244), .ZN(n18157) );
  OAI211_X1 U21279 ( .C1(n18159), .C2(n18192), .A(n18158), .B(n18157), .ZN(
        P3_U2978) );
  AOI22_X1 U21280 ( .A1(n18195), .A2(n18161), .B1(n18249), .B2(n18160), .ZN(
        n18164) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18162), .B1(
        n18251), .B2(n18252), .ZN(n18163) );
  OAI211_X1 U21282 ( .C1(n18200), .C2(n18192), .A(n18164), .B(n18163), .ZN(
        P3_U2979) );
  INV_X1 U21283 ( .A(n18165), .ZN(n18167) );
  NOR2_X1 U21284 ( .A1(n18166), .A2(n18167), .ZN(n18193) );
  AOI22_X1 U21285 ( .A1(n20659), .A2(n18193), .B1(n20658), .B2(n18194), .ZN(
        n18173) );
  NOR2_X1 U21286 ( .A1(n18194), .A2(n18235), .ZN(n18169) );
  OAI21_X1 U21287 ( .B1(n18169), .B2(n18168), .A(n18167), .ZN(n18170) );
  OAI211_X1 U21288 ( .C1(n18196), .C2(n18419), .A(n18171), .B(n18170), .ZN(
        n18197) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18197), .B1(
        n18206), .B2(n18196), .ZN(n18172) );
  OAI211_X1 U21290 ( .C1(n20665), .C2(n18257), .A(n18173), .B(n18172), .ZN(
        P3_U2980) );
  AOI22_X1 U21291 ( .A1(n18210), .A2(n18193), .B1(n18174), .B2(n18235), .ZN(
        n18176) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18212), .ZN(n18175) );
  OAI211_X1 U21293 ( .C1(n18177), .C2(n18192), .A(n18176), .B(n18175), .ZN(
        P3_U2981) );
  AOI22_X1 U21294 ( .A1(n18178), .A2(n18235), .B1(n18216), .B2(n18193), .ZN(
        n18180) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18218), .ZN(n18179) );
  OAI211_X1 U21296 ( .C1(n18181), .C2(n18192), .A(n18180), .B(n18179), .ZN(
        P3_U2982) );
  AOI22_X1 U21297 ( .A1(n18222), .A2(n18193), .B1(n18182), .B2(n18235), .ZN(
        n18184) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18224), .ZN(n18183) );
  OAI211_X1 U21299 ( .C1(n18185), .C2(n18192), .A(n18184), .B(n18183), .ZN(
        P3_U2983) );
  AOI22_X1 U21300 ( .A1(n18229), .A2(n18235), .B1(n18228), .B2(n18193), .ZN(
        n18187) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18230), .ZN(n18186) );
  OAI211_X1 U21302 ( .C1(n18233), .C2(n18192), .A(n18187), .B(n18186), .ZN(
        P3_U2984) );
  AOI22_X1 U21303 ( .A1(n18236), .A2(n18194), .B1(n18234), .B2(n18193), .ZN(
        n18189) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18237), .ZN(n18188) );
  OAI211_X1 U21305 ( .C1(n18240), .C2(n18257), .A(n18189), .B(n18188), .ZN(
        P3_U2985) );
  AOI22_X1 U21306 ( .A1(n18243), .A2(n18235), .B1(n18242), .B2(n18193), .ZN(
        n18191) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18244), .ZN(n18190) );
  OAI211_X1 U21308 ( .C1(n18247), .C2(n18192), .A(n18191), .B(n18190), .ZN(
        P3_U2986) );
  AOI22_X1 U21309 ( .A1(n18195), .A2(n18194), .B1(n18249), .B2(n18193), .ZN(
        n18199) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18252), .ZN(n18198) );
  OAI211_X1 U21311 ( .C1(n18200), .C2(n18257), .A(n18199), .B(n18198), .ZN(
        P3_U2987) );
  AND2_X1 U21312 ( .A1(n18324), .A2(n18202), .ZN(n18248) );
  AOI22_X1 U21313 ( .A1(n18201), .A2(n18251), .B1(n20659), .B2(n18248), .ZN(
        n18208) );
  AOI22_X1 U21314 ( .A1(n18205), .A2(n18204), .B1(n18203), .B2(n18202), .ZN(
        n18254) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18254), .B1(
        n18206), .B2(n18253), .ZN(n18207) );
  OAI211_X1 U21316 ( .C1(n18209), .C2(n18257), .A(n18208), .B(n18207), .ZN(
        P3_U2988) );
  AOI22_X1 U21317 ( .A1(n18211), .A2(n18235), .B1(n18210), .B2(n18248), .ZN(
        n18214) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18254), .B1(
        n18253), .B2(n18212), .ZN(n18213) );
  OAI211_X1 U21319 ( .C1(n18241), .C2(n18215), .A(n18214), .B(n18213), .ZN(
        P3_U2989) );
  AOI22_X1 U21320 ( .A1(n18217), .A2(n18235), .B1(n18216), .B2(n18248), .ZN(
        n18220) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18254), .B1(
        n18253), .B2(n18218), .ZN(n18219) );
  OAI211_X1 U21322 ( .C1(n18241), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        P3_U2990) );
  AOI22_X1 U21323 ( .A1(n18223), .A2(n18235), .B1(n18222), .B2(n18248), .ZN(
        n18226) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18254), .B1(
        n18253), .B2(n18224), .ZN(n18225) );
  OAI211_X1 U21325 ( .C1(n18241), .C2(n18227), .A(n18226), .B(n18225), .ZN(
        P3_U2991) );
  AOI22_X1 U21326 ( .A1(n18251), .A2(n18229), .B1(n18228), .B2(n18248), .ZN(
        n18232) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18254), .B1(
        n18253), .B2(n18230), .ZN(n18231) );
  OAI211_X1 U21328 ( .C1(n18233), .C2(n18257), .A(n18232), .B(n18231), .ZN(
        P3_U2992) );
  AOI22_X1 U21329 ( .A1(n18236), .A2(n18235), .B1(n18234), .B2(n18248), .ZN(
        n18239) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18254), .B1(
        n18253), .B2(n18237), .ZN(n18238) );
  OAI211_X1 U21331 ( .C1(n18241), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        P3_U2993) );
  AOI22_X1 U21332 ( .A1(n18251), .A2(n18243), .B1(n18242), .B2(n18248), .ZN(
        n18246) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18254), .B1(
        n18253), .B2(n18244), .ZN(n18245) );
  OAI211_X1 U21334 ( .C1(n18247), .C2(n18257), .A(n18246), .B(n18245), .ZN(
        P3_U2994) );
  AOI22_X1 U21335 ( .A1(n18251), .A2(n18250), .B1(n18249), .B2(n18248), .ZN(
        n18256) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18254), .B1(
        n18253), .B2(n18252), .ZN(n18255) );
  OAI211_X1 U21337 ( .C1(n18258), .C2(n18257), .A(n18256), .B(n18255), .ZN(
        P3_U2995) );
  OAI22_X1 U21338 ( .A1(n18262), .A2(n18261), .B1(n18260), .B2(n18259), .ZN(
        n18263) );
  AOI221_X1 U21339 ( .B1(n18266), .B2(n18265), .C1(n18264), .C2(n18265), .A(
        n18263), .ZN(n18464) );
  AOI211_X1 U21340 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18304), .A(
        n18268), .B(n18267), .ZN(n18314) );
  NAND2_X1 U21341 ( .A1(n18270), .A2(n18269), .ZN(n18272) );
  NOR2_X1 U21342 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18294), .ZN(
        n18300) );
  INV_X1 U21343 ( .A(n18300), .ZN(n18271) );
  AOI22_X1 U21344 ( .A1(n18440), .A2(n18272), .B1(n18443), .B2(n18271), .ZN(
        n18437) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18294), .B1(
        n18272), .B2(n18450), .ZN(n18444) );
  AOI222_X1 U21346 ( .A1(n18437), .A2(n18444), .B1(n18437), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18444), .C2(n18273), .ZN(
        n18275) );
  INV_X1 U21347 ( .A(n18304), .ZN(n18291) );
  AOI21_X1 U21348 ( .B1(n18275), .B2(n18291), .A(n18274), .ZN(n18293) );
  AND3_X1 U21349 ( .A1(n18277), .A2(n18299), .A3(n18276), .ZN(n18290) );
  AOI21_X1 U21350 ( .B1(n18280), .B2(n18279), .A(n18278), .ZN(n18297) );
  NOR3_X1 U21351 ( .A1(n18281), .A2(n18297), .A3(n18436), .ZN(n18289) );
  NAND2_X1 U21352 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18282), .ZN(
        n18284) );
  AOI21_X1 U21353 ( .B1(n9600), .B2(n18284), .A(n18283), .ZN(n18288) );
  OAI22_X1 U21354 ( .A1(n9600), .A2(n18285), .B1(n18432), .B2(n18301), .ZN(
        n18287) );
  NOR4_X1 U21355 ( .A1(n18290), .A2(n18289), .A3(n18288), .A4(n18287), .ZN(
        n18428) );
  MUX2_X1 U21356 ( .A(n18436), .B(n18428), .S(n18291), .Z(n18306) );
  OR2_X1 U21357 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18306), .ZN(
        n18292) );
  AOI221_X1 U21358 ( .B1(n18293), .B2(n18292), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18306), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18310) );
  NAND2_X1 U21359 ( .A1(n18299), .A2(n18294), .ZN(n18296) );
  INV_X1 U21360 ( .A(n18302), .ZN(n18295) );
  OAI211_X1 U21361 ( .C1(n18298), .C2(n18297), .A(n18296), .B(n18295), .ZN(
        n18424) );
  NOR2_X1 U21362 ( .A1(n18424), .A2(n18304), .ZN(n18305) );
  OAI22_X1 U21363 ( .A1(n18302), .A2(n18301), .B1(n18300), .B2(n18299), .ZN(
        n18303) );
  NAND2_X1 U21364 ( .A1(n18425), .A2(n18303), .ZN(n18421) );
  OAI22_X1 U21365 ( .A1(n18425), .A2(n18305), .B1(n18304), .B2(n18421), .ZN(
        n18309) );
  OAI21_X1 U21366 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18306), .ZN(n18307) );
  AOI222_X1 U21367 ( .A1(n18310), .A2(n18309), .B1(n18310), .B2(n18308), .C1(
        n18309), .C2(n18307), .ZN(n18313) );
  OAI21_X1 U21368 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18311), .ZN(n18312) );
  NAND4_X1 U21369 ( .A1(n18464), .A2(n18314), .A3(n18313), .A4(n18312), .ZN(
        n18321) );
  AOI211_X1 U21370 ( .C1(n18317), .C2(n18316), .A(n18315), .B(n18321), .ZN(
        n18417) );
  AOI21_X1 U21371 ( .B1(n18473), .B2(n18485), .A(n18417), .ZN(n18325) );
  NAND2_X1 U21372 ( .A1(n18473), .A2(n18467), .ZN(n18329) );
  INV_X1 U21373 ( .A(n18329), .ZN(n18318) );
  AOI211_X1 U21374 ( .C1(n18445), .C2(n18478), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18318), .ZN(n18319) );
  AOI211_X1 U21375 ( .C1(n18470), .C2(n18321), .A(n18320), .B(n18319), .ZN(
        n18322) );
  OAI221_X1 U21376 ( .B1(n18475), .B2(n18325), .C1(n18475), .C2(n18323), .A(
        n18322), .ZN(P3_U2996) );
  NOR4_X1 U21377 ( .A1(n18475), .A2(n18429), .A3(n18466), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18332) );
  INV_X1 U21378 ( .A(n18332), .ZN(n18328) );
  NAND3_X1 U21379 ( .A1(n18326), .A2(n18325), .A3(n18324), .ZN(n18327) );
  NAND4_X1 U21380 ( .A1(n18330), .A2(n18329), .A3(n18328), .A4(n18327), .ZN(
        P3_U2997) );
  OAI21_X1 U21381 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18331), .ZN(n18333) );
  AOI21_X1 U21382 ( .B1(n18334), .B2(n18333), .A(n18332), .ZN(P3_U2998) );
  AND2_X1 U21383 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18335), .ZN(
        P3_U2999) );
  AND2_X1 U21384 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18335), .ZN(
        P3_U3000) );
  AND2_X1 U21385 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18335), .ZN(
        P3_U3001) );
  AND2_X1 U21386 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18335), .ZN(
        P3_U3002) );
  AND2_X1 U21387 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18335), .ZN(
        P3_U3003) );
  AND2_X1 U21388 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18335), .ZN(
        P3_U3004) );
  AND2_X1 U21389 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18335), .ZN(
        P3_U3005) );
  AND2_X1 U21390 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18335), .ZN(
        P3_U3006) );
  AND2_X1 U21391 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18335), .ZN(
        P3_U3007) );
  AND2_X1 U21392 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18335), .ZN(
        P3_U3008) );
  AND2_X1 U21393 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18335), .ZN(
        P3_U3009) );
  AND2_X1 U21394 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18335), .ZN(
        P3_U3010) );
  AND2_X1 U21395 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18335), .ZN(
        P3_U3011) );
  AND2_X1 U21396 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18335), .ZN(
        P3_U3012) );
  AND2_X1 U21397 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18335), .ZN(
        P3_U3013) );
  AND2_X1 U21398 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18335), .ZN(
        P3_U3014) );
  AND2_X1 U21399 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18335), .ZN(
        P3_U3015) );
  AND2_X1 U21400 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18335), .ZN(
        P3_U3016) );
  AND2_X1 U21401 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18335), .ZN(
        P3_U3017) );
  AND2_X1 U21402 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18335), .ZN(
        P3_U3018) );
  AND2_X1 U21403 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18335), .ZN(
        P3_U3019) );
  AND2_X1 U21404 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18335), .ZN(
        P3_U3020) );
  AND2_X1 U21405 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18335), .ZN(P3_U3021) );
  AND2_X1 U21406 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18335), .ZN(P3_U3022) );
  AND2_X1 U21407 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18335), .ZN(P3_U3023) );
  AND2_X1 U21408 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18335), .ZN(P3_U3024) );
  AND2_X1 U21409 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18335), .ZN(P3_U3025) );
  AND2_X1 U21410 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18335), .ZN(P3_U3026) );
  AND2_X1 U21411 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18335), .ZN(P3_U3027) );
  AND2_X1 U21412 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18335), .ZN(P3_U3028) );
  OAI21_X1 U21413 ( .B1(n18336), .B2(n20407), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18337) );
  AOI22_X1 U21414 ( .A1(n18347), .A2(n18349), .B1(n18483), .B2(n18337), .ZN(
        n18338) );
  INV_X1 U21415 ( .A(NA), .ZN(n20413) );
  OR3_X1 U21416 ( .A1(n20413), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18342) );
  OAI211_X1 U21417 ( .C1(n18466), .C2(n18339), .A(n18338), .B(n18342), .ZN(
        P3_U3029) );
  NOR2_X1 U21418 ( .A1(n18349), .A2(n20407), .ZN(n18345) );
  INV_X1 U21419 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18480) );
  OAI22_X1 U21420 ( .A1(n18345), .A2(n18480), .B1(n20407), .B2(n18339), .ZN(
        n18340) );
  AOI21_X1 U21421 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n18340), .A(n18471), 
        .ZN(n18341) );
  NAND2_X1 U21422 ( .A1(n18473), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18343) );
  NAND2_X1 U21423 ( .A1(n18341), .A2(n18343), .ZN(P3_U3030) );
  AOI22_X1 U21424 ( .A1(n18473), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18347), 
        .B2(n18342), .ZN(n18348) );
  OAI22_X1 U21425 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18343), .ZN(n18344) );
  OAI22_X1 U21426 ( .A1(n18345), .A2(n18344), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18346) );
  OAI22_X1 U21427 ( .A1(n18348), .A2(n18349), .B1(n18347), .B2(n18346), .ZN(
        P3_U3031) );
  OAI222_X1 U21428 ( .A1(n18452), .A2(n9595), .B1(n18350), .B2(n18482), .C1(
        n18351), .C2(n18395), .ZN(P3_U3032) );
  OAI222_X1 U21429 ( .A1(n18395), .A2(n18353), .B1(n18352), .B2(n18482), .C1(
        n18351), .C2(n9595), .ZN(P3_U3033) );
  OAI222_X1 U21430 ( .A1(n18395), .A2(n18356), .B1(n18354), .B2(n18482), .C1(
        n18353), .C2(n9595), .ZN(P3_U3034) );
  INV_X1 U21431 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18359) );
  OAI222_X1 U21432 ( .A1(n18395), .A2(n18359), .B1(n18357), .B2(n18482), .C1(
        n18356), .C2(n9595), .ZN(P3_U3035) );
  OAI222_X1 U21433 ( .A1(n18359), .A2(n9595), .B1(n18358), .B2(n18482), .C1(
        n18360), .C2(n18395), .ZN(P3_U3036) );
  OAI222_X1 U21434 ( .A1(n18395), .A2(n18362), .B1(n18361), .B2(n18482), .C1(
        n18360), .C2(n9595), .ZN(P3_U3037) );
  OAI222_X1 U21435 ( .A1(n18395), .A2(n20608), .B1(n18363), .B2(n18482), .C1(
        n18362), .C2(n9595), .ZN(P3_U3038) );
  OAI222_X1 U21436 ( .A1(n20608), .A2(n9595), .B1(n18364), .B2(n18482), .C1(
        n18365), .C2(n18395), .ZN(P3_U3039) );
  OAI222_X1 U21437 ( .A1(n18395), .A2(n18367), .B1(n18366), .B2(n18482), .C1(
        n18365), .C2(n9595), .ZN(P3_U3040) );
  OAI222_X1 U21438 ( .A1(n18395), .A2(n18369), .B1(n18368), .B2(n18482), .C1(
        n18367), .C2(n9595), .ZN(P3_U3041) );
  OAI222_X1 U21439 ( .A1(n18395), .A2(n18371), .B1(n18370), .B2(n18482), .C1(
        n18369), .C2(n9595), .ZN(P3_U3042) );
  OAI222_X1 U21440 ( .A1(n18395), .A2(n18373), .B1(n18372), .B2(n18482), .C1(
        n18371), .C2(n9595), .ZN(P3_U3043) );
  OAI222_X1 U21441 ( .A1(n18395), .A2(n18376), .B1(n18374), .B2(n18482), .C1(
        n18373), .C2(n9595), .ZN(P3_U3044) );
  OAI222_X1 U21442 ( .A1(n18376), .A2(n9595), .B1(n18375), .B2(n18482), .C1(
        n18377), .C2(n18395), .ZN(P3_U3045) );
  INV_X1 U21443 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18379) );
  OAI222_X1 U21444 ( .A1(n18395), .A2(n18379), .B1(n18378), .B2(n18482), .C1(
        n18377), .C2(n9595), .ZN(P3_U3046) );
  OAI222_X1 U21445 ( .A1(n18395), .A2(n18381), .B1(n18380), .B2(n18482), .C1(
        n18379), .C2(n9595), .ZN(P3_U3047) );
  OAI222_X1 U21446 ( .A1(n18395), .A2(n18383), .B1(n18382), .B2(n18482), .C1(
        n18381), .C2(n9595), .ZN(P3_U3048) );
  INV_X1 U21447 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18384) );
  OAI222_X1 U21448 ( .A1(n18395), .A2(n18384), .B1(n20576), .B2(n18482), .C1(
        n18383), .C2(n9595), .ZN(P3_U3049) );
  OAI222_X1 U21449 ( .A1(n18395), .A2(n18387), .B1(n18385), .B2(n18482), .C1(
        n18384), .C2(n9595), .ZN(P3_U3050) );
  OAI222_X1 U21450 ( .A1(n18387), .A2(n9595), .B1(n18386), .B2(n18482), .C1(
        n18388), .C2(n18395), .ZN(P3_U3051) );
  OAI222_X1 U21451 ( .A1(n18395), .A2(n18390), .B1(n18389), .B2(n18482), .C1(
        n18388), .C2(n9595), .ZN(P3_U3052) );
  INV_X1 U21452 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18393) );
  OAI222_X1 U21453 ( .A1(n18395), .A2(n18393), .B1(n18391), .B2(n18482), .C1(
        n18390), .C2(n9595), .ZN(P3_U3053) );
  OAI222_X1 U21454 ( .A1(n18393), .A2(n9595), .B1(n18392), .B2(n18482), .C1(
        n20587), .C2(n18395), .ZN(P3_U3054) );
  INV_X1 U21455 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18396) );
  OAI222_X1 U21456 ( .A1(n18395), .A2(n18396), .B1(n18394), .B2(n18482), .C1(
        n20587), .C2(n9595), .ZN(P3_U3055) );
  OAI222_X1 U21457 ( .A1(n18395), .A2(n18398), .B1(n18397), .B2(n18482), .C1(
        n18396), .C2(n9595), .ZN(P3_U3056) );
  OAI222_X1 U21458 ( .A1(n18395), .A2(n18400), .B1(n18399), .B2(n18482), .C1(
        n18398), .C2(n9595), .ZN(P3_U3057) );
  INV_X1 U21459 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18403) );
  OAI222_X1 U21460 ( .A1(n18395), .A2(n18403), .B1(n18401), .B2(n18482), .C1(
        n18400), .C2(n9595), .ZN(P3_U3058) );
  OAI222_X1 U21461 ( .A1(n18403), .A2(n9595), .B1(n18402), .B2(n18482), .C1(
        n18404), .C2(n18395), .ZN(P3_U3059) );
  OAI222_X1 U21462 ( .A1(n18395), .A2(n18408), .B1(n18405), .B2(n18482), .C1(
        n18404), .C2(n9595), .ZN(P3_U3060) );
  OAI222_X1 U21463 ( .A1(n9595), .A2(n18408), .B1(n18407), .B2(n18482), .C1(
        n18406), .C2(n18395), .ZN(P3_U3061) );
  OAI22_X1 U21464 ( .A1(n18483), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18482), .ZN(n18409) );
  INV_X1 U21465 ( .A(n18409), .ZN(P3_U3274) );
  OAI22_X1 U21466 ( .A1(n18483), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18482), .ZN(n18410) );
  INV_X1 U21467 ( .A(n18410), .ZN(P3_U3275) );
  OAI22_X1 U21468 ( .A1(n18483), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18482), .ZN(n18411) );
  INV_X1 U21469 ( .A(n18411), .ZN(P3_U3276) );
  OAI22_X1 U21470 ( .A1(n18483), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18482), .ZN(n18412) );
  INV_X1 U21471 ( .A(n18412), .ZN(P3_U3277) );
  OAI21_X1 U21472 ( .B1(n18416), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18414), 
        .ZN(n18413) );
  INV_X1 U21473 ( .A(n18413), .ZN(P3_U3280) );
  OAI21_X1 U21474 ( .B1(n18416), .B2(n18415), .A(n18414), .ZN(P3_U3281) );
  NOR2_X1 U21475 ( .A1(n18417), .A2(n18475), .ZN(n18420) );
  OAI21_X1 U21476 ( .B1(n18420), .B2(n18419), .A(n18418), .ZN(P3_U3282) );
  INV_X1 U21477 ( .A(n18421), .ZN(n18423) );
  AOI22_X1 U21478 ( .A1(n18486), .A2(n18423), .B1(n18445), .B2(n18422), .ZN(
        n18427) );
  AOI21_X1 U21479 ( .B1(n18486), .B2(n18424), .A(n18451), .ZN(n18426) );
  OAI22_X1 U21480 ( .A1(n18451), .A2(n18427), .B1(n18426), .B2(n18425), .ZN(
        P3_U3285) );
  INV_X1 U21481 ( .A(n18428), .ZN(n18434) );
  NOR2_X1 U21482 ( .A1(n18429), .A2(n18447), .ZN(n18438) );
  OAI22_X1 U21483 ( .A1(n18431), .A2(n18430), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18439) );
  INV_X1 U21484 ( .A(n18439), .ZN(n18433) );
  AOI222_X1 U21485 ( .A1(n18434), .A2(n18486), .B1(n18438), .B2(n18433), .C1(
        n18445), .C2(n18432), .ZN(n18435) );
  AOI22_X1 U21486 ( .A1(n18451), .A2(n18436), .B1(n18435), .B2(n18448), .ZN(
        P3_U3288) );
  INV_X1 U21487 ( .A(n18437), .ZN(n18441) );
  AOI222_X1 U21488 ( .A1(n18441), .A2(n18486), .B1(n18445), .B2(n18440), .C1(
        n18439), .C2(n18438), .ZN(n18442) );
  AOI22_X1 U21489 ( .A1(n18451), .A2(n18443), .B1(n18442), .B2(n18448), .ZN(
        P3_U3289) );
  INV_X1 U21490 ( .A(n18444), .ZN(n18446) );
  AOI222_X1 U21491 ( .A1(n18447), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18486), 
        .B2(n18446), .C1(n18450), .C2(n18445), .ZN(n18449) );
  AOI22_X1 U21492 ( .A1(n18451), .A2(n18450), .B1(n18449), .B2(n18448), .ZN(
        P3_U3290) );
  AOI21_X1 U21493 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18453) );
  AOI22_X1 U21494 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18453), .B2(n18452), .ZN(n18455) );
  INV_X1 U21495 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U21496 ( .A1(n18456), .A2(n18455), .B1(n18454), .B2(n18459), .ZN(
        P3_U3292) );
  INV_X1 U21497 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18460) );
  NOR2_X1 U21498 ( .A1(n18459), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18457) );
  AOI22_X1 U21499 ( .A1(n18460), .A2(n18459), .B1(n18458), .B2(n18457), .ZN(
        P3_U3293) );
  INV_X1 U21500 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18489) );
  OAI22_X1 U21501 ( .A1(n18483), .A2(n18489), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18482), .ZN(n18461) );
  INV_X1 U21502 ( .A(n18461), .ZN(P3_U3294) );
  INV_X1 U21503 ( .A(n18462), .ZN(n18465) );
  NAND2_X1 U21504 ( .A1(n18465), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18463) );
  OAI21_X1 U21505 ( .B1(n18465), .B2(n18464), .A(n18463), .ZN(P3_U3295) );
  AOI21_X1 U21506 ( .B1(n18467), .B2(n18466), .A(n18488), .ZN(n18468) );
  OAI21_X1 U21507 ( .B1(n18470), .B2(n18469), .A(n18468), .ZN(n18481) );
  OAI21_X1 U21508 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18472), .A(n18471), 
        .ZN(n18474) );
  AOI211_X1 U21509 ( .C1(n18487), .C2(n18474), .A(n18473), .B(n18485), .ZN(
        n18476) );
  NOR2_X1 U21510 ( .A1(n18476), .A2(n18475), .ZN(n18477) );
  OAI21_X1 U21511 ( .B1(n18478), .B2(n18477), .A(n18481), .ZN(n18479) );
  OAI21_X1 U21512 ( .B1(n18481), .B2(n18480), .A(n18479), .ZN(P3_U3296) );
  OAI22_X1 U21513 ( .A1(n18483), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18482), .ZN(n18484) );
  INV_X1 U21514 ( .A(n18484), .ZN(P3_U3297) );
  AOI21_X1 U21515 ( .B1(n18486), .B2(n18485), .A(n18488), .ZN(n18492) );
  AOI22_X1 U21516 ( .A1(n18492), .A2(n18489), .B1(n18488), .B2(n18487), .ZN(
        P3_U3298) );
  INV_X1 U21517 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18491) );
  AOI21_X1 U21518 ( .B1(n18492), .B2(n18491), .A(n18490), .ZN(P3_U3299) );
  INV_X1 U21519 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18496) );
  NAND2_X1 U21520 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19485), .ZN(n19476) );
  NAND2_X1 U21521 ( .A1(n18496), .A2(n18493), .ZN(n19473) );
  OAI21_X1 U21522 ( .B1(n18496), .B2(n19476), .A(n19473), .ZN(n19542) );
  AOI21_X1 U21523 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19542), .ZN(n18494) );
  INV_X1 U21524 ( .A(n18494), .ZN(P2_U2815) );
  INV_X1 U21525 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18497) );
  NAND2_X1 U21526 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18495), .ZN(n19459) );
  OAI22_X1 U21527 ( .A1(n19600), .A2(n18497), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19459), .ZN(P2_U2816) );
  INV_X1 U21528 ( .A(n19468), .ZN(n19480) );
  NAND2_X1 U21529 ( .A1(n18496), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19607) );
  INV_X2 U21530 ( .A(n19607), .ZN(n19606) );
  AOI22_X1 U21531 ( .A1(n19606), .A2(n18497), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19607), .ZN(n18498) );
  OAI21_X1 U21532 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19480), .A(n18498), 
        .ZN(P2_U2817) );
  OAI21_X1 U21533 ( .B1(n19468), .B2(BS16), .A(n19542), .ZN(n19540) );
  OAI21_X1 U21534 ( .B1(n19542), .B2(n19072), .A(n19540), .ZN(P2_U2818) );
  NOR4_X1 U21535 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18502) );
  NOR4_X1 U21536 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18501) );
  NOR4_X1 U21537 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18500) );
  NOR4_X1 U21538 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18499) );
  NAND4_X1 U21539 ( .A1(n18502), .A2(n18501), .A3(n18500), .A4(n18499), .ZN(
        n18508) );
  NOR4_X1 U21540 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18506) );
  AOI211_X1 U21541 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_21__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18505) );
  NOR4_X1 U21542 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18504) );
  NOR4_X1 U21543 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18503) );
  NAND4_X1 U21544 ( .A1(n18506), .A2(n18505), .A3(n18504), .A4(n18503), .ZN(
        n18507) );
  NOR2_X1 U21545 ( .A1(n18508), .A2(n18507), .ZN(n18518) );
  INV_X1 U21546 ( .A(n18518), .ZN(n18516) );
  NOR2_X1 U21547 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18516), .ZN(n18511) );
  INV_X1 U21548 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U21549 ( .A1(n18511), .A2(n18680), .B1(n18516), .B2(n18509), .ZN(
        P2_U2820) );
  OR3_X1 U21550 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18515) );
  INV_X1 U21551 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18510) );
  AOI22_X1 U21552 ( .A1(n18511), .A2(n18515), .B1(n18516), .B2(n18510), .ZN(
        P2_U2821) );
  INV_X1 U21553 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19541) );
  NAND2_X1 U21554 ( .A1(n18511), .A2(n19541), .ZN(n18514) );
  OAI21_X1 U21555 ( .B1(n19486), .B2(n18680), .A(n18518), .ZN(n18512) );
  OAI21_X1 U21556 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18518), .A(n18512), 
        .ZN(n18513) );
  OAI221_X1 U21557 ( .B1(n18514), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18514), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18513), .ZN(P2_U2822) );
  INV_X1 U21558 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18517) );
  OAI221_X1 U21559 ( .B1(n18518), .B2(n18517), .C1(n18516), .C2(n18515), .A(
        n18514), .ZN(P2_U2823) );
  NAND2_X1 U21560 ( .A1(n18519), .A2(n18689), .ZN(n18521) );
  AOI22_X1 U21561 ( .A1(n18563), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18667), .ZN(n18520) );
  OAI211_X1 U21562 ( .C1(n18663), .C2(n18522), .A(n18521), .B(n18520), .ZN(
        n18523) );
  AOI21_X1 U21563 ( .B1(n18524), .B2(n18639), .A(n18523), .ZN(n18530) );
  INV_X1 U21564 ( .A(n18528), .ZN(n18526) );
  OAI221_X1 U21565 ( .B1(n18528), .B2(n18527), .C1(n18526), .C2(n18525), .A(
        n18678), .ZN(n18529) );
  OAI211_X1 U21566 ( .C1(n18676), .C2(n18531), .A(n18530), .B(n18529), .ZN(
        P2_U2834) );
  NAND2_X1 U21567 ( .A1(n18669), .A2(n18532), .ZN(n18533) );
  XOR2_X1 U21568 ( .A(n18534), .B(n18533), .Z(n18543) );
  AOI22_X1 U21569 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18677), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n18667), .ZN(n18535) );
  OAI21_X1 U21570 ( .B1(n18536), .B2(n18687), .A(n18535), .ZN(n18537) );
  AOI211_X1 U21571 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18563), .A(n18815), .B(
        n18537), .ZN(n18542) );
  OAI22_X1 U21572 ( .A1(n18539), .A2(n18656), .B1(n18676), .B2(n18538), .ZN(
        n18540) );
  INV_X1 U21573 ( .A(n18540), .ZN(n18541) );
  OAI211_X1 U21574 ( .C1(n19465), .C2(n18543), .A(n18542), .B(n18541), .ZN(
        P2_U2836) );
  NOR2_X1 U21575 ( .A1(n18653), .A2(n18544), .ZN(n18546) );
  XOR2_X1 U21576 ( .A(n18546), .B(n18545), .Z(n18556) );
  INV_X1 U21577 ( .A(n18547), .ZN(n18549) );
  AOI22_X1 U21578 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18677), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18667), .ZN(n18548) );
  OAI21_X1 U21579 ( .B1(n18549), .B2(n18687), .A(n18548), .ZN(n18550) );
  AOI211_X1 U21580 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n18563), .A(n18815), .B(
        n18550), .ZN(n18555) );
  OAI22_X1 U21581 ( .A1(n18552), .A2(n18656), .B1(n18551), .B2(n18676), .ZN(
        n18553) );
  INV_X1 U21582 ( .A(n18553), .ZN(n18554) );
  OAI211_X1 U21583 ( .C1(n19465), .C2(n18556), .A(n18555), .B(n18554), .ZN(
        P2_U2837) );
  NAND2_X1 U21584 ( .A1(n18669), .A2(n18557), .ZN(n18558) );
  XOR2_X1 U21585 ( .A(n18559), .B(n18558), .Z(n18569) );
  AOI22_X1 U21586 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n18667), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18677), .ZN(n18560) );
  OAI21_X1 U21587 ( .B1(n18561), .B2(n18687), .A(n18560), .ZN(n18562) );
  AOI211_X1 U21588 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18563), .A(n18815), .B(
        n18562), .ZN(n18568) );
  OAI22_X1 U21589 ( .A1(n18565), .A2(n18656), .B1(n18564), .B2(n18676), .ZN(
        n18566) );
  INV_X1 U21590 ( .A(n18566), .ZN(n18567) );
  OAI211_X1 U21591 ( .C1(n19465), .C2(n18569), .A(n18568), .B(n18567), .ZN(
        P2_U2838) );
  NOR2_X1 U21592 ( .A1(n18653), .A2(n18570), .ZN(n18572) );
  XOR2_X1 U21593 ( .A(n18572), .B(n18571), .Z(n18579) );
  AOI22_X1 U21594 ( .A1(n18573), .A2(n18639), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18677), .ZN(n18574) );
  OAI211_X1 U21595 ( .C1(n18679), .C2(n9804), .A(n18574), .B(n18662), .ZN(
        n18575) );
  AOI21_X1 U21596 ( .B1(P2_REIP_REG_16__SCAN_IN), .B2(n18667), .A(n18575), 
        .ZN(n18578) );
  AOI22_X1 U21597 ( .A1(n18576), .A2(n18689), .B1(n18684), .B2(n18704), .ZN(
        n18577) );
  OAI211_X1 U21598 ( .C1(n19465), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P2_U2839) );
  NAND2_X1 U21599 ( .A1(n18669), .A2(n18580), .ZN(n18582) );
  XOR2_X1 U21600 ( .A(n18582), .B(n18581), .Z(n18589) );
  AOI22_X1 U21601 ( .A1(n18583), .A2(n18639), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18677), .ZN(n18584) );
  OAI211_X1 U21602 ( .C1(n18679), .C2(n12071), .A(n18584), .B(n18662), .ZN(
        n18587) );
  OAI22_X1 U21603 ( .A1(n18585), .A2(n18656), .B1(n18676), .B2(n18710), .ZN(
        n18586) );
  AOI211_X1 U21604 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18667), .A(n18587), 
        .B(n18586), .ZN(n18588) );
  OAI21_X1 U21605 ( .B1(n18589), .B2(n19465), .A(n18588), .ZN(P2_U2840) );
  OAI21_X1 U21606 ( .B1(n18679), .B2(n12064), .A(n18662), .ZN(n18594) );
  INV_X1 U21607 ( .A(n18590), .ZN(n18592) );
  OAI22_X1 U21608 ( .A1(n18592), .A2(n18687), .B1(n18663), .B2(n18591), .ZN(
        n18593) );
  AOI211_X1 U21609 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18667), .A(n18594), 
        .B(n18593), .ZN(n18601) );
  NAND2_X1 U21610 ( .A1(n18669), .A2(n18595), .ZN(n18596) );
  XNOR2_X1 U21611 ( .A(n18597), .B(n18596), .ZN(n18599) );
  AOI22_X1 U21612 ( .A1(n18599), .A2(n18678), .B1(n18689), .B2(n18598), .ZN(
        n18600) );
  OAI211_X1 U21613 ( .C1(n18715), .C2(n18676), .A(n18601), .B(n18600), .ZN(
        P2_U2842) );
  OAI21_X1 U21614 ( .B1(n18679), .B2(n12059), .A(n18662), .ZN(n18605) );
  OAI22_X1 U21615 ( .A1(n18603), .A2(n18687), .B1(n18663), .B2(n18602), .ZN(
        n18604) );
  AOI211_X1 U21616 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n18667), .A(n18605), 
        .B(n18604), .ZN(n18612) );
  NAND2_X1 U21617 ( .A1(n18669), .A2(n18606), .ZN(n18607) );
  XNOR2_X1 U21618 ( .A(n18608), .B(n18607), .ZN(n18610) );
  AOI22_X1 U21619 ( .A1(n18610), .A2(n18678), .B1(n18689), .B2(n18609), .ZN(
        n18611) );
  OAI211_X1 U21620 ( .C1(n18721), .C2(n18676), .A(n18612), .B(n18611), .ZN(
        P2_U2844) );
  NOR2_X1 U21621 ( .A1(n18653), .A2(n18613), .ZN(n18614) );
  XOR2_X1 U21622 ( .A(n18615), .B(n18614), .Z(n18623) );
  AOI22_X1 U21623 ( .A1(n18616), .A2(n18639), .B1(P2_REIP_REG_10__SCAN_IN), 
        .B2(n18667), .ZN(n18617) );
  OAI211_X1 U21624 ( .C1(n18679), .C2(n12026), .A(n18617), .B(n18662), .ZN(
        n18621) );
  INV_X1 U21625 ( .A(n18618), .ZN(n18619) );
  OAI22_X1 U21626 ( .A1(n18619), .A2(n18656), .B1(n18676), .B2(n18724), .ZN(
        n18620) );
  AOI211_X1 U21627 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18677), .A(
        n18621), .B(n18620), .ZN(n18622) );
  OAI21_X1 U21628 ( .B1(n19465), .B2(n18623), .A(n18622), .ZN(P2_U2845) );
  OAI21_X1 U21629 ( .B1(n18679), .B2(n9978), .A(n18662), .ZN(n18628) );
  INV_X1 U21630 ( .A(n18624), .ZN(n18626) );
  OAI22_X1 U21631 ( .A1(n18626), .A2(n18687), .B1(n18663), .B2(n18625), .ZN(
        n18627) );
  AOI211_X1 U21632 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18667), .A(n18628), .B(
        n18627), .ZN(n18635) );
  NAND2_X1 U21633 ( .A1(n18669), .A2(n18629), .ZN(n18630) );
  XNOR2_X1 U21634 ( .A(n18631), .B(n18630), .ZN(n18633) );
  AOI22_X1 U21635 ( .A1(n18633), .A2(n18678), .B1(n18689), .B2(n18632), .ZN(
        n18634) );
  OAI211_X1 U21636 ( .C1(n18726), .C2(n18676), .A(n18635), .B(n18634), .ZN(
        P2_U2846) );
  NAND2_X1 U21637 ( .A1(n18669), .A2(n18636), .ZN(n18638) );
  XOR2_X1 U21638 ( .A(n18638), .B(n18637), .Z(n18646) );
  AOI22_X1 U21639 ( .A1(n18640), .A2(n18639), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18677), .ZN(n18641) );
  OAI211_X1 U21640 ( .C1(n18679), .C2(n12950), .A(n18641), .B(n18662), .ZN(
        n18644) );
  OAI22_X1 U21641 ( .A1(n18642), .A2(n18656), .B1(n18676), .B2(n18730), .ZN(
        n18643) );
  AOI211_X1 U21642 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n18667), .A(n18644), .B(
        n18643), .ZN(n18645) );
  OAI21_X1 U21643 ( .B1(n18646), .B2(n19465), .A(n18645), .ZN(P2_U2848) );
  OAI22_X1 U21644 ( .A1(n18647), .A2(n18687), .B1(n18663), .B2(n10008), .ZN(
        n18648) );
  INV_X1 U21645 ( .A(n18648), .ZN(n18649) );
  OAI211_X1 U21646 ( .C1(n18650), .C2(n18679), .A(n18662), .B(n18649), .ZN(
        n18651) );
  INV_X1 U21647 ( .A(n18651), .ZN(n18661) );
  NOR2_X1 U21648 ( .A1(n18653), .A2(n18652), .ZN(n18654) );
  XNOR2_X1 U21649 ( .A(n18655), .B(n18654), .ZN(n18659) );
  OAI22_X1 U21650 ( .A1(n18657), .A2(n18656), .B1(n18676), .B2(n18731), .ZN(
        n18658) );
  AOI21_X1 U21651 ( .B1(n18659), .B2(n18678), .A(n18658), .ZN(n18660) );
  OAI211_X1 U21652 ( .C1(n19495), .C2(n18681), .A(n18661), .B(n18660), .ZN(
        P2_U2849) );
  OAI21_X1 U21653 ( .B1(n18679), .B2(n12045), .A(n18662), .ZN(n18666) );
  OAI22_X1 U21654 ( .A1(n18664), .A2(n18687), .B1(n18663), .B2(n15822), .ZN(
        n18665) );
  AOI211_X1 U21655 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18667), .A(n18666), .B(
        n18665), .ZN(n18675) );
  NAND2_X1 U21656 ( .A1(n18669), .A2(n18668), .ZN(n18670) );
  XNOR2_X1 U21657 ( .A(n18671), .B(n18670), .ZN(n18673) );
  AOI22_X1 U21658 ( .A1(n18673), .A2(n18678), .B1(n18689), .B2(n18672), .ZN(
        n18674) );
  OAI211_X1 U21659 ( .C1(n18676), .C2(n18738), .A(n18675), .B(n18674), .ZN(
        P2_U2850) );
  NOR2_X1 U21660 ( .A1(n18678), .A2(n18677), .ZN(n18695) );
  INV_X1 U21661 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18694) );
  OAI22_X1 U21662 ( .A1(n18681), .A2(n18680), .B1(n18679), .B2(n12203), .ZN(
        n18682) );
  AOI21_X1 U21663 ( .B1(n18684), .B2(n18683), .A(n18682), .ZN(n18685) );
  OAI21_X1 U21664 ( .B1(n18687), .B2(n18686), .A(n18685), .ZN(n18688) );
  AOI21_X1 U21665 ( .B1(n18690), .B2(n18689), .A(n18688), .ZN(n18693) );
  NAND2_X1 U21666 ( .A1(n18691), .A2(n19127), .ZN(n18692) );
  OAI211_X1 U21667 ( .C1(n18695), .C2(n18694), .A(n18693), .B(n18692), .ZN(
        P2_U2855) );
  INV_X1 U21668 ( .A(n18696), .ZN(n18697) );
  AOI22_X1 U21669 ( .A1(n18697), .A2(n18757), .B1(n18702), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18699) );
  AOI22_X1 U21670 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n18756), .B1(n18703), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n18698) );
  NAND2_X1 U21671 ( .A1(n18699), .A2(n18698), .ZN(P2_U2888) );
  INV_X1 U21672 ( .A(n18866), .ZN(n18700) );
  AOI22_X1 U21673 ( .A1(n18701), .A2(n18700), .B1(n18756), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n18708) );
  AOI22_X1 U21674 ( .A1(n18703), .A2(BUF1_REG_16__SCAN_IN), .B1(n18702), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18707) );
  AOI22_X1 U21675 ( .A1(n18705), .A2(n18761), .B1(n18757), .B2(n18704), .ZN(
        n18706) );
  NAND3_X1 U21676 ( .A1(n18708), .A2(n18707), .A3(n18706), .ZN(P2_U2903) );
  OAI222_X1 U21677 ( .A1(n18710), .A2(n18739), .B1(n12224), .B2(n18755), .C1(
        n18709), .C2(n18765), .ZN(P2_U2904) );
  AOI22_X1 U21678 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n18756), .B1(n18711), 
        .B2(n18747), .ZN(n18712) );
  OAI21_X1 U21679 ( .B1(n18739), .B2(n18713), .A(n18712), .ZN(P2_U2905) );
  INV_X1 U21680 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18771) );
  OAI222_X1 U21681 ( .A1(n18715), .A2(n18739), .B1(n18771), .B2(n18755), .C1(
        n18765), .C2(n18714), .ZN(P2_U2906) );
  INV_X1 U21682 ( .A(n18716), .ZN(n18719) );
  AOI22_X1 U21683 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n18756), .B1(n18717), 
        .B2(n18747), .ZN(n18718) );
  OAI21_X1 U21684 ( .B1(n18739), .B2(n18719), .A(n18718), .ZN(P2_U2907) );
  INV_X1 U21685 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18775) );
  OAI222_X1 U21686 ( .A1(n18721), .A2(n18739), .B1(n18775), .B2(n18755), .C1(
        n18765), .C2(n18720), .ZN(P2_U2908) );
  AOI22_X1 U21687 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n18756), .B1(n18722), 
        .B2(n18747), .ZN(n18723) );
  OAI21_X1 U21688 ( .B1(n18739), .B2(n18724), .A(n18723), .ZN(P2_U2909) );
  INV_X1 U21689 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18779) );
  OAI222_X1 U21690 ( .A1(n18726), .A2(n18739), .B1(n18779), .B2(n18755), .C1(
        n18765), .C2(n18725), .ZN(P2_U2910) );
  INV_X1 U21691 ( .A(n18727), .ZN(n18729) );
  INV_X1 U21692 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18781) );
  OAI222_X1 U21693 ( .A1(n18729), .A2(n18739), .B1(n18781), .B2(n18755), .C1(
        n18765), .C2(n18728), .ZN(P2_U2911) );
  OAI222_X1 U21694 ( .A1(n18730), .A2(n18739), .B1(n18783), .B2(n18755), .C1(
        n18765), .C2(n18911), .ZN(P2_U2912) );
  OAI222_X1 U21695 ( .A1(n18731), .A2(n18739), .B1(n18785), .B2(n18755), .C1(
        n18765), .C2(n18902), .ZN(P2_U2913) );
  INV_X1 U21696 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18787) );
  OAI22_X1 U21697 ( .A1(n18787), .A2(n18755), .B1(n18897), .B2(n18765), .ZN(
        n18732) );
  INV_X1 U21698 ( .A(n18732), .ZN(n18737) );
  OR3_X1 U21699 ( .A1(n18735), .A2(n18734), .A3(n18733), .ZN(n18736) );
  OAI211_X1 U21700 ( .C1(n18739), .C2(n18738), .A(n18737), .B(n18736), .ZN(
        P2_U2914) );
  INV_X1 U21701 ( .A(n19546), .ZN(n18740) );
  AOI22_X1 U21702 ( .A1(n18740), .A2(n18757), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n18756), .ZN(n18746) );
  OAI21_X1 U21703 ( .B1(n18743), .B2(n18742), .A(n18741), .ZN(n18744) );
  NAND2_X1 U21704 ( .A1(n18744), .A2(n18761), .ZN(n18745) );
  OAI211_X1 U21705 ( .C1(n18887), .C2(n18765), .A(n18746), .B(n18745), .ZN(
        P2_U2916) );
  AOI22_X1 U21706 ( .A1(n19558), .A2(n18757), .B1(n18748), .B2(n18747), .ZN(
        n18754) );
  OAI21_X1 U21707 ( .B1(n18751), .B2(n18750), .A(n18749), .ZN(n18752) );
  NAND2_X1 U21708 ( .A1(n18752), .A2(n18761), .ZN(n18753) );
  OAI211_X1 U21709 ( .C1(n18755), .C2(n18793), .A(n18754), .B(n18753), .ZN(
        P2_U2917) );
  AOI22_X1 U21710 ( .A1(n18757), .A2(n19568), .B1(n18756), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n18764) );
  OAI21_X1 U21711 ( .B1(n18760), .B2(n18759), .A(n18758), .ZN(n18762) );
  NAND2_X1 U21712 ( .A1(n18762), .A2(n18761), .ZN(n18763) );
  OAI211_X1 U21713 ( .C1(n18878), .C2(n18765), .A(n18764), .B(n18763), .ZN(
        P2_U2918) );
  AND2_X1 U21714 ( .A1(n18796), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U21715 ( .A1(n19603), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18767) );
  OAI21_X1 U21716 ( .B1(n12224), .B2(n18799), .A(n18767), .ZN(P2_U2936) );
  AOI22_X1 U21717 ( .A1(n19603), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18768) );
  OAI21_X1 U21718 ( .B1(n18769), .B2(n18799), .A(n18768), .ZN(P2_U2937) );
  AOI22_X1 U21719 ( .A1(n19603), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18770) );
  OAI21_X1 U21720 ( .B1(n18771), .B2(n18799), .A(n18770), .ZN(P2_U2938) );
  AOI22_X1 U21721 ( .A1(n19603), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18772) );
  OAI21_X1 U21722 ( .B1(n18773), .B2(n18799), .A(n18772), .ZN(P2_U2939) );
  AOI22_X1 U21723 ( .A1(n19603), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18774) );
  OAI21_X1 U21724 ( .B1(n18775), .B2(n18799), .A(n18774), .ZN(P2_U2940) );
  AOI22_X1 U21725 ( .A1(n19603), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18776) );
  OAI21_X1 U21726 ( .B1(n18777), .B2(n18799), .A(n18776), .ZN(P2_U2941) );
  AOI22_X1 U21727 ( .A1(n19603), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18778) );
  OAI21_X1 U21728 ( .B1(n18779), .B2(n18799), .A(n18778), .ZN(P2_U2942) );
  AOI22_X1 U21729 ( .A1(n19603), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18780) );
  OAI21_X1 U21730 ( .B1(n18781), .B2(n18799), .A(n18780), .ZN(P2_U2943) );
  AOI22_X1 U21731 ( .A1(n18797), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18782) );
  OAI21_X1 U21732 ( .B1(n18783), .B2(n18799), .A(n18782), .ZN(P2_U2944) );
  AOI22_X1 U21733 ( .A1(n18797), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18784) );
  OAI21_X1 U21734 ( .B1(n18785), .B2(n18799), .A(n18784), .ZN(P2_U2945) );
  AOI22_X1 U21735 ( .A1(n18797), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18786) );
  OAI21_X1 U21736 ( .B1(n18787), .B2(n18799), .A(n18786), .ZN(P2_U2946) );
  INV_X1 U21737 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18789) );
  AOI22_X1 U21738 ( .A1(n18797), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18788) );
  OAI21_X1 U21739 ( .B1(n18789), .B2(n18799), .A(n18788), .ZN(P2_U2947) );
  INV_X1 U21740 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18791) );
  AOI22_X1 U21741 ( .A1(n18797), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18790) );
  OAI21_X1 U21742 ( .B1(n18791), .B2(n18799), .A(n18790), .ZN(P2_U2948) );
  AOI22_X1 U21743 ( .A1(n18797), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18792) );
  OAI21_X1 U21744 ( .B1(n18793), .B2(n18799), .A(n18792), .ZN(P2_U2949) );
  AOI22_X1 U21745 ( .A1(n18797), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18794) );
  OAI21_X1 U21746 ( .B1(n18795), .B2(n18799), .A(n18794), .ZN(P2_U2950) );
  AOI22_X1 U21747 ( .A1(n18797), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18796), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18798) );
  OAI21_X1 U21748 ( .B1(n12221), .B2(n18799), .A(n18798), .ZN(P2_U2951) );
  AOI22_X1 U21749 ( .A1(n18810), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n18815), .ZN(n18804) );
  AOI222_X1 U21750 ( .A1(n18802), .A2(n18811), .B1(n18819), .B2(n18801), .C1(
        n18800), .C2(n18814), .ZN(n18803) );
  OAI211_X1 U21751 ( .C1(n18817), .C2(n18805), .A(n18804), .B(n18803), .ZN(
        P2_U3010) );
  OAI21_X1 U21752 ( .B1(n18808), .B2(n18807), .A(n18806), .ZN(n18809) );
  XOR2_X1 U21753 ( .A(n18809), .B(n18850), .Z(n18843) );
  AOI22_X1 U21754 ( .A1(n18843), .A2(n18811), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18810), .ZN(n18821) );
  AOI21_X1 U21755 ( .B1(n18850), .B2(n18813), .A(n18812), .ZN(n18845) );
  NAND2_X1 U21756 ( .A1(n18845), .A2(n18814), .ZN(n18816) );
  NAND2_X1 U21757 ( .A1(n18815), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n18848) );
  OAI211_X1 U21758 ( .C1(n18817), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18816), .B(n18848), .ZN(n18818) );
  AOI21_X1 U21759 ( .B1(n12719), .B2(n18819), .A(n18818), .ZN(n18820) );
  NAND2_X1 U21760 ( .A1(n18821), .A2(n18820), .ZN(P2_U3013) );
  INV_X1 U21761 ( .A(n19558), .ZN(n18833) );
  NAND2_X1 U21762 ( .A1(n18823), .A2(n18822), .ZN(n18828) );
  NAND3_X1 U21763 ( .A1(n18825), .A2(n18844), .A3(n18824), .ZN(n18826) );
  NAND3_X1 U21764 ( .A1(n18828), .A2(n18827), .A3(n18826), .ZN(n18829) );
  AOI21_X1 U21765 ( .B1(n18853), .B2(n18830), .A(n18829), .ZN(n18831) );
  OAI21_X1 U21766 ( .B1(n18833), .B2(n18832), .A(n18831), .ZN(n18834) );
  AOI21_X1 U21767 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18835), .A(
        n18834), .ZN(n18840) );
  OAI21_X1 U21768 ( .B1(n18838), .B2(n18837), .A(n18836), .ZN(n18839) );
  OAI211_X1 U21769 ( .C1(n18842), .C2(n18841), .A(n18840), .B(n18839), .ZN(
        P2_U3044) );
  AOI22_X1 U21770 ( .A1(n18846), .A2(n18845), .B1(n18844), .B2(n18843), .ZN(
        n18858) );
  NAND2_X1 U21771 ( .A1(n18847), .A2(n19568), .ZN(n18849) );
  OAI211_X1 U21772 ( .C1(n18851), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        n18852) );
  AOI21_X1 U21773 ( .B1(n12719), .B2(n18853), .A(n18852), .ZN(n18857) );
  OAI211_X1 U21774 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n18855), .B(n18854), .ZN(n18856) );
  NAND3_X1 U21775 ( .A1(n18858), .A2(n18857), .A3(n18856), .ZN(P2_U3045) );
  NAND2_X1 U21776 ( .A1(n19355), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19566) );
  NAND2_X1 U21777 ( .A1(n19158), .A2(n19068), .ZN(n18906) );
  NAND2_X1 U21778 ( .A1(n19554), .A2(n19560), .ZN(n18978) );
  NOR2_X1 U21779 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18978), .ZN(
        n18927) );
  INV_X1 U21780 ( .A(n18927), .ZN(n18923) );
  NOR2_X1 U21781 ( .A1(n18923), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18914) );
  INV_X1 U21782 ( .A(n18914), .ZN(n18862) );
  AND2_X1 U21783 ( .A1(n18863), .A2(n18862), .ZN(n18865) );
  OAI21_X1 U21784 ( .B1(n18869), .B2(n18914), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n18864) );
  OAI21_X1 U21785 ( .B1(n18865), .B2(n19550), .A(n18864), .ZN(n18915) );
  NOR2_X2 U21786 ( .A1(n18868), .A2(n18898), .ZN(n19399) );
  AOI22_X1 U21787 ( .A1(n18915), .A2(n18867), .B1(n19399), .B2(n18914), .ZN(
        n18877) );
  INV_X1 U21788 ( .A(n18869), .ZN(n18874) );
  INV_X1 U21789 ( .A(n19297), .ZN(n18870) );
  OAI21_X1 U21790 ( .B1(n19436), .B2(n18944), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n18871) );
  INV_X1 U21791 ( .A(n18871), .ZN(n18872) );
  OAI21_X1 U21792 ( .B1(n19448), .B2(n18872), .A(n19571), .ZN(n18873) );
  AOI21_X1 U21793 ( .B1(n18874), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n18873), 
        .ZN(n18875) );
  OAI21_X1 U21794 ( .B1(n18875), .B2(n18914), .A(n19405), .ZN(n18918) );
  AOI22_X1 U21795 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18916), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n18917), .ZN(n19367) );
  AOI22_X1 U21796 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18918), .B1(
        n19436), .B2(n19407), .ZN(n18876) );
  OAI211_X1 U21797 ( .C1(n19410), .C2(n18906), .A(n18877), .B(n18876), .ZN(
        P2_U3048) );
  AOI22_X1 U21798 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18916), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n18917), .ZN(n19415) );
  NOR2_X2 U21799 ( .A1(n13275), .A2(n18898), .ZN(n19411) );
  AOI22_X1 U21800 ( .A1(n18915), .A2(n18879), .B1(n19411), .B2(n18914), .ZN(
        n18881) );
  AOI22_X1 U21801 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18916), .ZN(n19371) );
  INV_X1 U21802 ( .A(n19371), .ZN(n19412) );
  AOI22_X1 U21803 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18918), .B1(
        n18944), .B2(n19412), .ZN(n18880) );
  OAI211_X1 U21804 ( .C1(n19415), .C2(n19456), .A(n18881), .B(n18880), .ZN(
        P2_U3049) );
  AOI22_X1 U21805 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18916), .ZN(n19322) );
  NOR2_X2 U21806 ( .A1(n18884), .A2(n18898), .ZN(n19416) );
  AOI22_X1 U21807 ( .A1(n18915), .A2(n18883), .B1(n19416), .B2(n18914), .ZN(
        n18886) );
  AOI22_X1 U21808 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18916), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n18917), .ZN(n19420) );
  AOI22_X1 U21809 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18918), .B1(
        n19436), .B2(n19319), .ZN(n18885) );
  OAI211_X1 U21810 ( .C1(n19322), .C2(n18906), .A(n18886), .B(n18885), .ZN(
        P2_U3050) );
  AOI22_X1 U21811 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18916), .ZN(n19426) );
  NOR2_X2 U21812 ( .A1(n18887), .A2(n19162), .ZN(n19422) );
  INV_X1 U21813 ( .A(n18898), .ZN(n18912) );
  AOI22_X1 U21814 ( .A1(n18915), .A2(n19422), .B1(n19421), .B2(n18914), .ZN(
        n18890) );
  AOI22_X1 U21815 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18916), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n18917), .ZN(n19377) );
  AOI22_X1 U21816 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18918), .B1(
        n19436), .B2(n19423), .ZN(n18889) );
  OAI211_X1 U21817 ( .C1(n19426), .C2(n18906), .A(n18890), .B(n18889), .ZN(
        P2_U3051) );
  AOI22_X1 U21818 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18916), .ZN(n19432) );
  NOR2_X2 U21819 ( .A1(n18891), .A2(n19162), .ZN(n19428) );
  NOR2_X2 U21820 ( .A1(n18892), .A2(n18898), .ZN(n19427) );
  AOI22_X1 U21821 ( .A1(n18915), .A2(n19428), .B1(n19427), .B2(n18914), .ZN(
        n18894) );
  AOI22_X1 U21822 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18916), .ZN(n19381) );
  INV_X1 U21823 ( .A(n19381), .ZN(n19429) );
  AOI22_X1 U21824 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18918), .B1(
        n18944), .B2(n19429), .ZN(n18893) );
  OAI211_X1 U21825 ( .C1(n19432), .C2(n19456), .A(n18894), .B(n18893), .ZN(
        P2_U3052) );
  INV_X1 U21826 ( .A(n18917), .ZN(n18909) );
  INV_X1 U21827 ( .A(n18916), .ZN(n18907) );
  INV_X1 U21828 ( .A(n19382), .ZN(n19440) );
  NOR2_X2 U21829 ( .A1(n18897), .A2(n19162), .ZN(n19434) );
  NOR2_X2 U21830 ( .A1(n18899), .A2(n18898), .ZN(n19433) );
  AOI22_X1 U21831 ( .A1(n18915), .A2(n19434), .B1(n19433), .B2(n18914), .ZN(
        n18901) );
  AOI22_X1 U21832 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18916), .ZN(n19385) );
  AOI22_X1 U21833 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18918), .B1(
        n18944), .B2(n19435), .ZN(n18900) );
  OAI211_X1 U21834 ( .C1(n19440), .C2(n19456), .A(n18901), .B(n18900), .ZN(
        P2_U3053) );
  AOI22_X2 U21835 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n18916), .ZN(n19446) );
  NOR2_X2 U21836 ( .A1(n18902), .A2(n19162), .ZN(n19442) );
  AND2_X1 U21837 ( .A1(n18903), .A2(n18912), .ZN(n19441) );
  AOI22_X1 U21838 ( .A1(n18915), .A2(n19442), .B1(n19441), .B2(n18914), .ZN(
        n18905) );
  AOI22_X1 U21839 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18916), .ZN(n19390) );
  AOI22_X1 U21840 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18918), .B1(
        n19436), .B2(n19443), .ZN(n18904) );
  OAI211_X1 U21841 ( .C1(n19446), .C2(n18906), .A(n18905), .B(n18904), .ZN(
        P2_U3054) );
  OAI22_X2 U21842 ( .A1(n18910), .A2(n18909), .B1(n18908), .B2(n18907), .ZN(
        n19451) );
  INV_X1 U21843 ( .A(n19451), .ZN(n19263) );
  NOR2_X2 U21844 ( .A1(n18911), .A2(n19162), .ZN(n19449) );
  AND2_X1 U21845 ( .A1(n18913), .A2(n18912), .ZN(n19447) );
  AOI22_X1 U21846 ( .A1(n18915), .A2(n19449), .B1(n19447), .B2(n18914), .ZN(
        n18920) );
  AOI22_X1 U21847 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n18917), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18916), .ZN(n19457) );
  INV_X1 U21848 ( .A(n19457), .ZN(n19291) );
  AOI22_X1 U21849 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18918), .B1(
        n18944), .B2(n19291), .ZN(n18919) );
  OAI211_X1 U21850 ( .C1(n19263), .C2(n19456), .A(n18920), .B(n18919), .ZN(
        P2_U3055) );
  NOR2_X1 U21851 ( .A1(n19159), .A2(n18978), .ZN(n18942) );
  NOR3_X1 U21852 ( .A1(n18922), .A2(n18942), .A3(n18921), .ZN(n18924) );
  AOI211_X2 U21853 ( .C1(n18923), .C2(n18921), .A(n19011), .B(n18924), .ZN(
        n18943) );
  AOI22_X1 U21854 ( .A1(n18943), .A2(n18867), .B1(n19399), .B2(n18942), .ZN(
        n18929) );
  AND2_X1 U21855 ( .A1(n19160), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19100) );
  INV_X1 U21856 ( .A(n18942), .ZN(n18925) );
  AOI211_X1 U21857 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n18925), .A(n19162), 
        .B(n18924), .ZN(n18926) );
  OAI221_X1 U21858 ( .B1(n18927), .B2(n19158), .C1(n18927), .C2(n19100), .A(
        n18926), .ZN(n18945) );
  AOI22_X1 U21859 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19407), .ZN(n18928) );
  OAI211_X1 U21860 ( .C1(n19410), .C2(n18956), .A(n18929), .B(n18928), .ZN(
        P2_U3056) );
  AOI22_X1 U21861 ( .A1(n18943), .A2(n18879), .B1(n19411), .B2(n18942), .ZN(
        n18931) );
  INV_X1 U21862 ( .A(n19415), .ZN(n19368) );
  AOI22_X1 U21863 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19368), .ZN(n18930) );
  OAI211_X1 U21864 ( .C1(n19371), .C2(n18956), .A(n18931), .B(n18930), .ZN(
        P2_U3057) );
  AOI22_X1 U21865 ( .A1(n18943), .A2(n18883), .B1(n19416), .B2(n18942), .ZN(
        n18933) );
  AOI22_X1 U21866 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19319), .ZN(n18932) );
  OAI211_X1 U21867 ( .C1(n19322), .C2(n18956), .A(n18933), .B(n18932), .ZN(
        P2_U3058) );
  AOI22_X1 U21868 ( .A1(n18943), .A2(n19422), .B1(n19421), .B2(n18942), .ZN(
        n18935) );
  AOI22_X1 U21869 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19423), .ZN(n18934) );
  OAI211_X1 U21870 ( .C1(n19426), .C2(n18956), .A(n18935), .B(n18934), .ZN(
        P2_U3059) );
  AOI22_X1 U21871 ( .A1(n18943), .A2(n19428), .B1(n19427), .B2(n18942), .ZN(
        n18937) );
  AOI22_X1 U21872 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19378), .ZN(n18936) );
  OAI211_X1 U21873 ( .C1(n19381), .C2(n18956), .A(n18937), .B(n18936), .ZN(
        P2_U3060) );
  AOI22_X1 U21874 ( .A1(n18943), .A2(n19434), .B1(n19433), .B2(n18942), .ZN(
        n18939) );
  AOI22_X1 U21875 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19382), .ZN(n18938) );
  OAI211_X1 U21876 ( .C1(n19385), .C2(n18956), .A(n18939), .B(n18938), .ZN(
        P2_U3061) );
  AOI22_X1 U21877 ( .A1(n18943), .A2(n19442), .B1(n19441), .B2(n18942), .ZN(
        n18941) );
  AOI22_X1 U21878 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19443), .ZN(n18940) );
  OAI211_X1 U21879 ( .C1(n19446), .C2(n18956), .A(n18941), .B(n18940), .ZN(
        P2_U3062) );
  AOI22_X1 U21880 ( .A1(n18943), .A2(n19449), .B1(n19447), .B2(n18942), .ZN(
        n18947) );
  AOI22_X1 U21881 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18945), .B1(
        n18944), .B2(n19451), .ZN(n18946) );
  OAI211_X1 U21882 ( .C1(n19457), .C2(n18956), .A(n18947), .B(n18946), .ZN(
        P2_U3063) );
  NOR3_X2 U21883 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19570), .A3(
        n18978), .ZN(n18971) );
  OAI21_X1 U21884 ( .B1(n18950), .B2(n18971), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n18949) );
  NOR2_X1 U21885 ( .A1(n19192), .A2(n18978), .ZN(n18951) );
  INV_X1 U21886 ( .A(n18951), .ZN(n18948) );
  NAND2_X1 U21887 ( .A1(n18949), .A2(n18948), .ZN(n18972) );
  AOI22_X1 U21888 ( .A1(n18972), .A2(n18867), .B1(n19399), .B2(n18971), .ZN(
        n18958) );
  AOI21_X1 U21889 ( .B1(n18950), .B2(n19571), .A(n18971), .ZN(n18954) );
  AOI21_X1 U21890 ( .B1(n19007), .B2(n18956), .A(n19072), .ZN(n18952) );
  NOR2_X1 U21891 ( .A1(n18952), .A2(n18951), .ZN(n18953) );
  MUX2_X1 U21892 ( .A(n18954), .B(n18953), .S(n19355), .Z(n18955) );
  AOI22_X1 U21893 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19407), .ZN(n18957) );
  OAI211_X1 U21894 ( .C1(n19410), .C2(n19007), .A(n18958), .B(n18957), .ZN(
        P2_U3064) );
  AOI22_X1 U21895 ( .A1(n18972), .A2(n18879), .B1(n19411), .B2(n18971), .ZN(
        n18960) );
  AOI22_X1 U21896 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19368), .ZN(n18959) );
  OAI211_X1 U21897 ( .C1(n19371), .C2(n19007), .A(n18960), .B(n18959), .ZN(
        P2_U3065) );
  AOI22_X1 U21898 ( .A1(n18972), .A2(n18883), .B1(n19416), .B2(n18971), .ZN(
        n18962) );
  AOI22_X1 U21899 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19319), .ZN(n18961) );
  OAI211_X1 U21900 ( .C1(n19322), .C2(n19007), .A(n18962), .B(n18961), .ZN(
        P2_U3066) );
  AOI22_X1 U21901 ( .A1(n18972), .A2(n19422), .B1(n19421), .B2(n18971), .ZN(
        n18964) );
  AOI22_X1 U21902 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19423), .ZN(n18963) );
  OAI211_X1 U21903 ( .C1(n19426), .C2(n19007), .A(n18964), .B(n18963), .ZN(
        P2_U3067) );
  AOI22_X1 U21904 ( .A1(n18972), .A2(n19428), .B1(n19427), .B2(n18971), .ZN(
        n18966) );
  AOI22_X1 U21905 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19378), .ZN(n18965) );
  OAI211_X1 U21906 ( .C1(n19381), .C2(n19007), .A(n18966), .B(n18965), .ZN(
        P2_U3068) );
  AOI22_X1 U21907 ( .A1(n18972), .A2(n19434), .B1(n19433), .B2(n18971), .ZN(
        n18968) );
  AOI22_X1 U21908 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19382), .ZN(n18967) );
  OAI211_X1 U21909 ( .C1(n19385), .C2(n19007), .A(n18968), .B(n18967), .ZN(
        P2_U3069) );
  AOI22_X1 U21910 ( .A1(n18972), .A2(n19442), .B1(n19441), .B2(n18971), .ZN(
        n18970) );
  AOI22_X1 U21911 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19443), .ZN(n18969) );
  OAI211_X1 U21912 ( .C1(n19446), .C2(n19007), .A(n18970), .B(n18969), .ZN(
        P2_U3070) );
  AOI22_X1 U21913 ( .A1(n18972), .A2(n19449), .B1(n19447), .B2(n18971), .ZN(
        n18976) );
  AOI22_X1 U21914 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19451), .ZN(n18975) );
  OAI211_X1 U21915 ( .C1(n19457), .C2(n19007), .A(n18976), .B(n18975), .ZN(
        P2_U3071) );
  INV_X1 U21916 ( .A(n19410), .ZN(n19354) );
  INV_X1 U21917 ( .A(n18978), .ZN(n18977) );
  AND2_X1 U21918 ( .A1(n19221), .A2(n18977), .ZN(n19002) );
  AOI22_X1 U21919 ( .A1(n19354), .A2(n19035), .B1(n19002), .B2(n19399), .ZN(
        n18988) );
  INV_X1 U21920 ( .A(n19100), .ZN(n19039) );
  OAI21_X1 U21921 ( .B1(n19039), .B2(n19235), .A(n19355), .ZN(n18986) );
  NOR2_X1 U21922 ( .A1(n19570), .A2(n18978), .ZN(n18982) );
  INV_X1 U21923 ( .A(n18983), .ZN(n18980) );
  INV_X1 U21924 ( .A(n19002), .ZN(n18979) );
  OAI211_X1 U21925 ( .C1(n18980), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n18979), 
        .B(n19550), .ZN(n18981) );
  OAI211_X1 U21926 ( .C1(n18986), .C2(n18982), .A(n19405), .B(n18981), .ZN(
        n19004) );
  INV_X1 U21927 ( .A(n18982), .ZN(n18985) );
  OAI21_X1 U21928 ( .B1(n18983), .B2(n19002), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n18984) );
  OAI21_X1 U21929 ( .B1(n18986), .B2(n18985), .A(n18984), .ZN(n19003) );
  AOI22_X1 U21930 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19004), .B1(
        n18867), .B2(n19003), .ZN(n18987) );
  OAI211_X1 U21931 ( .C1(n19367), .C2(n19007), .A(n18988), .B(n18987), .ZN(
        P2_U3072) );
  AOI22_X1 U21932 ( .A1(n19412), .A2(n19035), .B1(n19002), .B2(n19411), .ZN(
        n18990) );
  AOI22_X1 U21933 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19004), .B1(
        n18879), .B2(n19003), .ZN(n18989) );
  OAI211_X1 U21934 ( .C1(n19415), .C2(n19007), .A(n18990), .B(n18989), .ZN(
        P2_U3073) );
  INV_X1 U21935 ( .A(n19322), .ZN(n19417) );
  AOI22_X1 U21936 ( .A1(n19417), .A2(n19035), .B1(n19002), .B2(n19416), .ZN(
        n18992) );
  AOI22_X1 U21937 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19004), .B1(
        n18883), .B2(n19003), .ZN(n18991) );
  OAI211_X1 U21938 ( .C1(n19420), .C2(n19007), .A(n18992), .B(n18991), .ZN(
        P2_U3074) );
  INV_X1 U21939 ( .A(n19426), .ZN(n19374) );
  AOI22_X1 U21940 ( .A1(n19374), .A2(n19035), .B1(n19002), .B2(n19421), .ZN(
        n18994) );
  AOI22_X1 U21941 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19004), .B1(
        n19422), .B2(n19003), .ZN(n18993) );
  OAI211_X1 U21942 ( .C1(n19377), .C2(n19007), .A(n18994), .B(n18993), .ZN(
        P2_U3075) );
  INV_X1 U21943 ( .A(n19035), .ZN(n19013) );
  INV_X1 U21944 ( .A(n19007), .ZN(n18995) );
  AOI22_X1 U21945 ( .A1(n19378), .A2(n18995), .B1(n19002), .B2(n19427), .ZN(
        n18997) );
  AOI22_X1 U21946 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19004), .B1(
        n19428), .B2(n19003), .ZN(n18996) );
  OAI211_X1 U21947 ( .C1(n19381), .C2(n19013), .A(n18997), .B(n18996), .ZN(
        P2_U3076) );
  AOI22_X1 U21948 ( .A1(n19435), .A2(n19035), .B1(n19002), .B2(n19433), .ZN(
        n18999) );
  AOI22_X1 U21949 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19004), .B1(
        n19434), .B2(n19003), .ZN(n18998) );
  OAI211_X1 U21950 ( .C1(n19440), .C2(n19007), .A(n18999), .B(n18998), .ZN(
        P2_U3077) );
  INV_X1 U21951 ( .A(n19446), .ZN(n19386) );
  AOI22_X1 U21952 ( .A1(n19386), .A2(n19035), .B1(n19002), .B2(n19441), .ZN(
        n19001) );
  AOI22_X1 U21953 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19004), .B1(
        n19442), .B2(n19003), .ZN(n19000) );
  OAI211_X1 U21954 ( .C1(n19390), .C2(n19007), .A(n19001), .B(n19000), .ZN(
        P2_U3078) );
  AOI22_X1 U21955 ( .A1(n19291), .A2(n19035), .B1(n19002), .B2(n19447), .ZN(
        n19006) );
  AOI22_X1 U21956 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19004), .B1(
        n19449), .B2(n19003), .ZN(n19005) );
  OAI211_X1 U21957 ( .C1(n19263), .C2(n19007), .A(n19006), .B(n19005), .ZN(
        P2_U3079) );
  INV_X1 U21958 ( .A(n19296), .ZN(n19304) );
  NOR2_X1 U21959 ( .A1(n19009), .A2(n19008), .ZN(n19264) );
  NAND2_X1 U21960 ( .A1(n19264), .A2(n19554), .ZN(n19012) );
  NOR3_X1 U21961 ( .A1(n19560), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19043) );
  NAND2_X1 U21962 ( .A1(n19578), .A2(n19043), .ZN(n19015) );
  INV_X1 U21963 ( .A(n19015), .ZN(n19033) );
  NOR3_X1 U21964 ( .A1(n19010), .A2(n19033), .A3(n18921), .ZN(n19014) );
  AOI211_X2 U21965 ( .C1(n19012), .C2(n18921), .A(n19011), .B(n19014), .ZN(
        n19034) );
  AOI22_X1 U21966 ( .A1(n19034), .A2(n18867), .B1(n19399), .B2(n19033), .ZN(
        n19020) );
  INV_X1 U21967 ( .A(n19012), .ZN(n19018) );
  AOI21_X1 U21968 ( .B1(n19013), .B2(n19056), .A(n19072), .ZN(n19017) );
  AOI211_X1 U21969 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19015), .A(n19162), 
        .B(n19014), .ZN(n19016) );
  AOI22_X1 U21970 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19407), .ZN(n19019) );
  OAI211_X1 U21971 ( .C1(n19410), .C2(n19056), .A(n19020), .B(n19019), .ZN(
        P2_U3080) );
  AOI22_X1 U21972 ( .A1(n19034), .A2(n18879), .B1(n19411), .B2(n19033), .ZN(
        n19022) );
  AOI22_X1 U21973 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19368), .ZN(n19021) );
  OAI211_X1 U21974 ( .C1(n19371), .C2(n19056), .A(n19022), .B(n19021), .ZN(
        P2_U3081) );
  AOI22_X1 U21975 ( .A1(n19034), .A2(n18883), .B1(n19416), .B2(n19033), .ZN(
        n19024) );
  AOI22_X1 U21976 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19319), .ZN(n19023) );
  OAI211_X1 U21977 ( .C1(n19322), .C2(n19056), .A(n19024), .B(n19023), .ZN(
        P2_U3082) );
  AOI22_X1 U21978 ( .A1(n19034), .A2(n19422), .B1(n19421), .B2(n19033), .ZN(
        n19026) );
  AOI22_X1 U21979 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19423), .ZN(n19025) );
  OAI211_X1 U21980 ( .C1(n19426), .C2(n19056), .A(n19026), .B(n19025), .ZN(
        P2_U3083) );
  AOI22_X1 U21981 ( .A1(n19034), .A2(n19428), .B1(n19427), .B2(n19033), .ZN(
        n19028) );
  AOI22_X1 U21982 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19378), .ZN(n19027) );
  OAI211_X1 U21983 ( .C1(n19381), .C2(n19056), .A(n19028), .B(n19027), .ZN(
        P2_U3084) );
  AOI22_X1 U21984 ( .A1(n19034), .A2(n19434), .B1(n19433), .B2(n19033), .ZN(
        n19030) );
  AOI22_X1 U21985 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19382), .ZN(n19029) );
  OAI211_X1 U21986 ( .C1(n19385), .C2(n19056), .A(n19030), .B(n19029), .ZN(
        P2_U3085) );
  AOI22_X1 U21987 ( .A1(n19034), .A2(n19442), .B1(n19441), .B2(n19033), .ZN(
        n19032) );
  AOI22_X1 U21988 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19443), .ZN(n19031) );
  OAI211_X1 U21989 ( .C1(n19446), .C2(n19056), .A(n19032), .B(n19031), .ZN(
        P2_U3086) );
  AOI22_X1 U21990 ( .A1(n19034), .A2(n19449), .B1(n19447), .B2(n19033), .ZN(
        n19038) );
  AOI22_X1 U21991 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19451), .ZN(n19037) );
  OAI211_X1 U21992 ( .C1(n19457), .C2(n19056), .A(n19038), .B(n19037), .ZN(
        P2_U3087) );
  INV_X1 U21993 ( .A(n19043), .ZN(n19046) );
  NOR2_X1 U21994 ( .A1(n19578), .A2(n19046), .ZN(n19074) );
  AOI22_X1 U21995 ( .A1(n19354), .A2(n19094), .B1(n19399), .B2(n19074), .ZN(
        n19049) );
  OAI21_X1 U21996 ( .B1(n19039), .B2(n19296), .A(n19355), .ZN(n19047) );
  INV_X1 U21997 ( .A(n19044), .ZN(n19041) );
  INV_X1 U21998 ( .A(n19074), .ZN(n19040) );
  OAI211_X1 U21999 ( .C1(n19041), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19040), 
        .B(n19550), .ZN(n19042) );
  OAI211_X1 U22000 ( .C1(n19047), .C2(n19043), .A(n19405), .B(n19042), .ZN(
        n19065) );
  OAI21_X1 U22001 ( .B1(n19044), .B2(n19074), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19045) );
  OAI21_X1 U22002 ( .B1(n19047), .B2(n19046), .A(n19045), .ZN(n19064) );
  AOI22_X1 U22003 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19065), .B1(
        n18867), .B2(n19064), .ZN(n19048) );
  OAI211_X1 U22004 ( .C1(n19367), .C2(n19056), .A(n19049), .B(n19048), .ZN(
        P2_U3088) );
  AOI22_X1 U22005 ( .A1(n19368), .A2(n19063), .B1(n19411), .B2(n19074), .ZN(
        n19051) );
  AOI22_X1 U22006 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19065), .B1(
        n18879), .B2(n19064), .ZN(n19050) );
  OAI211_X1 U22007 ( .C1(n19371), .C2(n19089), .A(n19051), .B(n19050), .ZN(
        P2_U3089) );
  AOI22_X1 U22008 ( .A1(n19319), .A2(n19063), .B1(n19416), .B2(n19074), .ZN(
        n19053) );
  AOI22_X1 U22009 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19065), .B1(
        n18883), .B2(n19064), .ZN(n19052) );
  OAI211_X1 U22010 ( .C1(n19322), .C2(n19089), .A(n19053), .B(n19052), .ZN(
        P2_U3090) );
  AOI22_X1 U22011 ( .A1(n19374), .A2(n19094), .B1(n19421), .B2(n19074), .ZN(
        n19055) );
  AOI22_X1 U22012 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19065), .B1(
        n19422), .B2(n19064), .ZN(n19054) );
  OAI211_X1 U22013 ( .C1(n19377), .C2(n19056), .A(n19055), .B(n19054), .ZN(
        P2_U3091) );
  AOI22_X1 U22014 ( .A1(n19378), .A2(n19063), .B1(n19427), .B2(n19074), .ZN(
        n19058) );
  AOI22_X1 U22015 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19065), .B1(
        n19428), .B2(n19064), .ZN(n19057) );
  OAI211_X1 U22016 ( .C1(n19381), .C2(n19089), .A(n19058), .B(n19057), .ZN(
        P2_U3092) );
  AOI22_X1 U22017 ( .A1(n19382), .A2(n19063), .B1(n19433), .B2(n19074), .ZN(
        n19060) );
  AOI22_X1 U22018 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19065), .B1(
        n19434), .B2(n19064), .ZN(n19059) );
  OAI211_X1 U22019 ( .C1(n19385), .C2(n19089), .A(n19060), .B(n19059), .ZN(
        P2_U3093) );
  AOI22_X1 U22020 ( .A1(n19443), .A2(n19063), .B1(n19441), .B2(n19074), .ZN(
        n19062) );
  AOI22_X1 U22021 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19065), .B1(
        n19442), .B2(n19064), .ZN(n19061) );
  OAI211_X1 U22022 ( .C1(n19446), .C2(n19089), .A(n19062), .B(n19061), .ZN(
        P2_U3094) );
  AOI22_X1 U22023 ( .A1(n19451), .A2(n19063), .B1(n19447), .B2(n19074), .ZN(
        n19067) );
  AOI22_X1 U22024 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19065), .B1(
        n19449), .B2(n19064), .ZN(n19066) );
  OAI211_X1 U22025 ( .C1(n19457), .C2(n19089), .A(n19067), .B(n19066), .ZN(
        P2_U3095) );
  NAND3_X1 U22026 ( .A1(n19554), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19101) );
  NOR2_X1 U22027 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19101), .ZN(
        n19092) );
  NOR2_X1 U22028 ( .A1(n19074), .A2(n19092), .ZN(n19069) );
  OR2_X1 U22029 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19069), .ZN(n19071) );
  NOR3_X1 U22030 ( .A1(n19070), .A2(n19092), .A3(n18921), .ZN(n19075) );
  AOI21_X1 U22031 ( .B1(n18921), .B2(n19071), .A(n19075), .ZN(n19093) );
  AOI22_X1 U22032 ( .A1(n19093), .A2(n18867), .B1(n19399), .B2(n19092), .ZN(
        n19078) );
  AOI21_X1 U22033 ( .B1(n19089), .B2(n19126), .A(n19072), .ZN(n19073) );
  AOI221_X1 U22034 ( .B1(n19571), .B2(n19074), .C1(n19571), .C2(n19073), .A(
        n19092), .ZN(n19076) );
  OR3_X1 U22035 ( .A1(n19076), .A2(n19075), .A3(n19162), .ZN(n19095) );
  AOI22_X1 U22036 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19407), .ZN(n19077) );
  OAI211_X1 U22037 ( .C1(n19410), .C2(n19126), .A(n19078), .B(n19077), .ZN(
        P2_U3096) );
  AOI22_X1 U22038 ( .A1(n19093), .A2(n18879), .B1(n19411), .B2(n19092), .ZN(
        n19080) );
  AOI22_X1 U22039 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19368), .ZN(n19079) );
  OAI211_X1 U22040 ( .C1(n19371), .C2(n19126), .A(n19080), .B(n19079), .ZN(
        P2_U3097) );
  AOI22_X1 U22041 ( .A1(n19093), .A2(n18883), .B1(n19416), .B2(n19092), .ZN(
        n19082) );
  AOI22_X1 U22042 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19319), .ZN(n19081) );
  OAI211_X1 U22043 ( .C1(n19322), .C2(n19126), .A(n19082), .B(n19081), .ZN(
        P2_U3098) );
  AOI22_X1 U22044 ( .A1(n19093), .A2(n19422), .B1(n19421), .B2(n19092), .ZN(
        n19084) );
  INV_X1 U22045 ( .A(n19126), .ZN(n19119) );
  AOI22_X1 U22046 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19095), .B1(
        n19119), .B2(n19374), .ZN(n19083) );
  OAI211_X1 U22047 ( .C1(n19377), .C2(n19089), .A(n19084), .B(n19083), .ZN(
        P2_U3099) );
  AOI22_X1 U22048 ( .A1(n19093), .A2(n19428), .B1(n19427), .B2(n19092), .ZN(
        n19086) );
  AOI22_X1 U22049 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19378), .ZN(n19085) );
  OAI211_X1 U22050 ( .C1(n19381), .C2(n19126), .A(n19086), .B(n19085), .ZN(
        P2_U3100) );
  AOI22_X1 U22051 ( .A1(n19093), .A2(n19434), .B1(n19433), .B2(n19092), .ZN(
        n19088) );
  AOI22_X1 U22052 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19095), .B1(
        n19119), .B2(n19435), .ZN(n19087) );
  OAI211_X1 U22053 ( .C1(n19440), .C2(n19089), .A(n19088), .B(n19087), .ZN(
        P2_U3101) );
  AOI22_X1 U22054 ( .A1(n19093), .A2(n19442), .B1(n19441), .B2(n19092), .ZN(
        n19091) );
  AOI22_X1 U22055 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19443), .ZN(n19090) );
  OAI211_X1 U22056 ( .C1(n19446), .C2(n19126), .A(n19091), .B(n19090), .ZN(
        P2_U3102) );
  AOI22_X1 U22057 ( .A1(n19093), .A2(n19449), .B1(n19447), .B2(n19092), .ZN(
        n19097) );
  AOI22_X1 U22058 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19451), .ZN(n19096) );
  OAI211_X1 U22059 ( .C1(n19457), .C2(n19126), .A(n19097), .B(n19096), .ZN(
        P2_U3103) );
  NOR2_X1 U22060 ( .A1(n19578), .A2(n19101), .ZN(n19134) );
  OAI21_X1 U22061 ( .B1(n19102), .B2(n19134), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19099) );
  OAI21_X1 U22062 ( .B1(n19101), .B2(n19550), .A(n19099), .ZN(n19122) );
  AOI22_X1 U22063 ( .A1(n19122), .A2(n18867), .B1(n19399), .B2(n19134), .ZN(
        n19108) );
  NAND2_X1 U22064 ( .A1(n19100), .A2(n19544), .ZN(n19551) );
  INV_X1 U22065 ( .A(n19551), .ZN(n19106) );
  INV_X1 U22066 ( .A(n19101), .ZN(n19105) );
  INV_X1 U22067 ( .A(n19102), .ZN(n19103) );
  INV_X1 U22068 ( .A(n19134), .ZN(n19131) );
  OAI211_X1 U22069 ( .C1(n19103), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19131), 
        .B(n19550), .ZN(n19104) );
  OAI211_X1 U22070 ( .C1(n19106), .C2(n19105), .A(n19405), .B(n19104), .ZN(
        n19123) );
  AOI22_X1 U22071 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19123), .B1(
        n19119), .B2(n19407), .ZN(n19107) );
  OAI211_X1 U22072 ( .C1(n19410), .C2(n19157), .A(n19108), .B(n19107), .ZN(
        P2_U3104) );
  AOI22_X1 U22073 ( .A1(n19122), .A2(n18879), .B1(n19411), .B2(n19134), .ZN(
        n19110) );
  AOI22_X1 U22074 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19123), .B1(
        n19149), .B2(n19412), .ZN(n19109) );
  OAI211_X1 U22075 ( .C1(n19415), .C2(n19126), .A(n19110), .B(n19109), .ZN(
        P2_U3105) );
  AOI22_X1 U22076 ( .A1(n19122), .A2(n18883), .B1(n19416), .B2(n19134), .ZN(
        n19112) );
  AOI22_X1 U22077 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19123), .B1(
        n19149), .B2(n19417), .ZN(n19111) );
  OAI211_X1 U22078 ( .C1(n19420), .C2(n19126), .A(n19112), .B(n19111), .ZN(
        P2_U3106) );
  AOI22_X1 U22079 ( .A1(n19122), .A2(n19422), .B1(n19421), .B2(n19134), .ZN(
        n19114) );
  AOI22_X1 U22080 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19123), .B1(
        n19149), .B2(n19374), .ZN(n19113) );
  OAI211_X1 U22081 ( .C1(n19377), .C2(n19126), .A(n19114), .B(n19113), .ZN(
        P2_U3107) );
  AOI22_X1 U22082 ( .A1(n19122), .A2(n19428), .B1(n19427), .B2(n19134), .ZN(
        n19116) );
  AOI22_X1 U22083 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19123), .B1(
        n19149), .B2(n19429), .ZN(n19115) );
  OAI211_X1 U22084 ( .C1(n19432), .C2(n19126), .A(n19116), .B(n19115), .ZN(
        P2_U3108) );
  AOI22_X1 U22085 ( .A1(n19122), .A2(n19434), .B1(n19433), .B2(n19134), .ZN(
        n19118) );
  AOI22_X1 U22086 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19123), .B1(
        n19149), .B2(n19435), .ZN(n19117) );
  OAI211_X1 U22087 ( .C1(n19440), .C2(n19126), .A(n19118), .B(n19117), .ZN(
        P2_U3109) );
  AOI22_X1 U22088 ( .A1(n19122), .A2(n19442), .B1(n19441), .B2(n19134), .ZN(
        n19121) );
  AOI22_X1 U22089 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19123), .B1(
        n19119), .B2(n19443), .ZN(n19120) );
  OAI211_X1 U22090 ( .C1(n19446), .C2(n19157), .A(n19121), .B(n19120), .ZN(
        P2_U3110) );
  AOI22_X1 U22091 ( .A1(n19122), .A2(n19449), .B1(n19447), .B2(n19134), .ZN(
        n19125) );
  AOI22_X1 U22092 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19123), .B1(
        n19149), .B2(n19291), .ZN(n19124) );
  OAI211_X1 U22093 ( .C1(n19263), .C2(n19126), .A(n19125), .B(n19124), .ZN(
        P2_U3111) );
  INV_X1 U22094 ( .A(n19353), .ZN(n19128) );
  NAND2_X1 U22095 ( .A1(n19560), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19224) );
  NOR2_X1 U22096 ( .A1(n19224), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19166) );
  INV_X1 U22097 ( .A(n19166), .ZN(n19169) );
  NOR2_X1 U22098 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19169), .ZN(
        n19152) );
  AOI22_X1 U22099 ( .A1(n19407), .A2(n19149), .B1(n19152), .B2(n19399), .ZN(
        n19138) );
  NAND2_X1 U22100 ( .A1(n19183), .A2(n19157), .ZN(n19129) );
  AOI21_X1 U22101 ( .B1(n19129), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19550), 
        .ZN(n19133) );
  OAI21_X1 U22102 ( .B1(n13233), .B2(n18921), .A(n19571), .ZN(n19130) );
  AOI21_X1 U22103 ( .B1(n19133), .B2(n19131), .A(n19130), .ZN(n19132) );
  OAI21_X1 U22104 ( .B1(n19152), .B2(n19132), .A(n19405), .ZN(n19154) );
  OAI21_X1 U22105 ( .B1(n19134), .B2(n19152), .A(n19133), .ZN(n19136) );
  OAI21_X1 U22106 ( .B1(n13233), .B2(n19152), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19135) );
  NAND2_X1 U22107 ( .A1(n19136), .A2(n19135), .ZN(n19153) );
  AOI22_X1 U22108 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19154), .B1(
        n18867), .B2(n19153), .ZN(n19137) );
  OAI211_X1 U22109 ( .C1(n19410), .C2(n19183), .A(n19138), .B(n19137), .ZN(
        P2_U3112) );
  AOI22_X1 U22110 ( .A1(n19412), .A2(n19186), .B1(n19411), .B2(n19152), .ZN(
        n19140) );
  AOI22_X1 U22111 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n18879), .ZN(n19139) );
  OAI211_X1 U22112 ( .C1(n19415), .C2(n19157), .A(n19140), .B(n19139), .ZN(
        P2_U3113) );
  AOI22_X1 U22113 ( .A1(n19319), .A2(n19149), .B1(n19152), .B2(n19416), .ZN(
        n19142) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n18883), .ZN(n19141) );
  OAI211_X1 U22115 ( .C1(n19322), .C2(n19183), .A(n19142), .B(n19141), .ZN(
        P2_U3114) );
  AOI22_X1 U22116 ( .A1(n19423), .A2(n19149), .B1(n19152), .B2(n19421), .ZN(
        n19144) );
  AOI22_X1 U22117 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19422), .ZN(n19143) );
  OAI211_X1 U22118 ( .C1(n19426), .C2(n19183), .A(n19144), .B(n19143), .ZN(
        P2_U3115) );
  AOI22_X1 U22119 ( .A1(n19429), .A2(n19186), .B1(n19427), .B2(n19152), .ZN(
        n19146) );
  AOI22_X1 U22120 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19428), .ZN(n19145) );
  OAI211_X1 U22121 ( .C1(n19432), .C2(n19157), .A(n19146), .B(n19145), .ZN(
        P2_U3116) );
  AOI22_X1 U22122 ( .A1(n19435), .A2(n19186), .B1(n19433), .B2(n19152), .ZN(
        n19148) );
  AOI22_X1 U22123 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19434), .ZN(n19147) );
  OAI211_X1 U22124 ( .C1(n19440), .C2(n19157), .A(n19148), .B(n19147), .ZN(
        P2_U3117) );
  AOI22_X1 U22125 ( .A1(n19443), .A2(n19149), .B1(n19152), .B2(n19441), .ZN(
        n19151) );
  AOI22_X1 U22126 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19442), .ZN(n19150) );
  OAI211_X1 U22127 ( .C1(n19446), .C2(n19183), .A(n19151), .B(n19150), .ZN(
        P2_U3118) );
  AOI22_X1 U22128 ( .A1(n19291), .A2(n19186), .B1(n19447), .B2(n19152), .ZN(
        n19156) );
  AOI22_X1 U22129 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19449), .ZN(n19155) );
  OAI211_X1 U22130 ( .C1(n19263), .C2(n19157), .A(n19156), .B(n19155), .ZN(
        P2_U3119) );
  INV_X1 U22131 ( .A(n19158), .ZN(n19161) );
  NOR2_X1 U22132 ( .A1(n19159), .A2(n19224), .ZN(n19193) );
  AOI22_X1 U22133 ( .A1(n19407), .A2(n19186), .B1(n19399), .B2(n19193), .ZN(
        n19172) );
  INV_X1 U22134 ( .A(n19160), .ZN(n19548) );
  NAND2_X1 U22135 ( .A1(n19548), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19228) );
  OAI21_X1 U22136 ( .B1(n19228), .B2(n19161), .A(n19355), .ZN(n19170) );
  INV_X1 U22137 ( .A(n13217), .ZN(n19167) );
  OAI21_X1 U22138 ( .B1(n19167), .B2(n18921), .A(n19571), .ZN(n19164) );
  INV_X1 U22139 ( .A(n19193), .ZN(n19163) );
  AOI21_X1 U22140 ( .B1(n19164), .B2(n19163), .A(n19162), .ZN(n19165) );
  OAI21_X1 U22141 ( .B1(n19170), .B2(n19166), .A(n19165), .ZN(n19188) );
  OAI21_X1 U22142 ( .B1(n19167), .B2(n19193), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19168) );
  OAI21_X1 U22143 ( .B1(n19170), .B2(n19169), .A(n19168), .ZN(n19187) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19188), .B1(
        n18867), .B2(n19187), .ZN(n19171) );
  OAI211_X1 U22145 ( .C1(n19410), .C2(n19219), .A(n19172), .B(n19171), .ZN(
        P2_U3120) );
  AOI22_X1 U22146 ( .A1(n19368), .A2(n19186), .B1(n19411), .B2(n19193), .ZN(
        n19174) );
  AOI22_X1 U22147 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19188), .B1(
        n18879), .B2(n19187), .ZN(n19173) );
  OAI211_X1 U22148 ( .C1(n19371), .C2(n19219), .A(n19174), .B(n19173), .ZN(
        P2_U3121) );
  AOI22_X1 U22149 ( .A1(n19319), .A2(n19186), .B1(n19193), .B2(n19416), .ZN(
        n19176) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19188), .B1(
        n18883), .B2(n19187), .ZN(n19175) );
  OAI211_X1 U22151 ( .C1(n19322), .C2(n19219), .A(n19176), .B(n19175), .ZN(
        P2_U3122) );
  AOI22_X1 U22152 ( .A1(n19374), .A2(n19210), .B1(n19193), .B2(n19421), .ZN(
        n19178) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19188), .B1(
        n19422), .B2(n19187), .ZN(n19177) );
  OAI211_X1 U22154 ( .C1(n19377), .C2(n19183), .A(n19178), .B(n19177), .ZN(
        P2_U3123) );
  AOI22_X1 U22155 ( .A1(n19378), .A2(n19186), .B1(n19427), .B2(n19193), .ZN(
        n19180) );
  AOI22_X1 U22156 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19188), .B1(
        n19428), .B2(n19187), .ZN(n19179) );
  OAI211_X1 U22157 ( .C1(n19381), .C2(n19219), .A(n19180), .B(n19179), .ZN(
        P2_U3124) );
  AOI22_X1 U22158 ( .A1(n19435), .A2(n19210), .B1(n19433), .B2(n19193), .ZN(
        n19182) );
  AOI22_X1 U22159 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19188), .B1(
        n19434), .B2(n19187), .ZN(n19181) );
  OAI211_X1 U22160 ( .C1(n19440), .C2(n19183), .A(n19182), .B(n19181), .ZN(
        P2_U3125) );
  AOI22_X1 U22161 ( .A1(n19443), .A2(n19186), .B1(n19193), .B2(n19441), .ZN(
        n19185) );
  AOI22_X1 U22162 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19188), .B1(
        n19442), .B2(n19187), .ZN(n19184) );
  OAI211_X1 U22163 ( .C1(n19446), .C2(n19219), .A(n19185), .B(n19184), .ZN(
        P2_U3126) );
  AOI22_X1 U22164 ( .A1(n19451), .A2(n19186), .B1(n19447), .B2(n19193), .ZN(
        n19190) );
  AOI22_X1 U22165 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19188), .B1(
        n19449), .B2(n19187), .ZN(n19189) );
  OAI211_X1 U22166 ( .C1(n19457), .C2(n19219), .A(n19190), .B(n19189), .ZN(
        P2_U3127) );
  NOR3_X2 U22167 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19570), .A3(
        n19224), .ZN(n19213) );
  OAI21_X1 U22168 ( .B1(n13232), .B2(n19213), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19191) );
  OAI21_X1 U22169 ( .B1(n19224), .B2(n19192), .A(n19191), .ZN(n19214) );
  AOI22_X1 U22170 ( .A1(n19214), .A2(n18867), .B1(n19399), .B2(n19213), .ZN(
        n19199) );
  INV_X1 U22171 ( .A(n13232), .ZN(n19195) );
  AOI221_X1 U22172 ( .B1(n19215), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19210), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19193), .ZN(n19194) );
  MUX2_X1 U22173 ( .A(n19195), .B(n19194), .S(n18921), .Z(n19196) );
  NOR2_X1 U22174 ( .A1(n19196), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19197) );
  OAI21_X1 U22175 ( .B1(n19197), .B2(n19213), .A(n19405), .ZN(n19216) );
  AOI22_X1 U22176 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19216), .B1(
        n19210), .B2(n19407), .ZN(n19198) );
  OAI211_X1 U22177 ( .C1(n19410), .C2(n19262), .A(n19199), .B(n19198), .ZN(
        P2_U3128) );
  AOI22_X1 U22178 ( .A1(n19214), .A2(n18879), .B1(n19411), .B2(n19213), .ZN(
        n19201) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19216), .B1(
        n19215), .B2(n19412), .ZN(n19200) );
  OAI211_X1 U22180 ( .C1(n19415), .C2(n19219), .A(n19201), .B(n19200), .ZN(
        P2_U3129) );
  AOI22_X1 U22181 ( .A1(n19214), .A2(n18883), .B1(n19416), .B2(n19213), .ZN(
        n19203) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19216), .B1(
        n19210), .B2(n19319), .ZN(n19202) );
  OAI211_X1 U22183 ( .C1(n19322), .C2(n19262), .A(n19203), .B(n19202), .ZN(
        P2_U3130) );
  AOI22_X1 U22184 ( .A1(n19214), .A2(n19422), .B1(n19421), .B2(n19213), .ZN(
        n19205) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19216), .B1(
        n19210), .B2(n19423), .ZN(n19204) );
  OAI211_X1 U22186 ( .C1(n19426), .C2(n19262), .A(n19205), .B(n19204), .ZN(
        P2_U3131) );
  AOI22_X1 U22187 ( .A1(n19214), .A2(n19428), .B1(n19427), .B2(n19213), .ZN(
        n19207) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19216), .B1(
        n19215), .B2(n19429), .ZN(n19206) );
  OAI211_X1 U22189 ( .C1(n19432), .C2(n19219), .A(n19207), .B(n19206), .ZN(
        P2_U3132) );
  AOI22_X1 U22190 ( .A1(n19214), .A2(n19434), .B1(n19433), .B2(n19213), .ZN(
        n19209) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19216), .B1(
        n19215), .B2(n19435), .ZN(n19208) );
  OAI211_X1 U22192 ( .C1(n19440), .C2(n19219), .A(n19209), .B(n19208), .ZN(
        P2_U3133) );
  AOI22_X1 U22193 ( .A1(n19214), .A2(n19442), .B1(n19441), .B2(n19213), .ZN(
        n19212) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19216), .B1(
        n19210), .B2(n19443), .ZN(n19211) );
  OAI211_X1 U22195 ( .C1(n19446), .C2(n19262), .A(n19212), .B(n19211), .ZN(
        P2_U3134) );
  AOI22_X1 U22196 ( .A1(n19214), .A2(n19449), .B1(n19447), .B2(n19213), .ZN(
        n19218) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19216), .B1(
        n19215), .B2(n19291), .ZN(n19217) );
  OAI211_X1 U22198 ( .C1(n19263), .C2(n19219), .A(n19218), .B(n19217), .ZN(
        P2_U3135) );
  INV_X1 U22199 ( .A(n19224), .ZN(n19220) );
  AND2_X1 U22200 ( .A1(n19221), .A2(n19220), .ZN(n19234) );
  NOR2_X1 U22201 ( .A1(n19234), .A2(n18921), .ZN(n19222) );
  AND2_X1 U22202 ( .A1(n19223), .A2(n19222), .ZN(n19230) );
  OR2_X1 U22203 ( .A1(n19570), .A2(n19224), .ZN(n19231) );
  INV_X1 U22204 ( .A(n19231), .ZN(n19225) );
  AOI21_X1 U22205 ( .B1(n19571), .B2(n19225), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19226) );
  INV_X1 U22206 ( .A(n18867), .ZN(n19302) );
  INV_X1 U22207 ( .A(n19399), .ZN(n19301) );
  INV_X1 U22208 ( .A(n19234), .ZN(n19256) );
  OAI22_X1 U22209 ( .A1(n19257), .A2(n19302), .B1(n19301), .B2(n19256), .ZN(
        n19227) );
  INV_X1 U22210 ( .A(n19227), .ZN(n19237) );
  INV_X1 U22211 ( .A(n19228), .ZN(n19402) );
  NAND2_X1 U22212 ( .A1(n19402), .A2(n19229), .ZN(n19232) );
  AOI21_X1 U22213 ( .B1(n19232), .B2(n19231), .A(n19230), .ZN(n19233) );
  OAI211_X1 U22214 ( .C1(n19234), .C2(n19571), .A(n19233), .B(n19405), .ZN(
        n19259) );
  NOR2_X2 U22215 ( .A1(n19297), .A2(n19235), .ZN(n19290) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19354), .ZN(n19236) );
  OAI211_X1 U22217 ( .C1(n19367), .C2(n19262), .A(n19237), .B(n19236), .ZN(
        P2_U3136) );
  INV_X1 U22218 ( .A(n18879), .ZN(n19312) );
  INV_X1 U22219 ( .A(n19411), .ZN(n19311) );
  OAI22_X1 U22220 ( .A1(n19257), .A2(n19312), .B1(n19311), .B2(n19256), .ZN(
        n19238) );
  INV_X1 U22221 ( .A(n19238), .ZN(n19240) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19412), .ZN(n19239) );
  OAI211_X1 U22223 ( .C1(n19415), .C2(n19262), .A(n19240), .B(n19239), .ZN(
        P2_U3137) );
  INV_X1 U22224 ( .A(n18883), .ZN(n19317) );
  INV_X1 U22225 ( .A(n19416), .ZN(n19316) );
  OAI22_X1 U22226 ( .A1(n19257), .A2(n19317), .B1(n19316), .B2(n19256), .ZN(
        n19241) );
  INV_X1 U22227 ( .A(n19241), .ZN(n19243) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19417), .ZN(n19242) );
  OAI211_X1 U22229 ( .C1(n19420), .C2(n19262), .A(n19243), .B(n19242), .ZN(
        P2_U3138) );
  INV_X1 U22230 ( .A(n19422), .ZN(n19324) );
  INV_X1 U22231 ( .A(n19421), .ZN(n19323) );
  OAI22_X1 U22232 ( .A1(n19257), .A2(n19324), .B1(n19323), .B2(n19256), .ZN(
        n19244) );
  INV_X1 U22233 ( .A(n19244), .ZN(n19246) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19374), .ZN(n19245) );
  OAI211_X1 U22235 ( .C1(n19377), .C2(n19262), .A(n19246), .B(n19245), .ZN(
        P2_U3139) );
  INV_X1 U22236 ( .A(n19428), .ZN(n19329) );
  INV_X1 U22237 ( .A(n19427), .ZN(n19328) );
  OAI22_X1 U22238 ( .A1(n19257), .A2(n19329), .B1(n19328), .B2(n19256), .ZN(
        n19247) );
  INV_X1 U22239 ( .A(n19247), .ZN(n19249) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19429), .ZN(n19248) );
  OAI211_X1 U22241 ( .C1(n19432), .C2(n19262), .A(n19249), .B(n19248), .ZN(
        P2_U3140) );
  INV_X1 U22242 ( .A(n19434), .ZN(n19334) );
  INV_X1 U22243 ( .A(n19433), .ZN(n19333) );
  OAI22_X1 U22244 ( .A1(n19257), .A2(n19334), .B1(n19333), .B2(n19256), .ZN(
        n19250) );
  INV_X1 U22245 ( .A(n19250), .ZN(n19252) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19435), .ZN(n19251) );
  OAI211_X1 U22247 ( .C1(n19440), .C2(n19262), .A(n19252), .B(n19251), .ZN(
        P2_U3141) );
  INV_X1 U22248 ( .A(n19442), .ZN(n19339) );
  INV_X1 U22249 ( .A(n19441), .ZN(n19338) );
  OAI22_X1 U22250 ( .A1(n19257), .A2(n19339), .B1(n19338), .B2(n19256), .ZN(
        n19253) );
  INV_X1 U22251 ( .A(n19253), .ZN(n19255) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19386), .ZN(n19254) );
  OAI211_X1 U22253 ( .C1(n19390), .C2(n19262), .A(n19255), .B(n19254), .ZN(
        P2_U3142) );
  INV_X1 U22254 ( .A(n19449), .ZN(n19345) );
  INV_X1 U22255 ( .A(n19447), .ZN(n19344) );
  OAI22_X1 U22256 ( .A1(n19257), .A2(n19345), .B1(n19344), .B2(n19256), .ZN(
        n19258) );
  INV_X1 U22257 ( .A(n19258), .ZN(n19261) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19259), .B1(
        n19290), .B2(n19291), .ZN(n19260) );
  OAI211_X1 U22259 ( .C1(n19263), .C2(n19262), .A(n19261), .B(n19260), .ZN(
        P2_U3143) );
  NOR2_X2 U22260 ( .A1(n19353), .A2(n19296), .ZN(n19348) );
  OAI21_X1 U22261 ( .B1(n19290), .B2(n19348), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19269) );
  NAND2_X1 U22262 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19264), .ZN(
        n19270) );
  NAND3_X1 U22263 ( .A1(n19570), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19306) );
  NOR2_X1 U22264 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19306), .ZN(
        n19288) );
  INV_X1 U22265 ( .A(n19288), .ZN(n19265) );
  AND2_X1 U22266 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19265), .ZN(n19266) );
  NAND2_X1 U22267 ( .A1(n19267), .A2(n19266), .ZN(n19272) );
  OAI211_X1 U22268 ( .C1(n19288), .C2(n19571), .A(n19272), .B(n19405), .ZN(
        n19268) );
  INV_X1 U22269 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n19275) );
  OAI21_X1 U22270 ( .B1(n19270), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n18921), 
        .ZN(n19271) );
  AND2_X1 U22271 ( .A1(n19272), .A2(n19271), .ZN(n19289) );
  AOI22_X1 U22272 ( .A1(n19289), .A2(n18867), .B1(n19399), .B2(n19288), .ZN(
        n19274) );
  AOI22_X1 U22273 ( .A1(n19290), .A2(n19407), .B1(n19348), .B2(n19354), .ZN(
        n19273) );
  OAI211_X1 U22274 ( .C1(n19295), .C2(n19275), .A(n19274), .B(n19273), .ZN(
        P2_U3144) );
  AOI22_X1 U22275 ( .A1(n19289), .A2(n18879), .B1(n19411), .B2(n19288), .ZN(
        n19277) );
  AOI22_X1 U22276 ( .A1(n19348), .A2(n19412), .B1(n19290), .B2(n19368), .ZN(
        n19276) );
  OAI211_X1 U22277 ( .C1(n19295), .C2(n10608), .A(n19277), .B(n19276), .ZN(
        P2_U3145) );
  AOI22_X1 U22278 ( .A1(n19289), .A2(n18883), .B1(n19416), .B2(n19288), .ZN(
        n19279) );
  AOI22_X1 U22279 ( .A1(n19290), .A2(n19319), .B1(n19348), .B2(n19417), .ZN(
        n19278) );
  OAI211_X1 U22280 ( .C1(n19295), .C2(n10636), .A(n19279), .B(n19278), .ZN(
        P2_U3146) );
  AOI22_X1 U22281 ( .A1(n19289), .A2(n19422), .B1(n19421), .B2(n19288), .ZN(
        n19281) );
  AOI22_X1 U22282 ( .A1(n19290), .A2(n19423), .B1(n19348), .B2(n19374), .ZN(
        n19280) );
  OAI211_X1 U22283 ( .C1(n19295), .C2(n12758), .A(n19281), .B(n19280), .ZN(
        P2_U3147) );
  AOI22_X1 U22284 ( .A1(n19289), .A2(n19428), .B1(n19427), .B2(n19288), .ZN(
        n19283) );
  AOI22_X1 U22285 ( .A1(n19348), .A2(n19429), .B1(n19290), .B2(n19378), .ZN(
        n19282) );
  OAI211_X1 U22286 ( .C1(n19295), .C2(n10682), .A(n19283), .B(n19282), .ZN(
        P2_U3148) );
  AOI22_X1 U22287 ( .A1(n19289), .A2(n19434), .B1(n19433), .B2(n19288), .ZN(
        n19285) );
  AOI22_X1 U22288 ( .A1(n19348), .A2(n19435), .B1(n19290), .B2(n19382), .ZN(
        n19284) );
  OAI211_X1 U22289 ( .C1(n19295), .C2(n13225), .A(n19285), .B(n19284), .ZN(
        P2_U3149) );
  AOI22_X1 U22290 ( .A1(n19289), .A2(n19442), .B1(n19441), .B2(n19288), .ZN(
        n19287) );
  AOI22_X1 U22291 ( .A1(n19290), .A2(n19443), .B1(n19348), .B2(n19386), .ZN(
        n19286) );
  OAI211_X1 U22292 ( .C1(n19295), .C2(n13262), .A(n19287), .B(n19286), .ZN(
        P2_U3150) );
  INV_X1 U22293 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19294) );
  AOI22_X1 U22294 ( .A1(n19289), .A2(n19449), .B1(n19447), .B2(n19288), .ZN(
        n19293) );
  AOI22_X1 U22295 ( .A1(n19348), .A2(n19291), .B1(n19290), .B2(n19451), .ZN(
        n19292) );
  OAI211_X1 U22296 ( .C1(n19295), .C2(n19294), .A(n19293), .B(n19292), .ZN(
        P2_U3151) );
  NOR2_X1 U22297 ( .A1(n19578), .A2(n19306), .ZN(n19357) );
  INV_X1 U22298 ( .A(n19357), .ZN(n19343) );
  AND2_X1 U22299 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19343), .ZN(n19298) );
  AND2_X1 U22300 ( .A1(n12753), .A2(n19298), .ZN(n19305) );
  INV_X1 U22301 ( .A(n19306), .ZN(n19299) );
  AOI21_X1 U22302 ( .B1(n19571), .B2(n19299), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19300) );
  OAI22_X1 U22303 ( .A1(n19346), .A2(n19302), .B1(n19301), .B2(n19343), .ZN(
        n19303) );
  INV_X1 U22304 ( .A(n19303), .ZN(n19310) );
  NAND2_X1 U22305 ( .A1(n19402), .A2(n19304), .ZN(n19307) );
  AOI21_X1 U22306 ( .B1(n19307), .B2(n19306), .A(n19305), .ZN(n19308) );
  OAI211_X1 U22307 ( .C1(n19357), .C2(n19571), .A(n19308), .B(n19405), .ZN(
        n19349) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19407), .ZN(n19309) );
  OAI211_X1 U22309 ( .C1(n19410), .C2(n19389), .A(n19310), .B(n19309), .ZN(
        P2_U3152) );
  OAI22_X1 U22310 ( .A1(n19346), .A2(n19312), .B1(n19311), .B2(n19343), .ZN(
        n19313) );
  INV_X1 U22311 ( .A(n19313), .ZN(n19315) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19368), .ZN(n19314) );
  OAI211_X1 U22313 ( .C1(n19371), .C2(n19389), .A(n19315), .B(n19314), .ZN(
        P2_U3153) );
  OAI22_X1 U22314 ( .A1(n19346), .A2(n19317), .B1(n19316), .B2(n19343), .ZN(
        n19318) );
  INV_X1 U22315 ( .A(n19318), .ZN(n19321) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19319), .ZN(n19320) );
  OAI211_X1 U22317 ( .C1(n19322), .C2(n19389), .A(n19321), .B(n19320), .ZN(
        P2_U3154) );
  OAI22_X1 U22318 ( .A1(n19346), .A2(n19324), .B1(n19323), .B2(n19343), .ZN(
        n19325) );
  INV_X1 U22319 ( .A(n19325), .ZN(n19327) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19423), .ZN(n19326) );
  OAI211_X1 U22321 ( .C1(n19426), .C2(n19389), .A(n19327), .B(n19326), .ZN(
        P2_U3155) );
  OAI22_X1 U22322 ( .A1(n19346), .A2(n19329), .B1(n19328), .B2(n19343), .ZN(
        n19330) );
  INV_X1 U22323 ( .A(n19330), .ZN(n19332) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19378), .ZN(n19331) );
  OAI211_X1 U22325 ( .C1(n19381), .C2(n19389), .A(n19332), .B(n19331), .ZN(
        P2_U3156) );
  OAI22_X1 U22326 ( .A1(n19346), .A2(n19334), .B1(n19333), .B2(n19343), .ZN(
        n19335) );
  INV_X1 U22327 ( .A(n19335), .ZN(n19337) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19382), .ZN(n19336) );
  OAI211_X1 U22329 ( .C1(n19385), .C2(n19389), .A(n19337), .B(n19336), .ZN(
        P2_U3157) );
  OAI22_X1 U22330 ( .A1(n19346), .A2(n19339), .B1(n19338), .B2(n19343), .ZN(
        n19340) );
  INV_X1 U22331 ( .A(n19340), .ZN(n19342) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19443), .ZN(n19341) );
  OAI211_X1 U22333 ( .C1(n19446), .C2(n19389), .A(n19342), .B(n19341), .ZN(
        P2_U3158) );
  OAI22_X1 U22334 ( .A1(n19346), .A2(n19345), .B1(n19344), .B2(n19343), .ZN(
        n19347) );
  INV_X1 U22335 ( .A(n19347), .ZN(n19351) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19451), .ZN(n19350) );
  OAI211_X1 U22337 ( .C1(n19457), .C2(n19389), .A(n19351), .B(n19350), .ZN(
        P2_U3159) );
  NAND3_X1 U22338 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19400) );
  NOR2_X1 U22339 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19400), .ZN(
        n19391) );
  AOI22_X1 U22340 ( .A1(n19354), .A2(n19452), .B1(n19391), .B2(n19399), .ZN(
        n19366) );
  OAI21_X1 U22341 ( .B1(n19452), .B2(n19392), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19356) );
  NAND2_X1 U22342 ( .A1(n19356), .A2(n19355), .ZN(n19364) );
  NOR2_X1 U22343 ( .A1(n19391), .A2(n19357), .ZN(n19363) );
  INV_X1 U22344 ( .A(n19363), .ZN(n19360) );
  INV_X1 U22345 ( .A(n19391), .ZN(n19358) );
  OAI211_X1 U22346 ( .C1(n13224), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19358), 
        .B(n19550), .ZN(n19359) );
  OAI211_X1 U22347 ( .C1(n19364), .C2(n19360), .A(n19405), .B(n19359), .ZN(
        n19394) );
  INV_X1 U22348 ( .A(n13224), .ZN(n19361) );
  OAI21_X1 U22349 ( .B1(n19361), .B2(n19391), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19362) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19394), .B1(
        n18867), .B2(n19393), .ZN(n19365) );
  OAI211_X1 U22351 ( .C1(n19367), .C2(n19389), .A(n19366), .B(n19365), .ZN(
        P2_U3160) );
  AOI22_X1 U22352 ( .A1(n19368), .A2(n19392), .B1(n19411), .B2(n19391), .ZN(
        n19370) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19394), .B1(
        n18879), .B2(n19393), .ZN(n19369) );
  OAI211_X1 U22354 ( .C1(n19371), .C2(n19439), .A(n19370), .B(n19369), .ZN(
        P2_U3161) );
  AOI22_X1 U22355 ( .A1(n19417), .A2(n19452), .B1(n19391), .B2(n19416), .ZN(
        n19373) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19394), .B1(
        n18883), .B2(n19393), .ZN(n19372) );
  OAI211_X1 U22357 ( .C1(n19420), .C2(n19389), .A(n19373), .B(n19372), .ZN(
        P2_U3162) );
  AOI22_X1 U22358 ( .A1(n19374), .A2(n19452), .B1(n19391), .B2(n19421), .ZN(
        n19376) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19394), .B1(
        n19422), .B2(n19393), .ZN(n19375) );
  OAI211_X1 U22360 ( .C1(n19377), .C2(n19389), .A(n19376), .B(n19375), .ZN(
        P2_U3163) );
  AOI22_X1 U22361 ( .A1(n19378), .A2(n19392), .B1(n19391), .B2(n19427), .ZN(
        n19380) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19394), .B1(
        n19428), .B2(n19393), .ZN(n19379) );
  OAI211_X1 U22363 ( .C1(n19381), .C2(n19439), .A(n19380), .B(n19379), .ZN(
        P2_U3164) );
  AOI22_X1 U22364 ( .A1(n19382), .A2(n19392), .B1(n19391), .B2(n19433), .ZN(
        n19384) );
  AOI22_X1 U22365 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19394), .B1(
        n19434), .B2(n19393), .ZN(n19383) );
  OAI211_X1 U22366 ( .C1(n19385), .C2(n19439), .A(n19384), .B(n19383), .ZN(
        P2_U3165) );
  AOI22_X1 U22367 ( .A1(n19386), .A2(n19452), .B1(n19391), .B2(n19441), .ZN(
        n19388) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19394), .B1(
        n19442), .B2(n19393), .ZN(n19387) );
  OAI211_X1 U22369 ( .C1(n19390), .C2(n19389), .A(n19388), .B(n19387), .ZN(
        P2_U3166) );
  AOI22_X1 U22370 ( .A1(n19451), .A2(n19392), .B1(n19391), .B2(n19447), .ZN(
        n19396) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19394), .B1(
        n19449), .B2(n19393), .ZN(n19395) );
  OAI211_X1 U22372 ( .C1(n19457), .C2(n19439), .A(n19396), .B(n19395), .ZN(
        P2_U3167) );
  INV_X1 U22373 ( .A(n19404), .ZN(n19397) );
  OAI21_X1 U22374 ( .B1(n19397), .B2(n19448), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19398) );
  OAI21_X1 U22375 ( .B1(n19400), .B2(n19550), .A(n19398), .ZN(n19450) );
  AOI22_X1 U22376 ( .A1(n19450), .A2(n18867), .B1(n19448), .B2(n19399), .ZN(
        n19409) );
  INV_X1 U22377 ( .A(n19400), .ZN(n19401) );
  AOI21_X1 U22378 ( .B1(n19402), .B2(n19544), .A(n19401), .ZN(n19403) );
  AOI211_X1 U22379 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19404), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19403), .ZN(n19406) );
  OAI21_X1 U22380 ( .B1(n19448), .B2(n19406), .A(n19405), .ZN(n19453) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19453), .B1(
        n19452), .B2(n19407), .ZN(n19408) );
  OAI211_X1 U22382 ( .C1(n19410), .C2(n19456), .A(n19409), .B(n19408), .ZN(
        P2_U3168) );
  AOI22_X1 U22383 ( .A1(n19450), .A2(n18879), .B1(n19448), .B2(n19411), .ZN(
        n19414) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19453), .B1(
        n19436), .B2(n19412), .ZN(n19413) );
  OAI211_X1 U22385 ( .C1(n19415), .C2(n19439), .A(n19414), .B(n19413), .ZN(
        P2_U3169) );
  AOI22_X1 U22386 ( .A1(n19450), .A2(n18883), .B1(n19448), .B2(n19416), .ZN(
        n19419) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19453), .B1(
        n19436), .B2(n19417), .ZN(n19418) );
  OAI211_X1 U22388 ( .C1(n19420), .C2(n19439), .A(n19419), .B(n19418), .ZN(
        P2_U3170) );
  AOI22_X1 U22389 ( .A1(n19450), .A2(n19422), .B1(n19448), .B2(n19421), .ZN(
        n19425) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19453), .B1(
        n19452), .B2(n19423), .ZN(n19424) );
  OAI211_X1 U22391 ( .C1(n19426), .C2(n19456), .A(n19425), .B(n19424), .ZN(
        P2_U3171) );
  AOI22_X1 U22392 ( .A1(n19450), .A2(n19428), .B1(n19448), .B2(n19427), .ZN(
        n19431) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19453), .B1(
        n19436), .B2(n19429), .ZN(n19430) );
  OAI211_X1 U22394 ( .C1(n19432), .C2(n19439), .A(n19431), .B(n19430), .ZN(
        P2_U3172) );
  AOI22_X1 U22395 ( .A1(n19450), .A2(n19434), .B1(n19448), .B2(n19433), .ZN(
        n19438) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19453), .B1(
        n19436), .B2(n19435), .ZN(n19437) );
  OAI211_X1 U22397 ( .C1(n19440), .C2(n19439), .A(n19438), .B(n19437), .ZN(
        P2_U3173) );
  AOI22_X1 U22398 ( .A1(n19450), .A2(n19442), .B1(n19448), .B2(n19441), .ZN(
        n19445) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19453), .B1(
        n19452), .B2(n19443), .ZN(n19444) );
  OAI211_X1 U22400 ( .C1(n19446), .C2(n19456), .A(n19445), .B(n19444), .ZN(
        P2_U3174) );
  AOI22_X1 U22401 ( .A1(n19450), .A2(n19449), .B1(n19448), .B2(n19447), .ZN(
        n19455) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19453), .B1(
        n19452), .B2(n19451), .ZN(n19454) );
  OAI211_X1 U22403 ( .C1(n19457), .C2(n19456), .A(n19455), .B(n19454), .ZN(
        P2_U3175) );
  OAI21_X1 U22404 ( .B1(n19595), .B2(n19459), .A(n19458), .ZN(n19463) );
  NAND2_X1 U22405 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19595), .ZN(n19460) );
  AOI21_X1 U22406 ( .B1(n19461), .B2(n19464), .A(n19460), .ZN(n19462) );
  AOI21_X1 U22407 ( .B1(n19464), .B2(n19463), .A(n19462), .ZN(n19466) );
  NAND2_X1 U22408 ( .A1(n19466), .A2(n19465), .ZN(P2_U3177) );
  AND2_X1 U22409 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19467), .ZN(
        P2_U3179) );
  AND2_X1 U22410 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19467), .ZN(
        P2_U3180) );
  AND2_X1 U22411 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19467), .ZN(
        P2_U3181) );
  AND2_X1 U22412 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19467), .ZN(
        P2_U3182) );
  AND2_X1 U22413 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19467), .ZN(
        P2_U3183) );
  AND2_X1 U22414 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19467), .ZN(
        P2_U3184) );
  AND2_X1 U22415 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19467), .ZN(
        P2_U3185) );
  AND2_X1 U22416 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19467), .ZN(
        P2_U3186) );
  AND2_X1 U22417 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19467), .ZN(
        P2_U3187) );
  AND2_X1 U22418 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19467), .ZN(
        P2_U3188) );
  INV_X1 U22419 ( .A(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20602) );
  NOR2_X1 U22420 ( .A1(n20602), .A2(n19542), .ZN(P2_U3189) );
  AND2_X1 U22421 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19467), .ZN(
        P2_U3190) );
  AND2_X1 U22422 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19467), .ZN(
        P2_U3191) );
  AND2_X1 U22423 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19467), .ZN(
        P2_U3192) );
  AND2_X1 U22424 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19467), .ZN(
        P2_U3193) );
  AND2_X1 U22425 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19467), .ZN(
        P2_U3194) );
  AND2_X1 U22426 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19467), .ZN(
        P2_U3195) );
  AND2_X1 U22427 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19467), .ZN(
        P2_U3196) );
  AND2_X1 U22428 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19467), .ZN(
        P2_U3197) );
  AND2_X1 U22429 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19467), .ZN(
        P2_U3198) );
  AND2_X1 U22430 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19467), .ZN(
        P2_U3199) );
  AND2_X1 U22431 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19467), .ZN(
        P2_U3200) );
  AND2_X1 U22432 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19467), .ZN(P2_U3201) );
  AND2_X1 U22433 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19467), .ZN(P2_U3202) );
  AND2_X1 U22434 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19467), .ZN(P2_U3203) );
  AND2_X1 U22435 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19467), .ZN(P2_U3204) );
  AND2_X1 U22436 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19467), .ZN(P2_U3205) );
  AND2_X1 U22437 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19467), .ZN(P2_U3206) );
  AND2_X1 U22438 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19467), .ZN(P2_U3207) );
  AND2_X1 U22439 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19467), .ZN(P2_U3208) );
  NAND2_X1 U22440 ( .A1(n19595), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19479) );
  NAND3_X1 U22441 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19479), .ZN(n19470) );
  AOI211_X1 U22442 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20407), .A(
        n19468), .B(n19606), .ZN(n19469) );
  NOR2_X1 U22443 ( .A1(n20413), .A2(n19473), .ZN(n19484) );
  AOI211_X1 U22444 ( .C1(n19485), .C2(n19470), .A(n19469), .B(n19484), .ZN(
        n19471) );
  INV_X1 U22445 ( .A(n19471), .ZN(P2_U3209) );
  INV_X1 U22446 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19472) );
  AOI21_X1 U22447 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20407), .A(n19485), 
        .ZN(n19477) );
  NOR2_X1 U22448 ( .A1(n19472), .A2(n19477), .ZN(n19474) );
  AOI21_X1 U22449 ( .B1(n19474), .B2(n19473), .A(n19591), .ZN(n19475) );
  OAI211_X1 U22450 ( .C1(n20407), .C2(n19476), .A(n19475), .B(n19479), .ZN(
        P2_U3210) );
  AOI21_X1 U22451 ( .B1(n19478), .B2(n19595), .A(n19477), .ZN(n19483) );
  OAI22_X1 U22452 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19480), .B1(NA), 
        .B2(n19479), .ZN(n19481) );
  OAI211_X1 U22453 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19481), .ZN(n19482) );
  OAI21_X1 U22454 ( .B1(n19484), .B2(n19483), .A(n19482), .ZN(P2_U3211) );
  OAI222_X1 U22455 ( .A1(n19534), .A2(n19488), .B1(n19487), .B2(n19606), .C1(
        n19486), .C2(n19531), .ZN(P2_U3212) );
  OAI222_X1 U22456 ( .A1(n19534), .A2(n19489), .B1(n20527), .B2(n19606), .C1(
        n19488), .C2(n19531), .ZN(P2_U3213) );
  OAI222_X1 U22457 ( .A1(n19534), .A2(n19491), .B1(n19490), .B2(n19606), .C1(
        n19489), .C2(n19531), .ZN(P2_U3214) );
  INV_X1 U22458 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19493) );
  OAI222_X1 U22459 ( .A1(n19534), .A2(n19493), .B1(n19492), .B2(n19606), .C1(
        n19491), .C2(n19531), .ZN(P2_U3215) );
  OAI222_X1 U22460 ( .A1(n19534), .A2(n19495), .B1(n19494), .B2(n19606), .C1(
        n19493), .C2(n19531), .ZN(P2_U3216) );
  OAI222_X1 U22461 ( .A1(n19534), .A2(n19497), .B1(n19496), .B2(n19606), .C1(
        n19495), .C2(n19531), .ZN(P2_U3217) );
  INV_X1 U22462 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19498) );
  OAI222_X1 U22463 ( .A1(n19534), .A2(n19498), .B1(n20544), .B2(n19606), .C1(
        n19497), .C2(n19531), .ZN(P2_U3218) );
  OAI222_X1 U22464 ( .A1(n19534), .A2(n19499), .B1(n20555), .B2(n19606), .C1(
        n19498), .C2(n19531), .ZN(P2_U3219) );
  OAI222_X1 U22465 ( .A1(n19534), .A2(n12029), .B1(n19500), .B2(n19606), .C1(
        n19499), .C2(n19531), .ZN(P2_U3220) );
  OAI222_X1 U22466 ( .A1(n19534), .A2(n19502), .B1(n19501), .B2(n19606), .C1(
        n12029), .C2(n19531), .ZN(P2_U3221) );
  OAI222_X1 U22467 ( .A1(n19534), .A2(n12062), .B1(n19503), .B2(n19606), .C1(
        n19502), .C2(n19531), .ZN(P2_U3222) );
  OAI222_X1 U22468 ( .A1(n19534), .A2(n12067), .B1(n19504), .B2(n19606), .C1(
        n12062), .C2(n19531), .ZN(P2_U3223) );
  OAI222_X1 U22469 ( .A1(n19534), .A2(n19506), .B1(n19505), .B2(n19606), .C1(
        n12067), .C2(n19531), .ZN(P2_U3224) );
  OAI222_X1 U22470 ( .A1(n19534), .A2(n12074), .B1(n19507), .B2(n19606), .C1(
        n19506), .C2(n19531), .ZN(P2_U3225) );
  OAI222_X1 U22471 ( .A1(n19534), .A2(n12078), .B1(n19508), .B2(n19606), .C1(
        n12074), .C2(n19531), .ZN(P2_U3226) );
  OAI222_X1 U22472 ( .A1(n19534), .A2(n19510), .B1(n19509), .B2(n19606), .C1(
        n12078), .C2(n19531), .ZN(P2_U3227) );
  INV_X1 U22473 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19512) );
  OAI222_X1 U22474 ( .A1(n19534), .A2(n19512), .B1(n19511), .B2(n19606), .C1(
        n19510), .C2(n19531), .ZN(P2_U3228) );
  OAI222_X1 U22475 ( .A1(n19534), .A2(n12088), .B1(n19513), .B2(n19606), .C1(
        n19512), .C2(n19531), .ZN(P2_U3229) );
  OAI222_X1 U22476 ( .A1(n19534), .A2(n19515), .B1(n19514), .B2(n19606), .C1(
        n12088), .C2(n19531), .ZN(P2_U3230) );
  OAI222_X1 U22477 ( .A1(n19534), .A2(n19517), .B1(n19516), .B2(n19606), .C1(
        n19515), .C2(n19531), .ZN(P2_U3231) );
  OAI222_X1 U22478 ( .A1(n19534), .A2(n12099), .B1(n19518), .B2(n19606), .C1(
        n19517), .C2(n19531), .ZN(P2_U3232) );
  OAI222_X1 U22479 ( .A1(n19534), .A2(n12104), .B1(n19519), .B2(n19606), .C1(
        n12099), .C2(n19531), .ZN(P2_U3233) );
  OAI222_X1 U22480 ( .A1(n19534), .A2(n12108), .B1(n19520), .B2(n19606), .C1(
        n12104), .C2(n19531), .ZN(P2_U3234) );
  INV_X1 U22481 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19522) );
  OAI222_X1 U22482 ( .A1(n19534), .A2(n19522), .B1(n19521), .B2(n19606), .C1(
        n12108), .C2(n19531), .ZN(P2_U3235) );
  OAI222_X1 U22483 ( .A1(n19534), .A2(n19524), .B1(n19523), .B2(n19606), .C1(
        n19522), .C2(n19531), .ZN(P2_U3236) );
  INV_X1 U22484 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19527) );
  OAI222_X1 U22485 ( .A1(n19534), .A2(n19527), .B1(n19525), .B2(n19606), .C1(
        n19524), .C2(n19531), .ZN(P2_U3237) );
  OAI222_X1 U22486 ( .A1(n19531), .A2(n19527), .B1(n19526), .B2(n19606), .C1(
        n12122), .C2(n19534), .ZN(P2_U3238) );
  OAI222_X1 U22487 ( .A1(n19534), .A2(n19529), .B1(n19528), .B2(n19606), .C1(
        n12122), .C2(n19531), .ZN(P2_U3239) );
  OAI222_X1 U22488 ( .A1(n19534), .A2(n14436), .B1(n19530), .B2(n19606), .C1(
        n19529), .C2(n19531), .ZN(P2_U3240) );
  INV_X1 U22489 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19533) );
  OAI222_X1 U22490 ( .A1(n19534), .A2(n19533), .B1(n19532), .B2(n19606), .C1(
        n14436), .C2(n19531), .ZN(P2_U3241) );
  OAI22_X1 U22491 ( .A1(n19607), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19606), .ZN(n19535) );
  INV_X1 U22492 ( .A(n19535), .ZN(P2_U3585) );
  OAI22_X1 U22493 ( .A1(n19607), .A2(P2_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P2_BE_N_REG_2__SCAN_IN), .B2(n19606), .ZN(n19536) );
  INV_X1 U22494 ( .A(n19536), .ZN(P2_U3586) );
  OAI22_X1 U22495 ( .A1(n19607), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19606), .ZN(n19537) );
  INV_X1 U22496 ( .A(n19537), .ZN(P2_U3587) );
  OAI22_X1 U22497 ( .A1(n19607), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19606), .ZN(n19538) );
  INV_X1 U22498 ( .A(n19538), .ZN(P2_U3588) );
  OAI21_X1 U22499 ( .B1(n19542), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19540), 
        .ZN(n19539) );
  INV_X1 U22500 ( .A(n19539), .ZN(P2_U3591) );
  OAI21_X1 U22501 ( .B1(n19542), .B2(n19541), .A(n19540), .ZN(P2_U3592) );
  NAND3_X1 U22502 ( .A1(n19544), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19543), 
        .ZN(n19545) );
  AND2_X1 U22503 ( .A1(n19545), .A2(n19561), .ZN(n19557) );
  NOR2_X1 U22504 ( .A1(n19546), .A2(n19571), .ZN(n19547) );
  AOI21_X1 U22505 ( .B1(n19557), .B2(n19548), .A(n19547), .ZN(n19549) );
  OAI21_X1 U22506 ( .B1(n19551), .B2(n19550), .A(n19549), .ZN(n19552) );
  INV_X1 U22507 ( .A(n19552), .ZN(n19553) );
  AOI22_X1 U22508 ( .A1(n19579), .A2(n19554), .B1(n19553), .B2(n19576), .ZN(
        P2_U3602) );
  OAI21_X1 U22509 ( .B1(n19563), .B2(n19566), .A(n19555), .ZN(n19556) );
  AOI22_X1 U22510 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19558), .B1(n19557), 
        .B2(n19556), .ZN(n19559) );
  AOI22_X1 U22511 ( .A1(n19579), .A2(n19560), .B1(n19559), .B2(n19576), .ZN(
        P2_U3603) );
  INV_X1 U22512 ( .A(n19561), .ZN(n19572) );
  OR3_X1 U22513 ( .A1(n19563), .A2(n19572), .A3(n19562), .ZN(n19564) );
  OAI21_X1 U22514 ( .B1(n19566), .B2(n19565), .A(n19564), .ZN(n19567) );
  AOI21_X1 U22515 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19568), .A(n19567), 
        .ZN(n19569) );
  AOI22_X1 U22516 ( .A1(n19579), .A2(n19570), .B1(n19569), .B2(n19576), .ZN(
        P2_U3604) );
  OAI22_X1 U22517 ( .A1(n19573), .A2(n19572), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19571), .ZN(n19574) );
  AOI21_X1 U22518 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19575), .A(n19574), 
        .ZN(n19577) );
  AOI22_X1 U22519 ( .A1(n19579), .A2(n19578), .B1(n19577), .B2(n19576), .ZN(
        P2_U3605) );
  INV_X1 U22520 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19580) );
  AOI22_X1 U22521 ( .A1(n19606), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19580), 
        .B2(n19607), .ZN(P2_U3608) );
  INV_X1 U22522 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19590) );
  INV_X1 U22523 ( .A(n19581), .ZN(n19589) );
  AOI22_X1 U22524 ( .A1(n19585), .A2(n19584), .B1(n19583), .B2(n19582), .ZN(
        n19588) );
  NOR2_X1 U22525 ( .A1(n19589), .A2(n19586), .ZN(n19587) );
  AOI22_X1 U22526 ( .A1(n19590), .A2(n19589), .B1(n19588), .B2(n19587), .ZN(
        P2_U3609) );
  OAI21_X1 U22527 ( .B1(n19592), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19591), 
        .ZN(n19593) );
  NAND3_X1 U22528 ( .A1(n19594), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19593), 
        .ZN(n19598) );
  OAI22_X1 U22529 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19596), .B1(n19595), 
        .B2(n18921), .ZN(n19597) );
  NAND2_X1 U22530 ( .A1(n19598), .A2(n19597), .ZN(n19605) );
  AOI21_X1 U22531 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19599), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19601) );
  AOI211_X1 U22532 ( .C1(n19603), .C2(n19602), .A(n19601), .B(n19600), .ZN(
        n19604) );
  MUX2_X1 U22533 ( .A(n19605), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19604), 
        .Z(P2_U3610) );
  OAI22_X1 U22534 ( .A1(n19607), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19606), .ZN(n19608) );
  INV_X1 U22535 ( .A(n19608), .ZN(P2_U3611) );
  AOI21_X1 U22536 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20422), .A(n20419), 
        .ZN(n19615) );
  INV_X1 U22537 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19609) );
  AOI21_X1 U22538 ( .B1(n19615), .B2(n19609), .A(n20487), .ZN(P1_U2802) );
  OAI21_X1 U22539 ( .B1(n19611), .B2(n19610), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19612) );
  OAI21_X1 U22540 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19613), .A(n19612), 
        .ZN(P1_U2803) );
  NOR2_X1 U22541 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19616) );
  OAI21_X1 U22542 ( .B1(n19616), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20502), .ZN(
        n19614) );
  OAI21_X1 U22543 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20502), .A(n19614), 
        .ZN(P1_U2804) );
  NOR2_X1 U22544 ( .A1(n20487), .A2(n19615), .ZN(n20475) );
  OAI21_X1 U22545 ( .B1(BS16), .B2(n19616), .A(n20475), .ZN(n20473) );
  OAI21_X1 U22546 ( .B1(n20475), .B2(n20291), .A(n20473), .ZN(P1_U2805) );
  OAI21_X1 U22547 ( .B1(n19618), .B2(n19617), .A(n19804), .ZN(P1_U2806) );
  NOR4_X1 U22548 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19622) );
  NOR4_X1 U22549 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19621) );
  NOR4_X1 U22550 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19620) );
  NOR4_X1 U22551 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19619) );
  NAND4_X1 U22552 ( .A1(n19622), .A2(n19621), .A3(n19620), .A4(n19619), .ZN(
        n19628) );
  NOR4_X1 U22553 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19626) );
  AOI211_X1 U22554 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_10__SCAN_IN), .B(
        P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n19625) );
  NOR4_X1 U22555 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19624) );
  NOR4_X1 U22556 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19623) );
  NAND4_X1 U22557 ( .A1(n19626), .A2(n19625), .A3(n19624), .A4(n19623), .ZN(
        n19627) );
  NOR2_X1 U22558 ( .A1(n19628), .A2(n19627), .ZN(n20480) );
  INV_X1 U22559 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19630) );
  NOR3_X1 U22560 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19631) );
  OAI21_X1 U22561 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19631), .A(n20480), .ZN(
        n19629) );
  OAI21_X1 U22562 ( .B1(n20480), .B2(n19630), .A(n19629), .ZN(P1_U2807) );
  INV_X1 U22563 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20474) );
  AOI21_X1 U22564 ( .B1(n20476), .B2(n20474), .A(n19631), .ZN(n19633) );
  INV_X1 U22565 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19632) );
  INV_X1 U22566 ( .A(n20480), .ZN(n20483) );
  AOI22_X1 U22567 ( .A1(n20480), .A2(n19633), .B1(n19632), .B2(n20483), .ZN(
        P1_U2808) );
  AOI22_X1 U22568 ( .A1(n19634), .A2(n20435), .B1(n19708), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19645) );
  OAI22_X1 U22569 ( .A1(n19636), .A2(n19686), .B1(n19673), .B2(n19635), .ZN(
        n19637) );
  AOI211_X1 U22570 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n19638), .A(n19650), .B(
        n19637), .ZN(n19644) );
  INV_X1 U22571 ( .A(n19639), .ZN(n19642) );
  AOI22_X1 U22572 ( .A1(n19642), .A2(n19667), .B1(n19641), .B2(n19640), .ZN(
        n19643) );
  NAND3_X1 U22573 ( .A1(n19645), .A2(n19644), .A3(n19643), .ZN(P1_U2831) );
  NAND2_X1 U22574 ( .A1(n19709), .A2(n19677), .ZN(n19684) );
  NAND2_X1 U22575 ( .A1(n19646), .A2(n19684), .ZN(n19699) );
  AOI21_X1 U22576 ( .B1(n19709), .B2(n19648), .A(n19699), .ZN(n19664) );
  NAND2_X1 U22577 ( .A1(n19647), .A2(n19667), .ZN(n19657) );
  NOR4_X1 U22578 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19678), .A3(n19677), .A4(
        n19648), .ZN(n19649) );
  AOI211_X1 U22579 ( .C1(n19710), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19650), .B(n19649), .ZN(n19656) );
  OAI22_X1 U22580 ( .A1(n19695), .A2(n19652), .B1(n19651), .B2(n19713), .ZN(
        n19653) );
  AOI21_X1 U22581 ( .B1(n19707), .B2(n19654), .A(n19653), .ZN(n19655) );
  AND3_X1 U22582 ( .A1(n19657), .A2(n19656), .A3(n19655), .ZN(n19658) );
  OAI21_X1 U22583 ( .B1(n19664), .B2(n20433), .A(n19658), .ZN(P1_U2833) );
  INV_X1 U22584 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19724) );
  NAND2_X1 U22585 ( .A1(n19710), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19659) );
  OAI211_X1 U22586 ( .C1(n19695), .C2(n19724), .A(n19659), .B(n19693), .ZN(
        n19660) );
  INV_X1 U22587 ( .A(n19660), .ZN(n19661) );
  OAI21_X1 U22588 ( .B1(n19673), .B2(n19662), .A(n19661), .ZN(n19666) );
  INV_X1 U22589 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20430) );
  INV_X1 U22590 ( .A(n19699), .ZN(n19663) );
  NAND2_X1 U22591 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19663), .ZN(n19679) );
  AOI21_X1 U22592 ( .B1(n20430), .B2(n19679), .A(n19664), .ZN(n19665) );
  AOI211_X1 U22593 ( .C1(n19667), .C2(n19722), .A(n19666), .B(n19665), .ZN(
        n19668) );
  OAI21_X1 U22594 ( .B1(n19669), .B2(n19713), .A(n19668), .ZN(P1_U2834) );
  OAI21_X1 U22595 ( .B1(n19686), .B2(n19670), .A(n19693), .ZN(n19671) );
  AOI21_X1 U22596 ( .B1(n19708), .B2(P1_EBX_REG_5__SCAN_IN), .A(n19671), .ZN(
        n19672) );
  OAI21_X1 U22597 ( .B1(n19674), .B2(n19673), .A(n19672), .ZN(n19675) );
  AOI21_X1 U22598 ( .B1(n19676), .B2(n19698), .A(n19675), .ZN(n19682) );
  NOR2_X1 U22599 ( .A1(n19678), .A2(n19677), .ZN(n19680) );
  OAI21_X1 U22600 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n19680), .A(n19679), .ZN(
        n19681) );
  OAI211_X1 U22601 ( .C1(n19713), .C2(n19683), .A(n19682), .B(n19681), .ZN(
        P1_U2835) );
  NAND3_X1 U22602 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19685) );
  OAI22_X1 U22603 ( .A1(n19687), .A2(n19686), .B1(n19685), .B2(n19684), .ZN(
        n19688) );
  INV_X1 U22604 ( .A(n19688), .ZN(n19703) );
  INV_X1 U22605 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19727) );
  NAND2_X1 U22606 ( .A1(n19690), .A2(n19689), .ZN(n19691) );
  AND2_X1 U22607 ( .A1(n19692), .A2(n19691), .ZN(n19814) );
  NAND2_X1 U22608 ( .A1(n19707), .A2(n19814), .ZN(n19694) );
  OAI211_X1 U22609 ( .C1(n19727), .C2(n19695), .A(n19694), .B(n19693), .ZN(
        n19696) );
  AOI21_X1 U22610 ( .B1(n19697), .B2(n19717), .A(n19696), .ZN(n19702) );
  NAND2_X1 U22611 ( .A1(n19793), .A2(n19698), .ZN(n19701) );
  NAND2_X1 U22612 ( .A1(n19699), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n19700) );
  AND4_X1 U22613 ( .A1(n19703), .A2(n19702), .A3(n19701), .A4(n19700), .ZN(
        n19704) );
  OAI21_X1 U22614 ( .B1(n19798), .B2(n19713), .A(n19704), .ZN(P1_U2836) );
  AOI21_X1 U22615 ( .B1(n19709), .B2(n20476), .A(n19705), .ZN(n19720) );
  INV_X1 U22616 ( .A(n19835), .ZN(n19706) );
  AOI22_X1 U22617 ( .A1(n19708), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n19707), .B2(
        n19706), .ZN(n19719) );
  INV_X1 U22618 ( .A(n20230), .ZN(n19860) );
  NAND3_X1 U22619 ( .A1(n19709), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n12916), 
        .ZN(n19712) );
  NAND2_X1 U22620 ( .A1(n19710), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19711) );
  OAI211_X1 U22621 ( .C1(n19809), .C2(n19713), .A(n19712), .B(n19711), .ZN(
        n19716) );
  NOR2_X1 U22622 ( .A1(n19805), .A2(n19714), .ZN(n19715) );
  AOI211_X1 U22623 ( .C1(n19717), .C2(n19860), .A(n19716), .B(n19715), .ZN(
        n19718) );
  OAI211_X1 U22624 ( .C1(n19720), .C2(n12916), .A(n19719), .B(n19718), .ZN(
        P1_U2838) );
  AOI22_X1 U22625 ( .A1(n19722), .A2(n11912), .B1(n19725), .B2(n19721), .ZN(
        n19723) );
  OAI21_X1 U22626 ( .B1(n19728), .B2(n19724), .A(n19723), .ZN(P1_U2866) );
  AOI22_X1 U22627 ( .A1(n19793), .A2(n11912), .B1(n19725), .B2(n19814), .ZN(
        n19726) );
  OAI21_X1 U22628 ( .B1(n19728), .B2(n19727), .A(n19726), .ZN(P1_U2868) );
  AOI22_X1 U22629 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19732), .B1(n19758), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19729) );
  OAI21_X1 U22630 ( .B1(n19731), .B2(n19730), .A(n19729), .ZN(P1_U2921) );
  INV_X1 U22631 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U22632 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19733) );
  OAI21_X1 U22633 ( .B1(n19734), .B2(n19761), .A(n19733), .ZN(P1_U2922) );
  INV_X1 U22634 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19736) );
  AOI22_X1 U22635 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19735) );
  OAI21_X1 U22636 ( .B1(n19736), .B2(n19761), .A(n19735), .ZN(P1_U2923) );
  INV_X1 U22637 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19738) );
  AOI22_X1 U22638 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19737) );
  OAI21_X1 U22639 ( .B1(n19738), .B2(n19761), .A(n19737), .ZN(P1_U2924) );
  INV_X1 U22640 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19740) );
  AOI22_X1 U22641 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19739) );
  OAI21_X1 U22642 ( .B1(n19740), .B2(n19761), .A(n19739), .ZN(P1_U2925) );
  AOI22_X1 U22643 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19741) );
  OAI21_X1 U22644 ( .B1(n20639), .B2(n19761), .A(n19741), .ZN(P1_U2926) );
  INV_X1 U22645 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U22646 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19742) );
  OAI21_X1 U22647 ( .B1(n19743), .B2(n19761), .A(n19742), .ZN(P1_U2927) );
  AOI22_X1 U22648 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19744) );
  OAI21_X1 U22649 ( .B1(n13081), .B2(n19761), .A(n19744), .ZN(P1_U2928) );
  AOI22_X1 U22650 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19745) );
  OAI21_X1 U22651 ( .B1(n11393), .B2(n19761), .A(n19745), .ZN(P1_U2929) );
  AOI22_X1 U22652 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19746) );
  OAI21_X1 U22653 ( .B1(n19747), .B2(n19761), .A(n19746), .ZN(P1_U2930) );
  AOI22_X1 U22654 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19748) );
  OAI21_X1 U22655 ( .B1(n19749), .B2(n19761), .A(n19748), .ZN(P1_U2931) );
  AOI22_X1 U22656 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19750) );
  OAI21_X1 U22657 ( .B1(n19751), .B2(n19761), .A(n19750), .ZN(P1_U2932) );
  AOI22_X1 U22658 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19752) );
  OAI21_X1 U22659 ( .B1(n19753), .B2(n19761), .A(n19752), .ZN(P1_U2933) );
  AOI22_X1 U22660 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19754) );
  OAI21_X1 U22661 ( .B1(n19755), .B2(n19761), .A(n19754), .ZN(P1_U2934) );
  AOI22_X1 U22662 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19756) );
  OAI21_X1 U22663 ( .B1(n19757), .B2(n19761), .A(n19756), .ZN(P1_U2935) );
  AOI22_X1 U22664 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19759), .B1(n19758), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19760) );
  OAI21_X1 U22665 ( .B1(n19762), .B2(n19761), .A(n19760), .ZN(P1_U2936) );
  AOI22_X1 U22666 ( .A1(n19786), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19767), .ZN(n19764) );
  NAND2_X1 U22667 ( .A1(n19773), .A2(n19763), .ZN(n19775) );
  NAND2_X1 U22668 ( .A1(n19764), .A2(n19775), .ZN(P1_U2945) );
  AOI22_X1 U22669 ( .A1(n19786), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n19785), .ZN(n19766) );
  NAND2_X1 U22670 ( .A1(n19773), .A2(n19765), .ZN(n19777) );
  NAND2_X1 U22671 ( .A1(n19766), .A2(n19777), .ZN(P1_U2946) );
  AOI22_X1 U22672 ( .A1(n19786), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n19767), .ZN(n19769) );
  NAND2_X1 U22673 ( .A1(n19773), .A2(n19768), .ZN(n19779) );
  NAND2_X1 U22674 ( .A1(n19769), .A2(n19779), .ZN(P1_U2948) );
  AOI22_X1 U22675 ( .A1(n19786), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19785), .ZN(n19771) );
  NAND2_X1 U22676 ( .A1(n19773), .A2(n19770), .ZN(n19781) );
  NAND2_X1 U22677 ( .A1(n19771), .A2(n19781), .ZN(P1_U2949) );
  AOI22_X1 U22678 ( .A1(n19786), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19785), .ZN(n19774) );
  NAND2_X1 U22679 ( .A1(n19773), .A2(n19772), .ZN(n19787) );
  NAND2_X1 U22680 ( .A1(n19774), .A2(n19787), .ZN(P1_U2951) );
  AOI22_X1 U22681 ( .A1(n19786), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19785), .ZN(n19776) );
  NAND2_X1 U22682 ( .A1(n19776), .A2(n19775), .ZN(P1_U2960) );
  AOI22_X1 U22683 ( .A1(n19786), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19767), .ZN(n19778) );
  NAND2_X1 U22684 ( .A1(n19778), .A2(n19777), .ZN(P1_U2961) );
  AOI22_X1 U22685 ( .A1(n19786), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19767), .ZN(n19780) );
  NAND2_X1 U22686 ( .A1(n19780), .A2(n19779), .ZN(P1_U2963) );
  AOI22_X1 U22687 ( .A1(n19786), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19785), .ZN(n19782) );
  NAND2_X1 U22688 ( .A1(n19782), .A2(n19781), .ZN(P1_U2964) );
  AOI22_X1 U22689 ( .A1(n19786), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19767), .ZN(n19784) );
  NAND2_X1 U22690 ( .A1(n19784), .A2(n19783), .ZN(P1_U2965) );
  AOI22_X1 U22691 ( .A1(n19786), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19785), .ZN(n19788) );
  NAND2_X1 U22692 ( .A1(n19788), .A2(n19787), .ZN(P1_U2966) );
  AOI22_X1 U22693 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19797) );
  OAI21_X1 U22694 ( .B1(n19791), .B2(n19790), .A(n19789), .ZN(n19792) );
  INV_X1 U22695 ( .A(n19792), .ZN(n19817) );
  AOI22_X1 U22696 ( .A1(n19817), .A2(n19795), .B1(n19794), .B2(n19793), .ZN(
        n19796) );
  OAI211_X1 U22697 ( .C1(n19810), .C2(n19798), .A(n19797), .B(n19796), .ZN(
        P1_U2995) );
  AOI22_X1 U22698 ( .A1(n19799), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12502), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n19808) );
  OR2_X1 U22699 ( .A1(n19801), .A2(n19800), .ZN(n19802) );
  NAND2_X1 U22700 ( .A1(n19803), .A2(n19802), .ZN(n19837) );
  OAI22_X1 U22701 ( .A1(n19805), .A2(n19851), .B1(n19837), .B2(n19804), .ZN(
        n19806) );
  INV_X1 U22702 ( .A(n19806), .ZN(n19807) );
  OAI211_X1 U22703 ( .C1(n19810), .C2(n19809), .A(n19808), .B(n19807), .ZN(
        P1_U2997) );
  NOR2_X1 U22704 ( .A1(n19812), .A2(n19811), .ZN(n19830) );
  NOR2_X1 U22705 ( .A1(n19830), .A2(n19813), .ZN(n19827) );
  AOI22_X1 U22706 ( .A1(n19814), .A2(n19825), .B1(n12502), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n19819) );
  AOI211_X1 U22707 ( .C1(n19820), .C2(n19828), .A(n19815), .B(n19829), .ZN(
        n19816) );
  AOI21_X1 U22708 ( .B1(n19817), .B2(n19823), .A(n19816), .ZN(n19818) );
  OAI211_X1 U22709 ( .C1(n19827), .C2(n19820), .A(n19819), .B(n19818), .ZN(
        P1_U3027) );
  INV_X1 U22710 ( .A(n19821), .ZN(n19822) );
  AOI222_X1 U22711 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n12502), .B1(n19825), 
        .B2(n19824), .C1(n19823), .C2(n19822), .ZN(n19826) );
  OAI221_X1 U22712 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19829), .C1(
        n19828), .C2(n19827), .A(n19826), .ZN(P1_U3028) );
  INV_X1 U22713 ( .A(n19830), .ZN(n19833) );
  NAND4_X1 U22714 ( .A1(n19831), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19832) );
  OAI211_X1 U22715 ( .C1(n19835), .C2(n19834), .A(n19833), .B(n19832), .ZN(
        n19836) );
  INV_X1 U22716 ( .A(n19836), .ZN(n19846) );
  OAI22_X1 U22717 ( .A1(n19839), .A2(n19841), .B1(n19838), .B2(n19837), .ZN(
        n19840) );
  INV_X1 U22718 ( .A(n19840), .ZN(n19845) );
  NAND2_X1 U22719 ( .A1(n12502), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n19844) );
  NAND3_X1 U22720 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19842), .A3(
        n19841), .ZN(n19843) );
  NAND4_X1 U22721 ( .A1(n19846), .A2(n19845), .A3(n19844), .A4(n19843), .ZN(
        P1_U3029) );
  NOR2_X1 U22722 ( .A1(n19848), .A2(n19847), .ZN(P1_U3032) );
  NOR2_X2 U22723 ( .A1(n19852), .A2(n19851), .ZN(n19894) );
  AOI22_X1 U22724 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19850), .B1(DATAI_16_), 
        .B2(n19894), .ZN(n20352) );
  INV_X1 U22725 ( .A(n19931), .ZN(n19853) );
  NAND2_X1 U22726 ( .A1(n19932), .A2(n19853), .ZN(n20201) );
  AOI22_X1 U22727 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19850), .B1(DATAI_24_), 
        .B2(n19894), .ZN(n20302) );
  INV_X1 U22728 ( .A(n20302), .ZN(n20349) );
  NOR2_X2 U22729 ( .A1(n19896), .A2(n19855), .ZN(n20340) );
  NOR3_X1 U22730 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19909) );
  NAND2_X1 U22731 ( .A1(n20259), .A2(n19909), .ZN(n19861) );
  INV_X1 U22732 ( .A(n19861), .ZN(n19897) );
  AOI22_X1 U22733 ( .A1(n19898), .A2(n20349), .B1(n20340), .B2(n19897), .ZN(
        n19870) );
  INV_X1 U22734 ( .A(n19856), .ZN(n20112) );
  INV_X1 U22735 ( .A(n20165), .ZN(n19857) );
  NOR2_X1 U22736 ( .A1(n20112), .A2(n19857), .ZN(n19866) );
  NAND2_X1 U22737 ( .A1(n19865), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20287) );
  AND2_X1 U22738 ( .A1(n20287), .A2(n19858), .ZN(n20167) );
  NAND2_X1 U22739 ( .A1(n19930), .A2(n20398), .ZN(n19859) );
  AOI21_X1 U22740 ( .B1(n19859), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20346), 
        .ZN(n19864) );
  NOR2_X1 U22741 ( .A1(n20110), .A2(n19860), .ZN(n19962) );
  NAND2_X1 U22742 ( .A1(n19962), .A2(n20111), .ZN(n19867) );
  AOI22_X1 U22743 ( .A1(n19864), .A2(n19867), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n19861), .ZN(n19862) );
  OAI211_X1 U22744 ( .C1(n19866), .C2(n11260), .A(n20167), .B(n19862), .ZN(
        n19901) );
  NOR2_X2 U22745 ( .A1(n19863), .A2(n19999), .ZN(n20339) );
  INV_X1 U22746 ( .A(n19864), .ZN(n19868) );
  NOR2_X1 U22747 ( .A1(n19865), .A2(n11260), .ZN(n20000) );
  INV_X1 U22748 ( .A(n20000), .ZN(n20170) );
  INV_X1 U22749 ( .A(n19866), .ZN(n19995) );
  OAI22_X1 U22750 ( .A1(n19868), .A2(n19867), .B1(n20170), .B2(n19995), .ZN(
        n19900) );
  AOI22_X1 U22751 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19901), .B1(
        n20339), .B2(n19900), .ZN(n19869) );
  OAI211_X1 U22752 ( .C1(n20352), .C2(n19930), .A(n19870), .B(n19869), .ZN(
        P1_U3033) );
  AOI22_X1 U22753 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19850), .B1(DATAI_17_), 
        .B2(n19894), .ZN(n20358) );
  AOI22_X1 U22754 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19850), .B1(DATAI_25_), 
        .B2(n19894), .ZN(n20306) );
  INV_X1 U22755 ( .A(n20306), .ZN(n20355) );
  NOR2_X2 U22756 ( .A1(n19896), .A2(n19871), .ZN(n20354) );
  AOI22_X1 U22757 ( .A1(n19898), .A2(n20355), .B1(n20354), .B2(n19897), .ZN(
        n19874) );
  NOR2_X2 U22758 ( .A1(n19872), .A2(n19999), .ZN(n20353) );
  AOI22_X1 U22759 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19901), .B1(
        n20353), .B2(n19900), .ZN(n19873) );
  OAI211_X1 U22760 ( .C1(n20358), .C2(n19930), .A(n19874), .B(n19873), .ZN(
        P1_U3034) );
  AOI22_X1 U22761 ( .A1(DATAI_18_), .A2(n19894), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n19850), .ZN(n20364) );
  AOI22_X1 U22762 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19850), .B1(DATAI_26_), 
        .B2(n19894), .ZN(n20310) );
  INV_X1 U22763 ( .A(n20310), .ZN(n20361) );
  NOR2_X2 U22764 ( .A1(n19896), .A2(n19875), .ZN(n20360) );
  AOI22_X1 U22765 ( .A1(n19898), .A2(n20361), .B1(n20360), .B2(n19897), .ZN(
        n19878) );
  NOR2_X2 U22766 ( .A1(n19876), .A2(n19999), .ZN(n20359) );
  AOI22_X1 U22767 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19901), .B1(
        n20359), .B2(n19900), .ZN(n19877) );
  OAI211_X1 U22768 ( .C1(n20364), .C2(n19930), .A(n19878), .B(n19877), .ZN(
        P1_U3035) );
  AOI22_X1 U22769 ( .A1(DATAI_19_), .A2(n19894), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n19850), .ZN(n20370) );
  AOI22_X1 U22770 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19850), .B1(DATAI_27_), 
        .B2(n19894), .ZN(n20314) );
  INV_X1 U22771 ( .A(n20314), .ZN(n20367) );
  NOR2_X2 U22772 ( .A1(n19896), .A2(n19879), .ZN(n20366) );
  AOI22_X1 U22773 ( .A1(n19898), .A2(n20367), .B1(n20366), .B2(n19897), .ZN(
        n19882) );
  NOR2_X2 U22774 ( .A1(n19880), .A2(n19999), .ZN(n20365) );
  AOI22_X1 U22775 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19901), .B1(
        n20365), .B2(n19900), .ZN(n19881) );
  OAI211_X1 U22776 ( .C1(n20370), .C2(n19930), .A(n19882), .B(n19881), .ZN(
        P1_U3036) );
  AOI22_X1 U22777 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19850), .B1(DATAI_20_), 
        .B2(n19894), .ZN(n20376) );
  AOI22_X1 U22778 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19850), .B1(DATAI_28_), 
        .B2(n19894), .ZN(n20318) );
  INV_X1 U22779 ( .A(n20318), .ZN(n20373) );
  NOR2_X2 U22780 ( .A1(n19896), .A2(n19883), .ZN(n20372) );
  AOI22_X1 U22781 ( .A1(n19898), .A2(n20373), .B1(n20372), .B2(n19897), .ZN(
        n19886) );
  NOR2_X2 U22782 ( .A1(n19884), .A2(n19999), .ZN(n20371) );
  AOI22_X1 U22783 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19901), .B1(
        n20371), .B2(n19900), .ZN(n19885) );
  OAI211_X1 U22784 ( .C1(n20376), .C2(n19930), .A(n19886), .B(n19885), .ZN(
        P1_U3037) );
  AOI22_X1 U22785 ( .A1(DATAI_21_), .A2(n19894), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n19850), .ZN(n20382) );
  AOI22_X1 U22786 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19850), .B1(DATAI_29_), 
        .B2(n19894), .ZN(n20322) );
  INV_X1 U22787 ( .A(n20322), .ZN(n20379) );
  NOR2_X2 U22788 ( .A1(n19896), .A2(n19887), .ZN(n20378) );
  AOI22_X1 U22789 ( .A1(n19898), .A2(n20379), .B1(n20378), .B2(n19897), .ZN(
        n19890) );
  NOR2_X2 U22790 ( .A1(n19888), .A2(n19999), .ZN(n20377) );
  AOI22_X1 U22791 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19901), .B1(
        n20377), .B2(n19900), .ZN(n19889) );
  OAI211_X1 U22792 ( .C1(n20382), .C2(n19930), .A(n19890), .B(n19889), .ZN(
        P1_U3038) );
  AOI22_X1 U22793 ( .A1(DATAI_22_), .A2(n19894), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n19850), .ZN(n20388) );
  AOI22_X1 U22794 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19850), .B1(DATAI_30_), 
        .B2(n19894), .ZN(n20326) );
  INV_X1 U22795 ( .A(n20326), .ZN(n20385) );
  AOI22_X1 U22796 ( .A1(n19898), .A2(n20385), .B1(n20384), .B2(n19897), .ZN(
        n19893) );
  NOR2_X2 U22797 ( .A1(n19891), .A2(n19999), .ZN(n20383) );
  AOI22_X1 U22798 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19901), .B1(
        n20383), .B2(n19900), .ZN(n19892) );
  OAI211_X1 U22799 ( .C1(n20388), .C2(n19930), .A(n19893), .B(n19892), .ZN(
        P1_U3039) );
  AOI22_X1 U22800 ( .A1(DATAI_23_), .A2(n19894), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n19850), .ZN(n20399) );
  AOI22_X1 U22801 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19850), .B1(DATAI_31_), 
        .B2(n19894), .ZN(n20334) );
  INV_X1 U22802 ( .A(n20334), .ZN(n20393) );
  NOR2_X2 U22803 ( .A1(n19896), .A2(n19895), .ZN(n20392) );
  AOI22_X1 U22804 ( .A1(n19898), .A2(n20393), .B1(n20392), .B2(n19897), .ZN(
        n19903) );
  NOR2_X2 U22805 ( .A1(n19899), .A2(n19999), .ZN(n20390) );
  AOI22_X1 U22806 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19901), .B1(
        n20390), .B2(n19900), .ZN(n19902) );
  OAI211_X1 U22807 ( .C1(n20399), .C2(n19930), .A(n19903), .B(n19902), .ZN(
        P1_U3040) );
  INV_X1 U22808 ( .A(n19909), .ZN(n19905) );
  NOR2_X1 U22809 ( .A1(n20259), .A2(n19905), .ZN(n19926) );
  INV_X1 U22810 ( .A(n19904), .ZN(n20261) );
  AOI21_X1 U22811 ( .B1(n19962), .B2(n20261), .A(n19926), .ZN(n19906) );
  OAI22_X1 U22812 ( .A1(n19906), .A2(n20346), .B1(n19905), .B2(n11260), .ZN(
        n19925) );
  AOI22_X1 U22813 ( .A1(n20340), .A2(n19926), .B1(n20339), .B2(n19925), .ZN(
        n19911) );
  INV_X1 U22814 ( .A(n19964), .ZN(n19907) );
  OAI211_X1 U22815 ( .C1(n19907), .C2(n20291), .A(n20348), .B(n19906), .ZN(
        n19908) );
  OAI211_X1 U22816 ( .C1(n20348), .C2(n19909), .A(n20344), .B(n19908), .ZN(
        n19927) );
  INV_X1 U22817 ( .A(n19930), .ZN(n19922) );
  AOI22_X1 U22818 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19927), .B1(
        n19922), .B2(n20349), .ZN(n19910) );
  OAI211_X1 U22819 ( .C1(n20352), .C2(n19959), .A(n19911), .B(n19910), .ZN(
        P1_U3041) );
  AOI22_X1 U22820 ( .A1(n20354), .A2(n19926), .B1(n20353), .B2(n19925), .ZN(
        n19913) );
  AOI22_X1 U22821 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19927), .B1(
        n19922), .B2(n20355), .ZN(n19912) );
  OAI211_X1 U22822 ( .C1(n20358), .C2(n19959), .A(n19913), .B(n19912), .ZN(
        P1_U3042) );
  AOI22_X1 U22823 ( .A1(n20360), .A2(n19926), .B1(n20359), .B2(n19925), .ZN(
        n19915) );
  AOI22_X1 U22824 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19927), .B1(
        n19922), .B2(n20361), .ZN(n19914) );
  OAI211_X1 U22825 ( .C1(n20364), .C2(n19959), .A(n19915), .B(n19914), .ZN(
        P1_U3043) );
  AOI22_X1 U22826 ( .A1(n20366), .A2(n19926), .B1(n20365), .B2(n19925), .ZN(
        n19917) );
  AOI22_X1 U22827 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19927), .B1(
        n19922), .B2(n20367), .ZN(n19916) );
  OAI211_X1 U22828 ( .C1(n20370), .C2(n19959), .A(n19917), .B(n19916), .ZN(
        P1_U3044) );
  AOI22_X1 U22829 ( .A1(n20372), .A2(n19926), .B1(n20371), .B2(n19925), .ZN(
        n19919) );
  INV_X1 U22830 ( .A(n19959), .ZN(n19951) );
  INV_X1 U22831 ( .A(n20376), .ZN(n20315) );
  AOI22_X1 U22832 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19927), .B1(
        n19951), .B2(n20315), .ZN(n19918) );
  OAI211_X1 U22833 ( .C1(n20318), .C2(n19930), .A(n19919), .B(n19918), .ZN(
        P1_U3045) );
  AOI22_X1 U22834 ( .A1(n20378), .A2(n19926), .B1(n20377), .B2(n19925), .ZN(
        n19921) );
  AOI22_X1 U22835 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19927), .B1(
        n19922), .B2(n20379), .ZN(n19920) );
  OAI211_X1 U22836 ( .C1(n20382), .C2(n19959), .A(n19921), .B(n19920), .ZN(
        P1_U3046) );
  AOI22_X1 U22837 ( .A1(n20384), .A2(n19926), .B1(n20383), .B2(n19925), .ZN(
        n19924) );
  AOI22_X1 U22838 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19927), .B1(
        n19922), .B2(n20385), .ZN(n19923) );
  OAI211_X1 U22839 ( .C1(n20388), .C2(n19959), .A(n19924), .B(n19923), .ZN(
        P1_U3047) );
  AOI22_X1 U22840 ( .A1(n20392), .A2(n19926), .B1(n20390), .B2(n19925), .ZN(
        n19929) );
  INV_X1 U22841 ( .A(n20399), .ZN(n20329) );
  AOI22_X1 U22842 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19927), .B1(
        n19951), .B2(n20329), .ZN(n19928) );
  OAI211_X1 U22843 ( .C1(n20334), .C2(n19930), .A(n19929), .B(n19928), .ZN(
        P1_U3048) );
  INV_X1 U22844 ( .A(n20352), .ZN(n20299) );
  NAND3_X1 U22845 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20626), .A3(
        n20226), .ZN(n19967) );
  NOR2_X1 U22846 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19967), .ZN(
        n19954) );
  AOI22_X1 U22847 ( .A1(n19980), .A2(n20299), .B1(n20340), .B2(n19954), .ZN(
        n19940) );
  NAND2_X1 U22848 ( .A1(n19991), .A2(n19959), .ZN(n19933) );
  AOI21_X1 U22849 ( .B1(n19933), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20346), 
        .ZN(n19936) );
  NAND2_X1 U22850 ( .A1(n19962), .A2(n20294), .ZN(n19937) );
  INV_X1 U22851 ( .A(n19954), .ZN(n19934) );
  AOI22_X1 U22852 ( .A1(n19936), .A2(n19937), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n19934), .ZN(n19935) );
  OR2_X1 U22853 ( .A1(n20165), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20051) );
  NAND2_X1 U22854 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20051), .ZN(n20048) );
  NAND3_X1 U22855 ( .A1(n20167), .A2(n19935), .A3(n20048), .ZN(n19956) );
  INV_X1 U22856 ( .A(n19936), .ZN(n19938) );
  OAI22_X1 U22857 ( .A1(n19938), .A2(n19937), .B1(n20170), .B2(n20051), .ZN(
        n19955) );
  AOI22_X1 U22858 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19956), .B1(
        n20339), .B2(n19955), .ZN(n19939) );
  OAI211_X1 U22859 ( .C1(n20302), .C2(n19959), .A(n19940), .B(n19939), .ZN(
        P1_U3049) );
  AOI22_X1 U22860 ( .A1(n19951), .A2(n20355), .B1(n20354), .B2(n19954), .ZN(
        n19942) );
  AOI22_X1 U22861 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19956), .B1(
        n20353), .B2(n19955), .ZN(n19941) );
  OAI211_X1 U22862 ( .C1(n20358), .C2(n19991), .A(n19942), .B(n19941), .ZN(
        P1_U3050) );
  INV_X1 U22863 ( .A(n20364), .ZN(n20307) );
  AOI22_X1 U22864 ( .A1(n19980), .A2(n20307), .B1(n20360), .B2(n19954), .ZN(
        n19944) );
  AOI22_X1 U22865 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19956), .B1(
        n20359), .B2(n19955), .ZN(n19943) );
  OAI211_X1 U22866 ( .C1(n20310), .C2(n19959), .A(n19944), .B(n19943), .ZN(
        P1_U3051) );
  INV_X1 U22867 ( .A(n20370), .ZN(n20311) );
  AOI22_X1 U22868 ( .A1(n19980), .A2(n20311), .B1(n20366), .B2(n19954), .ZN(
        n19946) );
  AOI22_X1 U22869 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19956), .B1(
        n20365), .B2(n19955), .ZN(n19945) );
  OAI211_X1 U22870 ( .C1(n20314), .C2(n19959), .A(n19946), .B(n19945), .ZN(
        P1_U3052) );
  AOI22_X1 U22871 ( .A1(n19951), .A2(n20373), .B1(n20372), .B2(n19954), .ZN(
        n19948) );
  AOI22_X1 U22872 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19956), .B1(
        n20371), .B2(n19955), .ZN(n19947) );
  OAI211_X1 U22873 ( .C1(n20376), .C2(n19991), .A(n19948), .B(n19947), .ZN(
        P1_U3053) );
  INV_X1 U22874 ( .A(n20382), .ZN(n20319) );
  AOI22_X1 U22875 ( .A1(n19980), .A2(n20319), .B1(n19954), .B2(n20378), .ZN(
        n19950) );
  AOI22_X1 U22876 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19956), .B1(
        n20377), .B2(n19955), .ZN(n19949) );
  OAI211_X1 U22877 ( .C1(n20322), .C2(n19959), .A(n19950), .B(n19949), .ZN(
        P1_U3054) );
  AOI22_X1 U22878 ( .A1(n19951), .A2(n20385), .B1(n20384), .B2(n19954), .ZN(
        n19953) );
  AOI22_X1 U22879 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19956), .B1(
        n20383), .B2(n19955), .ZN(n19952) );
  OAI211_X1 U22880 ( .C1(n20388), .C2(n19991), .A(n19953), .B(n19952), .ZN(
        P1_U3055) );
  AOI22_X1 U22881 ( .A1(n19980), .A2(n20329), .B1(n20392), .B2(n19954), .ZN(
        n19958) );
  AOI22_X1 U22882 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19956), .B1(
        n20390), .B2(n19955), .ZN(n19957) );
  OAI211_X1 U22883 ( .C1(n20334), .C2(n19959), .A(n19958), .B(n19957), .ZN(
        P1_U3056) );
  INV_X1 U22884 ( .A(n20018), .ZN(n19983) );
  NOR2_X1 U22885 ( .A1(n20194), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19986) );
  AOI22_X1 U22886 ( .A1(n19980), .A2(n20349), .B1(n19986), .B2(n20340), .ZN(
        n19971) );
  AND2_X1 U22887 ( .A1(n19961), .A2(n19960), .ZN(n20336) );
  AOI21_X1 U22888 ( .B1(n19962), .B2(n20336), .A(n19986), .ZN(n19968) );
  AOI21_X1 U22889 ( .B1(n19964), .B2(n19963), .A(n20346), .ZN(n19966) );
  AOI22_X1 U22890 ( .A1(n19968), .A2(n19966), .B1(n20346), .B2(n19967), .ZN(
        n19965) );
  NAND2_X1 U22891 ( .A1(n20344), .A2(n19965), .ZN(n19988) );
  INV_X1 U22892 ( .A(n19966), .ZN(n19969) );
  OAI22_X1 U22893 ( .A1(n19969), .A2(n19968), .B1(n11260), .B2(n19967), .ZN(
        n19987) );
  AOI22_X1 U22894 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19988), .B1(
        n20339), .B2(n19987), .ZN(n19970) );
  OAI211_X1 U22895 ( .C1(n20352), .C2(n19983), .A(n19971), .B(n19970), .ZN(
        P1_U3057) );
  INV_X1 U22896 ( .A(n20358), .ZN(n20303) );
  AOI22_X1 U22897 ( .A1(n20018), .A2(n20303), .B1(n20354), .B2(n19986), .ZN(
        n19973) );
  AOI22_X1 U22898 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19988), .B1(
        n20353), .B2(n19987), .ZN(n19972) );
  OAI211_X1 U22899 ( .C1(n20306), .C2(n19991), .A(n19973), .B(n19972), .ZN(
        P1_U3058) );
  AOI22_X1 U22900 ( .A1(n20018), .A2(n20307), .B1(n19986), .B2(n20360), .ZN(
        n19975) );
  AOI22_X1 U22901 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19988), .B1(
        n20359), .B2(n19987), .ZN(n19974) );
  OAI211_X1 U22902 ( .C1(n20310), .C2(n19991), .A(n19975), .B(n19974), .ZN(
        P1_U3059) );
  AOI22_X1 U22903 ( .A1(n20018), .A2(n20311), .B1(n19986), .B2(n20366), .ZN(
        n19977) );
  AOI22_X1 U22904 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19988), .B1(
        n20365), .B2(n19987), .ZN(n19976) );
  OAI211_X1 U22905 ( .C1(n20314), .C2(n19991), .A(n19977), .B(n19976), .ZN(
        P1_U3060) );
  AOI22_X1 U22906 ( .A1(n20018), .A2(n20315), .B1(n19986), .B2(n20372), .ZN(
        n19979) );
  AOI22_X1 U22907 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19988), .B1(
        n20371), .B2(n19987), .ZN(n19978) );
  OAI211_X1 U22908 ( .C1(n20318), .C2(n19991), .A(n19979), .B(n19978), .ZN(
        P1_U3061) );
  AOI22_X1 U22909 ( .A1(n19980), .A2(n20379), .B1(n19986), .B2(n20378), .ZN(
        n19982) );
  AOI22_X1 U22910 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19988), .B1(
        n20377), .B2(n19987), .ZN(n19981) );
  OAI211_X1 U22911 ( .C1(n20382), .C2(n19983), .A(n19982), .B(n19981), .ZN(
        P1_U3062) );
  INV_X1 U22912 ( .A(n20388), .ZN(n20323) );
  AOI22_X1 U22913 ( .A1(n20018), .A2(n20323), .B1(n19986), .B2(n20384), .ZN(
        n19985) );
  AOI22_X1 U22914 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19988), .B1(
        n20383), .B2(n19987), .ZN(n19984) );
  OAI211_X1 U22915 ( .C1(n20326), .C2(n19991), .A(n19985), .B(n19984), .ZN(
        P1_U3063) );
  AOI22_X1 U22916 ( .A1(n20018), .A2(n20329), .B1(n19986), .B2(n20392), .ZN(
        n19990) );
  AOI22_X1 U22917 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19988), .B1(
        n20390), .B2(n19987), .ZN(n19989) );
  OAI211_X1 U22918 ( .C1(n20334), .C2(n19991), .A(n19990), .B(n19989), .ZN(
        P1_U3064) );
  NOR3_X1 U22919 ( .A1(n20226), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20025) );
  INV_X1 U22920 ( .A(n20025), .ZN(n20022) );
  NOR2_X1 U22921 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20022), .ZN(
        n20017) );
  NOR2_X1 U22922 ( .A1(n20230), .A2(n19993), .ZN(n20078) );
  NAND3_X1 U22923 ( .A1(n20078), .A2(n20348), .A3(n20111), .ZN(n19994) );
  OAI21_X1 U22924 ( .B1(n20287), .B2(n19995), .A(n19994), .ZN(n20016) );
  AOI22_X1 U22925 ( .A1(n20340), .A2(n20017), .B1(n20339), .B2(n20016), .ZN(
        n20003) );
  INV_X1 U22926 ( .A(n20078), .ZN(n19998) );
  INV_X1 U22927 ( .A(n20045), .ZN(n19996) );
  OAI21_X1 U22928 ( .B1(n20018), .B2(n19996), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n19997) );
  OAI21_X1 U22929 ( .B1(n20294), .B2(n19998), .A(n19997), .ZN(n20001) );
  AOI22_X1 U22930 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20349), .ZN(n20002) );
  OAI211_X1 U22931 ( .C1(n20352), .C2(n20045), .A(n20003), .B(n20002), .ZN(
        P1_U3065) );
  AOI22_X1 U22932 ( .A1(n20354), .A2(n20017), .B1(n20353), .B2(n20016), .ZN(
        n20005) );
  AOI22_X1 U22933 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20355), .ZN(n20004) );
  OAI211_X1 U22934 ( .C1(n20358), .C2(n20045), .A(n20005), .B(n20004), .ZN(
        P1_U3066) );
  AOI22_X1 U22935 ( .A1(n20360), .A2(n20017), .B1(n20359), .B2(n20016), .ZN(
        n20007) );
  AOI22_X1 U22936 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20361), .ZN(n20006) );
  OAI211_X1 U22937 ( .C1(n20364), .C2(n20045), .A(n20007), .B(n20006), .ZN(
        P1_U3067) );
  AOI22_X1 U22938 ( .A1(n20366), .A2(n20017), .B1(n20365), .B2(n20016), .ZN(
        n20009) );
  AOI22_X1 U22939 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20367), .ZN(n20008) );
  OAI211_X1 U22940 ( .C1(n20370), .C2(n20045), .A(n20009), .B(n20008), .ZN(
        P1_U3068) );
  AOI22_X1 U22941 ( .A1(n20372), .A2(n20017), .B1(n20371), .B2(n20016), .ZN(
        n20011) );
  AOI22_X1 U22942 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20373), .ZN(n20010) );
  OAI211_X1 U22943 ( .C1(n20376), .C2(n20045), .A(n20011), .B(n20010), .ZN(
        P1_U3069) );
  AOI22_X1 U22944 ( .A1(n20378), .A2(n20017), .B1(n20377), .B2(n20016), .ZN(
        n20013) );
  AOI22_X1 U22945 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20379), .ZN(n20012) );
  OAI211_X1 U22946 ( .C1(n20382), .C2(n20045), .A(n20013), .B(n20012), .ZN(
        P1_U3070) );
  AOI22_X1 U22947 ( .A1(n9721), .A2(n20017), .B1(n20383), .B2(n20016), .ZN(
        n20015) );
  AOI22_X1 U22948 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20385), .ZN(n20014) );
  OAI211_X1 U22949 ( .C1(n20388), .C2(n20045), .A(n20015), .B(n20014), .ZN(
        P1_U3071) );
  AOI22_X1 U22950 ( .A1(n20392), .A2(n20017), .B1(n20390), .B2(n20016), .ZN(
        n20021) );
  AOI22_X1 U22951 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20393), .ZN(n20020) );
  OAI211_X1 U22952 ( .C1(n20399), .C2(n20045), .A(n20021), .B(n20020), .ZN(
        P1_U3072) );
  NOR2_X1 U22953 ( .A1(n20259), .A2(n20022), .ZN(n20041) );
  AOI21_X1 U22954 ( .B1(n20078), .B2(n20261), .A(n20041), .ZN(n20023) );
  OAI22_X1 U22955 ( .A1(n20023), .A2(n20346), .B1(n20022), .B2(n11260), .ZN(
        n20040) );
  AOI22_X1 U22956 ( .A1(n20340), .A2(n20041), .B1(n20339), .B2(n20040), .ZN(
        n20027) );
  OAI211_X1 U22957 ( .C1(n20081), .C2(n20291), .A(n20348), .B(n20023), .ZN(
        n20024) );
  OAI211_X1 U22958 ( .C1(n20348), .C2(n20025), .A(n20344), .B(n20024), .ZN(
        n20042) );
  AOI22_X1 U22959 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20299), .ZN(n20026) );
  OAI211_X1 U22960 ( .C1(n20302), .C2(n20045), .A(n20027), .B(n20026), .ZN(
        P1_U3073) );
  AOI22_X1 U22961 ( .A1(n20354), .A2(n20041), .B1(n20353), .B2(n20040), .ZN(
        n20029) );
  AOI22_X1 U22962 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20303), .ZN(n20028) );
  OAI211_X1 U22963 ( .C1(n20306), .C2(n20045), .A(n20029), .B(n20028), .ZN(
        P1_U3074) );
  AOI22_X1 U22964 ( .A1(n20360), .A2(n20041), .B1(n20359), .B2(n20040), .ZN(
        n20031) );
  AOI22_X1 U22965 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20307), .ZN(n20030) );
  OAI211_X1 U22966 ( .C1(n20310), .C2(n20045), .A(n20031), .B(n20030), .ZN(
        P1_U3075) );
  AOI22_X1 U22967 ( .A1(n20366), .A2(n20041), .B1(n20365), .B2(n20040), .ZN(
        n20033) );
  AOI22_X1 U22968 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20311), .ZN(n20032) );
  OAI211_X1 U22969 ( .C1(n20314), .C2(n20045), .A(n20033), .B(n20032), .ZN(
        P1_U3076) );
  AOI22_X1 U22970 ( .A1(n20372), .A2(n20041), .B1(n20371), .B2(n20040), .ZN(
        n20035) );
  AOI22_X1 U22971 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20315), .ZN(n20034) );
  OAI211_X1 U22972 ( .C1(n20318), .C2(n20045), .A(n20035), .B(n20034), .ZN(
        P1_U3077) );
  AOI22_X1 U22973 ( .A1(n20378), .A2(n20041), .B1(n20377), .B2(n20040), .ZN(
        n20037) );
  AOI22_X1 U22974 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20319), .ZN(n20036) );
  OAI211_X1 U22975 ( .C1(n20322), .C2(n20045), .A(n20037), .B(n20036), .ZN(
        P1_U3078) );
  AOI22_X1 U22976 ( .A1(n9721), .A2(n20041), .B1(n20383), .B2(n20040), .ZN(
        n20039) );
  AOI22_X1 U22977 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20323), .ZN(n20038) );
  OAI211_X1 U22978 ( .C1(n20326), .C2(n20045), .A(n20039), .B(n20038), .ZN(
        P1_U3079) );
  AOI22_X1 U22979 ( .A1(n20392), .A2(n20041), .B1(n20390), .B2(n20040), .ZN(
        n20044) );
  AOI22_X1 U22980 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20042), .B1(
        n20070), .B2(n20329), .ZN(n20043) );
  OAI211_X1 U22981 ( .C1(n20334), .C2(n20045), .A(n20044), .B(n20043), .ZN(
        P1_U3080) );
  NAND2_X1 U22982 ( .A1(n20259), .A2(n11291), .ZN(n20047) );
  INV_X1 U22983 ( .A(n20047), .ZN(n20069) );
  AOI22_X1 U22984 ( .A1(n20095), .A2(n20299), .B1(n20340), .B2(n20069), .ZN(
        n20055) );
  NAND2_X1 U22985 ( .A1(n20104), .A2(n20066), .ZN(n20046) );
  AOI21_X1 U22986 ( .B1(n20046), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20346), 
        .ZN(n20050) );
  NAND2_X1 U22987 ( .A1(n20078), .A2(n20294), .ZN(n20052) );
  AOI22_X1 U22988 ( .A1(n20050), .A2(n20052), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20047), .ZN(n20049) );
  NAND3_X1 U22989 ( .A1(n20297), .A2(n20049), .A3(n20048), .ZN(n20072) );
  INV_X1 U22990 ( .A(n20050), .ZN(n20053) );
  OAI22_X1 U22991 ( .A1(n20053), .A2(n20052), .B1(n20051), .B2(n20287), .ZN(
        n20071) );
  AOI22_X1 U22992 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20072), .B1(
        n20339), .B2(n20071), .ZN(n20054) );
  OAI211_X1 U22993 ( .C1(n20302), .C2(n20066), .A(n20055), .B(n20054), .ZN(
        P1_U3081) );
  AOI22_X1 U22994 ( .A1(n20095), .A2(n20303), .B1(n20354), .B2(n20069), .ZN(
        n20057) );
  AOI22_X1 U22995 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20072), .B1(
        n20353), .B2(n20071), .ZN(n20056) );
  OAI211_X1 U22996 ( .C1(n20306), .C2(n20066), .A(n20057), .B(n20056), .ZN(
        P1_U3082) );
  AOI22_X1 U22997 ( .A1(n20070), .A2(n20361), .B1(n20360), .B2(n20069), .ZN(
        n20059) );
  AOI22_X1 U22998 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20072), .B1(
        n20359), .B2(n20071), .ZN(n20058) );
  OAI211_X1 U22999 ( .C1(n20364), .C2(n20104), .A(n20059), .B(n20058), .ZN(
        P1_U3083) );
  AOI22_X1 U23000 ( .A1(n20070), .A2(n20367), .B1(n20366), .B2(n20069), .ZN(
        n20061) );
  AOI22_X1 U23001 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20072), .B1(
        n20365), .B2(n20071), .ZN(n20060) );
  OAI211_X1 U23002 ( .C1(n20370), .C2(n20104), .A(n20061), .B(n20060), .ZN(
        P1_U3084) );
  AOI22_X1 U23003 ( .A1(n20095), .A2(n20315), .B1(n20372), .B2(n20069), .ZN(
        n20063) );
  AOI22_X1 U23004 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20072), .B1(
        n20371), .B2(n20071), .ZN(n20062) );
  OAI211_X1 U23005 ( .C1(n20318), .C2(n20066), .A(n20063), .B(n20062), .ZN(
        P1_U3085) );
  AOI22_X1 U23006 ( .A1(n20095), .A2(n20319), .B1(n20378), .B2(n20069), .ZN(
        n20065) );
  AOI22_X1 U23007 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20072), .B1(
        n20377), .B2(n20071), .ZN(n20064) );
  OAI211_X1 U23008 ( .C1(n20322), .C2(n20066), .A(n20065), .B(n20064), .ZN(
        P1_U3086) );
  AOI22_X1 U23009 ( .A1(n20070), .A2(n20385), .B1(n20384), .B2(n20069), .ZN(
        n20068) );
  AOI22_X1 U23010 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20072), .B1(
        n20383), .B2(n20071), .ZN(n20067) );
  OAI211_X1 U23011 ( .C1(n20388), .C2(n20104), .A(n20068), .B(n20067), .ZN(
        P1_U3087) );
  AOI22_X1 U23012 ( .A1(n20070), .A2(n20393), .B1(n20392), .B2(n20069), .ZN(
        n20074) );
  AOI22_X1 U23013 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20072), .B1(
        n20390), .B2(n20071), .ZN(n20073) );
  OAI211_X1 U23014 ( .C1(n20399), .C2(n20104), .A(n20074), .B(n20073), .ZN(
        P1_U3088) );
  INV_X1 U23015 ( .A(n20077), .ZN(n20100) );
  AOI21_X1 U23016 ( .B1(n20078), .B2(n20336), .A(n20100), .ZN(n20080) );
  OAI22_X1 U23017 ( .A1(n20080), .A2(n20346), .B1(n20079), .B2(n11260), .ZN(
        n20099) );
  AOI22_X1 U23018 ( .A1(n20340), .A2(n20100), .B1(n20339), .B2(n20099), .ZN(
        n20084) );
  OAI211_X1 U23019 ( .C1(n20081), .C2(n20198), .A(n20348), .B(n20080), .ZN(
        n20082) );
  OAI211_X1 U23020 ( .C1(n11291), .C2(n20348), .A(n20344), .B(n20082), .ZN(
        n20101) );
  AOI22_X1 U23021 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20101), .B1(
        n20095), .B2(n20349), .ZN(n20083) );
  OAI211_X1 U23022 ( .C1(n20352), .C2(n20098), .A(n20084), .B(n20083), .ZN(
        P1_U3089) );
  AOI22_X1 U23023 ( .A1(n20354), .A2(n20100), .B1(n20353), .B2(n20099), .ZN(
        n20086) );
  AOI22_X1 U23024 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20101), .B1(
        n20095), .B2(n20355), .ZN(n20085) );
  OAI211_X1 U23025 ( .C1(n20358), .C2(n20098), .A(n20086), .B(n20085), .ZN(
        P1_U3090) );
  AOI22_X1 U23026 ( .A1(n20360), .A2(n20100), .B1(n20359), .B2(n20099), .ZN(
        n20088) );
  AOI22_X1 U23027 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20101), .B1(
        n20095), .B2(n20361), .ZN(n20087) );
  OAI211_X1 U23028 ( .C1(n20364), .C2(n20098), .A(n20088), .B(n20087), .ZN(
        P1_U3091) );
  AOI22_X1 U23029 ( .A1(n20366), .A2(n20100), .B1(n20365), .B2(n20099), .ZN(
        n20090) );
  AOI22_X1 U23030 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20101), .B1(
        n20133), .B2(n20311), .ZN(n20089) );
  OAI211_X1 U23031 ( .C1(n20314), .C2(n20104), .A(n20090), .B(n20089), .ZN(
        P1_U3092) );
  AOI22_X1 U23032 ( .A1(n20372), .A2(n20100), .B1(n20371), .B2(n20099), .ZN(
        n20092) );
  AOI22_X1 U23033 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20101), .B1(
        n20133), .B2(n20315), .ZN(n20091) );
  OAI211_X1 U23034 ( .C1(n20318), .C2(n20104), .A(n20092), .B(n20091), .ZN(
        P1_U3093) );
  AOI22_X1 U23035 ( .A1(n20378), .A2(n20100), .B1(n20377), .B2(n20099), .ZN(
        n20094) );
  AOI22_X1 U23036 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20101), .B1(
        n20095), .B2(n20379), .ZN(n20093) );
  OAI211_X1 U23037 ( .C1(n20382), .C2(n20098), .A(n20094), .B(n20093), .ZN(
        P1_U3094) );
  AOI22_X1 U23038 ( .A1(n9721), .A2(n20100), .B1(n20383), .B2(n20099), .ZN(
        n20097) );
  AOI22_X1 U23039 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20101), .B1(
        n20095), .B2(n20385), .ZN(n20096) );
  OAI211_X1 U23040 ( .C1(n20388), .C2(n20098), .A(n20097), .B(n20096), .ZN(
        P1_U3095) );
  AOI22_X1 U23041 ( .A1(n20392), .A2(n20100), .B1(n20390), .B2(n20099), .ZN(
        n20103) );
  AOI22_X1 U23042 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20101), .B1(
        n20133), .B2(n20329), .ZN(n20102) );
  OAI211_X1 U23043 ( .C1(n20334), .C2(n20104), .A(n20103), .B(n20102), .ZN(
        P1_U3096) );
  INV_X1 U23044 ( .A(n20105), .ZN(n20106) );
  INV_X1 U23045 ( .A(n20202), .ZN(n20109) );
  NOR3_X1 U23046 ( .A1(n20626), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20140) );
  INV_X1 U23047 ( .A(n20140), .ZN(n20137) );
  NOR2_X1 U23048 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20137), .ZN(
        n20132) );
  AND2_X1 U23049 ( .A1(n20110), .A2(n20230), .ZN(n20195) );
  AOI21_X1 U23050 ( .B1(n20195), .B2(n20111), .A(n20132), .ZN(n20114) );
  NAND2_X1 U23051 ( .A1(n20112), .A2(n20165), .ZN(n20234) );
  OAI22_X1 U23052 ( .A1(n20114), .A2(n20346), .B1(n20170), .B2(n20234), .ZN(
        n20131) );
  AOI22_X1 U23053 ( .A1(n20340), .A2(n20132), .B1(n20339), .B2(n20131), .ZN(
        n20118) );
  INV_X1 U23054 ( .A(n20161), .ZN(n20113) );
  OAI21_X1 U23055 ( .B1(n20113), .B2(n20133), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20115) );
  NAND2_X1 U23056 ( .A1(n20115), .A2(n20114), .ZN(n20116) );
  AOI22_X1 U23057 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20349), .ZN(n20117) );
  OAI211_X1 U23058 ( .C1(n20352), .C2(n20161), .A(n20118), .B(n20117), .ZN(
        P1_U3097) );
  AOI22_X1 U23059 ( .A1(n20354), .A2(n20132), .B1(n20353), .B2(n20131), .ZN(
        n20120) );
  AOI22_X1 U23060 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20355), .ZN(n20119) );
  OAI211_X1 U23061 ( .C1(n20358), .C2(n20161), .A(n20120), .B(n20119), .ZN(
        P1_U3098) );
  AOI22_X1 U23062 ( .A1(n20360), .A2(n20132), .B1(n20359), .B2(n20131), .ZN(
        n20122) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20361), .ZN(n20121) );
  OAI211_X1 U23064 ( .C1(n20364), .C2(n20161), .A(n20122), .B(n20121), .ZN(
        P1_U3099) );
  AOI22_X1 U23065 ( .A1(n20366), .A2(n20132), .B1(n20365), .B2(n20131), .ZN(
        n20124) );
  AOI22_X1 U23066 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20367), .ZN(n20123) );
  OAI211_X1 U23067 ( .C1(n20370), .C2(n20161), .A(n20124), .B(n20123), .ZN(
        P1_U3100) );
  AOI22_X1 U23068 ( .A1(n20372), .A2(n20132), .B1(n20371), .B2(n20131), .ZN(
        n20126) );
  AOI22_X1 U23069 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20373), .ZN(n20125) );
  OAI211_X1 U23070 ( .C1(n20376), .C2(n20161), .A(n20126), .B(n20125), .ZN(
        P1_U3101) );
  AOI22_X1 U23071 ( .A1(n20378), .A2(n20132), .B1(n20377), .B2(n20131), .ZN(
        n20128) );
  AOI22_X1 U23072 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20379), .ZN(n20127) );
  OAI211_X1 U23073 ( .C1(n20382), .C2(n20161), .A(n20128), .B(n20127), .ZN(
        P1_U3102) );
  AOI22_X1 U23074 ( .A1(n9721), .A2(n20132), .B1(n20383), .B2(n20131), .ZN(
        n20130) );
  AOI22_X1 U23075 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20385), .ZN(n20129) );
  OAI211_X1 U23076 ( .C1(n20388), .C2(n20161), .A(n20130), .B(n20129), .ZN(
        P1_U3103) );
  AOI22_X1 U23077 ( .A1(n20392), .A2(n20132), .B1(n20390), .B2(n20131), .ZN(
        n20136) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20134), .B1(
        n20133), .B2(n20393), .ZN(n20135) );
  OAI211_X1 U23079 ( .C1(n20399), .C2(n20161), .A(n20136), .B(n20135), .ZN(
        P1_U3104) );
  NOR2_X1 U23080 ( .A1(n20259), .A2(n20137), .ZN(n20157) );
  AOI21_X1 U23081 ( .B1(n20195), .B2(n20261), .A(n20157), .ZN(n20138) );
  OAI22_X1 U23082 ( .A1(n20138), .A2(n20346), .B1(n20137), .B2(n11260), .ZN(
        n20156) );
  AOI22_X1 U23083 ( .A1(n20340), .A2(n20157), .B1(n20339), .B2(n20156), .ZN(
        n20143) );
  OAI211_X1 U23084 ( .C1(n20202), .C2(n20291), .A(n20348), .B(n20138), .ZN(
        n20139) );
  OAI211_X1 U23085 ( .C1(n20348), .C2(n20140), .A(n20344), .B(n20139), .ZN(
        n20158) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20299), .ZN(n20142) );
  OAI211_X1 U23087 ( .C1(n20302), .C2(n20161), .A(n20143), .B(n20142), .ZN(
        P1_U3105) );
  AOI22_X1 U23088 ( .A1(n20354), .A2(n20157), .B1(n20353), .B2(n20156), .ZN(
        n20145) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20303), .ZN(n20144) );
  OAI211_X1 U23090 ( .C1(n20306), .C2(n20161), .A(n20145), .B(n20144), .ZN(
        P1_U3106) );
  AOI22_X1 U23091 ( .A1(n20360), .A2(n20157), .B1(n20359), .B2(n20156), .ZN(
        n20147) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20307), .ZN(n20146) );
  OAI211_X1 U23093 ( .C1(n20310), .C2(n20161), .A(n20147), .B(n20146), .ZN(
        P1_U3107) );
  AOI22_X1 U23094 ( .A1(n20366), .A2(n20157), .B1(n20365), .B2(n20156), .ZN(
        n20149) );
  AOI22_X1 U23095 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20311), .ZN(n20148) );
  OAI211_X1 U23096 ( .C1(n20314), .C2(n20161), .A(n20149), .B(n20148), .ZN(
        P1_U3108) );
  AOI22_X1 U23097 ( .A1(n20372), .A2(n20157), .B1(n20371), .B2(n20156), .ZN(
        n20151) );
  AOI22_X1 U23098 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20315), .ZN(n20150) );
  OAI211_X1 U23099 ( .C1(n20318), .C2(n20161), .A(n20151), .B(n20150), .ZN(
        P1_U3109) );
  AOI22_X1 U23100 ( .A1(n20378), .A2(n20157), .B1(n20377), .B2(n20156), .ZN(
        n20153) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20319), .ZN(n20152) );
  OAI211_X1 U23102 ( .C1(n20322), .C2(n20161), .A(n20153), .B(n20152), .ZN(
        P1_U3110) );
  AOI22_X1 U23103 ( .A1(n9721), .A2(n20157), .B1(n20383), .B2(n20156), .ZN(
        n20155) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20323), .ZN(n20154) );
  OAI211_X1 U23105 ( .C1(n20326), .C2(n20161), .A(n20155), .B(n20154), .ZN(
        P1_U3111) );
  AOI22_X1 U23106 ( .A1(n20392), .A2(n20157), .B1(n20390), .B2(n20156), .ZN(
        n20160) );
  AOI22_X1 U23107 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20158), .B1(
        n20177), .B2(n20329), .ZN(n20159) );
  OAI211_X1 U23108 ( .C1(n20334), .C2(n20161), .A(n20160), .B(n20159), .ZN(
        P1_U3112) );
  NOR3_X1 U23109 ( .A1(n20626), .A2(n20163), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20200) );
  INV_X1 U23110 ( .A(n20200), .ZN(n20196) );
  NOR2_X1 U23111 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20196), .ZN(
        n20188) );
  AOI22_X1 U23112 ( .A1(n20177), .A2(n20349), .B1(n20340), .B2(n20188), .ZN(
        n20174) );
  OAI21_X1 U23113 ( .B1(n20221), .B2(n20177), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20164) );
  NAND2_X1 U23114 ( .A1(n20164), .A2(n20348), .ZN(n20172) );
  AND2_X1 U23115 ( .A1(n20195), .A2(n20294), .ZN(n20169) );
  OR2_X1 U23116 ( .A1(n20165), .A2(n20626), .ZN(n20288) );
  NAND2_X1 U23117 ( .A1(n20288), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20296) );
  OAI21_X1 U23118 ( .B1(n20232), .B2(n20188), .A(n20296), .ZN(n20166) );
  INV_X1 U23119 ( .A(n20166), .ZN(n20168) );
  OAI211_X1 U23120 ( .C1(n20172), .C2(n20169), .A(n20168), .B(n20167), .ZN(
        n20190) );
  INV_X1 U23121 ( .A(n20169), .ZN(n20171) );
  AOI22_X1 U23122 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20190), .B1(
        n20339), .B2(n20189), .ZN(n20173) );
  OAI211_X1 U23123 ( .C1(n20352), .C2(n20218), .A(n20174), .B(n20173), .ZN(
        P1_U3113) );
  AOI22_X1 U23124 ( .A1(n20221), .A2(n20303), .B1(n20354), .B2(n20188), .ZN(
        n20176) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20190), .B1(
        n20353), .B2(n20189), .ZN(n20175) );
  OAI211_X1 U23126 ( .C1(n20306), .C2(n20193), .A(n20176), .B(n20175), .ZN(
        P1_U3114) );
  AOI22_X1 U23127 ( .A1(n20177), .A2(n20361), .B1(n20360), .B2(n20188), .ZN(
        n20179) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20190), .B1(
        n20359), .B2(n20189), .ZN(n20178) );
  OAI211_X1 U23129 ( .C1(n20364), .C2(n20218), .A(n20179), .B(n20178), .ZN(
        P1_U3115) );
  AOI22_X1 U23130 ( .A1(n20221), .A2(n20311), .B1(n20366), .B2(n20188), .ZN(
        n20181) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20190), .B1(
        n20365), .B2(n20189), .ZN(n20180) );
  OAI211_X1 U23132 ( .C1(n20314), .C2(n20193), .A(n20181), .B(n20180), .ZN(
        P1_U3116) );
  AOI22_X1 U23133 ( .A1(n20221), .A2(n20315), .B1(n20372), .B2(n20188), .ZN(
        n20183) );
  AOI22_X1 U23134 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20190), .B1(
        n20371), .B2(n20189), .ZN(n20182) );
  OAI211_X1 U23135 ( .C1(n20318), .C2(n20193), .A(n20183), .B(n20182), .ZN(
        P1_U3117) );
  AOI22_X1 U23136 ( .A1(n20221), .A2(n20319), .B1(n20378), .B2(n20188), .ZN(
        n20185) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20190), .B1(
        n20377), .B2(n20189), .ZN(n20184) );
  OAI211_X1 U23138 ( .C1(n20322), .C2(n20193), .A(n20185), .B(n20184), .ZN(
        P1_U3118) );
  AOI22_X1 U23139 ( .A1(n20221), .A2(n20323), .B1(n20384), .B2(n20188), .ZN(
        n20187) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20190), .B1(
        n20383), .B2(n20189), .ZN(n20186) );
  OAI211_X1 U23141 ( .C1(n20326), .C2(n20193), .A(n20187), .B(n20186), .ZN(
        P1_U3119) );
  AOI22_X1 U23142 ( .A1(n20221), .A2(n20329), .B1(n20392), .B2(n20188), .ZN(
        n20192) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20190), .B1(
        n20390), .B2(n20189), .ZN(n20191) );
  OAI211_X1 U23144 ( .C1(n20334), .C2(n20193), .A(n20192), .B(n20191), .ZN(
        P1_U3120) );
  NOR2_X1 U23145 ( .A1(n20194), .A2(n20626), .ZN(n20220) );
  AOI21_X1 U23146 ( .B1(n20195), .B2(n20336), .A(n20220), .ZN(n20197) );
  OAI22_X1 U23147 ( .A1(n20197), .A2(n20346), .B1(n20196), .B2(n11260), .ZN(
        n20219) );
  AOI22_X1 U23148 ( .A1(n20340), .A2(n20220), .B1(n20339), .B2(n20219), .ZN(
        n20204) );
  OAI211_X1 U23149 ( .C1(n20202), .C2(n20198), .A(n20348), .B(n20197), .ZN(
        n20199) );
  OAI211_X1 U23150 ( .C1(n20348), .C2(n20200), .A(n20344), .B(n20199), .ZN(
        n20222) );
  INV_X1 U23151 ( .A(n20256), .ZN(n20215) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20222), .B1(
        n20215), .B2(n20299), .ZN(n20203) );
  OAI211_X1 U23153 ( .C1(n20302), .C2(n20218), .A(n20204), .B(n20203), .ZN(
        P1_U3121) );
  AOI22_X1 U23154 ( .A1(n20354), .A2(n20220), .B1(n20353), .B2(n20219), .ZN(
        n20206) );
  AOI22_X1 U23155 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20222), .B1(
        n20215), .B2(n20303), .ZN(n20205) );
  OAI211_X1 U23156 ( .C1(n20306), .C2(n20218), .A(n20206), .B(n20205), .ZN(
        P1_U3122) );
  AOI22_X1 U23157 ( .A1(n20360), .A2(n20220), .B1(n20359), .B2(n20219), .ZN(
        n20208) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20222), .B1(
        n20215), .B2(n20307), .ZN(n20207) );
  OAI211_X1 U23159 ( .C1(n20310), .C2(n20218), .A(n20208), .B(n20207), .ZN(
        P1_U3123) );
  AOI22_X1 U23160 ( .A1(n20366), .A2(n20220), .B1(n20365), .B2(n20219), .ZN(
        n20210) );
  AOI22_X1 U23161 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20222), .B1(
        n20215), .B2(n20311), .ZN(n20209) );
  OAI211_X1 U23162 ( .C1(n20314), .C2(n20218), .A(n20210), .B(n20209), .ZN(
        P1_U3124) );
  AOI22_X1 U23163 ( .A1(n20372), .A2(n20220), .B1(n20371), .B2(n20219), .ZN(
        n20212) );
  AOI22_X1 U23164 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20222), .B1(
        n20215), .B2(n20315), .ZN(n20211) );
  OAI211_X1 U23165 ( .C1(n20318), .C2(n20218), .A(n20212), .B(n20211), .ZN(
        P1_U3125) );
  AOI22_X1 U23166 ( .A1(n20378), .A2(n20220), .B1(n20377), .B2(n20219), .ZN(
        n20214) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20222), .B1(
        n20221), .B2(n20379), .ZN(n20213) );
  OAI211_X1 U23168 ( .C1(n20382), .C2(n20256), .A(n20214), .B(n20213), .ZN(
        P1_U3126) );
  AOI22_X1 U23169 ( .A1(n9721), .A2(n20220), .B1(n20383), .B2(n20219), .ZN(
        n20217) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20222), .B1(
        n20215), .B2(n20323), .ZN(n20216) );
  OAI211_X1 U23171 ( .C1(n20326), .C2(n20218), .A(n20217), .B(n20216), .ZN(
        P1_U3127) );
  AOI22_X1 U23172 ( .A1(n20392), .A2(n20220), .B1(n20390), .B2(n20219), .ZN(
        n20224) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20222), .B1(
        n20221), .B2(n20393), .ZN(n20223) );
  OAI211_X1 U23174 ( .C1(n20399), .C2(n20256), .A(n20224), .B(n20223), .ZN(
        P1_U3128) );
  NOR3_X1 U23175 ( .A1(n20226), .A2(n20626), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20265) );
  INV_X1 U23176 ( .A(n20265), .ZN(n20262) );
  NOR2_X1 U23177 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20262), .ZN(
        n20251) );
  AOI22_X1 U23178 ( .A1(n20282), .A2(n20299), .B1(n20340), .B2(n20251), .ZN(
        n20238) );
  INV_X1 U23179 ( .A(n20282), .ZN(n20227) );
  AOI21_X1 U23180 ( .B1(n20227), .B2(n20256), .A(n20291), .ZN(n20228) );
  NOR2_X1 U23181 ( .A1(n20228), .A2(n20346), .ZN(n20233) );
  OR2_X1 U23182 ( .A1(n20230), .A2(n20229), .ZN(n20260) );
  OR2_X1 U23183 ( .A1(n20260), .A2(n20294), .ZN(n20235) );
  AOI22_X1 U23184 ( .A1(n20233), .A2(n20235), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20234), .ZN(n20231) );
  OAI211_X1 U23185 ( .C1(n20251), .C2(n20232), .A(n20297), .B(n20231), .ZN(
        n20253) );
  INV_X1 U23186 ( .A(n20233), .ZN(n20236) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20253), .B1(
        n20339), .B2(n20252), .ZN(n20237) );
  OAI211_X1 U23188 ( .C1(n20302), .C2(n20256), .A(n20238), .B(n20237), .ZN(
        P1_U3129) );
  AOI22_X1 U23189 ( .A1(n20282), .A2(n20303), .B1(n20354), .B2(n20251), .ZN(
        n20240) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20253), .B1(
        n20353), .B2(n20252), .ZN(n20239) );
  OAI211_X1 U23191 ( .C1(n20306), .C2(n20256), .A(n20240), .B(n20239), .ZN(
        P1_U3130) );
  AOI22_X1 U23192 ( .A1(n20282), .A2(n20307), .B1(n20360), .B2(n20251), .ZN(
        n20242) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20253), .B1(
        n20359), .B2(n20252), .ZN(n20241) );
  OAI211_X1 U23194 ( .C1(n20310), .C2(n20256), .A(n20242), .B(n20241), .ZN(
        P1_U3131) );
  AOI22_X1 U23195 ( .A1(n20282), .A2(n20311), .B1(n20366), .B2(n20251), .ZN(
        n20244) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20253), .B1(
        n20365), .B2(n20252), .ZN(n20243) );
  OAI211_X1 U23197 ( .C1(n20314), .C2(n20256), .A(n20244), .B(n20243), .ZN(
        P1_U3132) );
  AOI22_X1 U23198 ( .A1(n20282), .A2(n20315), .B1(n20372), .B2(n20251), .ZN(
        n20246) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20253), .B1(
        n20371), .B2(n20252), .ZN(n20245) );
  OAI211_X1 U23200 ( .C1(n20318), .C2(n20256), .A(n20246), .B(n20245), .ZN(
        P1_U3133) );
  AOI22_X1 U23201 ( .A1(n20282), .A2(n20319), .B1(n20378), .B2(n20251), .ZN(
        n20248) );
  AOI22_X1 U23202 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20253), .B1(
        n20377), .B2(n20252), .ZN(n20247) );
  OAI211_X1 U23203 ( .C1(n20322), .C2(n20256), .A(n20248), .B(n20247), .ZN(
        P1_U3134) );
  AOI22_X1 U23204 ( .A1(n20282), .A2(n20323), .B1(n20384), .B2(n20251), .ZN(
        n20250) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20253), .B1(
        n20383), .B2(n20252), .ZN(n20249) );
  OAI211_X1 U23206 ( .C1(n20326), .C2(n20256), .A(n20250), .B(n20249), .ZN(
        P1_U3135) );
  AOI22_X1 U23207 ( .A1(n20282), .A2(n20329), .B1(n20392), .B2(n20251), .ZN(
        n20255) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20253), .B1(
        n20390), .B2(n20252), .ZN(n20254) );
  OAI211_X1 U23209 ( .C1(n20334), .C2(n20256), .A(n20255), .B(n20254), .ZN(
        P1_U3136) );
  NOR2_X1 U23210 ( .A1(n20259), .A2(n20262), .ZN(n20281) );
  AOI21_X1 U23211 ( .B1(n20337), .B2(n20261), .A(n20281), .ZN(n20263) );
  OAI22_X1 U23212 ( .A1(n20263), .A2(n20346), .B1(n20262), .B2(n11260), .ZN(
        n20280) );
  AOI22_X1 U23213 ( .A1(n20340), .A2(n20281), .B1(n20339), .B2(n20280), .ZN(
        n20267) );
  NOR3_X1 U23214 ( .A1(n20290), .A2(n20346), .A3(n20291), .ZN(n20264) );
  OAI21_X1 U23215 ( .B1(n20265), .B2(n20264), .A(n20344), .ZN(n20283) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20349), .ZN(n20266) );
  OAI211_X1 U23217 ( .C1(n20352), .C2(n20333), .A(n20267), .B(n20266), .ZN(
        P1_U3137) );
  AOI22_X1 U23218 ( .A1(n20354), .A2(n20281), .B1(n20353), .B2(n20280), .ZN(
        n20269) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20355), .ZN(n20268) );
  OAI211_X1 U23220 ( .C1(n20358), .C2(n20333), .A(n20269), .B(n20268), .ZN(
        P1_U3138) );
  AOI22_X1 U23221 ( .A1(n20360), .A2(n20281), .B1(n20359), .B2(n20280), .ZN(
        n20271) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20361), .ZN(n20270) );
  OAI211_X1 U23223 ( .C1(n20364), .C2(n20333), .A(n20271), .B(n20270), .ZN(
        P1_U3139) );
  AOI22_X1 U23224 ( .A1(n20366), .A2(n20281), .B1(n20365), .B2(n20280), .ZN(
        n20273) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20367), .ZN(n20272) );
  OAI211_X1 U23226 ( .C1(n20370), .C2(n20333), .A(n20273), .B(n20272), .ZN(
        P1_U3140) );
  AOI22_X1 U23227 ( .A1(n20372), .A2(n20281), .B1(n20371), .B2(n20280), .ZN(
        n20275) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20373), .ZN(n20274) );
  OAI211_X1 U23229 ( .C1(n20376), .C2(n20333), .A(n20275), .B(n20274), .ZN(
        P1_U3141) );
  AOI22_X1 U23230 ( .A1(n20378), .A2(n20281), .B1(n20377), .B2(n20280), .ZN(
        n20277) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20379), .ZN(n20276) );
  OAI211_X1 U23232 ( .C1(n20382), .C2(n20333), .A(n20277), .B(n20276), .ZN(
        P1_U3142) );
  AOI22_X1 U23233 ( .A1(n9721), .A2(n20281), .B1(n20383), .B2(n20280), .ZN(
        n20279) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20385), .ZN(n20278) );
  OAI211_X1 U23235 ( .C1(n20388), .C2(n20333), .A(n20279), .B(n20278), .ZN(
        P1_U3143) );
  AOI22_X1 U23236 ( .A1(n20392), .A2(n20281), .B1(n20390), .B2(n20280), .ZN(
        n20285) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20283), .B1(
        n20282), .B2(n20393), .ZN(n20284) );
  OAI211_X1 U23238 ( .C1(n20399), .C2(n20333), .A(n20285), .B(n20284), .ZN(
        P1_U3144) );
  INV_X1 U23239 ( .A(n20347), .ZN(n20338) );
  NOR2_X1 U23240 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20338), .ZN(
        n20328) );
  NAND3_X1 U23241 ( .A1(n20337), .A2(n20294), .A3(n20348), .ZN(n20286) );
  OAI21_X1 U23242 ( .B1(n20288), .B2(n20287), .A(n20286), .ZN(n20327) );
  AOI22_X1 U23243 ( .A1(n20340), .A2(n20328), .B1(n20339), .B2(n20327), .ZN(
        n20301) );
  INV_X1 U23244 ( .A(n20394), .ZN(n20292) );
  AOI21_X1 U23245 ( .B1(n20292), .B2(n20333), .A(n20291), .ZN(n20293) );
  AOI21_X1 U23246 ( .B1(n20337), .B2(n20294), .A(n20293), .ZN(n20295) );
  NOR2_X1 U23247 ( .A1(n20295), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20298) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20299), .ZN(n20300) );
  OAI211_X1 U23249 ( .C1(n20302), .C2(n20333), .A(n20301), .B(n20300), .ZN(
        P1_U3145) );
  AOI22_X1 U23250 ( .A1(n20354), .A2(n20328), .B1(n20353), .B2(n20327), .ZN(
        n20305) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20303), .ZN(n20304) );
  OAI211_X1 U23252 ( .C1(n20306), .C2(n20333), .A(n20305), .B(n20304), .ZN(
        P1_U3146) );
  AOI22_X1 U23253 ( .A1(n20360), .A2(n20328), .B1(n20359), .B2(n20327), .ZN(
        n20309) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20307), .ZN(n20308) );
  OAI211_X1 U23255 ( .C1(n20310), .C2(n20333), .A(n20309), .B(n20308), .ZN(
        P1_U3147) );
  AOI22_X1 U23256 ( .A1(n20366), .A2(n20328), .B1(n20365), .B2(n20327), .ZN(
        n20313) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20311), .ZN(n20312) );
  OAI211_X1 U23258 ( .C1(n20314), .C2(n20333), .A(n20313), .B(n20312), .ZN(
        P1_U3148) );
  AOI22_X1 U23259 ( .A1(n20372), .A2(n20328), .B1(n20371), .B2(n20327), .ZN(
        n20317) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20315), .ZN(n20316) );
  OAI211_X1 U23261 ( .C1(n20318), .C2(n20333), .A(n20317), .B(n20316), .ZN(
        P1_U3149) );
  AOI22_X1 U23262 ( .A1(n20378), .A2(n20328), .B1(n20377), .B2(n20327), .ZN(
        n20321) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20319), .ZN(n20320) );
  OAI211_X1 U23264 ( .C1(n20322), .C2(n20333), .A(n20321), .B(n20320), .ZN(
        P1_U3150) );
  AOI22_X1 U23265 ( .A1(n9721), .A2(n20328), .B1(n20383), .B2(n20327), .ZN(
        n20325) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20323), .ZN(n20324) );
  OAI211_X1 U23267 ( .C1(n20326), .C2(n20333), .A(n20325), .B(n20324), .ZN(
        P1_U3151) );
  AOI22_X1 U23268 ( .A1(n20392), .A2(n20328), .B1(n20390), .B2(n20327), .ZN(
        n20332) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20330), .B1(
        n20394), .B2(n20329), .ZN(n20331) );
  OAI211_X1 U23270 ( .C1(n20334), .C2(n20333), .A(n20332), .B(n20331), .ZN(
        P1_U3152) );
  INV_X1 U23271 ( .A(n20335), .ZN(n20391) );
  AOI21_X1 U23272 ( .B1(n20337), .B2(n20336), .A(n20391), .ZN(n20342) );
  OAI22_X1 U23273 ( .A1(n20342), .A2(n20346), .B1(n20338), .B2(n11260), .ZN(
        n20389) );
  AOI22_X1 U23274 ( .A1(n20340), .A2(n20391), .B1(n20339), .B2(n20389), .ZN(
        n20351) );
  INV_X1 U23275 ( .A(n20341), .ZN(n20343) );
  NAND2_X1 U23276 ( .A1(n20343), .A2(n20342), .ZN(n20345) );
  OAI221_X1 U23277 ( .B1(n20348), .B2(n20347), .C1(n20346), .C2(n20345), .A(
        n20344), .ZN(n20395) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20349), .ZN(n20350) );
  OAI211_X1 U23279 ( .C1(n20352), .C2(n20398), .A(n20351), .B(n20350), .ZN(
        P1_U3153) );
  AOI22_X1 U23280 ( .A1(n20354), .A2(n20391), .B1(n20353), .B2(n20389), .ZN(
        n20357) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20355), .ZN(n20356) );
  OAI211_X1 U23282 ( .C1(n20358), .C2(n20398), .A(n20357), .B(n20356), .ZN(
        P1_U3154) );
  AOI22_X1 U23283 ( .A1(n20360), .A2(n20391), .B1(n20359), .B2(n20389), .ZN(
        n20363) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20361), .ZN(n20362) );
  OAI211_X1 U23285 ( .C1(n20364), .C2(n20398), .A(n20363), .B(n20362), .ZN(
        P1_U3155) );
  AOI22_X1 U23286 ( .A1(n20366), .A2(n20391), .B1(n20365), .B2(n20389), .ZN(
        n20369) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20367), .ZN(n20368) );
  OAI211_X1 U23288 ( .C1(n20370), .C2(n20398), .A(n20369), .B(n20368), .ZN(
        P1_U3156) );
  AOI22_X1 U23289 ( .A1(n20372), .A2(n20391), .B1(n20371), .B2(n20389), .ZN(
        n20375) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20373), .ZN(n20374) );
  OAI211_X1 U23291 ( .C1(n20376), .C2(n20398), .A(n20375), .B(n20374), .ZN(
        P1_U3157) );
  AOI22_X1 U23292 ( .A1(n20378), .A2(n20391), .B1(n20377), .B2(n20389), .ZN(
        n20381) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20379), .ZN(n20380) );
  OAI211_X1 U23294 ( .C1(n20382), .C2(n20398), .A(n20381), .B(n20380), .ZN(
        P1_U3158) );
  AOI22_X1 U23295 ( .A1(n9721), .A2(n20391), .B1(n20383), .B2(n20389), .ZN(
        n20387) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20385), .ZN(n20386) );
  OAI211_X1 U23297 ( .C1(n20388), .C2(n20398), .A(n20387), .B(n20386), .ZN(
        P1_U3159) );
  AOI22_X1 U23298 ( .A1(n20392), .A2(n20391), .B1(n20390), .B2(n20389), .ZN(
        n20397) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20393), .ZN(n20396) );
  OAI211_X1 U23300 ( .C1(n20399), .C2(n20398), .A(n20397), .B(n20396), .ZN(
        P1_U3160) );
  NOR2_X1 U23301 ( .A1(n20401), .A2(n20400), .ZN(n20404) );
  INV_X1 U23302 ( .A(n20402), .ZN(n20403) );
  OAI21_X1 U23303 ( .B1(n20404), .B2(n11260), .A(n20403), .ZN(P1_U3163) );
  AND2_X1 U23304 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20405), .ZN(
        P1_U3164) );
  AND2_X1 U23305 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20405), .ZN(
        P1_U3165) );
  AND2_X1 U23306 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20405), .ZN(
        P1_U3166) );
  AND2_X1 U23307 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20405), .ZN(
        P1_U3167) );
  AND2_X1 U23308 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20405), .ZN(
        P1_U3168) );
  AND2_X1 U23309 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20405), .ZN(
        P1_U3169) );
  AND2_X1 U23310 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20405), .ZN(
        P1_U3170) );
  AND2_X1 U23311 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20405), .ZN(
        P1_U3171) );
  AND2_X1 U23312 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20405), .ZN(
        P1_U3172) );
  INV_X1 U23313 ( .A(P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20571) );
  NOR2_X1 U23314 ( .A1(n20475), .A2(n20571), .ZN(P1_U3173) );
  AND2_X1 U23315 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20405), .ZN(
        P1_U3174) );
  AND2_X1 U23316 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20405), .ZN(
        P1_U3175) );
  AND2_X1 U23317 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20405), .ZN(
        P1_U3176) );
  AND2_X1 U23318 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20405), .ZN(
        P1_U3177) );
  AND2_X1 U23319 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20405), .ZN(
        P1_U3178) );
  INV_X1 U23320 ( .A(P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n20507) );
  NOR2_X1 U23321 ( .A1(n20475), .A2(n20507), .ZN(P1_U3179) );
  AND2_X1 U23322 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20405), .ZN(
        P1_U3180) );
  AND2_X1 U23323 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20405), .ZN(
        P1_U3181) );
  AND2_X1 U23324 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20405), .ZN(
        P1_U3182) );
  AND2_X1 U23325 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20405), .ZN(
        P1_U3183) );
  AND2_X1 U23326 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20405), .ZN(
        P1_U3184) );
  INV_X1 U23327 ( .A(P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20534) );
  NOR2_X1 U23328 ( .A1(n20475), .A2(n20534), .ZN(P1_U3185) );
  AND2_X1 U23329 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20405), .ZN(P1_U3186) );
  AND2_X1 U23330 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20405), .ZN(P1_U3187) );
  AND2_X1 U23331 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20405), .ZN(P1_U3188) );
  AND2_X1 U23332 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20405), .ZN(P1_U3189) );
  AND2_X1 U23333 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20405), .ZN(P1_U3190) );
  AND2_X1 U23334 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20405), .ZN(P1_U3191) );
  AND2_X1 U23335 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20405), .ZN(P1_U3192) );
  AND2_X1 U23336 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20405), .ZN(P1_U3193) );
  AND2_X1 U23337 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20406), .ZN(n20421) );
  NOR2_X1 U23338 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20408) );
  OAI21_X1 U23339 ( .B1(n20408), .B2(n20407), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20409) );
  AOI21_X1 U23340 ( .B1(NA), .B2(n20419), .A(n20409), .ZN(n20410) );
  OAI22_X1 U23341 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20421), .B1(n20487), 
        .B2(n20410), .ZN(P1_U3194) );
  INV_X1 U23342 ( .A(n20411), .ZN(n20414) );
  INV_X1 U23343 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20417) );
  NOR2_X1 U23344 ( .A1(n20419), .A2(n20417), .ZN(n20412) );
  OAI22_X1 U23345 ( .A1(n20414), .A2(n20413), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20412), .ZN(n20420) );
  OAI211_X1 U23346 ( .C1(NA), .C2(n20415), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20422), .ZN(n20416) );
  OAI211_X1 U23347 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20417), .A(HOLD), .B(
        n20416), .ZN(n20418) );
  OAI22_X1 U23348 ( .A1(n20421), .A2(n20420), .B1(n20419), .B2(n20418), .ZN(
        P1_U3196) );
  OR2_X1 U23349 ( .A1(n20485), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20462) );
  AOI222_X1 U23350 ( .A1(n20465), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20466), .ZN(n20423) );
  INV_X1 U23351 ( .A(n20423), .ZN(P1_U3197) );
  AOI222_X1 U23352 ( .A1(n20466), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20465), .ZN(n20424) );
  INV_X1 U23353 ( .A(n20424), .ZN(P1_U3198) );
  INV_X1 U23354 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20426) );
  INV_X1 U23355 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20428) );
  OAI222_X1 U23356 ( .A1(n20459), .A2(n20426), .B1(n20425), .B2(n20487), .C1(
        n20428), .C2(n20462), .ZN(P1_U3199) );
  AOI22_X1 U23357 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20465), .ZN(n20427) );
  OAI21_X1 U23358 ( .B1(n20428), .B2(n20459), .A(n20427), .ZN(P1_U3200) );
  AOI22_X1 U23359 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20466), .ZN(n20429) );
  OAI21_X1 U23360 ( .B1(n20430), .B2(n20462), .A(n20429), .ZN(P1_U3201) );
  AOI222_X1 U23361 ( .A1(n20466), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20465), .ZN(n20431) );
  INV_X1 U23362 ( .A(n20431), .ZN(P1_U3202) );
  AOI22_X1 U23363 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20465), .ZN(n20432) );
  OAI21_X1 U23364 ( .B1(n20433), .B2(n20459), .A(n20432), .ZN(P1_U3203) );
  AOI22_X1 U23365 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20466), .ZN(n20434) );
  OAI21_X1 U23366 ( .B1(n20435), .B2(n20462), .A(n20434), .ZN(P1_U3204) );
  AOI222_X1 U23367 ( .A1(n20466), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20465), .ZN(n20436) );
  INV_X1 U23368 ( .A(n20436), .ZN(P1_U3205) );
  AOI222_X1 U23369 ( .A1(n20466), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20465), .ZN(n20437) );
  INV_X1 U23370 ( .A(n20437), .ZN(P1_U3206) );
  AOI222_X1 U23371 ( .A1(n20466), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20465), .ZN(n20438) );
  INV_X1 U23372 ( .A(n20438), .ZN(P1_U3207) );
  AOI222_X1 U23373 ( .A1(n20466), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20465), .ZN(n20439) );
  INV_X1 U23374 ( .A(n20439), .ZN(P1_U3208) );
  AOI222_X1 U23375 ( .A1(n20466), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20465), .ZN(n20440) );
  INV_X1 U23376 ( .A(n20440), .ZN(P1_U3209) );
  AOI222_X1 U23377 ( .A1(n20465), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20502), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20466), .ZN(n20441) );
  INV_X1 U23378 ( .A(n20441), .ZN(P1_U3210) );
  AOI22_X1 U23379 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20465), .ZN(n20442) );
  OAI21_X1 U23380 ( .B1(n20443), .B2(n20459), .A(n20442), .ZN(P1_U3211) );
  AOI22_X1 U23381 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20466), .ZN(n20444) );
  OAI21_X1 U23382 ( .B1(n20445), .B2(n20462), .A(n20444), .ZN(P1_U3212) );
  AOI222_X1 U23383 ( .A1(n20466), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20465), .ZN(n20446) );
  INV_X1 U23384 ( .A(n20446), .ZN(P1_U3213) );
  AOI222_X1 U23385 ( .A1(n20466), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20465), .ZN(n20447) );
  INV_X1 U23386 ( .A(n20447), .ZN(P1_U3214) );
  AOI22_X1 U23387 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20465), .ZN(n20448) );
  OAI21_X1 U23388 ( .B1(n20449), .B2(n20459), .A(n20448), .ZN(P1_U3215) );
  AOI22_X1 U23389 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20502), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20466), .ZN(n20450) );
  OAI21_X1 U23390 ( .B1(n20451), .B2(n20462), .A(n20450), .ZN(P1_U3216) );
  AOI222_X1 U23391 ( .A1(n20465), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20466), .ZN(n20452) );
  INV_X1 U23392 ( .A(n20452), .ZN(P1_U3217) );
  AOI222_X1 U23393 ( .A1(n20466), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20465), .ZN(n20453) );
  INV_X1 U23394 ( .A(n20453), .ZN(P1_U3218) );
  AOI222_X1 U23395 ( .A1(n20466), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20465), .ZN(n20454) );
  INV_X1 U23396 ( .A(n20454), .ZN(P1_U3219) );
  AOI222_X1 U23397 ( .A1(n20466), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20465), .ZN(n20455) );
  INV_X1 U23398 ( .A(n20455), .ZN(P1_U3220) );
  AOI222_X1 U23399 ( .A1(n20466), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20465), .ZN(n20456) );
  INV_X1 U23400 ( .A(n20456), .ZN(P1_U3221) );
  AOI222_X1 U23401 ( .A1(n20466), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20465), .ZN(n20457) );
  INV_X1 U23402 ( .A(n20457), .ZN(P1_U3222) );
  AOI22_X1 U23403 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20465), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20485), .ZN(n20458) );
  OAI21_X1 U23404 ( .B1(n20460), .B2(n20459), .A(n20458), .ZN(P1_U3223) );
  AOI22_X1 U23405 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20466), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20485), .ZN(n20461) );
  OAI21_X1 U23406 ( .B1(n20463), .B2(n20462), .A(n20461), .ZN(P1_U3224) );
  AOI222_X1 U23407 ( .A1(n20466), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20465), .ZN(n20464) );
  INV_X1 U23408 ( .A(n20464), .ZN(P1_U3225) );
  AOI222_X1 U23409 ( .A1(n20466), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20485), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20465), .ZN(n20467) );
  INV_X1 U23410 ( .A(n20467), .ZN(P1_U3226) );
  OAI22_X1 U23411 ( .A1(n20502), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20487), .ZN(n20468) );
  INV_X1 U23412 ( .A(n20468), .ZN(P1_U3458) );
  OAI22_X1 U23413 ( .A1(n20485), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20487), .ZN(n20469) );
  INV_X1 U23414 ( .A(n20469), .ZN(P1_U3459) );
  OAI22_X1 U23415 ( .A1(n20502), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20487), .ZN(n20470) );
  INV_X1 U23416 ( .A(n20470), .ZN(P1_U3460) );
  OAI22_X1 U23417 ( .A1(n20502), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20487), .ZN(n20471) );
  INV_X1 U23418 ( .A(n20471), .ZN(P1_U3461) );
  OAI21_X1 U23419 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20475), .A(n20473), 
        .ZN(n20472) );
  INV_X1 U23420 ( .A(n20472), .ZN(P1_U3464) );
  OAI21_X1 U23421 ( .B1(n20475), .B2(n20474), .A(n20473), .ZN(P1_U3465) );
  AOI21_X1 U23422 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20477) );
  AOI22_X1 U23423 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20477), .B2(n20476), .ZN(n20479) );
  INV_X1 U23424 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20478) );
  AOI22_X1 U23425 ( .A1(n20480), .A2(n20479), .B1(n20478), .B2(n20483), .ZN(
        P1_U3481) );
  INV_X1 U23426 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20484) );
  NOR2_X1 U23427 ( .A1(n20483), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20481) );
  AOI22_X1 U23428 ( .A1(n20484), .A2(n20483), .B1(n20482), .B2(n20481), .ZN(
        P1_U3482) );
  AOI22_X1 U23429 ( .A1(n20487), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20486), 
        .B2(n20485), .ZN(P1_U3483) );
  AOI22_X1 U23430 ( .A1(n20490), .A2(n20489), .B1(P1_STATEBS16_REG_SCAN_IN), 
        .B2(n20488), .ZN(n20493) );
  NOR2_X1 U23431 ( .A1(n20491), .A2(n11260), .ZN(n20498) );
  INV_X1 U23432 ( .A(n20498), .ZN(n20492) );
  OAI21_X1 U23433 ( .B1(n20493), .B2(n20492), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n20495) );
  NAND2_X1 U23434 ( .A1(n20495), .A2(n20494), .ZN(n20501) );
  AOI211_X1 U23435 ( .C1(n20499), .C2(n20498), .A(n20497), .B(n20496), .ZN(
        n20500) );
  MUX2_X1 U23436 ( .A(n20501), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20500), 
        .Z(P1_U3485) );
  MUX2_X1 U23437 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20502), .Z(P1_U3486) );
  INV_X1 U23438 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n20504) );
  AOI22_X1 U23439 ( .A1(n20626), .A2(keyinput51), .B1(keyinput60), .B2(n20504), 
        .ZN(n20503) );
  OAI221_X1 U23440 ( .B1(n20626), .B2(keyinput51), .C1(n20504), .C2(keyinput60), .A(n20503), .ZN(n20515) );
  AOI22_X1 U23441 ( .A1(n20637), .A2(keyinput41), .B1(keyinput59), .B2(n20624), 
        .ZN(n20505) );
  OAI221_X1 U23442 ( .B1(n20637), .B2(keyinput41), .C1(n20624), .C2(keyinput59), .A(n20505), .ZN(n20514) );
  INV_X1 U23443 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n20508) );
  AOI22_X1 U23444 ( .A1(n20508), .A2(keyinput45), .B1(keyinput36), .B2(n20507), 
        .ZN(n20506) );
  OAI221_X1 U23445 ( .B1(n20508), .B2(keyinput45), .C1(n20507), .C2(keyinput36), .A(n20506), .ZN(n20513) );
  INV_X1 U23446 ( .A(DATAI_8_), .ZN(n20510) );
  AOI22_X1 U23447 ( .A1(n20511), .A2(keyinput17), .B1(keyinput53), .B2(n20510), 
        .ZN(n20509) );
  OAI221_X1 U23448 ( .B1(n20511), .B2(keyinput17), .C1(n20510), .C2(keyinput53), .A(n20509), .ZN(n20512) );
  NOR4_X1 U23449 ( .A1(n20515), .A2(n20514), .A3(n20513), .A4(n20512), .ZN(
        n20553) );
  AOI22_X1 U23450 ( .A1(n10720), .A2(keyinput37), .B1(n10684), .B2(keyinput25), 
        .ZN(n20516) );
  OAI221_X1 U23451 ( .B1(n10720), .B2(keyinput37), .C1(n10684), .C2(keyinput25), .A(n20516), .ZN(n20525) );
  AOI22_X1 U23452 ( .A1(n20627), .A2(keyinput63), .B1(keyinput31), .B2(n10030), 
        .ZN(n20517) );
  OAI221_X1 U23453 ( .B1(n20627), .B2(keyinput63), .C1(n10030), .C2(keyinput31), .A(n20517), .ZN(n20524) );
  AOI22_X1 U23454 ( .A1(n20519), .A2(keyinput4), .B1(n20638), .B2(keyinput58), 
        .ZN(n20518) );
  OAI221_X1 U23455 ( .B1(n20519), .B2(keyinput4), .C1(n20638), .C2(keyinput58), 
        .A(n20518), .ZN(n20523) );
  AOI22_X1 U23456 ( .A1(n20625), .A2(keyinput38), .B1(n20521), .B2(keyinput57), 
        .ZN(n20520) );
  OAI221_X1 U23457 ( .B1(n20625), .B2(keyinput38), .C1(n20521), .C2(keyinput57), .A(n20520), .ZN(n20522) );
  NOR4_X1 U23458 ( .A1(n20525), .A2(n20524), .A3(n20523), .A4(n20522), .ZN(
        n20552) );
  INV_X1 U23459 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20528) );
  AOI22_X1 U23460 ( .A1(n20528), .A2(keyinput27), .B1(keyinput61), .B2(n20527), 
        .ZN(n20526) );
  OAI221_X1 U23461 ( .B1(n20528), .B2(keyinput27), .C1(n20527), .C2(keyinput61), .A(n20526), .ZN(n20538) );
  INV_X1 U23462 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20530) );
  AOI22_X1 U23463 ( .A1(n20530), .A2(keyinput54), .B1(n12064), .B2(keyinput1), 
        .ZN(n20529) );
  OAI221_X1 U23464 ( .B1(n20530), .B2(keyinput54), .C1(n12064), .C2(keyinput1), 
        .A(n20529), .ZN(n20537) );
  XNOR2_X1 U23465 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput11), .ZN(
        n20533) );
  XNOR2_X1 U23466 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B(keyinput35), 
        .ZN(n20532) );
  XNOR2_X1 U23467 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B(keyinput55), .ZN(
        n20531) );
  NAND3_X1 U23468 ( .A1(n20533), .A2(n20532), .A3(n20531), .ZN(n20536) );
  XNOR2_X1 U23469 ( .A(n20534), .B(keyinput32), .ZN(n20535) );
  NOR4_X1 U23470 ( .A1(n20538), .A2(n20537), .A3(n20536), .A4(n20535), .ZN(
        n20551) );
  AOI22_X1 U23471 ( .A1(n20628), .A2(keyinput8), .B1(n20631), .B2(keyinput22), 
        .ZN(n20539) );
  OAI221_X1 U23472 ( .B1(n20628), .B2(keyinput8), .C1(n20631), .C2(keyinput22), 
        .A(n20539), .ZN(n20549) );
  INV_X1 U23473 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n20542) );
  INV_X1 U23474 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20541) );
  AOI22_X1 U23475 ( .A1(n20542), .A2(keyinput33), .B1(n20541), .B2(keyinput6), 
        .ZN(n20540) );
  OAI221_X1 U23476 ( .B1(n20542), .B2(keyinput33), .C1(n20541), .C2(keyinput6), 
        .A(n20540), .ZN(n20548) );
  AOI22_X1 U23477 ( .A1(n20544), .A2(keyinput47), .B1(keyinput40), .B2(n20633), 
        .ZN(n20543) );
  OAI221_X1 U23478 ( .B1(n20544), .B2(keyinput47), .C1(n20633), .C2(keyinput40), .A(n20543), .ZN(n20547) );
  INV_X1 U23479 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n20630) );
  AOI22_X1 U23480 ( .A1(n20629), .A2(keyinput9), .B1(n20630), .B2(keyinput0), 
        .ZN(n20545) );
  OAI221_X1 U23481 ( .B1(n20629), .B2(keyinput9), .C1(n20630), .C2(keyinput0), 
        .A(n20545), .ZN(n20546) );
  NOR4_X1 U23482 ( .A1(n20549), .A2(n20548), .A3(n20547), .A4(n20546), .ZN(
        n20550) );
  NAND4_X1 U23483 ( .A1(n20553), .A2(n20552), .A3(n20551), .A4(n20550), .ZN(
        n20619) );
  INV_X1 U23484 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20556) );
  AOI22_X1 U23485 ( .A1(n20556), .A2(keyinput14), .B1(keyinput10), .B2(n20555), 
        .ZN(n20554) );
  OAI221_X1 U23486 ( .B1(n20556), .B2(keyinput14), .C1(n20555), .C2(keyinput10), .A(n20554), .ZN(n20568) );
  AOI22_X1 U23487 ( .A1(n20640), .A2(keyinput44), .B1(n20558), .B2(keyinput50), 
        .ZN(n20557) );
  OAI221_X1 U23488 ( .B1(n20640), .B2(keyinput44), .C1(n20558), .C2(keyinput50), .A(n20557), .ZN(n20567) );
  INV_X1 U23489 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n20561) );
  INV_X1 U23490 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20560) );
  AOI22_X1 U23491 ( .A1(n20561), .A2(keyinput52), .B1(keyinput42), .B2(n20560), 
        .ZN(n20559) );
  OAI221_X1 U23492 ( .B1(n20561), .B2(keyinput52), .C1(n20560), .C2(keyinput42), .A(n20559), .ZN(n20566) );
  AOI22_X1 U23493 ( .A1(n20564), .A2(keyinput34), .B1(keyinput46), .B2(n20563), 
        .ZN(n20562) );
  OAI221_X1 U23494 ( .B1(n20564), .B2(keyinput34), .C1(n20563), .C2(keyinput46), .A(n20562), .ZN(n20565) );
  NOR4_X1 U23495 ( .A1(n20568), .A2(n20567), .A3(n20566), .A4(n20565), .ZN(
        n20617) );
  AOI22_X1 U23496 ( .A1(n20570), .A2(keyinput23), .B1(n14332), .B2(keyinput29), 
        .ZN(n20569) );
  OAI221_X1 U23497 ( .B1(n20570), .B2(keyinput23), .C1(n14332), .C2(keyinput29), .A(n20569), .ZN(n20574) );
  XOR2_X1 U23498 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B(keyinput18), .Z(
        n20573) );
  XNOR2_X1 U23499 ( .A(n20571), .B(keyinput39), .ZN(n20572) );
  OR3_X1 U23500 ( .A1(n20574), .A2(n20573), .A3(n20572), .ZN(n20582) );
  AOI22_X1 U23501 ( .A1(n13687), .A2(keyinput28), .B1(keyinput26), .B2(n20576), 
        .ZN(n20575) );
  OAI221_X1 U23502 ( .B1(n13687), .B2(keyinput28), .C1(n20576), .C2(keyinput26), .A(n20575), .ZN(n20581) );
  INV_X1 U23503 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n20578) );
  AOI22_X1 U23504 ( .A1(n20579), .A2(keyinput24), .B1(keyinput30), .B2(n20578), 
        .ZN(n20577) );
  OAI221_X1 U23505 ( .B1(n20579), .B2(keyinput24), .C1(n20578), .C2(keyinput30), .A(n20577), .ZN(n20580) );
  NOR3_X1 U23506 ( .A1(n20582), .A2(n20581), .A3(n20580), .ZN(n20616) );
  AOI22_X1 U23507 ( .A1(n20585), .A2(keyinput13), .B1(keyinput7), .B2(n20584), 
        .ZN(n20583) );
  OAI221_X1 U23508 ( .B1(n20585), .B2(keyinput13), .C1(n20584), .C2(keyinput7), 
        .A(n20583), .ZN(n20597) );
  INV_X1 U23509 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n20588) );
  AOI22_X1 U23510 ( .A1(n20588), .A2(keyinput62), .B1(n20587), .B2(keyinput56), 
        .ZN(n20586) );
  OAI221_X1 U23511 ( .B1(n20588), .B2(keyinput62), .C1(n20587), .C2(keyinput56), .A(n20586), .ZN(n20596) );
  INV_X1 U23512 ( .A(DATAI_22_), .ZN(n20590) );
  AOI22_X1 U23513 ( .A1(n20591), .A2(keyinput48), .B1(n20590), .B2(keyinput12), 
        .ZN(n20589) );
  OAI221_X1 U23514 ( .B1(n20591), .B2(keyinput48), .C1(n20590), .C2(keyinput12), .A(n20589), .ZN(n20595) );
  INV_X1 U23515 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n20593) );
  AOI22_X1 U23516 ( .A1(n20639), .A2(keyinput15), .B1(n20593), .B2(keyinput2), 
        .ZN(n20592) );
  OAI221_X1 U23517 ( .B1(n20639), .B2(keyinput15), .C1(n20593), .C2(keyinput2), 
        .A(n20592), .ZN(n20594) );
  NOR4_X1 U23518 ( .A1(n20597), .A2(n20596), .A3(n20595), .A4(n20594), .ZN(
        n20615) );
  AOI22_X1 U23519 ( .A1(n20600), .A2(keyinput21), .B1(keyinput19), .B2(n20599), 
        .ZN(n20598) );
  OAI221_X1 U23520 ( .B1(n20600), .B2(keyinput21), .C1(n20599), .C2(keyinput19), .A(n20598), .ZN(n20613) );
  AOI22_X1 U23521 ( .A1(n20603), .A2(keyinput20), .B1(keyinput5), .B2(n20602), 
        .ZN(n20601) );
  OAI221_X1 U23522 ( .B1(n20603), .B2(keyinput20), .C1(n20602), .C2(keyinput5), 
        .A(n20601), .ZN(n20612) );
  AOI22_X1 U23523 ( .A1(n20606), .A2(keyinput3), .B1(n20605), .B2(keyinput49), 
        .ZN(n20604) );
  OAI221_X1 U23524 ( .B1(n20606), .B2(keyinput3), .C1(n20605), .C2(keyinput49), 
        .A(n20604), .ZN(n20611) );
  AOI22_X1 U23525 ( .A1(n20609), .A2(keyinput43), .B1(keyinput16), .B2(n20608), 
        .ZN(n20607) );
  OAI221_X1 U23526 ( .B1(n20609), .B2(keyinput43), .C1(n20608), .C2(keyinput16), .A(n20607), .ZN(n20610) );
  NOR4_X1 U23527 ( .A1(n20613), .A2(n20612), .A3(n20611), .A4(n20610), .ZN(
        n20614) );
  NAND4_X1 U23528 ( .A1(n20617), .A2(n20616), .A3(n20615), .A4(n20614), .ZN(
        n20618) );
  NOR2_X1 U23529 ( .A1(n20619), .A2(n20618), .ZN(n20656) );
  NOR4_X1 U23530 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_EAX_REG_24__SCAN_IN), .A3(P2_DATAO_REG_29__SCAN_IN), .A4(
        P2_DATAO_REG_24__SCAN_IN), .ZN(n20623) );
  NOR4_X1 U23531 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_4__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_11__2__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n20622) );
  NOR4_X1 U23532 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(
        P2_EBX_REG_18__SCAN_IN), .A3(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n20621) );
  NOR4_X1 U23533 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(DATAI_22_), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A4(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n20620) );
  NAND4_X1 U23534 ( .A1(n20623), .A2(n20622), .A3(n20621), .A4(n20620), .ZN(
        n20654) );
  NAND4_X1 U23535 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(
        P2_LWORD_REG_14__SCAN_IN), .A3(P2_DATAO_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n20653) );
  NOR4_X1 U23536 ( .A1(n20627), .A2(n20626), .A3(n20625), .A4(n20624), .ZN(
        n20636) );
  NOR4_X1 U23537 ( .A1(n20631), .A2(n20630), .A3(n20629), .A4(n20628), .ZN(
        n20635) );
  INV_X1 U23538 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20632) );
  NOR4_X1 U23539 ( .A1(n20633), .A2(n20530), .A3(n20632), .A4(n12064), .ZN(
        n20634) );
  NAND3_X1 U23540 ( .A1(n20636), .A2(n20635), .A3(n20634), .ZN(n20652) );
  NOR4_X1 U23541 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_5__4__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), 
        .A4(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20650) );
  NOR4_X1 U23542 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__6__SCAN_IN), .A3(P3_INSTQUEUE_REG_0__6__SCAN_IN), 
        .A4(P3_DATAO_REG_3__SCAN_IN), .ZN(n20649) );
  NAND4_X1 U23543 ( .A1(n20640), .A2(n20639), .A3(n20638), .A4(n20637), .ZN(
        n20641) );
  NOR4_X1 U23544 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(DATAI_8_), .A3(
        n20642), .A4(n20641), .ZN(n20648) );
  NAND4_X1 U23545 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(
        P1_EBX_REG_16__SCAN_IN), .A3(P1_REIP_REG_10__SCAN_IN), .A4(
        P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20646) );
  NAND4_X1 U23546 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(P2_ADDRESS_REG_7__SCAN_IN), .A3(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A4(P1_DATAWIDTH_REG_22__SCAN_IN), 
        .ZN(n20645) );
  NAND4_X1 U23547 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(P3_REIP_REG_8__SCAN_IN), .A4(
        P3_EAX_REG_28__SCAN_IN), .ZN(n20644) );
  NAND4_X1 U23548 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        P1_EAX_REG_29__SCAN_IN), .A3(BUF1_REG_28__SCAN_IN), .A4(
        P3_REIP_REG_24__SCAN_IN), .ZN(n20643) );
  NOR4_X1 U23549 ( .A1(n20646), .A2(n20645), .A3(n20644), .A4(n20643), .ZN(
        n20647) );
  NAND4_X1 U23550 ( .A1(n20650), .A2(n20649), .A3(n20648), .A4(n20647), .ZN(
        n20651) );
  NOR4_X1 U23551 ( .A1(n20654), .A2(n20653), .A3(n20652), .A4(n20651), .ZN(
        n20655) );
  XNOR2_X1 U23552 ( .A(n20656), .B(n20655), .ZN(n20670) );
  AOI22_X1 U23553 ( .A1(n20660), .A2(n20659), .B1(n20658), .B2(n20657), .ZN(
        n20661) );
  INV_X1 U23554 ( .A(n20661), .ZN(n20667) );
  OAI22_X1 U23555 ( .A1(n20665), .A2(n20664), .B1(n20663), .B2(n20662), .ZN(
        n20666) );
  AOI211_X1 U23556 ( .C1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .C2(n20668), .A(
        n20667), .B(n20666), .ZN(n20669) );
  XOR2_X1 U23557 ( .A(n20670), .B(n20669), .Z(P3_U2900) );
  INV_X2 U11115 ( .A(n19592), .ZN(n13275) );
  AND2_X2 U13212 ( .A1(n10753), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10546) );
  BUF_X2 U11033 ( .A(n15274), .Z(n16763) );
  CLKBUF_X2 U11058 ( .A(n11634), .Z(n11615) );
  CLKBUF_X1 U11060 ( .A(n11073), .Z(n11817) );
  CLKBUF_X1 U11067 ( .A(n11150), .Z(n11165) );
  CLKBUF_X1 U11071 ( .A(n12125), .Z(n12119) );
  NAND2_X1 U11074 ( .A1(n10317), .A2(n10316), .ZN(n10347) );
  NAND2_X1 U11104 ( .A1(n12728), .A2(n12705), .ZN(n19404) );
  CLKBUF_X1 U11124 ( .A(n11148), .Z(n12470) );
  CLKBUF_X1 U11126 ( .A(n10271), .Z(n18868) );
  CLKBUF_X1 U11252 ( .A(n11921), .Z(n13471) );
  CLKBUF_X1 U11261 ( .A(n17047), .Z(n17057) );
  CLKBUF_X1 U11273 ( .A(n17477), .Z(n9601) );
  INV_X1 U11490 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19571) );
  CLKBUF_X1 U12218 ( .A(n16130), .Z(n16138) );
endmodule

