

module b21_C_SARLock_k_128_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4417, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10377;

  BUF_X2 U4923 ( .A(n6588), .Z(n6782) );
  CLKBUF_X2 U4924 ( .A(n6347), .Z(n6356) );
  BUF_X2 U4925 ( .A(n6779), .Z(n4424) );
  INV_X1 U4926 ( .A(n5389), .ZN(n5596) );
  BUF_X2 U4927 ( .A(n5376), .Z(n5594) );
  AND2_X1 U4928 ( .A1(n5947), .A2(n5946), .ZN(n5998) );
  CLKBUF_X2 U4929 ( .A(n5999), .Z(n6347) );
  INV_X1 U4930 ( .A(n10377), .ZN(n4417) );
  INV_X2 U4931 ( .A(n4417), .ZN(P1_U3084) );
  INV_X1 U4932 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10377) );
  INV_X1 U4934 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n4420) );
  INV_X1 U4935 ( .A(n5777), .ZN(n5762) );
  NAND2_X1 U4937 ( .A1(n5013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5010) );
  INV_X2 U4938 ( .A(n6786), .ZN(n6693) );
  BUF_X1 U4939 ( .A(n5937), .Z(n5939) );
  OR2_X1 U4940 ( .A1(n5195), .A2(n5194), .ZN(n4766) );
  INV_X1 U4941 ( .A(n5597), .ZN(n5459) );
  INV_X1 U4942 ( .A(n9399), .ZN(n9361) );
  NAND2_X1 U4944 ( .A1(n6535), .A2(n6526), .ZN(n6063) );
  NAND2_X1 U4945 ( .A1(n8283), .A2(n6433), .ZN(n8280) );
  INV_X1 U4946 ( .A(n7719), .ZN(n9861) );
  NAND2_X1 U4947 ( .A1(n5388), .A2(n5387), .ZN(n9061) );
  INV_X1 U4948 ( .A(n6063), .ZN(n7110) );
  AOI21_X1 U4949 ( .B1(n9390), .B2(n9397), .A(n8492), .ZN(n9375) );
  NAND2_X1 U4950 ( .A1(n6394), .A2(n6449), .ZN(n9519) );
  AND3_X1 U4951 ( .A1(n5104), .A2(n5103), .A3(n5102), .ZN(n10344) );
  INV_X1 U4952 ( .A(n5860), .ZN(n8929) );
  AOI21_X2 U4953 ( .B1(n9325), .B2(n6779), .A(n6557), .ZN(n7151) );
  AND2_X2 U4954 ( .A1(n4520), .A2(n6554), .ZN(n6779) );
  NAND2_X4 U4955 ( .A1(n4534), .A2(n4535), .ZN(n9323) );
  XNOR2_X2 U4956 ( .A(n5010), .B(n5009), .ZN(n5015) );
  OAI211_X2 U4957 ( .C1(n6354), .C2(n6353), .A(n6363), .B(n6352), .ZN(n6367)
         );
  NAND2_X2 U4958 ( .A1(n6692), .A2(n9294), .ZN(n9208) );
  NAND2_X1 U4959 ( .A1(n5709), .A2(n5708), .ZN(n8258) );
  INV_X1 U4960 ( .A(n9452), .ZN(n9256) );
  CLKBUF_X1 U4961 ( .A(n7548), .Z(n4422) );
  INV_X1 U4962 ( .A(n7456), .ZN(n7266) );
  INV_X2 U4963 ( .A(n8453), .ZN(n8448) );
  XNOR2_X1 U4964 ( .A(n5973), .B(n5966), .ZN(n6482) );
  CLKBUF_X2 U4965 ( .A(n6025), .Z(n6344) );
  NAND2_X2 U4966 ( .A1(n6913), .A2(n6912), .ZN(n6893) );
  INV_X2 U4967 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OR2_X1 U4968 ( .A1(n4719), .A2(n9901), .ZN(n4713) );
  NAND2_X1 U4969 ( .A1(n6749), .A2(n6748), .ZN(n9251) );
  NOR2_X1 U4970 ( .A1(n8610), .A2(n8609), .ZN(n8612) );
  AND2_X1 U4971 ( .A1(n8550), .A2(n4596), .ZN(n8610) );
  NAND2_X1 U4972 ( .A1(n9501), .A2(n4739), .ZN(n9482) );
  NAND2_X1 U4973 ( .A1(n5427), .A2(n5734), .ZN(n8891) );
  NAND2_X1 U4974 ( .A1(n4928), .A2(n4927), .ZN(n9170) );
  NAND2_X1 U4975 ( .A1(n8213), .A2(n4899), .ZN(n8222) );
  NAND2_X1 U4976 ( .A1(n6224), .A2(n6223), .ZN(n9610) );
  OR2_X1 U4977 ( .A1(n7737), .A2(n5192), .ZN(n7735) );
  OAI21_X1 U4978 ( .B1(n5385), .B2(n4780), .A(n5384), .ZN(n5396) );
  NAND2_X1 U4979 ( .A1(n5365), .A2(n5364), .ZN(n5385) );
  NAND2_X1 U4980 ( .A1(n6147), .A2(n6146), .ZN(n8158) );
  AND2_X1 U4981 ( .A1(n5689), .A2(n5686), .ZN(n7935) );
  NAND2_X1 U4982 ( .A1(n9477), .A2(n7415), .ZN(n9533) );
  AND2_X1 U4983 ( .A1(n7152), .A2(n6559), .ZN(n6567) );
  NAND2_X1 U4984 ( .A1(n5202), .A2(n5201), .ZN(n9929) );
  INV_X2 U4985 ( .A(n9477), .ZN(n4421) );
  NAND2_X1 U4986 ( .A1(n5217), .A2(n5216), .ZN(n7961) );
  NAND2_X1 U4987 ( .A1(n6087), .A2(n6086), .ZN(n9871) );
  CLKBUF_X2 U4988 ( .A(n6779), .Z(n4423) );
  INV_X2 U4989 ( .A(n6786), .ZN(n6778) );
  INV_X1 U4990 ( .A(n6572), .ZN(n6786) );
  INV_X2 U4991 ( .A(n9489), .ZN(n9530) );
  AND2_X1 U4992 ( .A1(n6545), .A2(n7116), .ZN(n6554) );
  AND2_X1 U4993 ( .A1(n6546), .A2(n6545), .ZN(n6588) );
  NAND2_X1 U4994 ( .A1(n5065), .A2(n4973), .ZN(n5660) );
  NAND2_X1 U4995 ( .A1(n4452), .A2(n6023), .ZN(n9322) );
  NAND2_X1 U4996 ( .A1(n4634), .A2(n5148), .ZN(n5167) );
  INV_X1 U4997 ( .A(n6553), .ZN(n6544) );
  INV_X1 U4998 ( .A(n7436), .ZN(n4823) );
  BUF_X1 U4999 ( .A(n6558), .Z(n9325) );
  NAND4_X1 U5000 ( .A1(n6050), .A2(n6049), .A3(n6048), .A4(n6047), .ZN(n9320)
         );
  NAND2_X1 U5001 ( .A1(n5136), .A2(n5135), .ZN(n5145) );
  AND2_X1 U5002 ( .A1(n6380), .A2(n5969), .ZN(n5971) );
  OR2_X1 U5003 ( .A1(n7192), .A2(n5810), .ZN(n7194) );
  NAND2_X1 U5004 ( .A1(n5968), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6380) );
  NAND4_X2 U5005 ( .A1(n5081), .A2(n5080), .A3(n5079), .A4(n5078), .ZN(n10348)
         );
  AND3_X1 U5006 ( .A1(n5064), .A2(n5063), .A3(n5062), .ZN(n9962) );
  NAND4_X1 U5007 ( .A1(n5054), .A2(n5053), .A3(n5052), .A4(n5051), .ZN(n8705)
         );
  BUF_X4 U5008 ( .A(n6000), .Z(n6355) );
  INV_X2 U5010 ( .A(n6054), .ZN(n6342) );
  AND3_X1 U5011 ( .A1(n5036), .A2(n5035), .A3(n5034), .ZN(n7408) );
  NAND2_X1 U5012 ( .A1(n6793), .A2(n6534), .ZN(n7116) );
  AND2_X2 U5013 ( .A1(n5015), .A2(n5016), .ZN(n5597) );
  INV_X1 U5014 ( .A(n5016), .ZN(n9166) );
  INV_X2 U5015 ( .A(n6893), .ZN(n5401) );
  OR2_X1 U5016 ( .A1(n9641), .A2(n6127), .ZN(n5938) );
  XNOR2_X1 U5017 ( .A(n5788), .B(n5787), .ZN(n8343) );
  NAND2_X1 U5018 ( .A1(n5939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5940) );
  INV_X1 U5019 ( .A(n5015), .ZN(n9161) );
  NAND2_X1 U5020 ( .A1(n5014), .A2(n5013), .ZN(n5016) );
  NAND2_X2 U5021 ( .A1(n6837), .A2(P1_U3084), .ZN(n9651) );
  NAND2_X2 U5022 ( .A1(n5032), .A2(n4420), .ZN(n9163) );
  INV_X4 U5023 ( .A(n5032), .ZN(n4538) );
  INV_X2 U5024 ( .A(n5032), .ZN(n6837) );
  OR2_X1 U5025 ( .A1(n4450), .A2(n4753), .ZN(n4436) );
  NOR2_X1 U5026 ( .A1(n4988), .A2(n4987), .ZN(n4992) );
  INV_X1 U5027 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6064) );
  NOR2_X1 U5028 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5917) );
  INV_X1 U5029 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6479) );
  NOR2_X1 U5030 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5962) );
  INV_X1 U5031 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6235) );
  NOR2_X2 U5032 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6005) );
  INV_X1 U5033 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4993) );
  INV_X1 U5034 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8376) );
  OAI21_X2 U5035 ( .B1(n6521), .B2(n4753), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6529) );
  NAND2_X2 U5036 ( .A1(n6108), .A2(n4731), .ZN(n6521) );
  NOR2_X2 U5037 ( .A1(n6142), .A2(n5963), .ZN(n6200) );
  AOI211_X2 U5038 ( .C1(n6323), .C2(n8493), .A(n9363), .B(n6322), .ZN(n6354)
         );
  OAI21_X2 U5039 ( .B1(n6629), .B2(n4431), .A(n4930), .ZN(n7977) );
  OAI211_X1 U5040 ( .C1(n6848), .C2(n6054), .A(n6016), .B(n6015), .ZN(n7548)
         );
  OAI21_X2 U5041 ( .B1(n7531), .B2(n6619), .A(n6618), .ZN(n7701) );
  XNOR2_X2 U5042 ( .A(n5971), .B(n5970), .ZN(n6553) );
  AND2_X1 U5043 ( .A1(n4768), .A2(n4975), .ZN(n4767) );
  NAND2_X1 U5044 ( .A1(n5194), .A2(n5193), .ZN(n4768) );
  OR2_X1 U5045 ( .A1(n7088), .A2(n7087), .ZN(n7090) );
  NAND2_X1 U5046 ( .A1(n8391), .A2(n8390), .ZN(n8392) );
  INV_X1 U5047 ( .A(n8974), .ZN(n5360) );
  OR2_X1 U5048 ( .A1(n9027), .A2(n8822), .ZN(n5633) );
  AND2_X1 U5049 ( .A1(n5007), .A2(n4479), .ZN(n5011) );
  INV_X1 U5050 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4855) );
  INV_X1 U5051 ( .A(n8531), .ZN(n4919) );
  AOI21_X1 U5052 ( .B1(n4798), .B2(n4800), .A(n4513), .ZN(n4795) );
  AND2_X1 U5053 ( .A1(n5925), .A2(n5920), .ZN(n4731) );
  NOR2_X1 U5054 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  INV_X1 U5055 ( .A(n5083), .ZN(n5574) );
  NAND2_X2 U5056 ( .A1(n9161), .A2(n5016), .ZN(n5376) );
  AND2_X1 U5057 ( .A1(n5558), .A2(n5903), .ZN(n8458) );
  AND2_X1 U5058 ( .A1(n6063), .A2(n5032), .ZN(n6025) );
  NAND2_X1 U5059 ( .A1(n6063), .A2(n4538), .ZN(n6054) );
  NOR2_X1 U5060 ( .A1(n8794), .A2(n8814), .ZN(n4604) );
  INV_X1 U5061 ( .A(n6668), .ZN(n4926) );
  AOI21_X1 U5062 ( .B1(n4780), .B2(n5384), .A(n5395), .ZN(n4779) );
  NAND2_X1 U5063 ( .A1(n5212), .A2(n5211), .ZN(n5229) );
  OAI21_X1 U5064 ( .B1(n4664), .B2(n8877), .A(n4502), .ZN(n4662) );
  OR2_X1 U5065 ( .A1(n9087), .A2(n8322), .ZN(n5709) );
  INV_X1 U5066 ( .A(n4836), .ZN(n4835) );
  NAND2_X1 U5067 ( .A1(n4836), .A2(n4834), .ZN(n4833) );
  INV_X1 U5068 ( .A(n4837), .ZN(n4834) );
  NAND2_X1 U5069 ( .A1(n7092), .A2(n7408), .ZN(n5662) );
  OR2_X1 U5070 ( .A1(n9131), .A2(n8893), .ZN(n5740) );
  OR2_X1 U5071 ( .A1(n9049), .A2(n8892), .ZN(n5734) );
  OR2_X1 U5072 ( .A1(n4949), .A2(n9220), .ZN(n4945) );
  OR2_X1 U5073 ( .A1(n4950), .A2(n4947), .ZN(n4946) );
  INV_X1 U5074 ( .A(n4512), .ZN(n4949) );
  INV_X1 U5075 ( .A(n7722), .ZN(n4710) );
  AOI21_X1 U5076 ( .B1(n4814), .B2(n4816), .A(n4813), .ZN(n4812) );
  INV_X1 U5077 ( .A(n5461), .ZN(n4813) );
  NAND2_X1 U5078 ( .A1(n5431), .A2(n5430), .ZN(n5444) );
  NAND2_X1 U5079 ( .A1(n5429), .A2(n5428), .ZN(n5431) );
  AND2_X1 U5080 ( .A1(n5364), .A2(n5345), .ZN(n5362) );
  NOR2_X1 U5081 ( .A1(n5320), .A2(n4810), .ZN(n4809) );
  INV_X1 U5082 ( .A(n5296), .ZN(n4810) );
  NAND2_X1 U5083 ( .A1(n5339), .A2(n5325), .ZN(n5340) );
  XNOR2_X1 U5084 ( .A(n5317), .B(SI_14_), .ZN(n5316) );
  NAND2_X1 U5085 ( .A1(n5295), .A2(n4974), .ZN(n5297) );
  OAI21_X1 U5086 ( .B1(n5276), .B2(n5275), .A(n5274), .ZN(n5295) );
  NAND2_X1 U5087 ( .A1(n5172), .A2(n5171), .ZN(n5193) );
  NAND2_X1 U5088 ( .A1(n8222), .A2(n8221), .ZN(n8391) );
  INV_X1 U5089 ( .A(n8464), .ZN(n4887) );
  NAND2_X1 U5090 ( .A1(n7357), .A2(n4585), .ZN(n4583) );
  NAND2_X1 U5091 ( .A1(n4591), .A2(n8645), .ZN(n8642) );
  NAND2_X1 U5092 ( .A1(n8646), .A2(n7233), .ZN(n4591) );
  OR2_X1 U5093 ( .A1(n8343), .A2(n8929), .ZN(n5864) );
  INV_X1 U5094 ( .A(n7803), .ZN(n7087) );
  AND4_X1 U5095 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n7859)
         );
  NOR2_X1 U5096 ( .A1(n7655), .A2(n7656), .ZN(n7678) );
  INV_X1 U5097 ( .A(n4555), .ZN(n8769) );
  AND2_X1 U5098 ( .A1(n5529), .A2(n5528), .ZN(n8802) );
  AND2_X1 U5099 ( .A1(n5547), .A2(n5546), .ZN(n8823) );
  AOI21_X1 U5100 ( .B1(n4700), .B2(n5360), .A(n4495), .ZN(n4699) );
  NAND2_X1 U5101 ( .A1(n8233), .A2(n5827), .ZN(n8259) );
  NAND2_X1 U5102 ( .A1(n5826), .A2(n4695), .ZN(n4694) );
  NOR2_X1 U5103 ( .A1(n8075), .A2(n4696), .ZN(n4695) );
  NAND2_X1 U5104 ( .A1(n8703), .A2(n7440), .ZN(n7444) );
  AND2_X1 U5105 ( .A1(n5655), .A2(n7444), .ZN(n7384) );
  NAND2_X1 U5106 ( .A1(n7600), .A2(n7604), .ZN(n7599) );
  INV_X1 U5107 ( .A(n5901), .ZN(n4829) );
  OR2_X1 U5108 ( .A1(n8689), .A2(n9027), .ZN(n4689) );
  INV_X1 U5109 ( .A(n4690), .ZN(n4687) );
  CLKBUF_X3 U5110 ( .A(n5071), .Z(n5328) );
  AND2_X1 U5111 ( .A1(n6893), .A2(n4538), .ZN(n5071) );
  MUX2_X1 U5112 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5012), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5014) );
  NAND2_X1 U5113 ( .A1(n5023), .A2(n5022), .ZN(n6913) );
  MUX2_X1 U5114 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5021), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5023) );
  NAND2_X1 U5115 ( .A1(n5026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U5116 ( .A1(n9200), .A2(n4920), .ZN(n4917) );
  NAND2_X1 U5117 ( .A1(n9250), .A2(n9253), .ZN(n6750) );
  AND2_X1 U5118 ( .A1(n9646), .A2(n5946), .ZN(n6000) );
  OR2_X1 U5119 ( .A1(n7166), .A2(n7165), .ZN(n4548) );
  AND2_X1 U5120 ( .A1(n5932), .A2(n5931), .ZN(n8499) );
  INV_X1 U5121 ( .A(n9347), .ZN(n8496) );
  AND2_X1 U5122 ( .A1(n9565), .A2(n9399), .ZN(n4705) );
  NAND2_X1 U5123 ( .A1(n4651), .A2(n4659), .ZN(n4650) );
  INV_X1 U5124 ( .A(n4654), .ZN(n4651) );
  AOI21_X1 U5125 ( .B1(n4656), .B2(n4658), .A(n4655), .ZN(n4654) );
  INV_X1 U5126 ( .A(n9519), .ZN(n4655) );
  NAND2_X1 U5127 ( .A1(n4656), .A2(n4659), .ZN(n4652) );
  OR2_X1 U5128 ( .A1(n9621), .A2(n8309), .ZN(n4970) );
  OR2_X1 U5129 ( .A1(n8303), .A2(n9313), .ZN(n8301) );
  AND2_X1 U5130 ( .A1(n7463), .A2(n6564), .ZN(n7288) );
  MUX2_X1 U5131 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5926), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5928) );
  INV_X1 U5132 ( .A(n6140), .ZN(n6128) );
  NOR3_X1 U5133 ( .A1(n6481), .A2(n4794), .A3(n6536), .ZN(n4792) );
  OR2_X1 U5134 ( .A1(n5660), .A2(n5663), .ZN(n4673) );
  OAI21_X1 U5135 ( .B1(n4569), .B2(n4568), .A(n5673), .ZN(n5688) );
  NOR2_X1 U5136 ( .A1(n5658), .A2(n5762), .ZN(n4568) );
  OAI21_X1 U5137 ( .B1(n5659), .B2(n5777), .A(n5669), .ZN(n4569) );
  AND2_X1 U5138 ( .A1(n5717), .A2(n5360), .ZN(n4567) );
  NOR2_X1 U5139 ( .A1(n5719), .A2(n5777), .ZN(n4566) );
  OAI21_X1 U5140 ( .B1(n4454), .B2(n4576), .A(n5760), .ZN(n4575) );
  NAND2_X1 U5141 ( .A1(n5753), .A2(n5752), .ZN(n4576) );
  NAND2_X1 U5142 ( .A1(n4574), .A2(n5895), .ZN(n4573) );
  AOI22_X1 U5143 ( .A1(n5763), .A2(n5762), .B1(n5761), .B2(n5777), .ZN(n4574)
         );
  NAND2_X1 U5144 ( .A1(n4528), .A2(n4525), .ZN(n6319) );
  AND2_X1 U5145 ( .A1(n4818), .A2(n4817), .ZN(n6363) );
  INV_X1 U5146 ( .A(n5362), .ZN(n4803) );
  NAND2_X1 U5147 ( .A1(n5323), .A2(n5322), .ZN(n5339) );
  INV_X1 U5148 ( .A(n4976), .ZN(n4760) );
  NAND2_X1 U5149 ( .A1(n5197), .A2(n10123), .ZN(n5209) );
  INV_X1 U5150 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5916) );
  INV_X1 U5151 ( .A(n7478), .ZN(n4877) );
  AND2_X1 U5152 ( .A1(n8405), .A2(n8400), .ZN(n4901) );
  INV_X1 U5153 ( .A(n8603), .ZN(n8405) );
  OR2_X1 U5154 ( .A1(n5602), .A2(n5900), .ZN(n5764) );
  INV_X1 U5155 ( .A(n4848), .ZN(n4847) );
  OAI21_X1 U5156 ( .B1(n4850), .B2(n4849), .A(n8840), .ZN(n4848) );
  INV_X1 U5157 ( .A(n5748), .ZN(n4849) );
  NOR2_X1 U5158 ( .A1(n8904), .A2(n9049), .ZN(n4607) );
  INV_X1 U5159 ( .A(n4870), .ZN(n4865) );
  NOR2_X1 U5160 ( .A1(n8958), .A2(n4871), .ZN(n4870) );
  INV_X1 U5161 ( .A(n5719), .ZN(n4871) );
  NOR2_X1 U5162 ( .A1(n8940), .A2(n4868), .ZN(n4867) );
  INV_X1 U5163 ( .A(n5641), .ZN(n4868) );
  NAND2_X1 U5164 ( .A1(n5305), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5332) );
  NOR2_X1 U5165 ( .A1(n9092), .A2(n8087), .ZN(n4613) );
  OR2_X1 U5166 ( .A1(n8814), .A2(n8823), .ZN(n5754) );
  NOR2_X1 U5167 ( .A1(n9115), .A2(n8834), .ZN(n8826) );
  OR2_X1 U5168 ( .A1(n9115), .A2(n8802), .ZN(n5635) );
  INV_X1 U5169 ( .A(n8258), .ZN(n8265) );
  NOR2_X1 U5170 ( .A1(n7488), .A2(n7632), .ZN(n7746) );
  INV_X1 U5171 ( .A(n5662), .ZN(n5048) );
  INV_X1 U5172 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5298) );
  NOR2_X1 U5173 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4982) );
  NOR2_X1 U5174 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4983) );
  INV_X1 U5175 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5115) );
  NOR2_X1 U5176 ( .A1(n4854), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U5177 ( .A1(n5346), .A2(n4902), .ZN(n4996) );
  AND2_X1 U5178 ( .A1(n4488), .A2(n4993), .ZN(n4902) );
  INV_X1 U5179 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4903) );
  AND2_X1 U5180 ( .A1(n5100), .A2(n4992), .ZN(n5346) );
  INV_X1 U5181 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n10294) );
  OR2_X1 U5182 ( .A1(n5215), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5256) );
  NOR2_X1 U5183 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4990) );
  NOR2_X1 U5184 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4989) );
  INV_X1 U5185 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4821) );
  AOI21_X1 U5186 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n4921) );
  INV_X1 U5187 ( .A(n6664), .ZN(n4923) );
  INV_X1 U5188 ( .A(n8134), .ZN(n4922) );
  OR2_X1 U5189 ( .A1(n8474), .A2(n8476), .ZN(n6741) );
  NOR2_X1 U5190 ( .A1(n9561), .A2(n4617), .ZN(n4616) );
  INV_X1 U5191 ( .A(n4618), .ZN(n4617) );
  OR2_X1 U5192 ( .A1(n9565), .A2(n9399), .ZN(n8493) );
  NOR2_X1 U5193 ( .A1(n9565), .A2(n9570), .ZN(n4618) );
  INV_X1 U5194 ( .A(n4749), .ZN(n4748) );
  AND2_X1 U5195 ( .A1(n6316), .A2(n9410), .ZN(n8515) );
  NAND2_X1 U5196 ( .A1(n9406), .A2(n9439), .ZN(n4644) );
  NOR2_X1 U5197 ( .A1(n9436), .A2(n4750), .ZN(n4749) );
  INV_X1 U5198 ( .A(n8513), .ZN(n4750) );
  NOR2_X1 U5199 ( .A1(n9592), .A2(n9595), .ZN(n4633) );
  NAND2_X1 U5200 ( .A1(n6269), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6280) );
  OR2_X1 U5201 ( .A1(n9592), .A2(n6286), .ZN(n8512) );
  OAI21_X1 U5202 ( .B1(n4650), .B2(n4435), .A(n4472), .ZN(n4649) );
  NAND2_X1 U5203 ( .A1(n9605), .A2(n9540), .ZN(n4659) );
  NAND2_X1 U5204 ( .A1(n9600), .A2(n9278), .ZN(n8509) );
  OR2_X1 U5205 ( .A1(n9617), .A2(n9302), .ZN(n6445) );
  OR2_X1 U5206 ( .A1(n8183), .A2(n8158), .ZN(n4628) );
  OR2_X1 U5207 ( .A1(n9319), .A2(n9867), .ZN(n7867) );
  OR2_X1 U5208 ( .A1(n9323), .A2(n9848), .ZN(n6421) );
  OR2_X1 U5209 ( .A1(n6573), .A2(n7566), .ZN(n6492) );
  NAND2_X1 U5210 ( .A1(n7266), .A2(n6564), .ZN(n6490) );
  NAND2_X1 U5211 ( .A1(n5535), .A2(n5534), .ZN(n5551) );
  NAND2_X1 U5212 ( .A1(n4783), .A2(n4781), .ZN(n5535) );
  AOI21_X1 U5213 ( .B1(n4784), .B2(n4506), .A(n4782), .ZN(n4781) );
  NOR2_X1 U5214 ( .A1(n5498), .A2(n4789), .ZN(n4788) );
  INV_X1 U5215 ( .A(n5482), .ZN(n4789) );
  AND2_X1 U5216 ( .A1(n5482), .A2(n5469), .ZN(n5480) );
  NAND2_X1 U5217 ( .A1(n4774), .A2(n4772), .ZN(n5429) );
  AOI21_X1 U5218 ( .B1(n4501), .B2(n4776), .A(n4773), .ZN(n4772) );
  INV_X1 U5219 ( .A(n5413), .ZN(n4773) );
  NAND2_X1 U5220 ( .A1(n5279), .A2(n5278), .ZN(n5296) );
  OAI21_X1 U5221 ( .B1(n5248), .B2(n5247), .A(n5246), .ZN(n5276) );
  AOI21_X1 U5222 ( .B1(n4767), .B2(n4764), .A(n4763), .ZN(n4762) );
  INV_X1 U5223 ( .A(n5209), .ZN(n4763) );
  INV_X1 U5224 ( .A(n5193), .ZN(n4764) );
  INV_X1 U5225 ( .A(n4767), .ZN(n4765) );
  NAND2_X1 U5226 ( .A1(n5193), .A2(n5174), .ZN(n5194) );
  NAND2_X1 U5227 ( .A1(n5170), .A2(n5169), .ZN(n5195) );
  CLKBUF_X1 U5228 ( .A(n6036), .Z(n6037) );
  OAI21_X1 U5229 ( .B1(n4538), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4539), .ZN(
        n5088) );
  NAND2_X1 U5230 ( .A1(n6837), .A2(n6843), .ZN(n4539) );
  NAND2_X1 U5231 ( .A1(n8431), .A2(n8430), .ZN(n8436) );
  INV_X1 U5232 ( .A(n7837), .ZN(n7839) );
  NAND2_X1 U5233 ( .A1(n4874), .A2(n4872), .ZN(n7836) );
  AOI21_X1 U5234 ( .B1(n4451), .B2(n4875), .A(n4873), .ZN(n4872) );
  INV_X1 U5235 ( .A(n8454), .ZN(n4893) );
  NAND2_X1 U5236 ( .A1(n4587), .A2(n4515), .ZN(n4584) );
  NOR2_X1 U5237 ( .A1(n8436), .A2(n8435), .ZN(n8609) );
  INV_X1 U5238 ( .A(n8434), .ZN(n8435) );
  NAND2_X1 U5239 ( .A1(n8556), .A2(n8412), .ZN(n8557) );
  NAND2_X1 U5240 ( .A1(n8029), .A2(n8028), .ZN(n8213) );
  INV_X1 U5241 ( .A(n4901), .ZN(n4595) );
  NAND2_X1 U5242 ( .A1(n8473), .A2(n4901), .ZN(n8654) );
  INV_X1 U5243 ( .A(n4584), .ZN(n4582) );
  NAND2_X1 U5244 ( .A1(n8392), .A2(n8393), .ZN(n8671) );
  NAND2_X1 U5245 ( .A1(n8395), .A2(n8394), .ZN(n8672) );
  INV_X1 U5246 ( .A(n8343), .ZN(n5805) );
  NAND2_X1 U5247 ( .A1(n5864), .A2(n7102), .ZN(n7088) );
  AND2_X1 U5248 ( .A1(n5479), .A2(n5478), .ZN(n8634) );
  AND4_X1 U5249 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), .ZN(n7377)
         );
  OAI211_X1 U5250 ( .C1(n8709), .C2(P2_REG2_REG_1__SCAN_IN), .A(n4564), .B(
        n4563), .ZN(n8711) );
  NOR2_X1 U5251 ( .A1(n8708), .A2(n6908), .ZN(n4564) );
  NAND2_X1 U5252 ( .A1(n8709), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4563) );
  INV_X1 U5253 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U5254 ( .A1(n9115), .A2(n8802), .ZN(n8799) );
  AOI21_X1 U5255 ( .B1(n8589), .B2(n5574), .A(n5510), .ZN(n8822) );
  NOR2_X1 U5256 ( .A1(n5616), .A2(n4851), .ZN(n4850) );
  INV_X1 U5257 ( .A(n5744), .ZN(n4851) );
  OR2_X1 U5258 ( .A1(n8858), .A2(n8690), .ZN(n5748) );
  NAND2_X1 U5259 ( .A1(n4859), .A2(n5740), .ZN(n4857) );
  AND2_X1 U5260 ( .A1(n5745), .A2(n5744), .ZN(n8865) );
  NAND2_X1 U5261 ( .A1(n4861), .A2(n4862), .ZN(n4860) );
  INV_X1 U5262 ( .A(n8891), .ZN(n4861) );
  NAND2_X1 U5263 ( .A1(n5408), .A2(n5407), .ZN(n5422) );
  INV_X1 U5264 ( .A(n5406), .ZN(n5408) );
  NAND2_X1 U5265 ( .A1(n5361), .A2(n5360), .ZN(n8976) );
  NOR2_X1 U5266 ( .A1(n4702), .A2(n4701), .ZN(n4700) );
  INV_X1 U5267 ( .A(n4505), .ZN(n4701) );
  OR2_X1 U5268 ( .A1(n8969), .A2(n5360), .ZN(n4703) );
  AND4_X1 U5269 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n8956)
         );
  NAND2_X1 U5270 ( .A1(n4839), .A2(n4840), .ZN(n8320) );
  AOI21_X1 U5271 ( .B1(n5315), .B2(n8235), .A(n4841), .ZN(n4840) );
  INV_X1 U5272 ( .A(n5709), .ZN(n4841) );
  AND4_X1 U5273 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n8978)
         );
  NOR2_X1 U5274 ( .A1(n5294), .A2(n4693), .ZN(n4692) );
  INV_X1 U5275 ( .A(n4697), .ZN(n4693) );
  NAND2_X1 U5276 ( .A1(n4842), .A2(n5294), .ZN(n8267) );
  INV_X1 U5277 ( .A(n8234), .ZN(n4842) );
  AND4_X1 U5278 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n8237)
         );
  OR2_X1 U5279 ( .A1(n5237), .A2(n7858), .ZN(n5264) );
  AND2_X1 U5280 ( .A1(n5689), .A2(n5682), .ZN(n4837) );
  NAND2_X1 U5281 ( .A1(n4474), .A2(n5689), .ZN(n4836) );
  NAND2_X1 U5282 ( .A1(n7735), .A2(n5821), .ZN(n7805) );
  NAND2_X1 U5283 ( .A1(n5164), .A2(n5163), .ZN(n7495) );
  INV_X1 U5284 ( .A(n7491), .ZN(n5163) );
  INV_X1 U5285 ( .A(n5837), .ZN(n5885) );
  AND2_X1 U5286 ( .A1(n5562), .A2(n5756), .ZN(n5837) );
  NAND2_X1 U5287 ( .A1(n4679), .A2(n4677), .ZN(n5886) );
  AOI21_X1 U5288 ( .B1(n4442), .B2(n4680), .A(n4678), .ZN(n4677) );
  NOR2_X1 U5289 ( .A1(n8814), .A2(n8687), .ZN(n4678) );
  NAND2_X1 U5290 ( .A1(n5505), .A2(n5504), .ZN(n9027) );
  NOR2_X1 U5291 ( .A1(n8858), .A2(n4691), .ZN(n4690) );
  INV_X1 U5292 ( .A(n5616), .ZN(n8852) );
  AOI21_X1 U5293 ( .B1(n4667), .B2(n4665), .A(n4496), .ZN(n4664) );
  INV_X1 U5294 ( .A(n8914), .ZN(n4665) );
  OR2_X1 U5295 ( .A1(n9143), .A2(n8946), .ZN(n5833) );
  NAND2_X1 U5296 ( .A1(n5372), .A2(n5371), .ZN(n8960) );
  NAND2_X1 U5297 ( .A1(n5304), .A2(n5303), .ZN(n9087) );
  NAND2_X1 U5298 ( .A1(n4676), .A2(n5816), .ZN(n7453) );
  NOR2_X1 U5299 ( .A1(n5817), .A2(n4675), .ZN(n4674) );
  INV_X1 U5300 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5301 ( .A1(n5346), .A2(n4993), .ZN(n5366) );
  NOR2_X1 U5302 ( .A1(n4468), .A2(n4440), .ZN(n4913) );
  INV_X1 U5303 ( .A(n6723), .ZN(n4939) );
  OR2_X1 U5304 ( .A1(n9192), .A2(n4939), .ZN(n4937) );
  OR2_X1 U5305 ( .A1(n6754), .A2(n4958), .ZN(n4957) );
  INV_X1 U5306 ( .A(n9183), .ZN(n4958) );
  INV_X1 U5307 ( .A(n4931), .ZN(n4930) );
  OAI21_X1 U5308 ( .B1(n4449), .B2(n4431), .A(n4933), .ZN(n4931) );
  INV_X1 U5309 ( .A(n7979), .ZN(n4933) );
  NAND2_X1 U5310 ( .A1(n7701), .A2(n7702), .ZN(n6629) );
  INV_X1 U5311 ( .A(n6579), .ZN(n6582) );
  INV_X1 U5312 ( .A(n6580), .ZN(n6581) );
  NAND2_X1 U5313 ( .A1(n4941), .A2(n4521), .ZN(n9275) );
  AND2_X1 U5314 ( .A1(n4944), .A2(n4438), .ZN(n4521) );
  NAND2_X1 U5315 ( .A1(n6608), .A2(n6611), .ZN(n4963) );
  AND2_X1 U5316 ( .A1(n6617), .A2(n6616), .ZN(n7528) );
  XNOR2_X1 U5317 ( .A(n5930), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6526) );
  OR2_X1 U5318 ( .A1(n6080), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6083) );
  NOR2_X1 U5319 ( .A1(n9781), .A2(n4549), .ZN(n7166) );
  AND2_X1 U5320 ( .A1(n9787), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U5321 ( .A1(n9799), .A2(n9800), .ZN(n7253) );
  INV_X1 U5322 ( .A(n9679), .ZN(n9339) );
  OAI21_X1 U5323 ( .B1(n9382), .B2(n4744), .A(n4743), .ZN(n9351) );
  NAND2_X1 U5324 ( .A1(n8521), .A2(n8519), .ZN(n4744) );
  NAND2_X1 U5325 ( .A1(n9363), .A2(n8521), .ZN(n4743) );
  NOR2_X1 U5326 ( .A1(n9383), .A2(n9384), .ZN(n9382) );
  NOR2_X1 U5327 ( .A1(n9570), .A2(n9414), .ZN(n8492) );
  OR2_X1 U5328 ( .A1(n9586), .A2(n9462), .ZN(n8488) );
  NAND2_X1 U5329 ( .A1(n9482), .A2(n8511), .ZN(n9461) );
  OR2_X1 U5330 ( .A1(n9479), .A2(n9194), .ZN(n4971) );
  OR2_X1 U5331 ( .A1(n9595), .A2(n9504), .ZN(n8485) );
  NOR2_X1 U5332 ( .A1(n9495), .A2(n9595), .ZN(n9476) );
  AND2_X1 U5333 ( .A1(n6393), .A2(n8509), .ZN(n9503) );
  AND2_X1 U5334 ( .A1(n4533), .A2(n4489), .ZN(n4656) );
  NAND2_X1 U5335 ( .A1(n4657), .A2(n4432), .ZN(n4533) );
  OR2_X1 U5336 ( .A1(n4447), .A2(n9617), .ZN(n9529) );
  AND2_X1 U5337 ( .A1(n9517), .A2(n6246), .ZN(n9535) );
  NAND2_X1 U5338 ( .A1(n6191), .A2(n6190), .ZN(n8303) );
  AOI21_X1 U5339 ( .B1(n8281), .B2(n8280), .A(n8279), .ZN(n8302) );
  NAND2_X1 U5340 ( .A1(n8010), .A2(n8009), .ZN(n8012) );
  AOI21_X1 U5341 ( .B1(n8008), .B2(n8007), .A(n8006), .ZN(n8050) );
  AOI21_X1 U5342 ( .B1(n4710), .B2(n7818), .A(n4463), .ZN(n4709) );
  INV_X1 U5343 ( .A(n7818), .ZN(n4711) );
  NAND2_X1 U5344 ( .A1(n7821), .A2(n6401), .ZN(n7869) );
  AND2_X1 U5345 ( .A1(n7869), .A2(n7864), .ZN(n7818) );
  AND2_X1 U5346 ( .A1(n7502), .A2(n7505), .ZN(n4721) );
  NAND2_X1 U5347 ( .A1(n7542), .A2(n7422), .ZN(n7423) );
  CLKBUF_X1 U5348 ( .A(n7419), .Z(n4530) );
  INV_X1 U5349 ( .A(n6383), .ZN(n7412) );
  OR2_X1 U5350 ( .A1(n7296), .A2(n4727), .ZN(n9380) );
  OAI211_X1 U5351 ( .C1(n8348), .C2(n4728), .A(n4726), .B(n4725), .ZN(n7456)
         );
  AND2_X1 U5352 ( .A1(n4730), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U5353 ( .A1(n4723), .A2(n4727), .ZN(n4726) );
  NOR2_X1 U5354 ( .A1(n4436), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4752) );
  OAI21_X1 U5355 ( .B1(n5607), .B2(n5606), .A(n5605), .ZN(n5611) );
  XNOR2_X1 U5356 ( .A(n5607), .B(n5606), .ZN(n9160) );
  OAI21_X1 U5357 ( .B1(n5483), .B2(n4506), .A(n4784), .ZN(n5533) );
  OAI21_X1 U5358 ( .B1(n5444), .B2(n4816), .A(n5448), .ZN(n5463) );
  OAI21_X1 U5359 ( .B1(n5385), .B2(n4778), .A(n4776), .ZN(n5415) );
  OAI21_X1 U5360 ( .B1(n5297), .B2(n4807), .A(n4805), .ZN(n5363) );
  CLKBUF_X1 U5361 ( .A(n6142), .Z(n6143) );
  OR2_X1 U5362 ( .A1(n6083), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6091) );
  XNOR2_X1 U5363 ( .A(n5133), .B(SI_5_), .ZN(n5131) );
  NAND2_X1 U5364 ( .A1(n7376), .A2(n7375), .ZN(n7480) );
  OAI21_X1 U5365 ( .B1(n8663), .B2(n8662), .A(n8447), .ZN(n8541) );
  AND4_X1 U5366 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n8269)
         );
  XNOR2_X1 U5367 ( .A(n8436), .B(n8434), .ZN(n8550) );
  INV_X1 U5368 ( .A(n7239), .ZN(n7240) );
  OAI22_X1 U5369 ( .A1(n4888), .A2(n4883), .B1(n4891), .B2(n4882), .ZN(n4881)
         );
  INV_X1 U5370 ( .A(n8457), .ZN(n4883) );
  NAND2_X1 U5371 ( .A1(n4892), .A2(n4887), .ZN(n4882) );
  NOR2_X1 U5372 ( .A1(n4891), .A2(n4889), .ZN(n4888) );
  NOR2_X1 U5373 ( .A1(n4889), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U5374 ( .A1(n4893), .A2(n4887), .ZN(n4886) );
  NAND2_X1 U5375 ( .A1(n4892), .A2(n4893), .ZN(n4890) );
  OAI21_X1 U5376 ( .B1(n8556), .B2(n4897), .A(n4894), .ZN(n8422) );
  AOI21_X1 U5377 ( .B1(n4896), .B2(n4898), .A(n4895), .ZN(n4894) );
  INV_X1 U5378 ( .A(n4898), .ZN(n4897) );
  NAND2_X1 U5379 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U5380 ( .A1(n5785), .A2(n5784), .ZN(n4571) );
  AOI21_X1 U5381 ( .B1(n8458), .B2(n5574), .A(n5561), .ZN(n8803) );
  NOR2_X1 U5382 ( .A1(n7067), .A2(n7066), .ZN(n7065) );
  OAI21_X1 U5383 ( .B1(n7065), .B2(n7047), .A(n7046), .ZN(n7049) );
  NOR2_X1 U5384 ( .A1(n7680), .A2(n7681), .ZN(n7684) );
  NAND2_X1 U5385 ( .A1(n7684), .A2(n7683), .ZN(n7776) );
  NAND2_X1 U5386 ( .A1(n8771), .A2(n4558), .ZN(n4557) );
  INV_X1 U5387 ( .A(n4559), .ZN(n4558) );
  OAI21_X1 U5388 ( .B1(n8772), .B2(n9906), .A(n9905), .ZN(n4559) );
  XNOR2_X1 U5389 ( .A(n8783), .B(n9103), .ZN(n9010) );
  AND2_X1 U5390 ( .A1(n4825), .A2(n4829), .ZN(n8378) );
  NAND2_X1 U5391 ( .A1(n5556), .A2(n5555), .ZN(n8794) );
  INV_X1 U5392 ( .A(n9081), .ZN(n9071) );
  AOI22_X1 U5393 ( .A1(n6343), .A2(n5117), .B1(n5328), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n9103) );
  AOI21_X1 U5394 ( .B1(n9010), .B2(n9959), .A(n9009), .ZN(n9100) );
  NAND2_X1 U5395 ( .A1(n4825), .A2(n4824), .ZN(n8382) );
  AND2_X1 U5396 ( .A1(n8377), .A2(n4829), .ZN(n4824) );
  AND2_X1 U5397 ( .A1(n9155), .A2(n9093), .ZN(n9142) );
  NAND2_X1 U5398 ( .A1(n4911), .A2(n4430), .ZN(n4910) );
  AOI21_X1 U5399 ( .B1(n9201), .B2(n4913), .A(n4908), .ZN(n4907) );
  NAND2_X1 U5400 ( .A1(n4912), .A2(n4909), .ZN(n4908) );
  NAND2_X1 U5401 ( .A1(n4913), .A2(n4915), .ZN(n4909) );
  OR2_X1 U5402 ( .A1(n9200), .A2(n4916), .ZN(n4915) );
  OAI211_X1 U5403 ( .C1(n6851), .C2(n6054), .A(n6029), .B(n6028), .ZN(n7504)
         );
  INV_X1 U5404 ( .A(n9309), .ZN(n9264) );
  XNOR2_X1 U5405 ( .A(n6745), .B(n7510), .ZN(n9253) );
  INV_X1 U5406 ( .A(n8004), .ZN(n8199) );
  NAND2_X1 U5407 ( .A1(n6132), .A2(n6131), .ZN(n8207) );
  OR2_X1 U5408 ( .A1(n6816), .A2(n4727), .ZN(n9301) );
  OAI21_X1 U5409 ( .B1(n4793), .B2(n6536), .A(n6539), .ZN(n4791) );
  INV_X1 U5410 ( .A(n6524), .ZN(n4793) );
  INV_X1 U5411 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5986) );
  AOI21_X1 U5412 ( .B1(n8373), .B2(n9816), .A(n4553), .ZN(n4552) );
  NAND2_X1 U5413 ( .A1(n9828), .A2(n9420), .ZN(n4553) );
  NAND2_X1 U5414 ( .A1(n4716), .A2(n4712), .ZN(n9554) );
  OR2_X1 U5415 ( .A1(n9344), .A2(n4717), .ZN(n4716) );
  INV_X1 U5416 ( .A(n8524), .ZN(n4717) );
  NAND2_X1 U5417 ( .A1(n9903), .A2(n9887), .ZN(n4714) );
  INV_X1 U5418 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4718) );
  AND2_X1 U5419 ( .A1(n9553), .A2(n4524), .ZN(n4719) );
  AOI21_X1 U5420 ( .B1(n9552), .B2(n9873), .A(n4499), .ZN(n4524) );
  NAND2_X1 U5421 ( .A1(n4719), .A2(n4531), .ZN(n4625) );
  NAND2_X1 U5422 ( .A1(n4532), .A2(n9887), .ZN(n4531) );
  INV_X1 U5423 ( .A(n9554), .ZN(n4532) );
  INV_X1 U5424 ( .A(n9710), .ZN(n8348) );
  CLKBUF_X1 U5425 ( .A(n6540), .Z(n6383) );
  OR2_X1 U5426 ( .A1(n5972), .A2(n6127), .ZN(n5973) );
  OR2_X1 U5427 ( .A1(n5660), .A2(n5665), .ZN(n4671) );
  NAND2_X1 U5428 ( .A1(n5688), .A2(n4461), .ZN(n5691) );
  OAI21_X1 U5429 ( .B1(n6217), .B2(n6216), .A(n6215), .ZN(n6233) );
  MUX2_X1 U5430 ( .A(n6185), .B(n6184), .S(n6371), .Z(n6217) );
  AND2_X1 U5431 ( .A1(n6393), .A2(n6394), .ZN(n4536) );
  OAI21_X1 U5432 ( .B1(n4565), .B2(n8958), .A(n5720), .ZN(n5730) );
  AOI21_X1 U5433 ( .B1(n5718), .B2(n4567), .A(n4566), .ZN(n4565) );
  NAND2_X1 U5434 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  AND2_X1 U5435 ( .A1(n8516), .A2(n4477), .ZN(n4526) );
  OR2_X1 U5436 ( .A1(n6317), .A2(n8514), .ZN(n4527) );
  INV_X1 U5437 ( .A(n5414), .ZN(n4775) );
  NAND2_X1 U5438 ( .A1(n4433), .A2(n4835), .ZN(n4830) );
  NOR2_X1 U5439 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4856) );
  INV_X1 U5440 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4636) );
  INV_X1 U5441 ( .A(n4799), .ZN(n4798) );
  OAI21_X1 U5442 ( .B1(n5550), .B2(n4800), .A(n5563), .ZN(n4799) );
  INV_X1 U5443 ( .A(n5552), .ZN(n4800) );
  INV_X1 U5444 ( .A(n5532), .ZN(n4782) );
  NOR2_X1 U5445 ( .A1(n5462), .A2(n4815), .ZN(n4814) );
  INV_X1 U5446 ( .A(n5448), .ZN(n4815) );
  NAND2_X1 U5447 ( .A1(n5250), .A2(n5249), .ZN(n5274) );
  INV_X1 U5448 ( .A(SI_9_), .ZN(n10123) );
  NOR2_X1 U5449 ( .A1(n5776), .A2(n5770), .ZN(n5773) );
  AOI21_X1 U5450 ( .B1(n4575), .B2(n4456), .A(n4573), .ZN(n5772) );
  NOR2_X1 U5451 ( .A1(n8871), .A2(n8858), .ZN(n8833) );
  OR2_X1 U5452 ( .A1(n9036), .A2(n8634), .ZN(n5745) );
  OR2_X1 U5453 ( .A1(n9080), .A2(n8978), .ZN(n5712) );
  NOR2_X1 U5454 ( .A1(n4612), .A2(n9087), .ZN(n4611) );
  INV_X1 U5455 ( .A(n4613), .ZN(n4612) );
  OR2_X1 U5456 ( .A1(n8087), .A2(n8237), .ZN(n5702) );
  OR2_X1 U5457 ( .A1(n7807), .A2(n9929), .ZN(n7806) );
  NAND2_X1 U5458 ( .A1(n4823), .A2(n4822), .ZN(n5653) );
  INV_X1 U5459 ( .A(n10348), .ZN(n4822) );
  NAND2_X1 U5460 ( .A1(n8826), .A2(n4604), .ZN(n5905) );
  NOR2_X1 U5461 ( .A1(n4603), .A2(n8383), .ZN(n4602) );
  INV_X1 U5462 ( .A(n4604), .ZN(n4603) );
  OR2_X1 U5463 ( .A1(n8383), .A2(n8460), .ZN(n5765) );
  OR2_X1 U5464 ( .A1(n8794), .A2(n8803), .ZN(n5562) );
  NAND2_X1 U5465 ( .A1(n8826), .A2(n9108), .ZN(n8811) );
  INV_X1 U5466 ( .A(n5815), .ZN(n4675) );
  OR2_X1 U5467 ( .A1(n4598), .A2(n8594), .ZN(n7488) );
  NOR2_X1 U5468 ( .A1(n9958), .A2(n7451), .ZN(n4599) );
  NAND2_X1 U5469 ( .A1(n5007), .A2(n4856), .ZN(n5026) );
  INV_X1 U5470 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5001) );
  INV_X1 U5471 ( .A(n7116), .ZN(n6548) );
  NOR2_X1 U5472 ( .A1(n9550), .A2(n9311), .ZN(n6370) );
  INV_X1 U5473 ( .A(n6389), .ZN(n6516) );
  NOR2_X1 U5474 ( .A1(n6370), .A2(n4425), .ZN(n6518) );
  NAND2_X1 U5475 ( .A1(n6347), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4518) );
  INV_X1 U5476 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5920) );
  NOR2_X1 U5477 ( .A1(n7916), .A2(n4550), .ZN(n7917) );
  AND2_X1 U5478 ( .A1(n7923), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4550) );
  OR2_X1 U5479 ( .A1(n9555), .A2(n8534), .ZN(n6469) );
  NAND2_X1 U5480 ( .A1(n9570), .A2(n9233), .ZN(n8517) );
  OR2_X1 U5481 ( .A1(n9570), .A2(n9233), .ZN(n8516) );
  NAND2_X1 U5482 ( .A1(n4633), .A2(n9448), .ZN(n4632) );
  NAND2_X1 U5483 ( .A1(n8175), .A2(n8172), .ZN(n4740) );
  NAND2_X1 U5484 ( .A1(n8183), .A2(n9177), .ZN(n8151) );
  OAI21_X1 U5485 ( .B1(n4737), .B2(n4710), .A(n7991), .ZN(n4735) );
  AND2_X1 U5486 ( .A1(n6113), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6133) );
  NOR2_X1 U5487 ( .A1(n6101), .A2(n6100), .ZN(n6113) );
  OR2_X1 U5488 ( .A1(n6074), .A2(n10095), .ZN(n6101) );
  NAND2_X1 U5489 ( .A1(n7575), .A2(n4441), .ZN(n4622) );
  NAND2_X1 U5490 ( .A1(n4730), .A2(n4729), .ZN(n4723) );
  NAND2_X1 U5491 ( .A1(n4724), .A2(n4538), .ZN(n4730) );
  AND2_X1 U5492 ( .A1(n8510), .A2(n8509), .ZN(n4739) );
  INV_X1 U5493 ( .A(n9485), .ZN(n8510) );
  NAND2_X1 U5494 ( .A1(n7286), .A2(n7287), .ZN(n7460) );
  INV_X1 U5495 ( .A(n5497), .ZN(n4786) );
  INV_X1 U5496 ( .A(n4785), .ZN(n4784) );
  OAI21_X1 U5497 ( .B1(n4788), .B2(n4506), .A(n5511), .ZN(n4785) );
  NAND2_X1 U5498 ( .A1(n6532), .A2(n4754), .ZN(n4753) );
  INV_X1 U5499 ( .A(n5445), .ZN(n4816) );
  INV_X1 U5500 ( .A(n4779), .ZN(n4778) );
  AOI21_X1 U5501 ( .B1(n4779), .B2(n4777), .A(n4500), .ZN(n4776) );
  INV_X1 U5502 ( .A(n5384), .ZN(n4777) );
  INV_X1 U5503 ( .A(n5381), .ZN(n4780) );
  AOI21_X1 U5504 ( .B1(n4805), .B2(n4807), .A(n4803), .ZN(n4802) );
  INV_X1 U5505 ( .A(n4806), .ZN(n4805) );
  OAI21_X1 U5506 ( .B1(n4809), .B2(n4807), .A(n5339), .ZN(n4806) );
  NAND2_X1 U5507 ( .A1(n4808), .A2(n5319), .ZN(n4807) );
  INV_X1 U5508 ( .A(n5340), .ZN(n4808) );
  XNOR2_X1 U5509 ( .A(n5244), .B(SI_11_), .ZN(n5243) );
  NAND2_X1 U5510 ( .A1(n5230), .A2(n5229), .ZN(n5248) );
  NAND2_X1 U5511 ( .A1(n4761), .A2(n4759), .ZN(n5230) );
  AOI21_X1 U5512 ( .B1(n4762), .B2(n4765), .A(n4760), .ZN(n4759) );
  XNOR2_X1 U5513 ( .A(n5168), .B(SI_7_), .ZN(n5165) );
  NAND2_X1 U5514 ( .A1(n5147), .A2(SI_6_), .ZN(n5148) );
  INV_X1 U5515 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U5516 ( .A1(n6834), .A2(n4537), .ZN(n5030) );
  NOR2_X1 U5517 ( .A1(n5038), .A2(n5028), .ZN(n4537) );
  INV_X1 U5518 ( .A(n8412), .ZN(n4896) );
  INV_X1 U5519 ( .A(n8421), .ZN(n4895) );
  NAND2_X1 U5520 ( .A1(n5352), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5373) );
  INV_X1 U5521 ( .A(n7639), .ZN(n4878) );
  AND2_X1 U5522 ( .A1(n4876), .A2(n7644), .ZN(n4875) );
  NAND2_X1 U5523 ( .A1(n7639), .A2(n4877), .ZN(n4876) );
  AND2_X1 U5524 ( .A1(n8621), .A2(n8416), .ZN(n4898) );
  NOR2_X1 U5525 ( .A1(n8253), .A2(n4900), .ZN(n4899) );
  INV_X1 U5526 ( .A(n8212), .ZN(n4900) );
  NAND3_X1 U5527 ( .A1(n7841), .A2(n7846), .A3(n7840), .ZN(n7955) );
  OR3_X1 U5528 ( .A1(n6890), .A2(n5855), .A3(n5854), .ZN(n7077) );
  AND4_X1 U5529 ( .A1(n5112), .A2(n5111), .A3(n5110), .A4(n5109), .ZN(n10342)
         );
  OR2_X1 U5530 ( .A1(n5083), .A2(n5049), .ZN(n5053) );
  OR2_X1 U5531 ( .A1(n5376), .A2(n8710), .ZN(n5017) );
  OR2_X1 U5532 ( .A1(n5389), .A2(n6895), .ZN(n5019) );
  OR2_X1 U5533 ( .A1(n5149), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5175) );
  NOR2_X1 U5534 ( .A1(n5175), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5178) );
  XNOR2_X1 U5535 ( .A(n7678), .B(n7679), .ZN(n7657) );
  OR2_X1 U5536 ( .A1(n8749), .A2(n8752), .ZN(n4555) );
  INV_X1 U5537 ( .A(n8777), .ZN(n8784) );
  NAND2_X1 U5538 ( .A1(n5521), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5557) );
  INV_X1 U5539 ( .A(n5522), .ZN(n5521) );
  AOI21_X1 U5540 ( .B1(n4847), .B2(n4849), .A(n4845), .ZN(n4844) );
  INV_X1 U5541 ( .A(n5633), .ZN(n4845) );
  OR2_X1 U5542 ( .A1(n5506), .A2(n8587), .ZN(n5522) );
  NAND2_X1 U5543 ( .A1(n8833), .A2(n5868), .ZN(n8834) );
  NAND2_X1 U5544 ( .A1(n8927), .A2(n4605), .ZN(n8871) );
  AND2_X1 U5545 ( .A1(n4427), .A2(n8872), .ZN(n4605) );
  INV_X1 U5546 ( .A(n8833), .ZN(n8853) );
  INV_X1 U5547 ( .A(n4660), .ZN(n8868) );
  INV_X1 U5548 ( .A(n4662), .ZN(n4661) );
  NAND2_X1 U5549 ( .A1(n4667), .A2(n8879), .ZN(n4663) );
  NAND2_X1 U5550 ( .A1(n8927), .A2(n4607), .ZN(n8901) );
  NAND2_X1 U5551 ( .A1(n5435), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5455) );
  INV_X1 U5552 ( .A(n5437), .ZN(n5435) );
  AND3_X1 U5553 ( .A1(n5426), .A2(n5425), .A3(n5424), .ZN(n8892) );
  AND2_X1 U5554 ( .A1(n8936), .A2(n8926), .ZN(n8927) );
  AOI21_X1 U5555 ( .B1(n4867), .B2(n4865), .A(n4864), .ZN(n4863) );
  INV_X1 U5556 ( .A(n4867), .ZN(n4866) );
  INV_X1 U5557 ( .A(n5731), .ZN(n4864) );
  NAND2_X1 U5558 ( .A1(n8976), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U5559 ( .A1(n4869), .A2(n4867), .ZN(n8941) );
  OR2_X1 U5560 ( .A1(n8987), .A2(n8960), .ZN(n8961) );
  NOR2_X1 U5561 ( .A1(n8961), .A2(n9061), .ZN(n8936) );
  AND2_X1 U5562 ( .A1(n8082), .A2(n4609), .ZN(n8988) );
  NOR2_X1 U5563 ( .A1(n9080), .A2(n4610), .ZN(n4609) );
  INV_X1 U5564 ( .A(n4611), .ZN(n4610) );
  AND2_X1 U5565 ( .A1(n5712), .A2(n5713), .ZN(n8319) );
  NAND2_X1 U5566 ( .A1(n8082), .A2(n4613), .ZN(n8260) );
  AND4_X1 U5567 ( .A1(n5313), .A2(n5312), .A3(n5311), .A4(n5310), .ZN(n8322)
         );
  AND2_X1 U5568 ( .A1(n7969), .A2(n7973), .ZN(n8082) );
  NAND2_X1 U5569 ( .A1(n8082), .A2(n9980), .ZN(n8241) );
  NAND2_X1 U5570 ( .A1(n5222), .A2(n5221), .ZN(n5237) );
  INV_X1 U5571 ( .A(n5220), .ZN(n5222) );
  INV_X1 U5572 ( .A(n7936), .ZN(n5823) );
  NOR2_X1 U5573 ( .A1(n7806), .A2(n7961), .ZN(n7969) );
  AND2_X1 U5574 ( .A1(n4838), .A2(n4439), .ZN(n7940) );
  NAND2_X1 U5575 ( .A1(n7808), .A2(n5682), .ZN(n4838) );
  AND4_X1 U5576 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n7941)
         );
  INV_X1 U5577 ( .A(n7741), .ZN(n5192) );
  AND4_X1 U5578 ( .A1(n5191), .A2(n5190), .A3(n5189), .A4(n5188), .ZN(n7646)
         );
  AND4_X1 U5579 ( .A1(n5130), .A2(n5129), .A3(n5128), .A4(n5127), .ZN(n7493)
         );
  OR2_X1 U5580 ( .A1(n4597), .A2(n8594), .ZN(n7450) );
  NAND2_X1 U5581 ( .A1(n4507), .A2(n10344), .ZN(n4597) );
  NAND2_X1 U5582 ( .A1(n4507), .A2(n10344), .ZN(n7601) );
  AND2_X1 U5583 ( .A1(n7192), .A2(n7408), .ZN(n7622) );
  NAND2_X1 U5584 ( .A1(n5811), .A2(n7191), .ZN(n7190) );
  NAND2_X1 U5585 ( .A1(n4685), .A2(n4491), .ZN(n4682) );
  NAND2_X1 U5586 ( .A1(n4681), .A2(n4491), .ZN(n4680) );
  INV_X1 U5587 ( .A(n4684), .ZN(n4681) );
  AOI21_X1 U5588 ( .B1(n4685), .B2(n8840), .A(n5530), .ZN(n4684) );
  NOR2_X1 U5589 ( .A1(n5830), .A2(n9061), .ZN(n5831) );
  NAND2_X1 U5590 ( .A1(n5007), .A2(n5006), .ZN(n5024) );
  INV_X1 U5591 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4986) );
  INV_X1 U5592 ( .A(n4854), .ZN(n4852) );
  INV_X1 U5593 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4991) );
  INV_X1 U5594 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U5595 ( .A1(n4590), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U5596 ( .A1(n4994), .A2(n4589), .ZN(n4590) );
  AND2_X1 U5597 ( .A1(n4968), .A2(n5002), .ZN(n4589) );
  NOR2_X1 U5598 ( .A1(n5366), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5368) );
  AND2_X1 U5599 ( .A1(n5326), .A2(n5302), .ZN(n7660) );
  AND2_X1 U5600 ( .A1(n5259), .A2(n5258), .ZN(n5299) );
  INV_X1 U5601 ( .A(n9285), .ZN(n4916) );
  INV_X1 U5602 ( .A(n6681), .ZN(n4927) );
  AND2_X1 U5603 ( .A1(n5942), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6300) );
  AOI21_X1 U5604 ( .B1(n4430), .B2(n4914), .A(n4428), .ZN(n4912) );
  AND2_X1 U5605 ( .A1(n6737), .A2(n6738), .ZN(n8476) );
  NAND2_X1 U5606 ( .A1(n6133), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6148) );
  AND2_X1 U5607 ( .A1(n6699), .A2(n6700), .ZN(n9210) );
  INV_X1 U5608 ( .A(n9210), .ZN(n4947) );
  OR2_X1 U5609 ( .A1(n6207), .A2(n6206), .ZN(n6226) );
  NAND2_X1 U5610 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n6300), .ZN(n6299) );
  XNOR2_X1 U5611 ( .A(n4904), .B(n6782), .ZN(n6599) );
  NAND2_X1 U5612 ( .A1(n4905), .A2(n6592), .ZN(n4904) );
  NAND2_X1 U5613 ( .A1(n9322), .A2(n6585), .ZN(n4905) );
  AND2_X1 U5614 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6030) );
  NAND2_X1 U5615 ( .A1(n7793), .A2(n7794), .ZN(n4932) );
  AND2_X1 U5616 ( .A1(n6253), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6259) );
  AND2_X1 U5617 ( .A1(n6240), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6253) );
  AOI21_X1 U5618 ( .B1(n4944), .B2(n4950), .A(n4438), .ZN(n4942) );
  NAND2_X1 U5619 ( .A1(n6030), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6045) );
  NOR2_X1 U5620 ( .A1(n6045), .A2(n7532), .ZN(n6056) );
  OR2_X1 U5621 ( .A1(n6385), .A2(n6384), .ZN(n6389) );
  NAND2_X1 U5622 ( .A1(n6368), .A2(n9551), .ZN(n6376) );
  INV_X1 U5623 ( .A(n5998), .ZN(n6273) );
  NAND2_X1 U5624 ( .A1(n7142), .A2(n4459), .ZN(n7335) );
  NAND2_X1 U5625 ( .A1(n7336), .A2(n7335), .ZN(n7334) );
  AND2_X1 U5626 ( .A1(n7334), .A2(n4546), .ZN(n7125) );
  NAND2_X1 U5627 ( .A1(n7123), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4546) );
  NAND2_X1 U5628 ( .A1(n7160), .A2(n7159), .ZN(n9720) );
  NAND2_X1 U5629 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7325) );
  OAI22_X1 U5630 ( .A1(n9720), .A2(n4543), .B1(n9718), .B2(
        P1_REG2_REG_4__SCAN_IN), .ZN(n9732) );
  INV_X1 U5631 ( .A(n9721), .ZN(n4543) );
  AND2_X1 U5632 ( .A1(n4548), .A2(n4547), .ZN(n9799) );
  NAND2_X1 U5633 ( .A1(n7252), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4547) );
  XNOR2_X1 U5634 ( .A(n7917), .B(n9807), .ZN(n9811) );
  OR2_X1 U5635 ( .A1(n8097), .A2(n8096), .ZN(n4540) );
  NAND2_X1 U5636 ( .A1(n9555), .A2(n8534), .ZN(n8522) );
  NOR2_X1 U5637 ( .A1(n8496), .A2(n9551), .ZN(n9340) );
  INV_X1 U5638 ( .A(n9345), .ZN(n9352) );
  NAND2_X1 U5639 ( .A1(n9351), .A2(n9352), .ZN(n9350) );
  AND2_X1 U5640 ( .A1(n6357), .A2(n6331), .ZN(n9348) );
  AND2_X1 U5641 ( .A1(n9409), .A2(n4478), .ZN(n9347) );
  NAND2_X1 U5642 ( .A1(n9409), .A2(n4616), .ZN(n9368) );
  NAND2_X1 U5643 ( .A1(n6469), .A2(n8522), .ZN(n9345) );
  NAND2_X1 U5644 ( .A1(n8519), .A2(n6463), .ZN(n9384) );
  AOI21_X1 U5645 ( .B1(n9450), .B2(n4457), .A(n4745), .ZN(n9398) );
  NAND2_X1 U5646 ( .A1(n4747), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U5647 ( .A1(n8515), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U5648 ( .A1(n9409), .A2(n9396), .ZN(n9391) );
  NAND2_X1 U5649 ( .A1(n4643), .A2(n8491), .ZN(n9390) );
  NAND2_X1 U5650 ( .A1(n8516), .A2(n8517), .ZN(n9397) );
  OR2_X1 U5651 ( .A1(n9581), .A2(n9256), .ZN(n9410) );
  NOR2_X1 U5652 ( .A1(n9426), .A2(n9406), .ZN(n9409) );
  NAND2_X1 U5653 ( .A1(n9449), .A2(n4749), .ZN(n9433) );
  NAND2_X1 U5654 ( .A1(n9449), .A2(n8513), .ZN(n9435) );
  NAND2_X1 U5655 ( .A1(n9450), .A2(n9451), .ZN(n9449) );
  NOR2_X1 U5656 ( .A1(n9495), .A2(n4631), .ZN(n9465) );
  INV_X1 U5657 ( .A(n4633), .ZN(n4631) );
  AND2_X1 U5658 ( .A1(n6455), .A2(n8513), .ZN(n9451) );
  INV_X1 U5659 ( .A(n4649), .ZN(n4648) );
  OR2_X1 U5660 ( .A1(n9510), .A2(n9600), .ZN(n9495) );
  NOR2_X1 U5661 ( .A1(n9529), .A2(n9610), .ZN(n9528) );
  NAND2_X1 U5662 ( .A1(n9686), .A2(n4627), .ZN(n4626) );
  NOR2_X1 U5663 ( .A1(n4628), .A2(n8303), .ZN(n4627) );
  NAND2_X1 U5664 ( .A1(n4740), .A2(n8151), .ZN(n8152) );
  AND2_X1 U5665 ( .A1(n8161), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5666 ( .A1(n4642), .A2(n8051), .ZN(n4638) );
  NAND2_X1 U5667 ( .A1(n4722), .A2(n8051), .ZN(n4641) );
  OR2_X1 U5668 ( .A1(n6148), .A2(n10166), .ZN(n6170) );
  OR2_X1 U5669 ( .A1(n6170), .A2(n6169), .ZN(n6172) );
  NOR2_X1 U5670 ( .A1(n8058), .A2(n4628), .ZN(n8181) );
  NOR2_X1 U5671 ( .A1(n8053), .A2(n4742), .ZN(n4741) );
  NOR2_X1 U5672 ( .A1(n8058), .A2(n8158), .ZN(n8179) );
  NAND2_X1 U5673 ( .A1(n4639), .A2(n8051), .ZN(n8169) );
  NAND2_X1 U5674 ( .A1(n8050), .A2(n8049), .ZN(n4639) );
  OR2_X1 U5675 ( .A1(n8015), .A2(n8207), .ZN(n8058) );
  NAND2_X1 U5676 ( .A1(n4707), .A2(n4706), .ZN(n8008) );
  AOI21_X1 U5677 ( .B1(n4437), .B2(n4711), .A(n4467), .ZN(n4706) );
  NOR2_X1 U5678 ( .A1(n4622), .A2(n4621), .ZN(n7989) );
  NAND2_X1 U5679 ( .A1(n7868), .A2(n7820), .ZN(n7992) );
  NAND2_X1 U5680 ( .A1(n4738), .A2(n4710), .ZN(n7868) );
  INV_X1 U5681 ( .A(n7714), .ZN(n4738) );
  NAND2_X1 U5682 ( .A1(n7575), .A2(n4434), .ZN(n7878) );
  NAND2_X1 U5683 ( .A1(n7575), .A2(n9861), .ZN(n7724) );
  AND2_X1 U5684 ( .A1(n7582), .A2(n7581), .ZN(n7585) );
  AND2_X1 U5685 ( .A1(n7513), .A2(n7521), .ZN(n7575) );
  NOR2_X1 U5686 ( .A1(n7547), .A2(n7504), .ZN(n7513) );
  NAND2_X1 U5687 ( .A1(n6018), .A2(n6421), .ZN(n6072) );
  OR2_X1 U5688 ( .A1(n7545), .A2(n4422), .ZN(n7547) );
  NAND2_X1 U5689 ( .A1(n7421), .A2(n7420), .ZN(n7544) );
  NAND2_X1 U5690 ( .A1(n7543), .A2(n7544), .ZN(n7542) );
  NAND2_X1 U5691 ( .A1(n7566), .A2(n7300), .ZN(n7545) );
  OAI211_X1 U5692 ( .C1(n6846), .C2(n6054), .A(n6007), .B(n6006), .ZN(n7419)
         );
  NAND2_X1 U5693 ( .A1(n6025), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6007) );
  INV_X1 U5694 ( .A(n9431), .ZN(n9537) );
  NOR2_X1 U5695 ( .A1(n8524), .A2(n4429), .ZN(n4715) );
  INV_X1 U5696 ( .A(n8499), .ZN(n9551) );
  INV_X1 U5697 ( .A(n9881), .ZN(n9872) );
  OR2_X1 U5698 ( .A1(n7302), .A2(n6483), .ZN(n9883) );
  INV_X1 U5699 ( .A(n9883), .ZN(n9873) );
  OR2_X1 U5700 ( .A1(n7302), .A2(n6552), .ZN(n9881) );
  AND2_X1 U5701 ( .A1(n7017), .A2(n7016), .ZN(n7410) );
  AND2_X1 U5702 ( .A1(n7015), .A2(n7014), .ZN(n7055) );
  XNOR2_X1 U5703 ( .A(n5578), .B(n5567), .ZN(n9164) );
  NAND2_X1 U5704 ( .A1(n4797), .A2(n5552), .ZN(n5564) );
  NAND2_X1 U5705 ( .A1(n5551), .A2(n5550), .ZN(n4797) );
  XNOR2_X1 U5706 ( .A(n5551), .B(n5550), .ZN(n8276) );
  NAND2_X1 U5707 ( .A1(n4787), .A2(n5497), .ZN(n5513) );
  NAND2_X1 U5708 ( .A1(n5483), .A2(n4788), .ZN(n4787) );
  CLKBUF_X1 U5709 ( .A(n6521), .Z(n6522) );
  NAND2_X1 U5710 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U5711 ( .A1(n4804), .A2(n5319), .ZN(n5341) );
  NAND2_X1 U5712 ( .A1(n5297), .A2(n4809), .ZN(n4804) );
  NAND2_X1 U5713 ( .A1(n5297), .A2(n5296), .ZN(n5321) );
  INV_X1 U5714 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U5715 ( .A1(n4758), .A2(n4762), .ZN(n5228) );
  OR2_X1 U5716 ( .A1(n5195), .A2(n4765), .ZN(n4758) );
  CLKBUF_X1 U5717 ( .A(n6093), .Z(n6094) );
  NAND2_X1 U5718 ( .A1(n4766), .A2(n5193), .ZN(n5208) );
  XNOR2_X1 U5719 ( .A(n5146), .B(SI_6_), .ZN(n5144) );
  AND2_X1 U5720 ( .A1(n6041), .A2(n6040), .ZN(n7177) );
  XNOR2_X1 U5721 ( .A(n5119), .B(SI_4_), .ZN(n5118) );
  NAND2_X1 U5722 ( .A1(n5095), .A2(n5093), .ZN(n4770) );
  NOR2_X2 U5723 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4906) );
  NAND2_X1 U5724 ( .A1(n5066), .A2(n4635), .ZN(n5092) );
  XNOR2_X1 U5725 ( .A(n5067), .B(SI_2_), .ZN(n4635) );
  NAND2_X1 U5726 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5990) );
  INV_X1 U5727 ( .A(n8549), .ZN(n4596) );
  NAND2_X1 U5728 ( .A1(n7841), .A2(n7840), .ZN(n7957) );
  NAND2_X1 U5729 ( .A1(n8642), .A2(n7237), .ZN(n7238) );
  NAND2_X1 U5730 ( .A1(n4879), .A2(n7478), .ZN(n7640) );
  OR2_X1 U5731 ( .A1(n7480), .A2(n7479), .ZN(n4879) );
  XNOR2_X1 U5732 ( .A(n7230), .B(n7231), .ZN(n7093) );
  AND2_X1 U5733 ( .A1(n7091), .A2(n7131), .ZN(n7094) );
  AND4_X1 U5734 ( .A1(n5242), .A2(n5241), .A3(n5240), .A4(n5239), .ZN(n8081)
         );
  INV_X1 U5735 ( .A(n9027), .ZN(n5868) );
  OR2_X1 U5736 ( .A1(n8611), .A2(n8614), .ZN(n8439) );
  NAND2_X1 U5737 ( .A1(n4503), .A2(n8396), .ZN(n8473) );
  OAI211_X1 U5738 ( .C1(n7357), .C2(n4582), .A(n8596), .B(n4580), .ZN(n8595)
         );
  NAND2_X1 U5739 ( .A1(n4583), .A2(n4584), .ZN(n8597) );
  NAND2_X1 U5740 ( .A1(n4586), .A2(n4584), .ZN(n4580) );
  NAND2_X1 U5741 ( .A1(n8473), .A2(n8400), .ZN(n8604) );
  NAND2_X1 U5742 ( .A1(n7357), .A2(n7356), .ZN(n10338) );
  AND2_X1 U5743 ( .A1(n8557), .A2(n8416), .ZN(n8620) );
  NAND2_X1 U5744 ( .A1(n8213), .A2(n8212), .ZN(n8254) );
  NAND2_X1 U5745 ( .A1(n5284), .A2(n5283), .ZN(n9092) );
  INV_X1 U5746 ( .A(n8665), .ZN(n10349) );
  AND3_X1 U5747 ( .A1(n5412), .A2(n5411), .A3(n5410), .ZN(n8658) );
  OR2_X1 U5748 ( .A1(n8637), .A2(n8979), .ZN(n10343) );
  AND2_X1 U5749 ( .A1(n4594), .A2(n8652), .ZN(n4593) );
  NAND2_X1 U5750 ( .A1(n4595), .A2(n8406), .ZN(n4594) );
  AOI21_X1 U5751 ( .B1(n4582), .B2(n8596), .A(n4581), .ZN(n4579) );
  INV_X1 U5752 ( .A(n7367), .ZN(n4581) );
  AND2_X1 U5753 ( .A1(n7098), .A2(n7086), .ZN(n8629) );
  CLKBUF_X1 U5754 ( .A(n7092), .Z(n8707) );
  OAI21_X1 U5755 ( .B1(n6909), .B2(n8710), .A(n8711), .ZN(n9665) );
  NAND2_X1 U5756 ( .A1(n9666), .A2(n9665), .ZN(n9664) );
  NAND2_X1 U5757 ( .A1(n7049), .A2(n4497), .ZN(n6961) );
  NAND2_X1 U5758 ( .A1(n6961), .A2(n6960), .ZN(n6966) );
  NOR2_X1 U5759 ( .A1(n9912), .A2(n7203), .ZN(n7205) );
  NOR2_X1 U5760 ( .A1(n7205), .A2(n7204), .ZN(n7655) );
  NAND2_X1 U5761 ( .A1(n7776), .A2(n7777), .ZN(n7779) );
  NAND2_X1 U5762 ( .A1(n7779), .A2(n7778), .ZN(n8747) );
  NOR2_X1 U5763 ( .A1(n8750), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U5764 ( .A1(n4555), .A2(n4554), .ZN(n8750) );
  NAND2_X1 U5765 ( .A1(n8749), .A2(n8752), .ZN(n4554) );
  OAI21_X1 U5766 ( .B1(n9658), .B2(n4637), .A(n8776), .ZN(n4561) );
  AOI21_X1 U5767 ( .B1(n5867), .B2(n8982), .A(n5866), .ZN(n8797) );
  AOI21_X1 U5768 ( .B1(n8805), .B2(n8982), .A(n8804), .ZN(n9017) );
  NAND2_X1 U5769 ( .A1(n4846), .A2(n5748), .ZN(n8841) );
  NAND2_X1 U5770 ( .A1(n8863), .A2(n4850), .ZN(n4846) );
  NAND2_X1 U5771 ( .A1(n8863), .A2(n5744), .ZN(n8846) );
  NAND2_X1 U5772 ( .A1(n4860), .A2(n4858), .ZN(n8881) );
  NAND2_X1 U5773 ( .A1(n5434), .A2(n5433), .ZN(n8904) );
  NAND2_X1 U5774 ( .A1(n8976), .A2(n5719), .ZN(n8952) );
  NAND2_X1 U5775 ( .A1(n4703), .A2(n4700), .ZN(n8957) );
  AND2_X1 U5776 ( .A1(n4703), .A2(n4505), .ZN(n8959) );
  NAND2_X1 U5777 ( .A1(n5351), .A2(n5350), .ZN(n8993) );
  NAND2_X1 U5778 ( .A1(n8267), .A2(n5315), .ZN(n8271) );
  NAND2_X1 U5779 ( .A1(n4694), .A2(n4697), .ZN(n8231) );
  NAND2_X1 U5780 ( .A1(n4832), .A2(n4836), .ZN(n7967) );
  NAND2_X1 U5781 ( .A1(n7808), .A2(n4837), .ZN(n4832) );
  NAND2_X1 U5782 ( .A1(n7495), .A2(n5674), .ZN(n7740) );
  NAND2_X1 U5783 ( .A1(n7599), .A2(n5815), .ZN(n7382) );
  INV_X1 U5784 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4828) );
  AND2_X1 U5785 ( .A1(n5590), .A2(n5589), .ZN(n9107) );
  NAND2_X1 U5786 ( .A1(n5520), .A2(n5519), .ZN(n9115) );
  NAND2_X1 U5787 ( .A1(n8145), .A2(n5568), .ZN(n5520) );
  NAND2_X1 U5788 ( .A1(n4683), .A2(n4685), .ZN(n8817) );
  NOR2_X1 U5789 ( .A1(n8850), .A2(n4690), .ZN(n8832) );
  OAI21_X1 U5790 ( .B1(n8907), .B2(n4666), .A(n4664), .ZN(n8878) );
  AND2_X1 U5791 ( .A1(n4668), .A2(n4670), .ZN(n8897) );
  NAND2_X1 U5792 ( .A1(n8907), .A2(n8914), .ZN(n4668) );
  NAND2_X1 U5793 ( .A1(n5403), .A2(n5402), .ZN(n9143) );
  AOI21_X1 U5794 ( .B1(n5328), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4469), .ZN(
        n4577) );
  INV_X1 U5795 ( .A(n9142), .ZN(n9152) );
  XNOR2_X1 U5796 ( .A(n5796), .B(P2_IR_REG_24__SCAN_IN), .ZN(n9949) );
  INV_X1 U5797 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U5798 ( .A1(n4588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4995) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6864) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10292) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6845) );
  INV_X1 U5802 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6852) );
  BUF_X1 U5803 ( .A(n6063), .Z(n7106) );
  NAND2_X1 U5804 ( .A1(n4956), .A2(n6754), .ZN(n9182) );
  NAND2_X1 U5805 ( .A1(n6750), .A2(n9251), .ZN(n4956) );
  OR2_X1 U5806 ( .A1(n6731), .A2(n4939), .ZN(n4938) );
  INV_X1 U5807 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5808 ( .B1(n6731), .B2(n4937), .A(n6730), .ZN(n4936) );
  INV_X1 U5809 ( .A(n4963), .ZN(n4962) );
  NAND2_X1 U5810 ( .A1(n6608), .A2(n6612), .ZN(n7519) );
  NAND2_X1 U5811 ( .A1(n4951), .A2(n9209), .ZN(n9222) );
  NAND2_X1 U5812 ( .A1(n4943), .A2(n4947), .ZN(n4951) );
  INV_X1 U5813 ( .A(n9208), .ZN(n4943) );
  OR2_X1 U5814 ( .A1(n9231), .A2(n4957), .ZN(n4954) );
  NOR2_X1 U5815 ( .A1(n9231), .A2(n4960), .ZN(n4955) );
  AND2_X1 U5816 ( .A1(n4953), .A2(n4957), .ZN(n9230) );
  INV_X1 U5817 ( .A(n9882), .ZN(n4621) );
  NAND2_X1 U5818 ( .A1(n4934), .A2(n6723), .ZN(n9241) );
  NAND2_X1 U5819 ( .A1(n9191), .A2(n9192), .ZN(n4934) );
  NAND2_X1 U5820 ( .A1(n6258), .A2(n6257), .ZN(n9595) );
  NAND2_X1 U5821 ( .A1(n6279), .A2(n6278), .ZN(n9586) );
  INV_X1 U5822 ( .A(n9301), .ZN(n9266) );
  AND2_X1 U5823 ( .A1(n6817), .A2(n4727), .ZN(n9298) );
  AOI21_X1 U5825 ( .B1(n9605), .B2(n6778), .A(n6714), .ZN(n9276) );
  NAND2_X1 U5826 ( .A1(n4963), .A2(n6612), .ZN(n7531) );
  INV_X1 U5827 ( .A(n9353), .ZN(n9381) );
  NAND2_X1 U5828 ( .A1(n5934), .A2(n5933), .ZN(n9565) );
  NAND2_X1 U5829 ( .A1(n8145), .A2(n6342), .ZN(n5934) );
  NAND2_X1 U5830 ( .A1(n6822), .A2(n6821), .ZN(n9306) );
  NAND2_X1 U5831 ( .A1(n6020), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U5832 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n7139) );
  NOR2_X1 U5833 ( .A1(n9747), .A2(n4545), .ZN(n9762) );
  AND2_X1 U5834 ( .A1(n9752), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U5835 ( .A1(n9762), .A2(n9761), .ZN(n9760) );
  AND2_X1 U5836 ( .A1(n6084), .A2(n6091), .ZN(n9769) );
  NAND2_X1 U5837 ( .A1(n9760), .A2(n4544), .ZN(n9774) );
  OR2_X1 U5838 ( .A1(n9756), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U5839 ( .A1(n9774), .A2(n9775), .ZN(n9773) );
  INV_X1 U5840 ( .A(n4548), .ZN(n7251) );
  NOR2_X1 U5841 ( .A1(n7398), .A2(n4511), .ZN(n7402) );
  NOR2_X1 U5842 ( .A1(n7402), .A2(n7401), .ZN(n7916) );
  NAND2_X1 U5843 ( .A1(n4540), .A2(n8365), .ZN(n9334) );
  AND2_X1 U5844 ( .A1(n6338), .A2(n6337), .ZN(n9679) );
  NOR2_X1 U5845 ( .A1(n9364), .A2(n9363), .ZN(n9362) );
  NAND2_X1 U5846 ( .A1(n4647), .A2(n4650), .ZN(n9494) );
  OR2_X1 U5847 ( .A1(n8484), .A2(n4652), .ZN(n4647) );
  NAND2_X1 U5848 ( .A1(n8484), .A2(n4657), .ZN(n4653) );
  AOI21_X1 U5849 ( .B1(n8484), .B2(n8500), .A(n4432), .ZN(n9527) );
  NAND2_X1 U5850 ( .A1(n8012), .A2(n8011), .ZN(n8052) );
  NAND2_X1 U5851 ( .A1(n4708), .A2(n4709), .ZN(n7988) );
  OR2_X1 U5852 ( .A1(n7723), .A2(n4711), .ZN(n4708) );
  NAND2_X1 U5853 ( .A1(n7819), .A2(n7818), .ZN(n7865) );
  NAND2_X1 U5854 ( .A1(n7506), .A2(n7505), .ZN(n7508) );
  NAND2_X1 U5855 ( .A1(n9653), .A2(n6063), .ZN(n5985) );
  AND2_X1 U5856 ( .A1(n9467), .A2(n9873), .ZN(n9545) );
  AND2_X2 U5857 ( .A1(n7055), .A2(n7410), .ZN(n9891) );
  INV_X1 U5858 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10244) );
  INV_X1 U5859 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6873) );
  INV_X1 U5860 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6866) );
  INV_X1 U5861 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6839) );
  INV_X1 U5862 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6843) );
  AOI21_X1 U5863 ( .B1(n4890), .B2(n8457), .A(n4885), .ZN(n4884) );
  INV_X1 U5864 ( .A(n4561), .ZN(n4560) );
  NAND2_X1 U5865 ( .A1(n4557), .A2(n5860), .ZN(n4556) );
  NAND2_X1 U5866 ( .A1(n8775), .A2(n8929), .ZN(n4562) );
  INV_X1 U5867 ( .A(n5913), .ZN(n5914) );
  OAI21_X1 U5868 ( .B1(n9100), .B2(n9994), .A(n4600), .ZN(P2_U3551) );
  INV_X1 U5869 ( .A(n4601), .ZN(n4600) );
  OAI22_X1 U5870 ( .A1(n9103), .A2(n9071), .B1(n9996), .B2(n9011), .ZN(n4601)
         );
  AOI21_X1 U5871 ( .B1(n8382), .B2(n9996), .A(n4826), .ZN(n8385) );
  OR2_X1 U5872 ( .A1(n8384), .A2(n4827), .ZN(n4826) );
  NOR2_X1 U5873 ( .A1(n9996), .A2(n4828), .ZN(n4827) );
  AND2_X1 U5874 ( .A1(n5871), .A2(n4965), .ZN(n5872) );
  NOR2_X1 U5875 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  AND2_X1 U5876 ( .A1(n8383), .A2(n9142), .ZN(n8379) );
  MUX2_X1 U5877 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8382), .S(n9155), .Z(n8380)
         );
  AND2_X1 U5878 ( .A1(n4910), .A2(n4907), .ZN(n8537) );
  NOR2_X1 U5879 ( .A1(n6388), .A2(n6387), .ZN(n4529) );
  NAND2_X1 U5880 ( .A1(n6386), .A2(n4492), .ZN(n4519) );
  OAI21_X1 U5881 ( .B1(n8374), .B2(n9420), .A(n4551), .ZN(n8375) );
  OAI21_X1 U5882 ( .B1(n8370), .B2(n8371), .A(n4552), .ZN(n4551) );
  OAI21_X1 U5883 ( .B1(n9554), .B2(n9547), .A(n4755), .ZN(P1_U3355) );
  AOI21_X1 U5884 ( .B1(n8528), .B2(n9477), .A(n4756), .ZN(n4755) );
  INV_X1 U5885 ( .A(n4757), .ZN(n4756) );
  AOI21_X1 U5886 ( .B1(n9552), .B2(n9545), .A(n8529), .ZN(n4757) );
  NAND2_X1 U5887 ( .A1(n4713), .A2(n4522), .ZN(P1_U3552) );
  INV_X1 U5888 ( .A(n4523), .ZN(n4522) );
  OAI21_X1 U5889 ( .B1(n9554), .B2(n4714), .A(n4508), .ZN(n4523) );
  NAND2_X1 U5890 ( .A1(n4625), .A2(n9891), .ZN(n4624) );
  INV_X1 U5891 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U5892 ( .A1(n4542), .A2(n4541), .ZN(P1_U3353) );
  NAND2_X1 U5893 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4541) );
  NAND2_X1 U5894 ( .A1(n9653), .A2(P1_U3084), .ZN(n4542) );
  OAI21_X1 U5895 ( .B1(n4425), .B2(n6384), .A(n6385), .ZN(n4818) );
  INV_X2 U5896 ( .A(n5032), .ZN(n6834) );
  AND2_X1 U5897 ( .A1(n9679), .A2(n9312), .ZN(n4425) );
  OR2_X1 U5898 ( .A1(n9581), .A2(n9452), .ZN(n4426) );
  AND2_X1 U5899 ( .A1(n4607), .A2(n4606), .ZN(n4427) );
  AND2_X1 U5900 ( .A1(n4919), .A2(n4918), .ZN(n4428) );
  AND2_X1 U5901 ( .A1(n9555), .A2(n9367), .ZN(n4429) );
  INV_X1 U5902 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6127) );
  AND2_X1 U5903 ( .A1(n4471), .A2(n4917), .ZN(n4430) );
  NOR2_X1 U5904 ( .A1(n7793), .A2(n7794), .ZN(n4431) );
  AND2_X1 U5905 ( .A1(n9617), .A2(n9538), .ZN(n4432) );
  INV_X1 U5906 ( .A(n7838), .ZN(n4873) );
  AND2_X1 U5907 ( .A1(n4833), .A2(n7966), .ZN(n4433) );
  NAND2_X1 U5908 ( .A1(n5485), .A2(n5484), .ZN(n8858) );
  AND2_X1 U5909 ( .A1(n9861), .A2(n9867), .ZN(n4434) );
  OR2_X1 U5910 ( .A1(n9561), .A2(n9381), .ZN(n8521) );
  AND2_X1 U5911 ( .A1(n9600), .A2(n9521), .ZN(n4435) );
  OR2_X1 U5912 ( .A1(n7961), .A2(n7859), .ZN(n5689) );
  INV_X1 U5913 ( .A(n8011), .ZN(n4742) );
  AND2_X1 U5914 ( .A1(n4709), .A2(n4462), .ZN(n4437) );
  NAND2_X1 U5915 ( .A1(n4720), .A2(n8488), .ZN(n9424) );
  XOR2_X1 U5916 ( .A(n6713), .B(n7510), .Z(n4438) );
  NAND2_X1 U5917 ( .A1(n9501), .A2(n8509), .ZN(n9481) );
  NAND2_X1 U5918 ( .A1(n9929), .A2(n7941), .ZN(n4439) );
  INV_X1 U5919 ( .A(n8840), .ZN(n4688) );
  AND2_X1 U5920 ( .A1(n5633), .A2(n5639), .ZN(n8840) );
  AND2_X1 U5921 ( .A1(n9285), .A2(n4914), .ZN(n4440) );
  XNOR2_X1 U5922 ( .A(n8453), .B(n7408), .ZN(n7230) );
  AND2_X1 U5923 ( .A1(n4434), .A2(n4620), .ZN(n4441) );
  NAND2_X1 U5924 ( .A1(n4796), .A2(n4795), .ZN(n5578) );
  AND2_X1 U5925 ( .A1(n6346), .A2(n6345), .ZN(n9550) );
  AND2_X1 U5926 ( .A1(n4682), .A2(n8806), .ZN(n4442) );
  AND2_X1 U5927 ( .A1(n9049), .A2(n8924), .ZN(n5835) );
  INV_X1 U5928 ( .A(n8877), .ZN(n8879) );
  AND2_X1 U5929 ( .A1(n5740), .A2(n5727), .ZN(n8877) );
  NAND2_X1 U5930 ( .A1(n6290), .A2(n6289), .ZN(n9406) );
  INV_X1 U5931 ( .A(n4686), .ZN(n4685) );
  OAI21_X1 U5932 ( .B1(n8840), .B2(n4687), .A(n4689), .ZN(n4686) );
  NAND2_X1 U5933 ( .A1(n6252), .A2(n6251), .ZN(n9600) );
  INV_X1 U5934 ( .A(n4493), .ZN(n4918) );
  AND2_X1 U5935 ( .A1(n4680), .A2(n8806), .ZN(n4443) );
  AND2_X1 U5936 ( .A1(n5192), .A2(n5674), .ZN(n4444) );
  INV_X1 U5937 ( .A(n7466), .ZN(n9477) );
  INV_X1 U5938 ( .A(n8958), .ZN(n4702) );
  INV_X1 U5939 ( .A(n8893), .ZN(n4669) );
  INV_X1 U5940 ( .A(n9131), .ZN(n4606) );
  INV_X1 U5941 ( .A(n9555), .ZN(n4615) );
  AND2_X1 U5942 ( .A1(n8451), .A2(n8450), .ZN(n4445) );
  AND4_X1 U5943 ( .A1(n6335), .A2(n6334), .A3(n6333), .A4(n6332), .ZN(n8534)
         );
  AND2_X1 U5944 ( .A1(n6389), .A2(n6483), .ZN(n4446) );
  NAND2_X1 U5945 ( .A1(n5660), .A2(n4455), .ZN(n7316) );
  INV_X1 U5946 ( .A(n6025), .ZN(n6062) );
  NAND2_X1 U5947 ( .A1(n8705), .A2(n9962), .ZN(n4672) );
  OR2_X1 U5948 ( .A1(n8058), .A2(n4626), .ZN(n4447) );
  OR2_X1 U5949 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4448) );
  AND2_X1 U5950 ( .A1(n6628), .A2(n4932), .ZN(n4449) );
  OR3_X1 U5951 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .A3(
        P1_IR_REG_27__SCAN_IN), .ZN(n4450) );
  OR2_X1 U5952 ( .A1(n4878), .A2(n7479), .ZN(n4451) );
  AND3_X1 U5953 ( .A1(n6021), .A2(n6024), .A3(n6022), .ZN(n4452) );
  NAND2_X1 U5954 ( .A1(n6715), .A2(n9275), .ZN(n9191) );
  AND2_X1 U5955 ( .A1(n6893), .A2(n5032), .ZN(n5117) );
  INV_X1 U5956 ( .A(n5117), .ZN(n5419) );
  AND2_X1 U5957 ( .A1(n5098), .A2(n4991), .ZN(n5100) );
  NAND2_X1 U5958 ( .A1(n5542), .A2(n5541), .ZN(n8814) );
  NOR2_X1 U5959 ( .A1(n6218), .A2(n5965), .ZN(n5972) );
  AND2_X1 U5960 ( .A1(n4990), .A2(n4989), .ZN(n5098) );
  OR2_X1 U5961 ( .A1(n6522), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4453) );
  AND3_X1 U5962 ( .A1(n8840), .A2(n5751), .A3(n5750), .ZN(n4454) );
  INV_X1 U5963 ( .A(n7440), .ZN(n8594) );
  AND2_X1 U5964 ( .A1(n5122), .A2(n4577), .ZN(n7440) );
  AND3_X1 U5965 ( .A1(n5653), .A2(n5648), .A3(n4672), .ZN(n4455) );
  NOR2_X1 U5966 ( .A1(n5759), .A2(n5761), .ZN(n4456) );
  NAND2_X1 U5967 ( .A1(n6298), .A2(n6297), .ZN(n9581) );
  AND2_X1 U5968 ( .A1(n8515), .A2(n9451), .ZN(n4457) );
  NAND2_X1 U5969 ( .A1(n6005), .A2(n4906), .ZN(n6026) );
  NOR2_X1 U5970 ( .A1(n9134), .A2(n8633), .ZN(n4458) );
  INV_X1 U5971 ( .A(n4658), .ZN(n4657) );
  OAI21_X1 U5972 ( .B1(n8500), .B2(n4432), .A(n4460), .ZN(n4658) );
  NAND2_X1 U5973 ( .A1(n5977), .A2(n5976), .ZN(n9561) );
  NAND2_X1 U5974 ( .A1(n5330), .A2(n5329), .ZN(n9080) );
  NAND2_X1 U5975 ( .A1(n6268), .A2(n6267), .ZN(n9592) );
  NAND2_X1 U5976 ( .A1(n5421), .A2(n5420), .ZN(n9049) );
  OR2_X1 U5977 ( .A1(n7147), .A2(n7122), .ZN(n4459) );
  NAND2_X1 U5978 ( .A1(n5262), .A2(n5261), .ZN(n8087) );
  INV_X1 U5979 ( .A(n9570), .ZN(n9396) );
  NAND2_X1 U5980 ( .A1(n5936), .A2(n5935), .ZN(n9570) );
  NAND2_X1 U5981 ( .A1(n9409), .A2(n4618), .ZN(n4619) );
  OR2_X1 U5982 ( .A1(n9610), .A2(n9522), .ZN(n4460) );
  AND2_X1 U5983 ( .A1(n5192), .A2(n5687), .ZN(n4461) );
  NAND2_X1 U5984 ( .A1(n7987), .A2(n7995), .ZN(n4462) );
  INV_X1 U5985 ( .A(n4950), .ZN(n4948) );
  NAND2_X1 U5986 ( .A1(n4512), .A2(n9209), .ZN(n4950) );
  AND2_X1 U5987 ( .A1(n9406), .A2(n8490), .ZN(n8514) );
  INV_X1 U5988 ( .A(n8514), .ZN(n4746) );
  AND2_X1 U5989 ( .A1(n9871), .A2(n9318), .ZN(n4463) );
  OR2_X1 U5990 ( .A1(n4652), .A2(n4435), .ZN(n4464) );
  NAND2_X1 U5991 ( .A1(n5635), .A2(n8799), .ZN(n8820) );
  AND2_X1 U5992 ( .A1(n8153), .A2(n8151), .ZN(n4465) );
  OR2_X1 U5993 ( .A1(n9565), .A2(n9361), .ZN(n8519) );
  INV_X1 U5994 ( .A(n5895), .ZN(n5887) );
  AND2_X1 U5995 ( .A1(n5765), .A2(n5766), .ZN(n5895) );
  NAND2_X1 U5996 ( .A1(n5570), .A2(n5569), .ZN(n8383) );
  NAND2_X1 U5997 ( .A1(n4860), .A2(n5737), .ZN(n4466) );
  NOR2_X1 U5998 ( .A1(n7987), .A2(n7995), .ZN(n4467) );
  OR2_X1 U5999 ( .A1(n4919), .A2(n4918), .ZN(n4468) );
  NAND2_X1 U6000 ( .A1(n5032), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4729) );
  AND2_X1 U6001 ( .A1(n5401), .A2(n8724), .ZN(n4469) );
  INV_X1 U6002 ( .A(n4960), .ZN(n4959) );
  NOR2_X1 U6003 ( .A1(n4961), .A2(n9183), .ZN(n4960) );
  NAND3_X1 U6004 ( .A1(n6750), .A2(n9251), .A3(n4961), .ZN(n4470) );
  INV_X1 U6005 ( .A(n4667), .ZN(n4666) );
  NOR2_X1 U6006 ( .A1(n4458), .A2(n5835), .ZN(n4667) );
  AND2_X1 U6007 ( .A1(n4919), .A2(n9285), .ZN(n4471) );
  OR2_X1 U6008 ( .A1(n9600), .A2(n9521), .ZN(n4472) );
  INV_X1 U6009 ( .A(n4925), .ZN(n4924) );
  OR2_X1 U6010 ( .A1(n8133), .A2(n4926), .ZN(n4925) );
  NAND2_X1 U6011 ( .A1(n4862), .A2(n5740), .ZN(n4473) );
  NAND2_X1 U6012 ( .A1(n7935), .A2(n4439), .ZN(n4474) );
  INV_X1 U6013 ( .A(n4859), .ZN(n4858) );
  NAND2_X1 U6014 ( .A1(n8877), .A2(n5737), .ZN(n4859) );
  INV_X1 U6015 ( .A(n8049), .ZN(n4722) );
  AND2_X1 U6016 ( .A1(n4771), .A2(n4770), .ZN(n4475) );
  NAND2_X1 U6017 ( .A1(n6168), .A2(n6167), .ZN(n8183) );
  AND2_X1 U6018 ( .A1(n8524), .A2(n4429), .ZN(n4476) );
  AND2_X1 U6019 ( .A1(n6316), .A2(n7007), .ZN(n4477) );
  AND2_X1 U6020 ( .A1(n4616), .A2(n4615), .ZN(n4478) );
  AND2_X1 U6021 ( .A1(n4856), .A2(n4855), .ZN(n4479) );
  AND2_X1 U6022 ( .A1(n4673), .A2(n4672), .ZN(n4480) );
  AND2_X1 U6023 ( .A1(n6419), .A2(n6397), .ZN(n4481) );
  INV_X1 U6024 ( .A(n7820), .ZN(n4737) );
  AND2_X1 U6025 ( .A1(n6392), .A2(n8509), .ZN(n4482) );
  OR2_X1 U6026 ( .A1(n9448), .A2(n9432), .ZN(n4483) );
  AND2_X1 U6027 ( .A1(n4830), .A2(n5272), .ZN(n4484) );
  AND2_X1 U6028 ( .A1(n8509), .A2(n6449), .ZN(n4485) );
  AND2_X1 U6029 ( .A1(n8468), .A2(n8406), .ZN(n4486) );
  AND2_X1 U6030 ( .A1(n7240), .A2(n7237), .ZN(n4487) );
  INV_X1 U6031 ( .A(n4980), .ZN(n4642) );
  NOR2_X1 U6032 ( .A1(n8160), .A2(n8159), .ZN(n4980) );
  AND2_X1 U6033 ( .A1(n5001), .A2(n4903), .ZN(n4488) );
  INV_X1 U6034 ( .A(n9036), .ZN(n8872) );
  NAND2_X1 U6035 ( .A1(n5471), .A2(n5470), .ZN(n9036) );
  OR2_X1 U6036 ( .A1(n9534), .A2(n9216), .ZN(n4489) );
  AND2_X1 U6037 ( .A1(n4946), .A2(n4945), .ZN(n4944) );
  INV_X1 U6038 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U6039 ( .A1(n8557), .A2(n4898), .ZN(n8567) );
  INV_X1 U6040 ( .A(n5007), .ZN(n5797) );
  AND2_X1 U6041 ( .A1(n8927), .A2(n8911), .ZN(n4490) );
  NAND2_X1 U6042 ( .A1(n5836), .A2(n8802), .ZN(n4491) );
  INV_X1 U6043 ( .A(n8806), .ZN(n8800) );
  NAND2_X1 U6044 ( .A1(n5754), .A2(n5755), .ZN(n8806) );
  NAND2_X1 U6045 ( .A1(n5454), .A2(n5453), .ZN(n9131) );
  NAND2_X1 U6046 ( .A1(n7722), .A2(n7723), .ZN(n7819) );
  NAND2_X1 U6047 ( .A1(n8110), .A2(n6668), .ZN(n8132) );
  NAND2_X1 U6048 ( .A1(n4653), .A2(n4656), .ZN(n9509) );
  NAND2_X1 U6049 ( .A1(n8200), .A2(n6664), .ZN(n8110) );
  AND2_X1 U6050 ( .A1(n4446), .A2(n7931), .ZN(n4492) );
  OR2_X1 U6051 ( .A1(n6767), .A2(n6766), .ZN(n4920) );
  INV_X1 U6052 ( .A(n4920), .ZN(n4914) );
  NOR3_X1 U6053 ( .A1(n9495), .A2(n9581), .A3(n4632), .ZN(n4629) );
  NAND2_X1 U6054 ( .A1(n6108), .A2(n5920), .ZN(n6140) );
  OR2_X1 U6055 ( .A1(n6771), .A2(n6770), .ZN(n4493) );
  AND2_X1 U6056 ( .A1(n4869), .A2(n5641), .ZN(n4494) );
  AND2_X1 U6057 ( .A1(n5493), .A2(n5492), .ZN(n8690) );
  INV_X1 U6058 ( .A(n8690), .ZN(n4691) );
  AND2_X1 U6059 ( .A1(n5829), .A2(n8980), .ZN(n4495) );
  INV_X1 U6060 ( .A(n4630), .ZN(n9444) );
  NOR2_X1 U6061 ( .A1(n9495), .A2(n4632), .ZN(n4630) );
  AND2_X1 U6062 ( .A1(n9134), .A2(n8633), .ZN(n4496) );
  OR2_X1 U6063 ( .A1(n6959), .A2(n6958), .ZN(n4497) );
  AND2_X1 U6064 ( .A1(n9581), .A2(n9452), .ZN(n4498) );
  AND2_X1 U6065 ( .A1(n9551), .A2(n9872), .ZN(n4499) );
  NAND2_X1 U6066 ( .A1(n6325), .A2(n6324), .ZN(n9555) );
  NAND2_X1 U6067 ( .A1(n8927), .A2(n4427), .ZN(n4608) );
  AND2_X1 U6068 ( .A1(n5397), .A2(SI_18_), .ZN(n4500) );
  AND2_X1 U6069 ( .A1(n4778), .A2(n4775), .ZN(n4501) );
  OR2_X1 U6070 ( .A1(n9131), .A2(n4669), .ZN(n4502) );
  AND2_X1 U6071 ( .A1(n8672), .A2(n8468), .ZN(n4503) );
  AND2_X1 U6072 ( .A1(n4776), .A2(n4775), .ZN(n4504) );
  NAND2_X1 U6073 ( .A1(n8993), .A2(n8692), .ZN(n4505) );
  INV_X1 U6074 ( .A(n5835), .ZN(n4670) );
  AND2_X1 U6075 ( .A1(n7413), .A2(n9489), .ZN(n7466) );
  INV_X1 U6076 ( .A(n7804), .ZN(n4704) );
  OR2_X1 U6077 ( .A1(n5512), .A2(n4786), .ZN(n4506) );
  NOR2_X1 U6078 ( .A1(n4823), .A2(n9958), .ZN(n4507) );
  OR2_X1 U6079 ( .A1(n9903), .A2(n4718), .ZN(n4508) );
  OAI21_X1 U6080 ( .B1(n7480), .B2(n4451), .A(n4875), .ZN(n7837) );
  NAND2_X1 U6081 ( .A1(n6629), .A2(n6628), .ZN(n7792) );
  NAND2_X1 U6082 ( .A1(n6553), .A2(n9420), .ZN(n7007) );
  NAND2_X1 U6083 ( .A1(n7506), .A2(n4721), .ZN(n7582) );
  OR3_X1 U6084 ( .A1(n8058), .A2(n9179), .A3(n4628), .ZN(n4509) );
  AND2_X1 U6085 ( .A1(n6612), .A2(n4962), .ZN(n4510) );
  AND2_X1 U6086 ( .A1(n7399), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U6087 ( .A1(n8082), .A2(n4611), .ZN(n4614) );
  NAND2_X1 U6088 ( .A1(n6710), .A2(n6709), .ZN(n4512) );
  AND2_X1 U6089 ( .A1(n5566), .A2(n5565), .ZN(n4513) );
  OR2_X1 U6090 ( .A1(n9891), .A2(n4623), .ZN(n4514) );
  AOI21_X1 U6091 ( .B1(n6629), .B2(n4449), .A(n4431), .ZN(n4929) );
  INV_X1 U6092 ( .A(n6535), .ZN(n4727) );
  INV_X1 U6093 ( .A(n9542), .ZN(n9484) );
  INV_X1 U6094 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4754) );
  INV_X1 U6095 ( .A(n9871), .ZN(n4620) );
  AND2_X1 U6096 ( .A1(n7359), .A2(n7358), .ZN(n4515) );
  INV_X1 U6097 ( .A(n4586), .ZN(n4585) );
  NAND2_X1 U6098 ( .A1(n4587), .A2(n7356), .ZN(n4586) );
  AND2_X1 U6099 ( .A1(n5660), .A2(n4672), .ZN(n4516) );
  NAND2_X1 U6100 ( .A1(n4517), .A2(n6451), .ZN(n6265) );
  NAND2_X1 U6101 ( .A1(n6264), .A2(n4485), .ZN(n4517) );
  MUX2_X1 U6102 ( .A(n6125), .B(n6124), .S(n7007), .Z(n6139) );
  OAI211_X1 U6103 ( .C1(n6121), .C2(n6120), .A(n7993), .B(n6401), .ZN(n6123)
         );
  NAND4_X1 U6104 ( .A1(n4518), .A2(n5989), .A3(n5987), .A4(n5988), .ZN(n6558)
         );
  NAND2_X1 U6105 ( .A1(n6044), .A2(n4481), .ZN(n6055) );
  OAI21_X1 U6106 ( .B1(n4519), .B2(n4529), .A(n4790), .ZN(P1_U3240) );
  NAND2_X1 U6107 ( .A1(n6263), .A2(n4482), .ZN(n6266) );
  AOI211_X2 U6108 ( .C1(n6307), .C2(n8515), .A(n6484), .B(n6462), .ZN(n6318)
         );
  AND3_X1 U6109 ( .A1(n6009), .A2(n6010), .A3(n6008), .ZN(n4534) );
  AOI211_X2 U6110 ( .C1(n9539), .C2(n9367), .A(n9366), .B(n9365), .ZN(n9563)
         );
  NAND2_X1 U6111 ( .A1(n7994), .A2(n7993), .ZN(n8010) );
  NAND2_X1 U6112 ( .A1(n8150), .A2(n8149), .ZN(n8175) );
  OAI21_X1 U6113 ( .B1(n8307), .B2(n8306), .A(n8305), .ZN(n8502) );
  AOI21_X1 U6114 ( .B1(n8508), .B2(n6431), .A(n8507), .ZN(n9502) );
  NAND2_X1 U6115 ( .A1(n7151), .A2(n7153), .ZN(n7152) );
  NAND2_X1 U6116 ( .A1(n6552), .A2(n6553), .ZN(n4520) );
  NAND2_X1 U6117 ( .A1(n9260), .A2(n9263), .ZN(n9261) );
  XNOR2_X2 U6118 ( .A(n6480), .B(n6479), .ZN(n4794) );
  NAND2_X1 U6119 ( .A1(n5059), .A2(n5058), .ZN(n5066) );
  XNOR2_X2 U6120 ( .A(n5208), .B(n4975), .ZN(n6872) );
  NAND2_X1 U6121 ( .A1(n4740), .A2(n4465), .ZN(n8284) );
  OAI21_X2 U6122 ( .B1(n7293), .B2(n7292), .A(n6492), .ZN(n7538) );
  NAND2_X1 U6123 ( .A1(n6318), .A2(n6371), .ZN(n4528) );
  INV_X1 U6124 ( .A(n7584), .ZN(n7583) );
  NOR2_X1 U6125 ( .A1(n6309), .A2(n6308), .ZN(n6313) );
  NAND3_X1 U6126 ( .A1(n6005), .A2(n4906), .A3(n5916), .ZN(n6036) );
  INV_X1 U6127 ( .A(n9424), .ZN(n4645) );
  NAND2_X1 U6128 ( .A1(n9404), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U6129 ( .A1(n4624), .A2(n4514), .ZN(P1_U3520) );
  AOI22_X1 U6130 ( .A1(n9359), .A2(n9363), .B1(n9381), .B2(n9360), .ZN(n9346)
         );
  MUX2_X1 U6131 ( .A(n6835), .B(n6847), .S(n5032), .Z(n5067) );
  AND2_X2 U6132 ( .A1(n4819), .A2(n4820), .ZN(n5032) );
  INV_X1 U6133 ( .A(n4646), .ZN(n9474) );
  NAND2_X1 U6134 ( .A1(n9443), .A2(n4483), .ZN(n4720) );
  XNOR2_X2 U6135 ( .A(n5938), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9646) );
  OAI21_X2 U6136 ( .B1(n6072), .B2(n6420), .A(n6423), .ZN(n7711) );
  NAND2_X1 U6137 ( .A1(n6355), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4535) );
  NAND2_X1 U6138 ( .A1(n6264), .A2(n4536), .ZN(n6263) );
  NAND2_X1 U6139 ( .A1(n6249), .A2(n6248), .ZN(n6264) );
  OAI21_X1 U6140 ( .B1(n5786), .B2(n4570), .A(n5793), .ZN(n5809) );
  INV_X1 U6141 ( .A(n8528), .ZN(n9553) );
  INV_X1 U6142 ( .A(n5794), .ZN(n4572) );
  XNOR2_X2 U6143 ( .A(n5321), .B(n5316), .ZN(n7004) );
  AOI21_X1 U6144 ( .B1(n6315), .B2(n6461), .A(n6314), .ZN(n6317) );
  NAND4_X1 U6145 ( .A1(n5917), .A2(n6064), .A3(n6038), .A4(n6081), .ZN(n5918)
         );
  AND2_X1 U6146 ( .A1(n6583), .A2(n6584), .ZN(n9263) );
  NAND2_X2 U6147 ( .A1(n7218), .A2(n7219), .ZN(n7274) );
  NAND2_X1 U6148 ( .A1(n9170), .A2(n9172), .ZN(n6689) );
  NAND2_X1 U6149 ( .A1(n4910), .A2(n4912), .ZN(n8530) );
  INV_X1 U6150 ( .A(n9201), .ZN(n4911) );
  NAND2_X1 U6151 ( .A1(n9208), .A2(n4948), .ZN(n4941) );
  INV_X1 U6152 ( .A(n5094), .ZN(n5095) );
  NOR2_X2 U6153 ( .A1(n6036), .A2(n5918), .ZN(n6093) );
  MUX2_X2 U6154 ( .A(n6266), .B(n6265), .S(n7007), .Z(n6309) );
  MUX2_X2 U6155 ( .A(n6090), .B(n6089), .S(n6371), .Z(n6121) );
  NAND2_X2 U6156 ( .A1(n6492), .A2(n6497), .ZN(n7292) );
  INV_X1 U6157 ( .A(n4540), .ZN(n8364) );
  NOR2_X1 U6158 ( .A1(n8094), .A2(n8095), .ZN(n8097) );
  NAND3_X1 U6159 ( .A1(n4562), .A2(n4560), .A3(n4556), .ZN(P2_U3264) );
  AND4_X2 U6160 ( .A1(n4853), .A2(n4992), .A3(n4969), .A4(n5100), .ZN(n5007)
         );
  NAND2_X1 U6161 ( .A1(n5783), .A2(n7733), .ZN(n5785) );
  NAND3_X1 U6162 ( .A1(n7357), .A2(n8596), .A3(n4585), .ZN(n4578) );
  NAND2_X1 U6163 ( .A1(n4579), .A2(n4578), .ZN(n7368) );
  INV_X1 U6164 ( .A(n10336), .ZN(n4587) );
  NAND2_X1 U6165 ( .A1(n8343), .A2(n7803), .ZN(n7102) );
  NAND2_X1 U6166 ( .A1(n4994), .A2(n4968), .ZN(n4588) );
  NAND2_X1 U6167 ( .A1(n7093), .A2(n7094), .ZN(n8646) );
  NAND3_X1 U6168 ( .A1(n8396), .A2(n8672), .A3(n4486), .ZN(n4592) );
  NAND2_X1 U6169 ( .A1(n4592), .A2(n4593), .ZN(n8556) );
  NAND3_X1 U6170 ( .A1(n10344), .A2(n4599), .A3(n7436), .ZN(n4598) );
  NAND2_X1 U6171 ( .A1(n8826), .A2(n4602), .ZN(n8777) );
  INV_X1 U6172 ( .A(n4608), .ZN(n8883) );
  INV_X1 U6173 ( .A(n4614), .ZN(n8323) );
  INV_X1 U6174 ( .A(n4619), .ZN(n9376) );
  INV_X1 U6175 ( .A(n4622), .ZN(n7877) );
  INV_X1 U6176 ( .A(n4629), .ZN(n9426) );
  INV_X1 U6177 ( .A(n7419), .ZN(n7566) );
  NAND2_X1 U6178 ( .A1(n5167), .A2(n5166), .ZN(n5170) );
  NAND2_X1 U6179 ( .A1(n5145), .A2(n5144), .ZN(n4634) );
  XNOR2_X1 U6180 ( .A(n5066), .B(n4635), .ZN(n6846) );
  NAND3_X1 U6181 ( .A1(n8376), .A2(n4637), .A3(n4636), .ZN(n4819) );
  OAI22_X1 U6182 ( .A1(n8050), .A2(n4638), .B1(n4640), .B2(n4980), .ZN(n8281)
         );
  AOI21_X2 U6183 ( .B1(n4645), .B2(n4426), .A(n4498), .ZN(n9404) );
  OAI21_X1 U6184 ( .B1(n4464), .B2(n8484), .A(n4648), .ZN(n4646) );
  OAI21_X1 U6185 ( .B1(n8907), .B2(n4663), .A(n4661), .ZN(n4660) );
  AND2_X1 U6186 ( .A1(n4973), .A2(n4672), .ZN(n7615) );
  NAND2_X1 U6187 ( .A1(n4671), .A2(n4672), .ZN(n5666) );
  NAND2_X1 U6188 ( .A1(n7599), .A2(n4674), .ZN(n4676) );
  NAND2_X1 U6189 ( .A1(n7453), .A2(n5818), .ZN(n5820) );
  OAI21_X1 U6190 ( .B1(n8850), .B2(n4682), .A(n4680), .ZN(n8807) );
  NAND2_X1 U6191 ( .A1(n8850), .A2(n4443), .ZN(n4679) );
  NAND2_X1 U6192 ( .A1(n8850), .A2(n4688), .ZN(n4683) );
  NAND2_X1 U6193 ( .A1(n4694), .A2(n4692), .ZN(n8233) );
  NAND2_X1 U6194 ( .A1(n5826), .A2(n5825), .ZN(n8076) );
  INV_X1 U6195 ( .A(n5825), .ZN(n4696) );
  OR2_X1 U6196 ( .A1(n8087), .A2(n8696), .ZN(n4697) );
  NAND2_X1 U6197 ( .A1(n8969), .A2(n4700), .ZN(n4698) );
  NAND2_X1 U6198 ( .A1(n4698), .A2(n4699), .ZN(n8935) );
  INV_X1 U6199 ( .A(n4703), .ZN(n8971) );
  OAI21_X1 U6200 ( .B1(n7805), .B2(n4704), .A(n5822), .ZN(n7936) );
  NAND2_X1 U6201 ( .A1(n7289), .A2(n7292), .ZN(n7421) );
  AOI21_X2 U6202 ( .B1(n9375), .B2(n8493), .A(n4705), .ZN(n9359) );
  NAND2_X1 U6203 ( .A1(n7723), .A2(n4437), .ZN(n4707) );
  AOI21_X1 U6204 ( .B1(n9344), .B2(n4715), .A(n4476), .ZN(n4712) );
  INV_X1 U6205 ( .A(n6841), .ZN(n4724) );
  NAND3_X1 U6206 ( .A1(n8348), .A2(n6535), .A3(n7121), .ZN(n4725) );
  AND2_X2 U6207 ( .A1(n6093), .A2(n5919), .ZN(n6108) );
  AOI21_X1 U6208 ( .B1(n9458), .B2(n9457), .A(n8487), .ZN(n9443) );
  NAND2_X1 U6209 ( .A1(n7585), .A2(n7584), .ZN(n7721) );
  NAND2_X1 U6210 ( .A1(n7423), .A2(n7424), .ZN(n7506) );
  NAND2_X1 U6211 ( .A1(n7456), .A2(n5996), .ZN(n6396) );
  AOI21_X1 U6212 ( .B1(n8935), .B2(n5832), .A(n5831), .ZN(n8920) );
  INV_X1 U6213 ( .A(n7317), .ZN(n7312) );
  OAI22_X1 U6214 ( .A1(n7487), .A2(n5163), .B1(n7632), .B2(n8701), .ZN(n7737)
         );
  NAND2_X1 U6215 ( .A1(n7934), .A2(n5824), .ZN(n7963) );
  OR2_X1 U6216 ( .A1(n8705), .A2(n9962), .ZN(n4973) );
  NAND2_X1 U6217 ( .A1(n5820), .A2(n5819), .ZN(n7487) );
  NAND2_X1 U6218 ( .A1(n6529), .A2(n5929), .ZN(n5930) );
  AOI21_X1 U6219 ( .B1(n7460), .B2(n7456), .A(n7288), .ZN(n7289) );
  INV_X1 U6220 ( .A(n4732), .ZN(n4733) );
  OR2_X1 U6221 ( .A1(n6558), .A2(n7022), .ZN(n4732) );
  NAND2_X1 U6222 ( .A1(n4732), .A2(n6489), .ZN(n7018) );
  NAND2_X1 U6223 ( .A1(n4732), .A2(n6396), .ZN(n5997) );
  XNOR2_X1 U6224 ( .A(n7286), .B(n4733), .ZN(n7464) );
  NAND2_X1 U6225 ( .A1(n4736), .A2(n4734), .ZN(n7994) );
  INV_X1 U6226 ( .A(n4735), .ZN(n4734) );
  NAND2_X1 U6227 ( .A1(n7714), .A2(n7820), .ZN(n4736) );
  NAND2_X1 U6228 ( .A1(n8012), .A2(n4741), .ZN(n8148) );
  NAND2_X1 U6229 ( .A1(n8148), .A2(n8147), .ZN(n8150) );
  NOR2_X1 U6230 ( .A1(n9382), .A2(n8520), .ZN(n9364) );
  INV_X1 U6231 ( .A(n6521), .ZN(n4751) );
  NAND2_X1 U6232 ( .A1(n4751), .A2(n4752), .ZN(n5937) );
  NOR2_X1 U6233 ( .A1(n6521), .A2(n4436), .ZN(n5927) );
  NAND2_X1 U6234 ( .A1(n5195), .A2(n4762), .ZN(n4761) );
  NAND2_X1 U6235 ( .A1(n5092), .A2(n5091), .ZN(n4771) );
  NAND2_X1 U6236 ( .A1(n4769), .A2(n5121), .ZN(n5132) );
  NAND3_X1 U6237 ( .A1(n4771), .A2(n4770), .A3(n5118), .ZN(n4769) );
  NAND2_X1 U6238 ( .A1(n5385), .A2(n4504), .ZN(n4774) );
  NAND2_X1 U6239 ( .A1(n5483), .A2(n4784), .ZN(n4783) );
  NAND2_X1 U6240 ( .A1(n5483), .A2(n5482), .ZN(n5499) );
  NOR2_X1 U6241 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U6242 ( .A1(n5551), .A2(n4798), .ZN(n4796) );
  NAND2_X1 U6243 ( .A1(n5297), .A2(n4805), .ZN(n4801) );
  NAND2_X1 U6244 ( .A1(n4801), .A2(n4802), .ZN(n5365) );
  NAND2_X1 U6245 ( .A1(n5444), .A2(n4814), .ZN(n4811) );
  NAND2_X1 U6246 ( .A1(n4811), .A2(n4812), .ZN(n5481) );
  INV_X1 U6247 ( .A(n6372), .ZN(n4817) );
  NAND3_X1 U6248 ( .A1(n4821), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U6249 ( .A1(n7316), .A2(n5653), .ZN(n7606) );
  AND2_X1 U6250 ( .A1(n5653), .A2(n5648), .ZN(n7317) );
  NAND2_X1 U6251 ( .A1(n5902), .A2(n8982), .ZN(n4825) );
  NAND2_X1 U6252 ( .A1(n4831), .A2(n4484), .ZN(n5273) );
  NAND2_X1 U6253 ( .A1(n7808), .A2(n4433), .ZN(n4831) );
  OAI21_X1 U6254 ( .B1(n7808), .B2(n4835), .A(n4433), .ZN(n7965) );
  NAND2_X1 U6255 ( .A1(n8234), .A2(n5315), .ZN(n4839) );
  NAND2_X1 U6256 ( .A1(n8863), .A2(n4847), .ZN(n4843) );
  NAND2_X1 U6257 ( .A1(n4843), .A2(n4844), .ZN(n8818) );
  NAND2_X1 U6258 ( .A1(n7495), .A2(n4444), .ZN(n7738) );
  NAND3_X1 U6259 ( .A1(n5004), .A2(n5005), .A3(n5003), .ZN(n4854) );
  NAND4_X1 U6260 ( .A1(n4992), .A2(n4969), .A3(n5100), .A4(n4852), .ZN(n5800)
         );
  OAI21_X2 U6261 ( .B1(n8891), .B2(n4473), .A(n4857), .ZN(n8864) );
  INV_X1 U6262 ( .A(n8896), .ZN(n4862) );
  OAI21_X1 U6263 ( .B1(n8976), .B2(n4866), .A(n4863), .ZN(n8922) );
  NAND2_X1 U6264 ( .A1(n7480), .A2(n4875), .ZN(n4874) );
  NAND2_X1 U6265 ( .A1(n8452), .A2(n4881), .ZN(n4880) );
  OAI211_X1 U6266 ( .C1(n8452), .C2(n4884), .A(n4880), .B(n8463), .ZN(P2_U3222) );
  INV_X1 U6267 ( .A(n4892), .ZN(n4889) );
  NOR2_X1 U6268 ( .A1(n4445), .A2(n8454), .ZN(n4891) );
  NAND2_X1 U6269 ( .A1(n4445), .A2(n8454), .ZN(n4892) );
  NAND2_X1 U6270 ( .A1(n7955), .A2(n7853), .ZN(n7855) );
  NAND2_X1 U6271 ( .A1(n8642), .A2(n4487), .ZN(n7357) );
  INV_X1 U6272 ( .A(n4996), .ZN(n4994) );
  OAI21_X1 U6273 ( .B1(n9201), .B2(n9200), .A(n4920), .ZN(n9287) );
  OAI21_X2 U6274 ( .B1(n8111), .B2(n4925), .A(n4921), .ZN(n6682) );
  INV_X1 U6275 ( .A(n6682), .ZN(n4928) );
  OAI21_X2 U6276 ( .B1(n9191), .B2(n4938), .A(n4935), .ZN(n8474) );
  NAND2_X1 U6277 ( .A1(n4940), .A2(n4942), .ZN(n9274) );
  NAND3_X1 U6278 ( .A1(n6692), .A2(n9294), .A3(n4944), .ZN(n4940) );
  NAND3_X1 U6279 ( .A1(n6750), .A2(n9251), .A3(n4955), .ZN(n4952) );
  NAND2_X1 U6280 ( .A1(n4952), .A2(n4954), .ZN(n9229) );
  NAND3_X1 U6281 ( .A1(n6750), .A2(n9251), .A3(n4959), .ZN(n4953) );
  INV_X1 U6282 ( .A(n6754), .ZN(n4961) );
  XNOR2_X1 U6283 ( .A(n5564), .B(n5563), .ZN(n8330) );
  NAND2_X1 U6284 ( .A1(n5481), .A2(n5480), .ZN(n5483) );
  OR2_X1 U6285 ( .A1(n8788), .A2(n5915), .ZN(n8796) );
  XNOR2_X1 U6286 ( .A(n5533), .B(n5532), .ZN(n8145) );
  XNOR2_X1 U6287 ( .A(n5513), .B(n5512), .ZN(n8188) );
  NAND2_X2 U6288 ( .A1(n5928), .A2(n5939), .ZN(n6535) );
  NAND4_X1 U6289 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n5017), .ZN(n7092)
         );
  AOI22_X1 U6290 ( .A1(n5886), .A2(n5885), .B1(n5884), .B2(n8803), .ZN(n5888)
         );
  CLKBUF_X1 U6291 ( .A(n8111), .Z(n8200) );
  NAND2_X1 U6292 ( .A1(n5617), .A2(n5662), .ZN(n5811) );
  NAND2_X1 U6293 ( .A1(n8922), .A2(n8923), .ZN(n8921) );
  AND2_X1 U6294 ( .A1(n5896), .A2(n5895), .ZN(n5894) );
  XNOR2_X1 U6295 ( .A(n8524), .B(n8523), .ZN(n8527) );
  AND4_X1 U6296 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n8980)
         );
  INV_X1 U6297 ( .A(n7007), .ZN(n6371) );
  OR2_X1 U6298 ( .A1(n5884), .A2(n9152), .ZN(n4964) );
  INV_X1 U6299 ( .A(n9439), .ZN(n8490) );
  INV_X1 U6300 ( .A(n6889), .ZN(n5793) );
  INV_X1 U6301 ( .A(n9414), .ZN(n9233) );
  OR2_X1 U6302 ( .A1(n5884), .A2(n9071), .ZN(n4965) );
  NOR2_X1 U6303 ( .A1(n6133), .A2(n6114), .ZN(n4966) );
  OR2_X1 U6304 ( .A1(n8926), .A2(n8658), .ZN(n4967) );
  AND2_X1 U6305 ( .A1(n5003), .A2(n4998), .ZN(n4968) );
  AND4_X1 U6306 ( .A1(n5002), .A2(n4993), .A3(n5787), .A4(n5001), .ZN(n4969)
         );
  NAND2_X2 U6307 ( .A1(n5908), .A2(n8989), .ZN(n9001) );
  OR2_X1 U6308 ( .A1(n8872), .A2(n8634), .ZN(n4972) );
  AND3_X1 U6309 ( .A1(n5394), .A2(n5393), .A3(n5392), .ZN(n8955) );
  INV_X1 U6310 ( .A(n8955), .ZN(n5830) );
  INV_X1 U6311 ( .A(n4794), .ZN(n6483) );
  AND2_X1 U6312 ( .A1(n5296), .A2(n5281), .ZN(n4974) );
  AND2_X1 U6313 ( .A1(n5209), .A2(n5199), .ZN(n4975) );
  INV_X1 U6314 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5966) );
  INV_X1 U6315 ( .A(n7502), .ZN(n7572) );
  AND2_X1 U6316 ( .A1(n5229), .A2(n5214), .ZN(n4976) );
  NAND2_X1 U6317 ( .A1(n8183), .A2(n9315), .ZN(n4977) );
  AND2_X1 U6318 ( .A1(n6760), .A2(n6759), .ZN(n4978) );
  AND4_X1 U6319 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9575), .ZN(n4979)
         );
  INV_X1 U6320 ( .A(n8960), .ZN(n5829) );
  OR4_X1 U6321 ( .A1(n9945), .A2(n6912), .A3(n5853), .A4(n8977), .ZN(n4981) );
  INV_X1 U6322 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4985) );
  INV_X1 U6323 ( .A(n6564), .ZN(n5996) );
  INV_X1 U6324 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5006) );
  AOI21_X1 U6325 ( .B1(n6373), .B2(n6372), .A(n6371), .ZN(n6374) );
  NAND2_X1 U6326 ( .A1(n6235), .A2(n6219), .ZN(n5965) );
  INV_X1 U6327 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5961) );
  INV_X1 U6328 ( .A(n5307), .ZN(n5305) );
  INV_X1 U6329 ( .A(n5184), .ZN(n5183) );
  INV_X1 U6330 ( .A(n5354), .ZN(n5352) );
  OR2_X1 U6331 ( .A1(n5332), .A2(n5331), .ZN(n5354) );
  INV_X1 U6332 ( .A(n5473), .ZN(n5472) );
  INV_X1 U6333 ( .A(n5288), .ZN(n5286) );
  INV_X1 U6334 ( .A(n8235), .ZN(n5294) );
  NAND2_X1 U6335 ( .A1(n6567), .A2(n6568), .ZN(n7262) );
  AND2_X1 U6336 ( .A1(n7276), .A2(n7273), .ZN(n6598) );
  XNOR2_X1 U6337 ( .A(n6576), .B(n6588), .ZN(n6579) );
  INV_X1 U6338 ( .A(n6280), .ZN(n5942) );
  INV_X1 U6339 ( .A(n5165), .ZN(n5166) );
  NAND2_X1 U6340 ( .A1(n5154), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6341 ( .A1(n7839), .A2(n4873), .ZN(n7840) );
  OR2_X1 U6342 ( .A1(n5264), .A2(n5263), .ZN(n5288) );
  OR2_X1 U6343 ( .A1(n5486), .A2(n10230), .ZN(n5506) );
  NAND2_X1 U6344 ( .A1(n5183), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5220) );
  INV_X1 U6345 ( .A(n7958), .ZN(n7846) );
  NAND2_X1 U6346 ( .A1(n5472), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6347 ( .A1(n5286), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5307) );
  OR2_X1 U6348 ( .A1(n9946), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5856) );
  INV_X1 U6349 ( .A(n5419), .ZN(n5568) );
  OR2_X1 U6350 ( .A1(n7529), .A2(n7528), .ZN(n6618) );
  NAND2_X1 U6351 ( .A1(n5952), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6330) );
  NOR2_X1 U6352 ( .A1(n6172), .A2(n9173), .ZN(n6192) );
  AND2_X1 U6353 ( .A1(n9592), .A2(n9488), .ZN(n8487) );
  INV_X1 U6354 ( .A(n6588), .ZN(n6562) );
  AND2_X1 U6355 ( .A1(n6482), .A2(n4794), .ZN(n6552) );
  OR2_X1 U6356 ( .A1(n6380), .A2(n6379), .ZN(n6382) );
  INV_X1 U6357 ( .A(n5316), .ZN(n5320) );
  INV_X1 U6358 ( .A(n5243), .ZN(n5247) );
  INV_X1 U6359 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6081) );
  INV_X1 U6360 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6038) );
  INV_X1 U6361 ( .A(n8627), .ZN(n8456) );
  OR2_X1 U6362 ( .A1(n5422), .A2(n8622), .ZN(n5437) );
  OR2_X1 U6363 ( .A1(n5455), .A2(n8635), .ZN(n5473) );
  OR2_X1 U6364 ( .A1(n5373), .A2(n7784), .ZN(n5406) );
  OR2_X1 U6365 ( .A1(n8637), .A2(n8977), .ZN(n8665) );
  OR3_X1 U6366 ( .A1(n5557), .A2(n8544), .A3(n8459), .ZN(n5903) );
  INV_X1 U6367 ( .A(n8865), .ZN(n8867) );
  OR2_X1 U6368 ( .A1(n9981), .A2(n8929), .ZN(n5892) );
  AND2_X1 U6369 ( .A1(n5857), .A2(n5856), .ZN(n7073) );
  INV_X1 U6370 ( .A(n8319), .ZN(n8317) );
  INV_X1 U6371 ( .A(n8945), .ZN(n8979) );
  OR2_X1 U6372 ( .A1(n7102), .A2(n7076), .ZN(n9981) );
  OR2_X1 U6373 ( .A1(n6890), .A2(n5804), .ZN(n9945) );
  NOR2_X1 U6374 ( .A1(n6226), .A2(n6225), .ZN(n6240) );
  NAND2_X1 U6375 ( .A1(n6544), .A2(n7412), .ZN(n7296) );
  AND2_X1 U6376 ( .A1(n6330), .A2(n5955), .ZN(n9377) );
  AND2_X1 U6377 ( .A1(n6259), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6269) );
  INV_X1 U6378 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7532) );
  INV_X1 U6379 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10095) );
  OR2_X1 U6380 ( .A1(n9832), .A2(n9831), .ZN(n9835) );
  AND2_X1 U6381 ( .A1(n6395), .A2(n8151), .ZN(n8172) );
  OR2_X1 U6382 ( .A1(n7296), .A2(n6525), .ZN(n7509) );
  INV_X1 U6383 ( .A(n6482), .ZN(n9420) );
  OR3_X1 U6384 ( .A1(n9876), .A2(n7412), .A3(n7411), .ZN(n9489) );
  INV_X1 U6385 ( .A(n7817), .ZN(n9867) );
  OR2_X1 U6386 ( .A1(n7296), .A2(n6535), .ZN(n9431) );
  OR2_X1 U6387 ( .A1(n7007), .A2(n6483), .ZN(n9876) );
  XNOR2_X1 U6388 ( .A(n5611), .B(n5610), .ZN(n6343) );
  AND2_X1 U6389 ( .A1(n5430), .A2(n5418), .ZN(n5428) );
  NAND2_X1 U6390 ( .A1(n5274), .A2(n5252), .ZN(n5275) );
  NOR2_X1 U6391 ( .A1(n8803), .A2(n8456), .ZN(n8457) );
  INV_X1 U6392 ( .A(n10343), .ZN(n8675) );
  AND2_X1 U6393 ( .A1(n5443), .A2(n5442), .ZN(n8633) );
  AND2_X1 U6394 ( .A1(n6915), .A2(n6914), .ZN(n9904) );
  OR2_X1 U6395 ( .A1(n9945), .A2(n5892), .ZN(n8989) );
  AND2_X1 U6396 ( .A1(n8383), .A2(n9081), .ZN(n8384) );
  NOR2_X1 U6397 ( .A1(n9994), .A2(n9979), .ZN(n9081) );
  INV_X1 U6398 ( .A(n8814), .ZN(n9108) );
  AND2_X1 U6399 ( .A1(n5733), .A2(n8912), .ZN(n8923) );
  OR2_X1 U6400 ( .A1(n7075), .A2(n5876), .ZN(n5889) );
  NAND2_X1 U6401 ( .A1(n9952), .A2(n5850), .ZN(n9946) );
  INV_X1 U6402 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5002) );
  INV_X1 U6403 ( .A(n9303), .ZN(n9291) );
  AND4_X1 U6404 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n6825)
         );
  NAND2_X1 U6405 ( .A1(n6355), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6023) );
  INV_X1 U6406 ( .A(n9833), .ZN(n9816) );
  INV_X1 U6407 ( .A(n9782), .ZN(n9823) );
  NAND2_X1 U6408 ( .A1(n8521), .A2(n6464), .ZN(n9363) );
  INV_X1 U6409 ( .A(n9380), .ZN(n9539) );
  AND2_X1 U6410 ( .A1(n7054), .A2(n7053), .ZN(n7056) );
  AND2_X1 U6411 ( .A1(n9672), .A2(n9876), .ZN(n9683) );
  INV_X1 U6412 ( .A(n9683), .ZN(n9887) );
  AND2_X1 U6413 ( .A1(n6795), .A2(n6794), .ZN(n7052) );
  INV_X1 U6414 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6187) );
  XNOR2_X1 U6415 ( .A(n5057), .B(n5031), .ZN(n5056) );
  AND2_X1 U6416 ( .A1(n9949), .A2(n5803), .ZN(n6890) );
  INV_X1 U6417 ( .A(n8904), .ZN(n9134) );
  INV_X1 U6418 ( .A(n8858), .ZN(n9123) );
  INV_X1 U6419 ( .A(n8668), .ZN(n10345) );
  INV_X1 U6420 ( .A(n8629), .ZN(n10351) );
  INV_X1 U6421 ( .A(n9001), .ZN(n8998) );
  INV_X1 U6422 ( .A(n9002), .ZN(n9937) );
  OR2_X1 U6423 ( .A1(n7075), .A2(n5858), .ZN(n9994) );
  AND2_X1 U6424 ( .A1(n5881), .A2(n4964), .ZN(n5882) );
  OR2_X1 U6425 ( .A1(n5889), .A2(n5878), .ZN(n9987) );
  AND2_X1 U6426 ( .A1(n5852), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9957) );
  OR2_X1 U6427 ( .A1(n5260), .A2(n5299), .ZN(n6986) );
  INV_X1 U6428 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6881) );
  INV_X1 U6429 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6849) );
  OR2_X1 U6430 ( .A1(n8530), .A2(n6808), .ZN(n6832) );
  OR2_X1 U6431 ( .A1(n9237), .A2(n9881), .ZN(n9303) );
  OR2_X1 U6432 ( .A1(n6815), .A2(n6819), .ZN(n9309) );
  NAND4_X1 U6433 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n9399)
         );
  OR2_X1 U6434 ( .A1(n9713), .A2(n9710), .ZN(n9833) );
  OR2_X1 U6435 ( .A1(n8371), .A2(n4727), .ZN(n9828) );
  NAND2_X1 U6436 ( .A1(n9477), .A2(n7511), .ZN(n9547) );
  INV_X1 U6437 ( .A(n9903), .ZN(n9901) );
  AND2_X2 U6438 ( .A1(n7056), .A2(n7055), .ZN(n9903) );
  OR3_X1 U6439 ( .A1(n9625), .A2(n9624), .A3(n9623), .ZN(n9640) );
  INV_X1 U6440 ( .A(n9891), .ZN(n9889) );
  AND2_X1 U6441 ( .A1(n7116), .A2(n6862), .ZN(n6860) );
  INV_X1 U6442 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10315) );
  INV_X1 U6443 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6879) );
  AND2_X1 U6444 ( .A1(n6890), .A2(n9957), .ZN(P2_U3966) );
  INV_X1 U6445 ( .A(n9324), .ZN(P1_U4006) );
  NOR2_X1 U6446 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4984) );
  NAND4_X1 U6447 ( .A1(n4984), .A2(n4983), .A3(n4982), .A4(n10294), .ZN(n4988)
         );
  NAND4_X1 U6448 ( .A1(n5298), .A2(n4986), .A3(n4985), .A4(n5115), .ZN(n4987)
         );
  INV_X1 U6449 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4998) );
  XNOR2_X1 U6450 ( .A(n4995), .B(n5002), .ZN(n7803) );
  NAND2_X1 U6451 ( .A1(n4996), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U6452 ( .A1(n5000), .A2(n5003), .ZN(n4997) );
  NAND2_X1 U6453 ( .A1(n4997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4999) );
  XNOR2_X1 U6454 ( .A(n4999), .B(n4998), .ZN(n7733) );
  XNOR2_X1 U6455 ( .A(n5000), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U6456 ( .A1(n7733), .A2(n8929), .ZN(n5853) );
  OR2_X1 U6457 ( .A1(n7102), .A2(n5853), .ZN(n8432) );
  INV_X1 U6458 ( .A(n7733), .ZN(n7076) );
  NAND2_X1 U6459 ( .A1(n7076), .A2(n7087), .ZN(n5863) );
  NOR2_X1 U6460 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5005) );
  NOR2_X1 U6461 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5004) );
  INV_X1 U6462 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6463 ( .A1(n5011), .A2(n5008), .ZN(n5013) );
  INV_X1 U6464 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5009) );
  INV_X1 U6465 ( .A(n5011), .ZN(n5022) );
  NAND2_X1 U6466 ( .A1(n5022), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5012) );
  NAND2_X4 U6467 ( .A1(n9161), .A2(n9166), .ZN(n5083) );
  INV_X1 U6468 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7594) );
  OR2_X1 U6469 ( .A1(n5083), .A2(n7594), .ZN(n5020) );
  NAND2_X2 U6470 ( .A1(n9166), .A2(n5015), .ZN(n5389) );
  INV_X1 U6471 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6895) );
  NAND2_X1 U6472 ( .A1(n5597), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5018) );
  INV_X1 U6473 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U6474 ( .A1(n5024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5025) );
  MUX2_X1 U6475 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5025), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5027) );
  NAND2_X1 U6476 ( .A1(n5027), .A2(n5026), .ZN(n6912) );
  INV_X1 U6477 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5028) );
  AND2_X1 U6478 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U6479 ( .A1(n5032), .A2(n5029), .ZN(n5039) );
  NAND2_X1 U6480 ( .A1(n5030), .A2(n5039), .ZN(n5057) );
  INV_X1 U6481 ( .A(SI_1_), .ZN(n5031) );
  MUX2_X1 U6482 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6834), .Z(n5055) );
  XNOR2_X1 U6483 ( .A(n5056), .B(n5055), .ZN(n6841) );
  NAND2_X1 U6484 ( .A1(n5117), .A2(n4724), .ZN(n5036) );
  NAND2_X1 U6485 ( .A1(n5071), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6486 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5033) );
  XNOR2_X1 U6487 ( .A(n5033), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U6488 ( .A1(n5401), .A2(n8709), .ZN(n5034) );
  INV_X1 U6489 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8708) );
  INV_X1 U6490 ( .A(SI_0_), .ZN(n5038) );
  INV_X1 U6491 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5037) );
  OAI21_X1 U6492 ( .B1(n4538), .B2(n5038), .A(n5037), .ZN(n5040) );
  NAND2_X1 U6493 ( .A1(n5040), .A2(n5039), .ZN(n9168) );
  MUX2_X1 U6494 ( .A(n8708), .B(n9168), .S(n6893), .Z(n7192) );
  INV_X1 U6495 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7135) );
  OR2_X1 U6496 ( .A1(n5083), .A2(n7135), .ZN(n5045) );
  NAND2_X1 U6497 ( .A1(n5597), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5044) );
  INV_X1 U6498 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5041) );
  OR2_X1 U6499 ( .A1(n5389), .A2(n5041), .ZN(n5043) );
  INV_X1 U6500 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6908) );
  OR2_X1 U6501 ( .A1(n5376), .A2(n6908), .ZN(n5042) );
  NAND4_X2 U6502 ( .A1(n5045), .A2(n5044), .A3(n5043), .A4(n5042), .ZN(n5810)
         );
  INV_X1 U6503 ( .A(n7092), .ZN(n5047) );
  INV_X1 U6504 ( .A(n7408), .ZN(n5046) );
  NAND2_X1 U6505 ( .A1(n5047), .A2(n5046), .ZN(n5617) );
  OAI21_X2 U6506 ( .B1(n5048), .B2(n7194), .A(n5617), .ZN(n7616) );
  INV_X1 U6507 ( .A(n7616), .ZN(n5065) );
  NAND2_X1 U6508 ( .A1(n5597), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5054) );
  INV_X1 U6509 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5049) );
  INV_X1 U6510 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9989) );
  OR2_X1 U6511 ( .A1(n5389), .A2(n9989), .ZN(n5052) );
  INV_X1 U6512 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5050) );
  OR2_X1 U6513 ( .A1(n5376), .A2(n5050), .ZN(n5051) );
  NAND2_X1 U6514 ( .A1(n5056), .A2(n5055), .ZN(n5059) );
  NAND2_X1 U6515 ( .A1(n5057), .A2(SI_1_), .ZN(n5058) );
  INV_X1 U6516 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6847) );
  INV_X1 U6517 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6835) );
  INV_X1 U6518 ( .A(n6846), .ZN(n5060) );
  NAND2_X1 U6519 ( .A1(n5117), .A2(n5060), .ZN(n5064) );
  NAND2_X1 U6520 ( .A1(n5071), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U6521 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4448), .ZN(n5061) );
  XNOR2_X1 U6522 ( .A(n5061), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U6523 ( .A1(n5401), .A2(n6907), .ZN(n5062) );
  INV_X1 U6524 ( .A(n5067), .ZN(n5068) );
  NAND2_X1 U6525 ( .A1(n5068), .A2(SI_2_), .ZN(n5090) );
  NAND2_X1 U6526 ( .A1(n5092), .A2(n5090), .ZN(n5069) );
  XNOR2_X1 U6527 ( .A(n5088), .B(SI_3_), .ZN(n5094) );
  XNOR2_X1 U6528 ( .A(n5069), .B(n5094), .ZN(n6848) );
  INV_X1 U6529 ( .A(n6848), .ZN(n5070) );
  NAND2_X1 U6530 ( .A1(n5117), .A2(n5070), .ZN(n5075) );
  NAND2_X1 U6531 ( .A1(n5328), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5074) );
  OAI21_X1 U6532 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n4448), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5072) );
  XNOR2_X1 U6533 ( .A(n5072), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6906) );
  NAND2_X1 U6534 ( .A1(n5401), .A2(n6906), .ZN(n5073) );
  AND3_X2 U6535 ( .A1(n5075), .A2(n5074), .A3(n5073), .ZN(n7436) );
  NAND2_X1 U6536 ( .A1(n5597), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5081) );
  OR2_X1 U6537 ( .A1(n5083), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5080) );
  INV_X1 U6538 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5076) );
  OR2_X1 U6539 ( .A1(n5594), .A2(n5076), .ZN(n5079) );
  INV_X1 U6540 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5077) );
  OR2_X1 U6541 ( .A1(n5389), .A2(n5077), .ZN(n5078) );
  NAND2_X1 U6542 ( .A1(n10348), .A2(n7436), .ZN(n5648) );
  NAND2_X1 U6543 ( .A1(n5596), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5087) );
  INV_X1 U6544 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5082) );
  OR2_X1 U6545 ( .A1(n5459), .A2(n5082), .ZN(n5086) );
  XNOR2_X1 U6546 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n10340) );
  OR2_X1 U6547 ( .A1(n5083), .A2(n10340), .ZN(n5085) );
  INV_X1 U6548 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6911) );
  OR2_X1 U6549 ( .A1(n5376), .A2(n6911), .ZN(n5084) );
  NAND4_X1 U6550 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n8704)
         );
  INV_X1 U6551 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6552 ( .A1(n5089), .A2(SI_3_), .ZN(n5093) );
  AND2_X1 U6553 ( .A1(n5090), .A2(n5093), .ZN(n5091) );
  MUX2_X1 U6554 ( .A(n6852), .B(n5096), .S(n4538), .Z(n5119) );
  XNOR2_X1 U6555 ( .A(n4475), .B(n5118), .ZN(n6851) );
  INV_X1 U6556 ( .A(n6851), .ZN(n5097) );
  NAND2_X1 U6557 ( .A1(n5097), .A2(n5117), .ZN(n5104) );
  NOR2_X1 U6558 ( .A1(n5098), .A2(n9157), .ZN(n5099) );
  MUX2_X1 U6559 ( .A(n9157), .B(n5099), .S(P2_IR_REG_4__SCAN_IN), .Z(n5101) );
  NOR2_X1 U6560 ( .A1(n5101), .A2(n5100), .ZN(n6950) );
  NAND2_X1 U6561 ( .A1(n5401), .A2(n6950), .ZN(n5103) );
  NAND2_X1 U6562 ( .A1(n5328), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6563 ( .A1(n8704), .A2(n10344), .ZN(n5649) );
  NOR2_X1 U6564 ( .A1(n8704), .A2(n10344), .ZN(n5618) );
  AOI21_X1 U6565 ( .B1(n7606), .B2(n5649), .A(n5618), .ZN(n7385) );
  NAND2_X1 U6566 ( .A1(n5596), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5112) );
  INV_X1 U6567 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5105) );
  OR2_X1 U6568 ( .A1(n5459), .A2(n5105), .ZN(n5111) );
  NAND3_X1 U6569 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5124) );
  INV_X1 U6570 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6571 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5106) );
  NAND2_X1 U6572 ( .A1(n5107), .A2(n5106), .ZN(n5108) );
  NAND2_X1 U6573 ( .A1(n5124), .A2(n5108), .ZN(n8592) );
  OR2_X1 U6574 ( .A1(n5083), .A2(n8592), .ZN(n5110) );
  INV_X1 U6575 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7760) );
  OR2_X1 U6576 ( .A1(n5594), .A2(n7760), .ZN(n5109) );
  NOR2_X1 U6577 ( .A1(n5100), .A2(n9157), .ZN(n5113) );
  MUX2_X1 U6578 ( .A(n9157), .B(n5113), .S(P2_IR_REG_5__SCAN_IN), .Z(n5114) );
  INV_X1 U6579 ( .A(n5114), .ZN(n5116) );
  NAND2_X1 U6580 ( .A1(n5100), .A2(n5115), .ZN(n5149) );
  AND2_X1 U6581 ( .A1(n5116), .A2(n5149), .ZN(n8724) );
  INV_X1 U6582 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6583 ( .A1(n5120), .A2(SI_4_), .ZN(n5121) );
  MUX2_X1 U6584 ( .A(n6845), .B(n6839), .S(n4538), .Z(n5133) );
  XNOR2_X1 U6585 ( .A(n5132), .B(n5131), .ZN(n6844) );
  OR2_X1 U6586 ( .A1(n5419), .A2(n6844), .ZN(n5122) );
  NAND2_X1 U6587 ( .A1(n10342), .A2(n8594), .ZN(n5655) );
  INV_X1 U6588 ( .A(n10342), .ZN(n8703) );
  NAND2_X1 U6589 ( .A1(n7385), .A2(n7384), .ZN(n7445) );
  NAND2_X1 U6590 ( .A1(n5597), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5130) );
  INV_X1 U6591 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6954) );
  OR2_X1 U6592 ( .A1(n5594), .A2(n6954), .ZN(n5129) );
  INV_X1 U6593 ( .A(n5124), .ZN(n5123) );
  NAND2_X1 U6594 ( .A1(n5123), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5156) );
  INV_X1 U6595 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U6596 ( .A1(n5124), .A2(n7370), .ZN(n5125) );
  NAND2_X1 U6597 ( .A1(n5156), .A2(n5125), .ZN(n7691) );
  OR2_X1 U6598 ( .A1(n5083), .A2(n7691), .ZN(n5128) );
  INV_X1 U6599 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5126) );
  OR2_X1 U6600 ( .A1(n5389), .A2(n5126), .ZN(n5127) );
  NAND2_X1 U6601 ( .A1(n5132), .A2(n5131), .ZN(n5136) );
  INV_X1 U6602 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6603 ( .A1(n5134), .A2(SI_5_), .ZN(n5135) );
  INV_X1 U6604 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5137) );
  MUX2_X1 U6605 ( .A(n10292), .B(n5137), .S(n4538), .Z(n5146) );
  XNOR2_X1 U6606 ( .A(n5145), .B(n5144), .ZN(n6850) );
  OR2_X1 U6607 ( .A1(n6850), .A2(n5419), .ZN(n5140) );
  NAND2_X1 U6608 ( .A1(n5149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5138) );
  XNOR2_X1 U6609 ( .A(n5138), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7032) );
  AOI22_X1 U6610 ( .A1(n5328), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5401), .B2(
        n7032), .ZN(n5139) );
  NAND2_X1 U6611 ( .A1(n5140), .A2(n5139), .ZN(n7451) );
  NAND2_X1 U6612 ( .A1(n7493), .A2(n7451), .ZN(n5671) );
  INV_X1 U6613 ( .A(n7451), .ZN(n7695) );
  INV_X1 U6614 ( .A(n7493), .ZN(n8702) );
  NAND2_X1 U6615 ( .A1(n7695), .A2(n8702), .ZN(n5670) );
  NAND2_X1 U6616 ( .A1(n5671), .A2(n5670), .ZN(n5818) );
  INV_X1 U6617 ( .A(n7444), .ZN(n5141) );
  NOR2_X1 U6618 ( .A1(n5818), .A2(n5141), .ZN(n5142) );
  NAND2_X1 U6619 ( .A1(n7445), .A2(n5142), .ZN(n5143) );
  NAND2_X1 U6620 ( .A1(n5143), .A2(n5671), .ZN(n7492) );
  INV_X1 U6621 ( .A(n7492), .ZN(n5164) );
  INV_X1 U6622 ( .A(n5146), .ZN(n5147) );
  MUX2_X1 U6623 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4538), .Z(n5168) );
  XNOR2_X1 U6624 ( .A(n5167), .B(n5165), .ZN(n6855) );
  NAND2_X1 U6625 ( .A1(n6855), .A2(n5117), .ZN(n5152) );
  NAND2_X1 U6626 ( .A1(n5175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5150) );
  XNOR2_X1 U6627 ( .A(n5150), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8737) );
  AOI22_X1 U6628 ( .A1(n5328), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5401), .B2(
        n8737), .ZN(n5151) );
  NAND2_X1 U6629 ( .A1(n5152), .A2(n5151), .ZN(n7632) );
  NAND2_X1 U6630 ( .A1(n5596), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5162) );
  INV_X1 U6631 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5153) );
  OR2_X1 U6632 ( .A1(n5459), .A2(n5153), .ZN(n5161) );
  INV_X1 U6633 ( .A(n5156), .ZN(n5154) );
  INV_X1 U6634 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6635 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U6636 ( .A1(n5184), .A2(n5157), .ZN(n7629) );
  OR2_X1 U6637 ( .A1(n5083), .A2(n7629), .ZN(n5160) );
  INV_X1 U6638 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5158) );
  OR2_X1 U6639 ( .A1(n5376), .A2(n5158), .ZN(n5159) );
  OR2_X1 U6640 ( .A1(n7632), .A2(n7377), .ZN(n5674) );
  NAND2_X1 U6641 ( .A1(n7632), .A2(n7377), .ZN(n5687) );
  NAND2_X1 U6642 ( .A1(n5674), .A2(n5687), .ZN(n7491) );
  NAND2_X1 U6643 ( .A1(n5168), .A2(SI_7_), .ZN(n5169) );
  MUX2_X1 U6644 ( .A(n6864), .B(n6866), .S(n4538), .Z(n5172) );
  INV_X1 U6645 ( .A(SI_8_), .ZN(n5171) );
  INV_X1 U6646 ( .A(n5172), .ZN(n5173) );
  NAND2_X1 U6647 ( .A1(n5173), .A2(SI_8_), .ZN(n5174) );
  XNOR2_X1 U6648 ( .A(n5195), .B(n5194), .ZN(n6863) );
  NAND2_X1 U6649 ( .A1(n6863), .A2(n5568), .ZN(n5182) );
  NOR2_X1 U6650 ( .A1(n5178), .A2(n9157), .ZN(n5176) );
  MUX2_X1 U6651 ( .A(n9157), .B(n5176), .S(P2_IR_REG_8__SCAN_IN), .Z(n5180) );
  INV_X1 U6652 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6653 ( .A1(n5178), .A2(n5177), .ZN(n5215) );
  INV_X1 U6654 ( .A(n5215), .ZN(n5179) );
  NOR2_X1 U6655 ( .A1(n5180), .A2(n5179), .ZN(n7070) );
  AOI22_X1 U6656 ( .A1(n5328), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5401), .B2(
        n7070), .ZN(n5181) );
  NAND2_X1 U6657 ( .A1(n5182), .A2(n5181), .ZN(n7771) );
  NAND2_X1 U6658 ( .A1(n5597), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5191) );
  INV_X1 U6659 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U6660 ( .A1(n5184), .A2(n10175), .ZN(n5185) );
  NAND2_X1 U6661 ( .A1(n5220), .A2(n5185), .ZN(n7483) );
  OR2_X1 U6662 ( .A1(n5083), .A2(n7483), .ZN(n5190) );
  INV_X1 U6663 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5186) );
  OR2_X1 U6664 ( .A1(n5594), .A2(n5186), .ZN(n5189) );
  INV_X1 U6665 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6666 ( .A1(n5389), .A2(n5187), .ZN(n5188) );
  OR2_X1 U6667 ( .A1(n7771), .A2(n7646), .ZN(n5679) );
  NAND2_X1 U6668 ( .A1(n7771), .A2(n7646), .ZN(n5676) );
  NAND2_X1 U6669 ( .A1(n5679), .A2(n5676), .ZN(n7741) );
  NAND2_X1 U6670 ( .A1(n7738), .A2(n5676), .ZN(n7808) );
  INV_X1 U6671 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5196) );
  MUX2_X1 U6672 ( .A(n5196), .B(n6873), .S(n4538), .Z(n5197) );
  INV_X1 U6673 ( .A(n5197), .ZN(n5198) );
  NAND2_X1 U6674 ( .A1(n5198), .A2(SI_9_), .ZN(n5199) );
  NAND2_X1 U6675 ( .A1(n6872), .A2(n5117), .ZN(n5202) );
  NAND2_X1 U6676 ( .A1(n5215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5200) );
  XNOR2_X1 U6677 ( .A(n5200), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7045) );
  AOI22_X1 U6678 ( .A1(n5328), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5401), .B2(
        n7045), .ZN(n5201) );
  NAND2_X1 U6679 ( .A1(n5597), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5207) );
  INV_X1 U6680 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6681 ( .A1(n5389), .A2(n5203), .ZN(n5206) );
  INV_X1 U6682 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7649) );
  XNOR2_X1 U6683 ( .A(n5220), .B(n7649), .ZN(n9932) );
  OR2_X1 U6684 ( .A1(n5083), .A2(n9932), .ZN(n5205) );
  INV_X1 U6685 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6958) );
  OR2_X1 U6686 ( .A1(n5594), .A2(n6958), .ZN(n5204) );
  OR2_X1 U6687 ( .A1(n9929), .A2(n7941), .ZN(n5682) );
  INV_X1 U6688 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5210) );
  MUX2_X1 U6689 ( .A(n5210), .B(n6879), .S(n6837), .Z(n5212) );
  INV_X1 U6690 ( .A(SI_10_), .ZN(n5211) );
  INV_X1 U6691 ( .A(n5212), .ZN(n5213) );
  NAND2_X1 U6692 ( .A1(n5213), .A2(SI_10_), .ZN(n5214) );
  XNOR2_X1 U6693 ( .A(n5228), .B(n4976), .ZN(n6875) );
  NAND2_X1 U6694 ( .A1(n6875), .A2(n5117), .ZN(n5217) );
  NAND2_X1 U6695 ( .A1(n5256), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6696 ( .A(n5231), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6972) );
  AOI22_X1 U6697 ( .A1(n5328), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5401), .B2(
        n6972), .ZN(n5216) );
  NAND2_X1 U6698 ( .A1(n5597), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5227) );
  INV_X1 U6699 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5218) );
  OR2_X1 U6700 ( .A1(n5389), .A2(n5218), .ZN(n5226) );
  INV_X1 U6701 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5219) );
  OAI21_X1 U6702 ( .B1(n5220), .B2(n7649), .A(n5219), .ZN(n5223) );
  AND2_X1 U6703 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n5221) );
  NAND2_X1 U6704 ( .A1(n5223), .A2(n5237), .ZN(n7954) );
  OR2_X1 U6705 ( .A1(n5083), .A2(n7954), .ZN(n5225) );
  INV_X1 U6706 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7945) );
  OR2_X1 U6707 ( .A1(n5376), .A2(n7945), .ZN(n5224) );
  NAND2_X1 U6708 ( .A1(n7961), .A2(n7859), .ZN(n5686) );
  MUX2_X1 U6709 ( .A(n6881), .B(n10244), .S(n6837), .Z(n5244) );
  XNOR2_X1 U6710 ( .A(n5248), .B(n5243), .ZN(n6880) );
  NAND2_X1 U6711 ( .A1(n6880), .A2(n5117), .ZN(n5235) );
  INV_X1 U6712 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6713 ( .A1(n5231), .A2(n5254), .ZN(n5232) );
  NAND2_X1 U6714 ( .A1(n5232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5233) );
  XNOR2_X1 U6715 ( .A(n5233), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6976) );
  AOI22_X1 U6716 ( .A1(n5328), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5401), .B2(
        n6976), .ZN(n5234) );
  NAND2_X1 U6717 ( .A1(n5235), .A2(n5234), .ZN(n8043) );
  NAND2_X1 U6718 ( .A1(n5596), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5242) );
  INV_X1 U6719 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5236) );
  OR2_X1 U6720 ( .A1(n5459), .A2(n5236), .ZN(n5241) );
  INV_X1 U6721 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U6722 ( .A1(n5237), .A2(n7858), .ZN(n5238) );
  NAND2_X1 U6723 ( .A1(n5264), .A2(n5238), .ZN(n8038) );
  OR2_X1 U6724 ( .A1(n5083), .A2(n8038), .ZN(n5240) );
  INV_X1 U6725 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8039) );
  OR2_X1 U6726 ( .A1(n5594), .A2(n8039), .ZN(n5239) );
  OR2_X1 U6727 ( .A1(n8043), .A2(n8081), .ZN(n5694) );
  NAND2_X1 U6728 ( .A1(n8043), .A2(n8081), .ZN(n8077) );
  NAND2_X1 U6729 ( .A1(n5694), .A2(n8077), .ZN(n7964) );
  INV_X1 U6730 ( .A(n5244), .ZN(n5245) );
  NAND2_X1 U6731 ( .A1(n5245), .A2(SI_11_), .ZN(n5246) );
  INV_X1 U6732 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6888) );
  INV_X1 U6733 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6886) );
  MUX2_X1 U6734 ( .A(n6888), .B(n6886), .S(n6837), .Z(n5250) );
  INV_X1 U6735 ( .A(SI_12_), .ZN(n5249) );
  INV_X1 U6736 ( .A(n5250), .ZN(n5251) );
  NAND2_X1 U6737 ( .A1(n5251), .A2(SI_12_), .ZN(n5252) );
  XNOR2_X1 U6738 ( .A(n5276), .B(n5275), .ZN(n6884) );
  NAND2_X1 U6739 ( .A1(n6884), .A2(n5117), .ZN(n5262) );
  INV_X1 U6740 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6741 ( .A1(n5254), .A2(n5253), .ZN(n5255) );
  NOR2_X1 U6742 ( .A1(n5256), .A2(n5255), .ZN(n5259) );
  NOR2_X1 U6743 ( .A1(n5259), .A2(n9157), .ZN(n5257) );
  MUX2_X1 U6744 ( .A(n9157), .B(n5257), .S(P2_IR_REG_12__SCAN_IN), .Z(n5260)
         );
  INV_X1 U6745 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5258) );
  INV_X1 U6746 ( .A(n6986), .ZN(n7209) );
  AOI22_X1 U6747 ( .A1(n7209), .A2(n5401), .B1(n5328), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6748 ( .A1(n5597), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5270) );
  INV_X1 U6749 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6977) );
  OR2_X1 U6750 ( .A1(n5389), .A2(n6977), .ZN(n5269) );
  INV_X1 U6751 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6752 ( .A1(n5264), .A2(n5263), .ZN(n5265) );
  NAND2_X1 U6753 ( .A1(n5288), .A2(n5265), .ZN(n8085) );
  OR2_X1 U6754 ( .A1(n5083), .A2(n8085), .ZN(n5268) );
  INV_X1 U6755 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6756 ( .A1(n5594), .A2(n5266), .ZN(n5267) );
  NAND2_X1 U6757 ( .A1(n8087), .A2(n8237), .ZN(n5701) );
  NAND2_X1 U6758 ( .A1(n5702), .A2(n5701), .ZN(n8078) );
  INV_X1 U6759 ( .A(n8077), .ZN(n5271) );
  NOR2_X1 U6760 ( .A1(n8078), .A2(n5271), .ZN(n5272) );
  NAND2_X1 U6761 ( .A1(n5273), .A2(n5702), .ZN(n8234) );
  INV_X1 U6762 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7003) );
  INV_X1 U6763 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5277) );
  MUX2_X1 U6764 ( .A(n7003), .B(n5277), .S(n4538), .Z(n5279) );
  INV_X1 U6765 ( .A(SI_13_), .ZN(n5278) );
  INV_X1 U6766 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6767 ( .A1(n5280), .A2(SI_13_), .ZN(n5281) );
  XNOR2_X1 U6768 ( .A(n5295), .B(n4974), .ZN(n6964) );
  NAND2_X1 U6769 ( .A1(n6964), .A2(n5568), .ZN(n5284) );
  OR2_X1 U6770 ( .A1(n5299), .A2(n9157), .ZN(n5282) );
  XNOR2_X1 U6771 ( .A(n5282), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9923) );
  AOI22_X1 U6772 ( .A1(n9923), .A2(n5401), .B1(n5328), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6773 ( .A1(n5597), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5293) );
  INV_X1 U6774 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6775 ( .A1(n5389), .A2(n5285), .ZN(n5292) );
  INV_X1 U6776 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6777 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  NAND2_X1 U6778 ( .A1(n5307), .A2(n5289), .ZN(n8251) );
  OR2_X1 U6779 ( .A1(n5083), .A2(n8251), .ZN(n5291) );
  INV_X1 U6780 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8243) );
  OR2_X1 U6781 ( .A1(n5376), .A2(n8243), .ZN(n5290) );
  OR2_X1 U6782 ( .A1(n9092), .A2(n8269), .ZN(n5705) );
  NAND2_X1 U6783 ( .A1(n9092), .A2(n8269), .ZN(n8266) );
  NAND2_X1 U6784 ( .A1(n5705), .A2(n8266), .ZN(n8235) );
  INV_X1 U6785 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7006) );
  MUX2_X1 U6786 ( .A(n7006), .B(n10315), .S(n4538), .Z(n5317) );
  NAND2_X1 U6787 ( .A1(n7004), .A2(n5568), .ZN(n5304) );
  NAND2_X1 U6788 ( .A1(n5299), .A2(n5298), .ZN(n5300) );
  NAND2_X1 U6789 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6790 ( .A1(n5301), .A2(n10294), .ZN(n5326) );
  OR2_X1 U6791 ( .A1(n5301), .A2(n10294), .ZN(n5302) );
  AOI22_X1 U6792 ( .A1(n7660), .A2(n5401), .B1(n5328), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5303) );
  INV_X1 U6793 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7206) );
  OR2_X1 U6794 ( .A1(n5389), .A2(n7206), .ZN(n5313) );
  INV_X1 U6795 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10156) );
  OR2_X1 U6796 ( .A1(n5459), .A2(n10156), .ZN(n5312) );
  INV_X1 U6797 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6798 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U6799 ( .A1(n5332), .A2(n5308), .ZN(n8261) );
  OR2_X1 U6800 ( .A1(n5083), .A2(n8261), .ZN(n5311) );
  INV_X1 U6801 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5309) );
  OR2_X1 U6802 ( .A1(n5594), .A2(n5309), .ZN(n5310) );
  NAND2_X1 U6803 ( .A1(n9087), .A2(n8322), .ZN(n5708) );
  INV_X1 U6804 ( .A(n8266), .ZN(n5314) );
  NOR2_X1 U6805 ( .A1(n8258), .A2(n5314), .ZN(n5315) );
  INV_X1 U6806 ( .A(n5317), .ZN(n5318) );
  NAND2_X1 U6807 ( .A1(n5318), .A2(SI_14_), .ZN(n5319) );
  INV_X1 U6808 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7187) );
  INV_X1 U6809 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7189) );
  MUX2_X1 U6810 ( .A(n7187), .B(n7189), .S(n6837), .Z(n5323) );
  INV_X1 U6811 ( .A(SI_15_), .ZN(n5322) );
  INV_X1 U6812 ( .A(n5323), .ZN(n5324) );
  NAND2_X1 U6813 ( .A1(n5324), .A2(SI_15_), .ZN(n5325) );
  XNOR2_X1 U6814 ( .A(n5341), .B(n5340), .ZN(n7186) );
  NAND2_X1 U6815 ( .A1(n7186), .A2(n5568), .ZN(n5330) );
  NAND2_X1 U6816 ( .A1(n5326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5327) );
  XNOR2_X1 U6817 ( .A(n5327), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7679) );
  AOI22_X1 U6818 ( .A1(n7679), .A2(n5401), .B1(n5328), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5329) );
  INV_X1 U6819 ( .A(n5594), .ZN(n5598) );
  NAND2_X1 U6820 ( .A1(n5598), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5337) );
  INV_X1 U6821 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9079) );
  OR2_X1 U6822 ( .A1(n5389), .A2(n9079), .ZN(n5336) );
  INV_X1 U6823 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10314) );
  OR2_X1 U6824 ( .A1(n5459), .A2(n10314), .ZN(n5335) );
  INV_X1 U6825 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6826 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  NAND2_X1 U6827 ( .A1(n5354), .A2(n5333), .ZN(n8324) );
  OR2_X1 U6828 ( .A1(n5083), .A2(n8324), .ZN(n5334) );
  NAND2_X1 U6829 ( .A1(n9080), .A2(n8978), .ZN(n5713) );
  NAND2_X1 U6830 ( .A1(n8320), .A2(n8319), .ZN(n5338) );
  NAND2_X1 U6831 ( .A1(n5338), .A2(n5712), .ZN(n8973) );
  INV_X1 U6832 ( .A(n8973), .ZN(n5361) );
  INV_X1 U6833 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7272) );
  INV_X1 U6834 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7285) );
  MUX2_X1 U6835 ( .A(n7272), .B(n7285), .S(n4538), .Z(n5343) );
  INV_X1 U6836 ( .A(SI_16_), .ZN(n5342) );
  NAND2_X1 U6837 ( .A1(n5343), .A2(n5342), .ZN(n5364) );
  INV_X1 U6838 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U6839 ( .A1(n5344), .A2(SI_16_), .ZN(n5345) );
  XNOR2_X1 U6840 ( .A(n5363), .B(n5362), .ZN(n7271) );
  NAND2_X1 U6841 ( .A1(n7271), .A2(n5568), .ZN(n5351) );
  INV_X1 U6842 ( .A(n5346), .ZN(n5347) );
  NAND2_X1 U6843 ( .A1(n5347), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5348) );
  MUX2_X1 U6844 ( .A(n5348), .B(P2_IR_REG_31__SCAN_IN), .S(n4993), .Z(n5349)
         );
  AND2_X1 U6845 ( .A1(n5349), .A2(n5366), .ZN(n7781) );
  AOI22_X1 U6846 ( .A1(n5328), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5401), .B2(
        n7781), .ZN(n5350) );
  NAND2_X1 U6847 ( .A1(n5597), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5359) );
  INV_X1 U6848 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7671) );
  OR2_X1 U6849 ( .A1(n5389), .A2(n7671), .ZN(n5358) );
  INV_X1 U6850 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6851 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6852 ( .A1(n5373), .A2(n5355), .ZN(n8990) );
  OR2_X1 U6853 ( .A1(n5083), .A2(n8990), .ZN(n5357) );
  INV_X1 U6854 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8991) );
  OR2_X1 U6855 ( .A1(n5594), .A2(n8991), .ZN(n5356) );
  OR2_X1 U6856 ( .A1(n8993), .A2(n8956), .ZN(n5642) );
  NAND2_X1 U6857 ( .A1(n8993), .A2(n8956), .ZN(n5719) );
  NAND2_X1 U6858 ( .A1(n5642), .A2(n5719), .ZN(n8974) );
  INV_X1 U6859 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7310) );
  INV_X1 U6860 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7343) );
  MUX2_X1 U6861 ( .A(n7310), .B(n7343), .S(n4538), .Z(n5382) );
  XNOR2_X1 U6862 ( .A(n5382), .B(SI_17_), .ZN(n5381) );
  XNOR2_X1 U6863 ( .A(n5385), .B(n5381), .ZN(n7309) );
  NAND2_X1 U6864 ( .A1(n7309), .A2(n5568), .ZN(n5372) );
  NAND2_X1 U6865 ( .A1(n5366), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5367) );
  MUX2_X1 U6866 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5367), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5370) );
  INV_X1 U6867 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6868 ( .A1(n5370), .A2(n5369), .ZN(n7791) );
  INV_X1 U6869 ( .A(n7791), .ZN(n8754) );
  AOI22_X1 U6870 ( .A1(n5328), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5401), .B2(
        n8754), .ZN(n5371) );
  INV_X1 U6871 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U6872 ( .A1(n5373), .A2(n7784), .ZN(n5374) );
  AND2_X1 U6873 ( .A1(n5406), .A2(n5374), .ZN(n8963) );
  NAND2_X1 U6874 ( .A1(n8963), .A2(n5574), .ZN(n5380) );
  NAND2_X1 U6875 ( .A1(n5597), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5379) );
  INV_X1 U6876 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9069) );
  OR2_X1 U6877 ( .A1(n5389), .A2(n9069), .ZN(n5378) );
  INV_X1 U6878 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n5375) );
  OR2_X1 U6879 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  XNOR2_X1 U6880 ( .A(n8960), .B(n8980), .ZN(n8958) );
  OR2_X1 U6881 ( .A1(n8960), .A2(n8980), .ZN(n5641) );
  INV_X1 U6882 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6883 ( .A1(n5383), .A2(SI_17_), .ZN(n5384) );
  MUX2_X1 U6884 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6837), .Z(n5397) );
  XNOR2_X1 U6885 ( .A(n5397), .B(SI_18_), .ZN(n5395) );
  XNOR2_X1 U6886 ( .A(n5396), .B(n5395), .ZN(n7473) );
  NAND2_X1 U6887 ( .A1(n7473), .A2(n5568), .ZN(n5388) );
  OR2_X1 U6888 ( .A1(n5368), .A2(n9157), .ZN(n5386) );
  XNOR2_X1 U6889 ( .A(n5386), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8752) );
  AOI22_X1 U6890 ( .A1(n5328), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5401), .B2(
        n8752), .ZN(n5387) );
  XNOR2_X1 U6891 ( .A(n5406), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U6892 ( .A1(n8937), .A2(n5574), .ZN(n5394) );
  INV_X1 U6893 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8763) );
  OR2_X1 U6894 ( .A1(n5389), .A2(n8763), .ZN(n5391) );
  INV_X1 U6895 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10317) );
  OR2_X1 U6896 ( .A1(n5459), .A2(n10317), .ZN(n5390) );
  AND2_X1 U6897 ( .A1(n5391), .A2(n5390), .ZN(n5393) );
  NAND2_X1 U6898 ( .A1(n5598), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5392) );
  OR2_X1 U6899 ( .A1(n9061), .A2(n8955), .ZN(n5729) );
  NAND2_X1 U6900 ( .A1(n9061), .A2(n8955), .ZN(n5731) );
  NAND2_X1 U6901 ( .A1(n5729), .A2(n5731), .ZN(n8940) );
  INV_X1 U6902 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7591) );
  INV_X1 U6903 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7589) );
  MUX2_X1 U6904 ( .A(n7591), .B(n7589), .S(n4538), .Z(n5398) );
  INV_X1 U6905 ( .A(SI_19_), .ZN(n10320) );
  NAND2_X1 U6906 ( .A1(n5398), .A2(n10320), .ZN(n5413) );
  INV_X1 U6907 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U6908 ( .A1(n5399), .A2(SI_19_), .ZN(n5400) );
  NAND2_X1 U6909 ( .A1(n5413), .A2(n5400), .ZN(n5414) );
  XNOR2_X1 U6910 ( .A(n5415), .B(n5414), .ZN(n7588) );
  NAND2_X1 U6911 ( .A1(n7588), .A2(n5568), .ZN(n5403) );
  AOI22_X1 U6912 ( .A1(n5328), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5401), .B2(
        n5860), .ZN(n5402) );
  AOI22_X1 U6913 ( .A1(n5596), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n5597), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5412) );
  INV_X1 U6914 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5405) );
  INV_X1 U6915 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5404) );
  OAI21_X1 U6916 ( .B1(n5406), .B2(n5405), .A(n5404), .ZN(n5409) );
  AND2_X1 U6917 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5407) );
  NAND2_X1 U6918 ( .A1(n5409), .A2(n5422), .ZN(n8931) );
  OR2_X1 U6919 ( .A1(n8931), .A2(n5083), .ZN(n5411) );
  NAND2_X1 U6920 ( .A1(n5598), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5410) );
  OR2_X1 U6921 ( .A1(n9143), .A2(n8658), .ZN(n5733) );
  NAND2_X1 U6922 ( .A1(n9143), .A2(n8658), .ZN(n8912) );
  INV_X1 U6923 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7734) );
  INV_X1 U6924 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7774) );
  MUX2_X1 U6925 ( .A(n7734), .B(n7774), .S(n4538), .Z(n5416) );
  INV_X1 U6926 ( .A(SI_20_), .ZN(n10118) );
  NAND2_X1 U6927 ( .A1(n5416), .A2(n10118), .ZN(n5430) );
  INV_X1 U6928 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U6929 ( .A1(n5417), .A2(SI_20_), .ZN(n5418) );
  XNOR2_X1 U6930 ( .A(n5429), .B(n5428), .ZN(n7732) );
  NAND2_X1 U6931 ( .A1(n7732), .A2(n5568), .ZN(n5421) );
  NAND2_X1 U6932 ( .A1(n5328), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5420) );
  INV_X1 U6933 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U6934 ( .A1(n5422), .A2(n8622), .ZN(n5423) );
  AND2_X1 U6935 ( .A1(n5437), .A2(n5423), .ZN(n8909) );
  NAND2_X1 U6936 ( .A1(n8909), .A2(n5574), .ZN(n5426) );
  AOI22_X1 U6937 ( .A1(n5596), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5597), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6938 ( .A1(n5598), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6939 ( .A1(n9049), .A2(n8892), .ZN(n5736) );
  AND2_X1 U6940 ( .A1(n5736), .A2(n8912), .ZN(n5722) );
  NAND2_X1 U6941 ( .A1(n8921), .A2(n5722), .ZN(n5427) );
  INV_X1 U6942 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n5432) );
  INV_X1 U6943 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7833) );
  MUX2_X1 U6944 ( .A(n5432), .B(n7833), .S(n6837), .Z(n5446) );
  XNOR2_X1 U6945 ( .A(n5446), .B(SI_21_), .ZN(n5445) );
  XNOR2_X1 U6946 ( .A(n5444), .B(n5445), .ZN(n7802) );
  NAND2_X1 U6947 ( .A1(n7802), .A2(n5568), .ZN(n5434) );
  NAND2_X1 U6948 ( .A1(n5328), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5433) );
  INV_X1 U6949 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6950 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  NAND2_X1 U6951 ( .A1(n5455), .A2(n5438), .ZN(n8899) );
  OR2_X1 U6952 ( .A1(n8899), .A2(n5083), .ZN(n5443) );
  INV_X1 U6953 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U6954 ( .A1(n5597), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6955 ( .A1(n5596), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5439) );
  OAI211_X1 U6956 ( .C1(n5594), .C2(n8900), .A(n5440), .B(n5439), .ZN(n5441)
         );
  INV_X1 U6957 ( .A(n5441), .ZN(n5442) );
  OR2_X1 U6958 ( .A1(n8904), .A2(n8633), .ZN(n5739) );
  NAND2_X1 U6959 ( .A1(n8904), .A2(n8633), .ZN(n5737) );
  NAND2_X1 U6960 ( .A1(n5739), .A2(n5737), .ZN(n8896) );
  INV_X1 U6961 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6962 ( .A1(n5447), .A2(SI_21_), .ZN(n5448) );
  INV_X1 U6963 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8344) );
  INV_X1 U6964 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8539) );
  MUX2_X1 U6965 ( .A(n8344), .B(n8539), .S(n4538), .Z(n5450) );
  INV_X1 U6966 ( .A(SI_22_), .ZN(n5449) );
  NAND2_X1 U6967 ( .A1(n5450), .A2(n5449), .ZN(n5461) );
  INV_X1 U6968 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U6969 ( .A1(n5451), .A2(SI_22_), .ZN(n5452) );
  NAND2_X1 U6970 ( .A1(n5461), .A2(n5452), .ZN(n5462) );
  XNOR2_X1 U6971 ( .A(n5463), .B(n5462), .ZN(n8342) );
  NAND2_X1 U6972 ( .A1(n8342), .A2(n5568), .ZN(n5454) );
  NAND2_X1 U6973 ( .A1(n5328), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5453) );
  INV_X1 U6974 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U6975 ( .A1(n5455), .A2(n8635), .ZN(n5456) );
  AND2_X1 U6976 ( .A1(n5473), .A2(n5456), .ZN(n8885) );
  INV_X1 U6977 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U6978 ( .A1(n5596), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6979 ( .A1(n5598), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5457) );
  OAI211_X1 U6980 ( .C1(n5459), .C2(n10232), .A(n5458), .B(n5457), .ZN(n5460)
         );
  AOI21_X1 U6981 ( .B1(n8885), .B2(n5574), .A(n5460), .ZN(n8893) );
  NAND2_X1 U6982 ( .A1(n9131), .A2(n8893), .ZN(n5727) );
  INV_X1 U6983 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5465) );
  INV_X1 U6984 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5464) );
  MUX2_X1 U6985 ( .A(n5465), .B(n5464), .S(n4538), .Z(n5467) );
  INV_X1 U6986 ( .A(SI_23_), .ZN(n5466) );
  NAND2_X1 U6987 ( .A1(n5467), .A2(n5466), .ZN(n5482) );
  INV_X1 U6988 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U6989 ( .A1(n5468), .A2(SI_23_), .ZN(n5469) );
  XNOR2_X1 U6990 ( .A(n5481), .B(n5480), .ZN(n7929) );
  NAND2_X1 U6991 ( .A1(n7929), .A2(n5568), .ZN(n5471) );
  NAND2_X1 U6992 ( .A1(n5328), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5470) );
  INV_X1 U6993 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U6994 ( .A1(n5473), .A2(n8551), .ZN(n5474) );
  NAND2_X1 U6995 ( .A1(n5486), .A2(n5474), .ZN(n8869) );
  OR2_X1 U6996 ( .A1(n8869), .A2(n5083), .ZN(n5479) );
  INV_X1 U6997 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U6998 ( .A1(n5597), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6999 ( .A1(n5596), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5475) );
  OAI211_X1 U7000 ( .C1(n8870), .C2(n5594), .A(n5476), .B(n5475), .ZN(n5477)
         );
  INV_X1 U7001 ( .A(n5477), .ZN(n5478) );
  NAND2_X1 U7002 ( .A1(n9036), .A2(n8634), .ZN(n5744) );
  NAND2_X1 U7003 ( .A1(n8864), .A2(n8865), .ZN(n8863) );
  INV_X1 U7004 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10187) );
  INV_X1 U7005 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8002) );
  MUX2_X1 U7006 ( .A(n10187), .B(n8002), .S(n6837), .Z(n5495) );
  XNOR2_X1 U7007 ( .A(n5495), .B(SI_24_), .ZN(n5494) );
  XNOR2_X1 U7008 ( .A(n5499), .B(n5494), .ZN(n8001) );
  NAND2_X1 U7009 ( .A1(n8001), .A2(n5568), .ZN(n5485) );
  NAND2_X1 U7010 ( .A1(n5328), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5484) );
  INV_X1 U7011 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U7012 ( .A1(n5486), .A2(n10230), .ZN(n5487) );
  NAND2_X1 U7013 ( .A1(n5506), .A2(n5487), .ZN(n8856) );
  OR2_X1 U7014 ( .A1(n8856), .A2(n5083), .ZN(n5493) );
  INV_X1 U7015 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7016 ( .A1(n5596), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7017 ( .A1(n5597), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5488) );
  OAI211_X1 U7018 ( .C1(n5490), .C2(n5594), .A(n5489), .B(n5488), .ZN(n5491)
         );
  INV_X1 U7019 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U7020 ( .A1(n8858), .A2(n8690), .ZN(n5749) );
  NAND2_X1 U7021 ( .A1(n5748), .A2(n5749), .ZN(n5616) );
  INV_X1 U7022 ( .A(n5494), .ZN(n5498) );
  INV_X1 U7023 ( .A(n5495), .ZN(n5496) );
  NAND2_X1 U7024 ( .A1(n5496), .A2(SI_24_), .ZN(n5497) );
  INV_X1 U7025 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10218) );
  INV_X1 U7026 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8192) );
  MUX2_X1 U7027 ( .A(n10218), .B(n8192), .S(n4538), .Z(n5501) );
  INV_X1 U7028 ( .A(SI_25_), .ZN(n5500) );
  NAND2_X1 U7029 ( .A1(n5501), .A2(n5500), .ZN(n5511) );
  INV_X1 U7030 ( .A(n5501), .ZN(n5502) );
  NAND2_X1 U7031 ( .A1(n5502), .A2(SI_25_), .ZN(n5503) );
  NAND2_X1 U7032 ( .A1(n5511), .A2(n5503), .ZN(n5512) );
  NAND2_X1 U7033 ( .A1(n8188), .A2(n5568), .ZN(n5505) );
  NAND2_X1 U7034 ( .A1(n5328), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5504) );
  INV_X1 U7035 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U7036 ( .A1(n5506), .A2(n8587), .ZN(n5507) );
  NAND2_X1 U7037 ( .A1(n5522), .A2(n5507), .ZN(n8836) );
  INV_X1 U7038 ( .A(n8836), .ZN(n8589) );
  INV_X1 U7039 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U7040 ( .A1(n5596), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7041 ( .A1(n5597), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5508) );
  OAI211_X1 U7042 ( .C1(n8837), .C2(n5594), .A(n5509), .B(n5508), .ZN(n5510)
         );
  NAND2_X1 U7043 ( .A1(n9027), .A2(n8822), .ZN(n5639) );
  INV_X1 U7044 ( .A(n8818), .ZN(n5531) );
  INV_X1 U7045 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5514) );
  INV_X1 U7046 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8193) );
  MUX2_X1 U7047 ( .A(n5514), .B(n8193), .S(n6837), .Z(n5516) );
  INV_X1 U7048 ( .A(SI_26_), .ZN(n5515) );
  NAND2_X1 U7049 ( .A1(n5516), .A2(n5515), .ZN(n5534) );
  INV_X1 U7050 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U7051 ( .A1(n5517), .A2(SI_26_), .ZN(n5518) );
  AND2_X1 U7052 ( .A1(n5534), .A2(n5518), .ZN(n5532) );
  NAND2_X1 U7053 ( .A1(n5328), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5519) );
  INV_X1 U7054 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U7055 ( .A1(n5522), .A2(n8664), .ZN(n5523) );
  NAND2_X1 U7056 ( .A1(n5557), .A2(n5523), .ZN(n8828) );
  OR2_X1 U7057 ( .A1(n8828), .A2(n5083), .ZN(n5529) );
  INV_X1 U7058 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7059 ( .A1(n5596), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7060 ( .A1(n5597), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5524) );
  OAI211_X1 U7061 ( .C1(n5526), .C2(n5594), .A(n5525), .B(n5524), .ZN(n5527)
         );
  INV_X1 U7062 ( .A(n5527), .ZN(n5528) );
  INV_X1 U7063 ( .A(n8820), .ZN(n5530) );
  NAND2_X1 U7064 ( .A1(n5531), .A2(n5530), .ZN(n8798) );
  INV_X1 U7065 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5536) );
  INV_X1 U7066 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8335) );
  MUX2_X1 U7067 ( .A(n5536), .B(n8335), .S(n6834), .Z(n5538) );
  INV_X1 U7068 ( .A(SI_27_), .ZN(n5537) );
  NAND2_X1 U7069 ( .A1(n5538), .A2(n5537), .ZN(n5552) );
  INV_X1 U7070 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U7071 ( .A1(n5539), .A2(SI_27_), .ZN(n5540) );
  AND2_X1 U7072 ( .A1(n5552), .A2(n5540), .ZN(n5550) );
  NAND2_X1 U7073 ( .A1(n8276), .A2(n5568), .ZN(n5542) );
  NAND2_X1 U7074 ( .A1(n5328), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5541) );
  XNOR2_X1 U7075 ( .A(n5557), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U7076 ( .A1(n8543), .A2(n5574), .ZN(n5547) );
  INV_X1 U7077 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U7078 ( .A1(n5596), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7079 ( .A1(n5597), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5543) );
  OAI211_X1 U7080 ( .C1(n8810), .C2(n5594), .A(n5544), .B(n5543), .ZN(n5545)
         );
  INV_X1 U7081 ( .A(n5545), .ZN(n5546) );
  NAND2_X1 U7082 ( .A1(n8814), .A2(n8823), .ZN(n5755) );
  INV_X1 U7083 ( .A(n8799), .ZN(n5636) );
  NOR2_X1 U7084 ( .A1(n8806), .A2(n5636), .ZN(n5548) );
  NAND2_X1 U7085 ( .A1(n8798), .A2(n5548), .ZN(n5549) );
  NAND2_X1 U7086 ( .A1(n5549), .A2(n5754), .ZN(n5862) );
  INV_X1 U7087 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5554) );
  INV_X1 U7088 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5553) );
  MUX2_X1 U7089 ( .A(n5554), .B(n5553), .S(n4538), .Z(n5566) );
  XNOR2_X1 U7090 ( .A(n5566), .B(SI_28_), .ZN(n5563) );
  NAND2_X1 U7091 ( .A1(n8330), .A2(n5568), .ZN(n5556) );
  NAND2_X1 U7092 ( .A1(n5328), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5555) );
  INV_X1 U7093 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8544) );
  INV_X1 U7094 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8459) );
  OAI21_X1 U7095 ( .B1(n5557), .B2(n8544), .A(n8459), .ZN(n5558) );
  INV_X1 U7096 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U7097 ( .A1(n5596), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7098 ( .A1(n5597), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5559) );
  OAI211_X1 U7099 ( .C1(n8790), .C2(n5594), .A(n5560), .B(n5559), .ZN(n5561)
         );
  NAND2_X1 U7100 ( .A1(n8794), .A2(n8803), .ZN(n5756) );
  INV_X1 U7101 ( .A(n5562), .ZN(n5761) );
  AOI21_X1 U7102 ( .B1(n5862), .B2(n5837), .A(n5761), .ZN(n5896) );
  INV_X1 U7103 ( .A(SI_28_), .ZN(n5565) );
  MUX2_X1 U7104 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4538), .Z(n5576) );
  INV_X1 U7105 ( .A(SI_29_), .ZN(n5579) );
  XNOR2_X1 U7106 ( .A(n5576), .B(n5579), .ZN(n5567) );
  NAND2_X1 U7107 ( .A1(n9164), .A2(n5568), .ZN(n5570) );
  NAND2_X1 U7108 ( .A1(n5328), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5569) );
  INV_X1 U7109 ( .A(n5903), .ZN(n5575) );
  INV_X1 U7110 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7111 ( .A1(n5597), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7112 ( .A1(n5596), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5571) );
  OAI211_X1 U7113 ( .C1(n5904), .C2(n5376), .A(n5572), .B(n5571), .ZN(n5573)
         );
  AOI21_X1 U7114 ( .B1(n5575), .B2(n5574), .A(n5573), .ZN(n8460) );
  NAND2_X1 U7115 ( .A1(n8383), .A2(n8460), .ZN(n5766) );
  NAND2_X1 U7116 ( .A1(n5578), .A2(n5579), .ZN(n5577) );
  NAND2_X1 U7117 ( .A1(n5577), .A2(n5576), .ZN(n5582) );
  INV_X1 U7118 ( .A(n5578), .ZN(n5580) );
  NAND2_X1 U7119 ( .A1(n5580), .A2(SI_29_), .ZN(n5581) );
  NAND2_X1 U7120 ( .A1(n5582), .A2(n5581), .ZN(n5607) );
  INV_X1 U7121 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5584) );
  INV_X1 U7122 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n5583) );
  MUX2_X1 U7123 ( .A(n5584), .B(n5583), .S(n6837), .Z(n5586) );
  INV_X1 U7124 ( .A(SI_30_), .ZN(n5585) );
  NAND2_X1 U7125 ( .A1(n5586), .A2(n5585), .ZN(n5605) );
  INV_X1 U7126 ( .A(n5586), .ZN(n5587) );
  NAND2_X1 U7127 ( .A1(n5587), .A2(SI_30_), .ZN(n5588) );
  NAND2_X1 U7128 ( .A1(n5605), .A2(n5588), .ZN(n5606) );
  NAND2_X1 U7129 ( .A1(n9160), .A2(n5568), .ZN(n5590) );
  NAND2_X1 U7130 ( .A1(n5328), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5589) );
  INV_X1 U7131 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7132 ( .A1(n5596), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7133 ( .A1(n5597), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7134 ( .C1(n5594), .C2(n5593), .A(n5592), .B(n5591), .ZN(n8779)
         );
  OR2_X1 U7135 ( .A1(n8779), .A2(n7803), .ZN(n5595) );
  OAI21_X1 U7136 ( .B1(n9107), .B2(n5595), .A(n5766), .ZN(n5604) );
  INV_X1 U7137 ( .A(n5595), .ZN(n5603) );
  INV_X1 U7138 ( .A(n9107), .ZN(n5602) );
  NAND2_X1 U7139 ( .A1(n5596), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7140 ( .A1(n5597), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7141 ( .A1(n5598), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5599) );
  AND3_X1 U7142 ( .A1(n5601), .A2(n5600), .A3(n5599), .ZN(n5900) );
  OAI22_X1 U7143 ( .A1(n5894), .A2(n5604), .B1(n5603), .B2(n5764), .ZN(n5612)
         );
  MUX2_X1 U7144 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6834), .Z(n5609) );
  INV_X1 U7145 ( .A(SI_31_), .ZN(n5608) );
  XNOR2_X1 U7146 ( .A(n5609), .B(n5608), .ZN(n5610) );
  AND2_X1 U7147 ( .A1(n9103), .A2(n8779), .ZN(n5776) );
  INV_X1 U7148 ( .A(n5900), .ZN(n8685) );
  NOR2_X1 U7149 ( .A1(n9107), .A2(n8685), .ZN(n5770) );
  NOR2_X1 U7150 ( .A1(n9103), .A2(n8779), .ZN(n5615) );
  AOI21_X1 U7151 ( .B1(n5612), .B2(n5773), .A(n5615), .ZN(n5613) );
  XNOR2_X1 U7152 ( .A(n5613), .B(n5860), .ZN(n5614) );
  AOI21_X1 U7153 ( .B1(n8432), .B2(n5863), .A(n5614), .ZN(n5794) );
  INV_X1 U7154 ( .A(n5615), .ZN(n5779) );
  NAND2_X1 U7155 ( .A1(n5779), .A2(n5764), .ZN(n5774) );
  INV_X1 U7156 ( .A(n5774), .ZN(n5630) );
  NAND2_X1 U7157 ( .A1(n5734), .A2(n5736), .ZN(n8914) );
  INV_X1 U7158 ( .A(n8078), .ZN(n8075) );
  INV_X1 U7159 ( .A(n7935), .ZN(n7939) );
  NAND2_X1 U7160 ( .A1(n5682), .A2(n4439), .ZN(n7804) );
  NAND2_X1 U7161 ( .A1(n5810), .A2(n7192), .ZN(n5661) );
  AND2_X1 U7162 ( .A1(n7194), .A2(n5661), .ZN(n7759) );
  INV_X1 U7163 ( .A(n5811), .ZN(n7196) );
  NAND4_X1 U7164 ( .A1(n7759), .A2(n7196), .A3(n7615), .A4(n7076), .ZN(n5620)
         );
  INV_X1 U7165 ( .A(n7384), .ZN(n5619) );
  INV_X1 U7166 ( .A(n5618), .ZN(n5654) );
  NAND2_X1 U7167 ( .A1(n5654), .A2(n5649), .ZN(n7604) );
  NOR4_X1 U7168 ( .A1(n5620), .A2(n5619), .A3(n7604), .A4(n7312), .ZN(n5621)
         );
  INV_X1 U7169 ( .A(n5818), .ZN(n7452) );
  NAND4_X1 U7170 ( .A1(n5621), .A2(n5192), .A3(n5163), .A4(n7452), .ZN(n5622)
         );
  NOR4_X1 U7171 ( .A1(n7964), .A2(n7939), .A3(n7804), .A4(n5622), .ZN(n5623)
         );
  NAND4_X1 U7172 ( .A1(n8265), .A2(n5294), .A3(n8075), .A4(n5623), .ZN(n5624)
         );
  NOR4_X1 U7173 ( .A1(n8940), .A2(n8974), .A3(n8317), .A4(n5624), .ZN(n5625)
         );
  NAND3_X1 U7174 ( .A1(n8923), .A2(n5625), .A3(n4702), .ZN(n5626) );
  NOR4_X1 U7175 ( .A1(n8879), .A2(n8896), .A3(n8914), .A4(n5626), .ZN(n5627)
         );
  NAND4_X1 U7176 ( .A1(n8840), .A2(n8852), .A3(n8865), .A4(n5627), .ZN(n5628)
         );
  NOR4_X1 U7177 ( .A1(n5885), .A2(n8806), .A3(n8820), .A4(n5628), .ZN(n5629)
         );
  NAND4_X1 U7178 ( .A1(n5630), .A2(n5773), .A3(n5895), .A4(n5629), .ZN(n5631)
         );
  XNOR2_X1 U7179 ( .A(n5631), .B(n8929), .ZN(n5632) );
  OAI22_X1 U7180 ( .A1(n5632), .A2(n7087), .B1(n7076), .B2(n5864), .ZN(n5784)
         );
  INV_X1 U7181 ( .A(n5756), .ZN(n5763) );
  OR2_X1 U7182 ( .A1(n7088), .A2(n8929), .ZN(n5777) );
  NAND2_X1 U7183 ( .A1(n5635), .A2(n5633), .ZN(n5634) );
  NAND2_X1 U7184 ( .A1(n5634), .A2(n5762), .ZN(n5752) );
  INV_X1 U7185 ( .A(n5635), .ZN(n5637) );
  AOI22_X1 U7186 ( .A1(n5752), .A2(n5637), .B1(n5636), .B2(n5762), .ZN(n5638)
         );
  AND2_X1 U7187 ( .A1(n5638), .A2(n8800), .ZN(n5760) );
  INV_X1 U7188 ( .A(n5639), .ZN(n5640) );
  OAI21_X1 U7189 ( .B1(n8820), .B2(n5640), .A(n5777), .ZN(n5753) );
  OAI211_X1 U7190 ( .C1(n8958), .C2(n5642), .A(n5641), .B(n5729), .ZN(n5644)
         );
  AND2_X1 U7191 ( .A1(n8960), .A2(n8980), .ZN(n5643) );
  MUX2_X1 U7192 ( .A(n5644), .B(n5643), .S(n5762), .Z(n5645) );
  INV_X1 U7193 ( .A(n5645), .ZN(n5720) );
  NAND2_X1 U7194 ( .A1(n5655), .A2(n5654), .ZN(n5647) );
  NAND2_X1 U7195 ( .A1(n7444), .A2(n5649), .ZN(n5646) );
  MUX2_X1 U7196 ( .A(n5647), .B(n5646), .S(n5777), .Z(n5652) );
  AND2_X1 U7197 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  OAI211_X1 U7198 ( .C1(n5652), .C2(n5650), .A(n5670), .B(n7444), .ZN(n5651)
         );
  INV_X1 U7199 ( .A(n5651), .ZN(n5659) );
  INV_X1 U7200 ( .A(n5652), .ZN(n5667) );
  NAND2_X1 U7201 ( .A1(n5654), .A2(n5653), .ZN(n5657) );
  NAND2_X1 U7202 ( .A1(n5671), .A2(n5655), .ZN(n5656) );
  AOI21_X1 U7203 ( .B1(n5667), .B2(n5657), .A(n5656), .ZN(n5658) );
  NAND2_X1 U7204 ( .A1(n5662), .A2(n5661), .ZN(n5664) );
  NOR2_X1 U7205 ( .A1(n5664), .A2(n7803), .ZN(n5663) );
  INV_X1 U7206 ( .A(n5664), .ZN(n5665) );
  MUX2_X1 U7207 ( .A(n4480), .B(n5666), .S(n5762), .Z(n5668) );
  NAND3_X1 U7208 ( .A1(n5668), .A2(n5667), .A3(n7317), .ZN(n5669) );
  MUX2_X1 U7209 ( .A(n5671), .B(n5670), .S(n5777), .Z(n5672) );
  AND2_X1 U7210 ( .A1(n5163), .A2(n5672), .ZN(n5673) );
  INV_X1 U7211 ( .A(n5674), .ZN(n5675) );
  NOR2_X1 U7212 ( .A1(n7741), .A2(n5675), .ZN(n5678) );
  INV_X1 U7213 ( .A(n5676), .ZN(n5677) );
  AOI21_X1 U7214 ( .B1(n5688), .B2(n5678), .A(n5677), .ZN(n5681) );
  AND2_X1 U7215 ( .A1(n5682), .A2(n5679), .ZN(n5680) );
  MUX2_X1 U7216 ( .A(n5681), .B(n5680), .S(n5777), .Z(n5685) );
  AND2_X1 U7217 ( .A1(n5689), .A2(n5682), .ZN(n5683) );
  MUX2_X1 U7218 ( .A(n4439), .B(n5683), .S(n5762), .Z(n5684) );
  NAND2_X1 U7219 ( .A1(n5684), .A2(n5686), .ZN(n5690) );
  AOI21_X1 U7220 ( .B1(n5685), .B2(n4439), .A(n5690), .ZN(n5700) );
  NAND2_X1 U7221 ( .A1(n8077), .A2(n5686), .ZN(n5693) );
  OAI211_X1 U7222 ( .C1(n5691), .C2(n5690), .A(n5694), .B(n5689), .ZN(n5692)
         );
  MUX2_X1 U7223 ( .A(n5693), .B(n5692), .S(n5777), .Z(n5699) );
  NAND2_X1 U7224 ( .A1(n5701), .A2(n8077), .ZN(n5696) );
  NAND2_X1 U7225 ( .A1(n5702), .A2(n5694), .ZN(n5695) );
  MUX2_X1 U7226 ( .A(n5696), .B(n5695), .S(n5762), .Z(n5697) );
  INV_X1 U7227 ( .A(n5697), .ZN(n5698) );
  OAI21_X1 U7228 ( .B1(n5700), .B2(n5699), .A(n5698), .ZN(n5704) );
  MUX2_X1 U7229 ( .A(n5702), .B(n5701), .S(n5762), .Z(n5703) );
  NAND3_X1 U7230 ( .A1(n5704), .A2(n5294), .A3(n5703), .ZN(n5707) );
  MUX2_X1 U7231 ( .A(n5705), .B(n8266), .S(n5777), .Z(n5706) );
  NAND3_X1 U7232 ( .A1(n5707), .A2(n8265), .A3(n5706), .ZN(n5711) );
  MUX2_X1 U7233 ( .A(n5709), .B(n5708), .S(n5762), .Z(n5710) );
  NAND3_X1 U7234 ( .A1(n5711), .A2(n8319), .A3(n5710), .ZN(n5718) );
  INV_X1 U7235 ( .A(n5712), .ZN(n5715) );
  INV_X1 U7236 ( .A(n5713), .ZN(n5714) );
  MUX2_X1 U7237 ( .A(n5715), .B(n5714), .S(n5777), .Z(n5716) );
  INV_X1 U7238 ( .A(n5716), .ZN(n5717) );
  INV_X1 U7239 ( .A(n5733), .ZN(n5721) );
  AOI21_X1 U7240 ( .B1(n5730), .B2(n5731), .A(n5721), .ZN(n5724) );
  INV_X1 U7241 ( .A(n5722), .ZN(n5723) );
  OAI211_X1 U7242 ( .C1(n5724), .C2(n5723), .A(n5739), .B(n5734), .ZN(n5725)
         );
  NAND3_X1 U7243 ( .A1(n5725), .A2(n5727), .A3(n5737), .ZN(n5726) );
  AND2_X1 U7244 ( .A1(n5726), .A2(n5740), .ZN(n5728) );
  MUX2_X1 U7245 ( .A(n5728), .B(n5727), .S(n5762), .Z(n5743) );
  NAND2_X1 U7246 ( .A1(n5730), .A2(n5729), .ZN(n5732) );
  NAND3_X1 U7247 ( .A1(n5732), .A2(n8912), .A3(n5731), .ZN(n5735) );
  NAND3_X1 U7248 ( .A1(n5735), .A2(n5734), .A3(n5733), .ZN(n5738) );
  NAND3_X1 U7249 ( .A1(n5738), .A2(n5737), .A3(n5736), .ZN(n5741) );
  NAND4_X1 U7250 ( .A1(n5741), .A2(n5740), .A3(n5762), .A4(n5739), .ZN(n5742)
         );
  NAND3_X1 U7251 ( .A1(n5743), .A2(n8865), .A3(n5742), .ZN(n5747) );
  MUX2_X1 U7252 ( .A(n5745), .B(n5744), .S(n5777), .Z(n5746) );
  NAND3_X1 U7253 ( .A1(n8852), .A2(n5747), .A3(n5746), .ZN(n5751) );
  MUX2_X1 U7254 ( .A(n5749), .B(n5748), .S(n5777), .Z(n5750) );
  INV_X1 U7255 ( .A(n5754), .ZN(n5758) );
  NAND2_X1 U7256 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  MUX2_X1 U7257 ( .A(n5758), .B(n5757), .S(n5777), .Z(n5759) );
  INV_X1 U7258 ( .A(n5764), .ZN(n5771) );
  INV_X1 U7259 ( .A(n5765), .ZN(n5768) );
  INV_X1 U7260 ( .A(n5766), .ZN(n5767) );
  MUX2_X1 U7261 ( .A(n5768), .B(n5767), .S(n5777), .Z(n5769) );
  NOR4_X1 U7262 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n5782)
         );
  INV_X1 U7263 ( .A(n5773), .ZN(n5775) );
  MUX2_X1 U7264 ( .A(n5775), .B(n5774), .S(n5777), .Z(n5781) );
  INV_X1 U7265 ( .A(n5776), .ZN(n5778) );
  MUX2_X1 U7266 ( .A(n5779), .B(n5778), .S(n5777), .Z(n5780) );
  OAI21_X1 U7267 ( .B1(n5782), .B2(n5781), .A(n5780), .ZN(n5783) );
  NOR2_X1 U7268 ( .A1(n5785), .A2(n7088), .ZN(n5786) );
  NAND2_X1 U7269 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  NAND2_X1 U7270 ( .A1(n5789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  INV_X1 U7271 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7272 ( .A1(n5791), .A2(n5790), .ZN(n5795) );
  OR2_X1 U7273 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  NAND2_X1 U7274 ( .A1(n5795), .A2(n5792), .ZN(n5852) );
  OR2_X1 U7275 ( .A1(n5852), .A2(n4420), .ZN(n6889) );
  NAND2_X1 U7276 ( .A1(n5795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7277 ( .A1(n5797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5798) );
  MUX2_X1 U7278 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5798), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5799) );
  AND2_X1 U7279 ( .A1(n5024), .A2(n5799), .ZN(n9952) );
  NAND2_X1 U7280 ( .A1(n5800), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5801) );
  MUX2_X1 U7281 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5801), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5802) );
  NAND2_X1 U7282 ( .A1(n5802), .A2(n5797), .ZN(n8189) );
  INV_X1 U7283 ( .A(n8189), .ZN(n9953) );
  AND2_X1 U7284 ( .A1(n9952), .A2(n9953), .ZN(n5803) );
  INV_X1 U7285 ( .A(n9957), .ZN(n5804) );
  NAND2_X1 U7286 ( .A1(n5805), .A2(n7087), .ZN(n7085) );
  OR2_X1 U7287 ( .A1(n6913), .A2(n7085), .ZN(n8977) );
  OAI21_X1 U7288 ( .B1(n6889), .B2(n5805), .A(P2_B_REG_SCAN_IN), .ZN(n5806) );
  INV_X1 U7289 ( .A(n5806), .ZN(n5807) );
  NAND2_X1 U7290 ( .A1(n4981), .A2(n5807), .ZN(n5808) );
  NAND2_X1 U7291 ( .A1(n5809), .A2(n5808), .ZN(P2_U3244) );
  INV_X1 U7292 ( .A(n7192), .ZN(n7754) );
  NAND2_X1 U7293 ( .A1(n5810), .A2(n7754), .ZN(n7191) );
  OR2_X1 U7294 ( .A1(n5046), .A2(n7092), .ZN(n5812) );
  NAND2_X1 U7295 ( .A1(n7190), .A2(n5812), .ZN(n7614) );
  INV_X1 U7296 ( .A(n7615), .ZN(n7613) );
  NAND2_X1 U7297 ( .A1(n7614), .A2(n7613), .ZN(n7612) );
  INV_X1 U7298 ( .A(n9962), .ZN(n7623) );
  OR2_X1 U7299 ( .A1(n7623), .A2(n8705), .ZN(n5813) );
  NAND2_X1 U7300 ( .A1(n7612), .A2(n5813), .ZN(n7313) );
  NAND2_X1 U7301 ( .A1(n7313), .A2(n7312), .ZN(n7311) );
  OR2_X1 U7302 ( .A1(n4823), .A2(n10348), .ZN(n5814) );
  NAND2_X1 U7303 ( .A1(n7311), .A2(n5814), .ZN(n7600) );
  INV_X1 U7304 ( .A(n8704), .ZN(n7227) );
  NAND2_X1 U7305 ( .A1(n7227), .A2(n10344), .ZN(n5815) );
  AND2_X1 U7306 ( .A1(n10342), .A2(n7440), .ZN(n5817) );
  NAND2_X1 U7307 ( .A1(n7384), .A2(n8594), .ZN(n5816) );
  OR2_X1 U7308 ( .A1(n7695), .A2(n7493), .ZN(n5819) );
  INV_X1 U7309 ( .A(n7377), .ZN(n8701) );
  INV_X1 U7310 ( .A(n7646), .ZN(n8700) );
  NAND2_X1 U7311 ( .A1(n7771), .A2(n8700), .ZN(n5821) );
  INV_X1 U7312 ( .A(n7941), .ZN(n8699) );
  OR2_X1 U7313 ( .A1(n9929), .A2(n8699), .ZN(n5822) );
  NAND2_X1 U7314 ( .A1(n5823), .A2(n7939), .ZN(n7934) );
  INV_X1 U7315 ( .A(n7859), .ZN(n8698) );
  NAND2_X1 U7316 ( .A1(n7961), .A2(n8698), .ZN(n5824) );
  NAND2_X1 U7317 ( .A1(n7963), .A2(n7964), .ZN(n5826) );
  INV_X1 U7318 ( .A(n8081), .ZN(n8697) );
  NAND2_X1 U7319 ( .A1(n8043), .A2(n8697), .ZN(n5825) );
  INV_X1 U7320 ( .A(n8237), .ZN(n8696) );
  INV_X1 U7321 ( .A(n8269), .ZN(n8695) );
  NAND2_X1 U7322 ( .A1(n9092), .A2(n8695), .ZN(n5827) );
  INV_X1 U7323 ( .A(n8322), .ZN(n8694) );
  OAI22_X1 U7324 ( .A1(n8259), .A2(n8265), .B1(n8694), .B2(n9087), .ZN(n8318)
         );
  NAND2_X1 U7325 ( .A1(n8318), .A2(n8317), .ZN(n8316) );
  INV_X1 U7326 ( .A(n8978), .ZN(n8693) );
  OR2_X1 U7327 ( .A1(n9080), .A2(n8693), .ZN(n5828) );
  NAND2_X1 U7328 ( .A1(n8316), .A2(n5828), .ZN(n8969) );
  INV_X1 U7329 ( .A(n8956), .ZN(n8692) );
  INV_X1 U7330 ( .A(n8980), .ZN(n8944) );
  NAND2_X1 U7331 ( .A1(n9061), .A2(n5830), .ZN(n5832) );
  INV_X1 U7332 ( .A(n9061), .ZN(n8939) );
  INV_X1 U7333 ( .A(n8658), .ZN(n8946) );
  NAND2_X1 U7334 ( .A1(n8920), .A2(n5833), .ZN(n5834) );
  INV_X1 U7335 ( .A(n9143), .ZN(n8926) );
  NAND2_X1 U7336 ( .A1(n5834), .A2(n4967), .ZN(n8907) );
  INV_X1 U7337 ( .A(n8892), .ZN(n8924) );
  INV_X1 U7338 ( .A(n8633), .ZN(n8915) );
  NAND2_X1 U7339 ( .A1(n8868), .A2(n8867), .ZN(n9034) );
  NAND2_X1 U7340 ( .A1(n9034), .A2(n4972), .ZN(n8851) );
  NOR2_X2 U7341 ( .A1(n8851), .A2(n8852), .ZN(n8850) );
  INV_X1 U7342 ( .A(n8822), .ZN(n8689) );
  INV_X1 U7343 ( .A(n9115), .ZN(n5836) );
  INV_X1 U7344 ( .A(n8823), .ZN(n8687) );
  XNOR2_X1 U7345 ( .A(n5886), .B(n5837), .ZN(n8788) );
  NOR4_X1 U7346 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5846) );
  NOR4_X1 U7347 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5845) );
  INV_X1 U7348 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10289) );
  INV_X1 U7349 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10140) );
  INV_X1 U7350 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10181) );
  INV_X1 U7351 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10105) );
  NAND4_X1 U7352 ( .A1(n10289), .A2(n10140), .A3(n10181), .A4(n10105), .ZN(
        n5843) );
  NOR4_X1 U7353 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5841) );
  NOR4_X1 U7354 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5840) );
  NOR4_X1 U7355 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5839) );
  NOR4_X1 U7356 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5838) );
  NAND4_X1 U7357 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n5842)
         );
  NOR4_X1 U7358 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5843), .A4(n5842), .ZN(n5844) );
  AND3_X1 U7359 ( .A1(n5846), .A2(n5845), .A3(n5844), .ZN(n5851) );
  INV_X1 U7360 ( .A(n9949), .ZN(n8023) );
  INV_X1 U7361 ( .A(P2_B_REG_SCAN_IN), .ZN(n5847) );
  AOI22_X1 U7362 ( .A1(P2_B_REG_SCAN_IN), .A2(n8023), .B1(n9949), .B2(n5847), 
        .ZN(n5848) );
  INV_X1 U7363 ( .A(n5848), .ZN(n5849) );
  NAND2_X1 U7364 ( .A1(n8189), .A2(n5849), .ZN(n5850) );
  NOR2_X1 U7365 ( .A1(n5851), .A2(n9946), .ZN(n7075) );
  INV_X1 U7366 ( .A(n5852), .ZN(n5855) );
  INV_X1 U7367 ( .A(n5853), .ZN(n7082) );
  NOR2_X1 U7368 ( .A1(n7085), .A2(n7082), .ZN(n5854) );
  NOR2_X1 U7369 ( .A1(n7077), .A2(n4420), .ZN(n5875) );
  OR2_X1 U7370 ( .A1(n9949), .A2(n9952), .ZN(n5857) );
  OAI22_X1 U7371 ( .A1(n9946), .A2(P2_D_REG_1__SCAN_IN), .B1(n9953), .B2(n9952), .ZN(n5890) );
  AND2_X1 U7372 ( .A1(n5892), .A2(n5890), .ZN(n5877) );
  NAND3_X1 U7373 ( .A1(n5875), .A2(n7073), .A3(n5877), .ZN(n5858) );
  INV_X2 U7374 ( .A(n9994), .ZN(n9996) );
  NAND2_X1 U7375 ( .A1(n7087), .A2(n7733), .ZN(n7089) );
  XNOR2_X1 U7376 ( .A(n7089), .B(n8343), .ZN(n5859) );
  OR2_X1 U7377 ( .A1(n5859), .A2(n5860), .ZN(n8972) );
  AND2_X1 U7378 ( .A1(n7733), .A2(n5860), .ZN(n5861) );
  NAND2_X1 U7379 ( .A1(n8343), .A2(n5861), .ZN(n9096) );
  NAND2_X1 U7380 ( .A1(n8972), .A2(n9096), .ZN(n9985) );
  NAND2_X1 U7381 ( .A1(n9996), .A2(n9985), .ZN(n9060) );
  OR2_X1 U7382 ( .A1(n8788), .A2(n9060), .ZN(n5873) );
  XNOR2_X1 U7383 ( .A(n5862), .B(n5885), .ZN(n5867) );
  NAND2_X1 U7384 ( .A1(n5864), .A2(n5863), .ZN(n8982) );
  INV_X1 U7385 ( .A(n6913), .ZN(n5865) );
  NOR2_X2 U7386 ( .A1(n7085), .A2(n5865), .ZN(n8945) );
  OAI22_X1 U7387 ( .A1(n8823), .A2(n8977), .B1(n8460), .B2(n8979), .ZN(n5866)
         );
  NAND2_X1 U7388 ( .A1(n7622), .A2(n9962), .ZN(n9958) );
  INV_X1 U7389 ( .A(n7771), .ZN(n7745) );
  NAND2_X1 U7390 ( .A1(n7746), .A2(n7745), .ZN(n7807) );
  INV_X1 U7391 ( .A(n8043), .ZN(n7973) );
  INV_X1 U7392 ( .A(n8087), .ZN(n9980) );
  INV_X1 U7393 ( .A(n9080), .ZN(n8678) );
  INV_X1 U7394 ( .A(n8993), .ZN(n9073) );
  NAND2_X1 U7395 ( .A1(n8988), .A2(n9073), .ZN(n8987) );
  INV_X1 U7396 ( .A(n9049), .ZN(n8911) );
  INV_X1 U7397 ( .A(n8811), .ZN(n5869) );
  INV_X1 U7398 ( .A(n8794), .ZN(n5884) );
  INV_X1 U7399 ( .A(n9981), .ZN(n9959) );
  OAI211_X1 U7400 ( .C1(n5869), .C2(n5884), .A(n9959), .B(n5905), .ZN(n8791)
         );
  NAND2_X1 U7401 ( .A1(n8797), .A2(n8791), .ZN(n5879) );
  MUX2_X1 U7402 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n5879), .S(n9996), .Z(n5870)
         );
  INV_X1 U7403 ( .A(n5870), .ZN(n5871) );
  OR2_X1 U7404 ( .A1(n7102), .A2(n7082), .ZN(n9979) );
  NAND2_X1 U7405 ( .A1(n5873), .A2(n5872), .ZN(P2_U3548) );
  INV_X1 U7406 ( .A(n7073), .ZN(n5874) );
  NAND2_X1 U7407 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  INV_X1 U7408 ( .A(n5877), .ZN(n5878) );
  INV_X2 U7409 ( .A(n9987), .ZN(n9155) );
  NAND2_X1 U7410 ( .A1(n9155), .A2(n9985), .ZN(n9146) );
  OR2_X1 U7411 ( .A1(n8788), .A2(n9146), .ZN(n5883) );
  MUX2_X1 U7412 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n5879), .S(n9155), .Z(n5880)
         );
  INV_X1 U7413 ( .A(n5880), .ZN(n5881) );
  INV_X1 U7414 ( .A(n9979), .ZN(n9093) );
  NAND2_X1 U7415 ( .A1(n5883), .A2(n5882), .ZN(P2_U3516) );
  XNOR2_X1 U7416 ( .A(n5888), .B(n5887), .ZN(n8386) );
  INV_X1 U7417 ( .A(n5889), .ZN(n5891) );
  INV_X1 U7418 ( .A(n5890), .ZN(n7072) );
  NAND2_X1 U7419 ( .A1(n5891), .A2(n7072), .ZN(n5908) );
  OR2_X1 U7420 ( .A1(n7089), .A2(n8929), .ZN(n7938) );
  AND2_X1 U7421 ( .A1(n8972), .A2(n7938), .ZN(n5893) );
  NOR2_X2 U7422 ( .A1(n9944), .A2(n5893), .ZN(n9940) );
  INV_X1 U7423 ( .A(n9940), .ZN(n5915) );
  INV_X1 U7424 ( .A(n5894), .ZN(n5898) );
  OR2_X1 U7425 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  NAND2_X1 U7426 ( .A1(n5898), .A2(n5897), .ZN(n5902) );
  INV_X1 U7427 ( .A(n6912), .ZN(n8277) );
  NAND2_X1 U7428 ( .A1(n8277), .A2(P2_B_REG_SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7429 ( .A1(n8945), .A2(n5899), .ZN(n8778) );
  OAI22_X1 U7430 ( .A1(n8803), .A2(n8977), .B1(n5900), .B2(n8778), .ZN(n5901)
         );
  OR2_X1 U7431 ( .A1(n7102), .A2(n7733), .ZN(n7096) );
  NOR2_X2 U7432 ( .A1(n8998), .A2(n7096), .ZN(n9002) );
  OAI22_X1 U7433 ( .A1(n9001), .A2(n5904), .B1(n5903), .B2(n8989), .ZN(n5911)
         );
  INV_X1 U7434 ( .A(n5905), .ZN(n5907) );
  INV_X1 U7435 ( .A(n8383), .ZN(n5906) );
  OAI211_X1 U7436 ( .C1(n5906), .C2(n5907), .A(n9959), .B(n8777), .ZN(n8377)
         );
  INV_X1 U7437 ( .A(n5908), .ZN(n5909) );
  NAND2_X1 U7438 ( .A1(n5909), .A2(n8929), .ZN(n8995) );
  NOR2_X1 U7439 ( .A1(n8377), .A2(n8995), .ZN(n5910) );
  AOI211_X1 U7440 ( .C1(n9002), .C2(n8383), .A(n5911), .B(n5910), .ZN(n5912)
         );
  OAI21_X1 U7441 ( .B1(n8378), .B2(n8998), .A(n5912), .ZN(n5913) );
  OAI21_X1 U7442 ( .B1(n8386), .B2(n5915), .A(n5914), .ZN(P2_U3267) );
  NOR2_X1 U7443 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5922) );
  NOR2_X1 U7444 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5921) );
  NAND4_X1 U7445 ( .A1(n5962), .A2(n5922), .A3(n5921), .A4(n5961), .ZN(n5924)
         );
  NAND4_X1 U7446 ( .A1(n6187), .A2(n6219), .A3(n6235), .A4(n6479), .ZN(n5923)
         );
  INV_X1 U7447 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6532) );
  OR2_X1 U7448 ( .A1(n5927), .A2(n6127), .ZN(n5926) );
  OAI21_X1 U7449 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7450 ( .A1(n9164), .A2(n6342), .ZN(n5932) );
  NAND2_X1 U7451 ( .A1(n6344), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7452 ( .A1(n6344), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7453 ( .A1(n8188), .A2(n6342), .ZN(n5936) );
  NAND2_X1 U7454 ( .A1(n6344), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5935) );
  NOR2_X2 U7455 ( .A1(n5937), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9641) );
  XNOR2_X2 U7456 ( .A(n5940), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5941) );
  INV_X1 U7457 ( .A(n5941), .ZN(n5946) );
  NAND2_X1 U7458 ( .A1(n6355), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5951) );
  INV_X1 U7459 ( .A(n9646), .ZN(n5947) );
  AND2_X2 U7460 ( .A1(n5947), .A2(n5941), .ZN(n5999) );
  NAND2_X1 U7461 ( .A1(n6356), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5950) );
  AND2_X4 U7462 ( .A1(n9646), .A2(n5941), .ZN(n6020) );
  NAND2_X1 U7463 ( .A1(n6056), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6074) );
  INV_X1 U7464 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6100) );
  INV_X1 U7465 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10166) );
  INV_X1 U7466 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6169) );
  INV_X1 U7467 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U7468 ( .A1(n6192), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6207) );
  INV_X1 U7469 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6206) );
  INV_X1 U7470 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6225) );
  INV_X1 U7471 ( .A(n6299), .ZN(n5943) );
  NAND2_X1 U7472 ( .A1(n5943), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6292) );
  INV_X1 U7473 ( .A(n6292), .ZN(n5944) );
  NAND2_X1 U7474 ( .A1(n5944), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5954) );
  INV_X1 U7475 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U7476 ( .A1(n6292), .A2(n9203), .ZN(n5945) );
  AND2_X1 U7477 ( .A1(n5954), .A2(n5945), .ZN(n9394) );
  NAND2_X1 U7478 ( .A1(n6020), .A2(n9394), .ZN(n5949) );
  INV_X4 U7479 ( .A(n6273), .ZN(n6358) );
  NAND2_X1 U7480 ( .A1(n6358), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5948) );
  NAND4_X1 U7481 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n9414)
         );
  NAND2_X1 U7482 ( .A1(n6355), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7483 ( .A1(n6358), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5958) );
  INV_X1 U7484 ( .A(n5954), .ZN(n5952) );
  INV_X1 U7485 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7486 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7487 ( .A1(n6020), .A2(n9377), .ZN(n5957) );
  NAND2_X1 U7488 ( .A1(n6356), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5956) );
  OAI21_X1 U7489 ( .B1(n9565), .B2(n8516), .A(n9361), .ZN(n5975) );
  NOR2_X1 U7490 ( .A1(n8517), .A2(n9399), .ZN(n5960) );
  OR2_X1 U7491 ( .A1(n9565), .A2(n5960), .ZN(n5974) );
  NAND2_X1 U7492 ( .A1(n6128), .A2(n5961), .ZN(n6142) );
  NAND2_X1 U7493 ( .A1(n5962), .A2(n6187), .ZN(n5963) );
  INV_X1 U7494 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7495 ( .A1(n6200), .A2(n5964), .ZN(n6218) );
  NAND2_X1 U7496 ( .A1(n5972), .A2(n5966), .ZN(n5967) );
  NAND2_X1 U7497 ( .A1(n6478), .A2(n6479), .ZN(n5968) );
  INV_X1 U7498 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6379) );
  OR2_X1 U7499 ( .A1(n6127), .A2(n6379), .ZN(n5969) );
  INV_X1 U7500 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5970) );
  MUX2_X1 U7501 ( .A(n5975), .B(n5974), .S(n7007), .Z(n6321) );
  INV_X1 U7502 ( .A(n6321), .ZN(n6323) );
  NAND2_X1 U7503 ( .A1(n8276), .A2(n6342), .ZN(n5977) );
  NAND2_X1 U7504 ( .A1(n6344), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7505 ( .A1(n6355), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7506 ( .A1(n6358), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5980) );
  XNOR2_X1 U7507 ( .A(n6330), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U7508 ( .A1(n6020), .A2(n9370), .ZN(n5979) );
  NAND2_X1 U7509 ( .A1(n6356), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5978) );
  NAND4_X1 U7510 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n9353)
         );
  NAND2_X1 U7511 ( .A1(n9561), .A2(n9381), .ZN(n6464) );
  NAND2_X1 U7512 ( .A1(n9565), .A2(n8516), .ZN(n5983) );
  NAND2_X1 U7513 ( .A1(n8517), .A2(n9399), .ZN(n5982) );
  MUX2_X1 U7514 ( .A(n5983), .B(n5982), .S(n7007), .Z(n6320) );
  NAND2_X1 U7515 ( .A1(n4538), .A2(SI_0_), .ZN(n5984) );
  XNOR2_X1 U7516 ( .A(n5984), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9653) );
  OAI21_X2 U7517 ( .B1(n6063), .B2(n5986), .A(n5985), .ZN(n7457) );
  INV_X1 U7518 ( .A(n7457), .ZN(n7022) );
  NAND2_X1 U7519 ( .A1(n6020), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7520 ( .A1(n6000), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7521 ( .A1(n5998), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7522 ( .A(n5990), .B(P1_IR_REG_1__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U7523 ( .A1(n5999), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7524 ( .A1(n5998), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5991) );
  AND2_X1 U7525 ( .A1(n5992), .A2(n5991), .ZN(n5994) );
  NAND2_X1 U7526 ( .A1(n6000), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5993) );
  NAND3_X2 U7527 ( .A1(n5995), .A2(n5994), .A3(n5993), .ZN(n6564) );
  NAND2_X1 U7528 ( .A1(n5997), .A2(n6490), .ZN(n7293) );
  NAND2_X1 U7529 ( .A1(n6020), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7530 ( .A1(n5998), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7531 ( .A1(n5999), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7532 ( .A1(n6000), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6001) );
  NAND4_X2 U7533 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n6573)
         );
  OR2_X1 U7534 ( .A1(n6005), .A2(n6127), .ZN(n6012) );
  XNOR2_X1 U7535 ( .A(n6012), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7123) );
  NAND2_X1 U7536 ( .A1(n7110), .A2(n7123), .ZN(n6006) );
  NAND2_X1 U7537 ( .A1(n6573), .A2(n7566), .ZN(n6497) );
  NAND2_X1 U7538 ( .A1(n5998), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7539 ( .A1(n5999), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6009) );
  INV_X1 U7540 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10165) );
  NAND2_X1 U7541 ( .A1(n6020), .A2(n10165), .ZN(n6008) );
  NAND2_X1 U7542 ( .A1(n6025), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6016) );
  INV_X1 U7543 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7544 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  NAND2_X1 U7545 ( .A1(n6013), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6014) );
  XNOR2_X1 U7546 ( .A(n6014), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U7547 ( .A1(n7110), .A2(n7175), .ZN(n6015) );
  INV_X1 U7548 ( .A(n7548), .ZN(n9848) );
  NAND2_X1 U7549 ( .A1(n9323), .A2(n9848), .ZN(n6417) );
  NAND2_X2 U7550 ( .A1(n6421), .A2(n6417), .ZN(n7543) );
  INV_X1 U7551 ( .A(n7543), .ZN(n6017) );
  NAND2_X1 U7552 ( .A1(n7538), .A2(n6017), .ZN(n6018) );
  NAND2_X1 U7553 ( .A1(n6358), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6024) );
  NOR2_X1 U7554 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6019) );
  NOR2_X1 U7555 ( .A1(n6030), .A2(n6019), .ZN(n7555) );
  NAND2_X1 U7556 ( .A1(n6020), .A2(n7555), .ZN(n6022) );
  NAND2_X1 U7557 ( .A1(n6347), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7558 ( .A1(n6025), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7559 ( .A1(n6026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6027) );
  XNOR2_X1 U7560 ( .A(n6027), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U7561 ( .A1(n7110), .A2(n9718), .ZN(n6028) );
  INV_X1 U7562 ( .A(n7504), .ZN(n7558) );
  NAND2_X1 U7563 ( .A1(n9322), .A2(n7558), .ZN(n6423) );
  NAND2_X1 U7564 ( .A1(n6072), .A2(n6423), .ZN(n6044) );
  NAND2_X1 U7565 ( .A1(n6358), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7566 ( .A1(n6355), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U7567 ( .B1(n6030), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6045), .ZN(
        n6031) );
  INV_X1 U7568 ( .A(n6031), .ZN(n7525) );
  NAND2_X1 U7569 ( .A1(n6020), .A2(n7525), .ZN(n6033) );
  NAND2_X1 U7570 ( .A1(n6347), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6032) );
  NAND4_X1 U7571 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n9321)
         );
  NAND2_X1 U7572 ( .A1(n6344), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7573 ( .A1(n6037), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6039) );
  MUX2_X1 U7574 ( .A(n6039), .B(P1_IR_REG_31__SCAN_IN), .S(n6038), .Z(n6041)
         );
  NOR2_X1 U7575 ( .A1(n6037), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6065) );
  INV_X1 U7576 ( .A(n6065), .ZN(n6040) );
  NAND2_X1 U7577 ( .A1(n7110), .A2(n7177), .ZN(n6042) );
  OAI211_X1 U7578 ( .C1(n6844), .C2(n6054), .A(n6043), .B(n6042), .ZN(n7580)
         );
  INV_X1 U7579 ( .A(n7580), .ZN(n7521) );
  OR2_X1 U7580 ( .A1(n9321), .A2(n7521), .ZN(n6419) );
  OR2_X1 U7581 ( .A1(n9322), .A2(n7558), .ZN(n6397) );
  NAND2_X1 U7582 ( .A1(n6358), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7583 ( .A1(n6355), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6049) );
  AND2_X1 U7584 ( .A1(n6045), .A2(n7532), .ZN(n6046) );
  NOR2_X1 U7585 ( .A1(n6056), .A2(n6046), .ZN(n7576) );
  NAND2_X1 U7586 ( .A1(n6020), .A2(n7576), .ZN(n6048) );
  NAND2_X1 U7587 ( .A1(n6347), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7588 ( .A1(n6344), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6053) );
  OR2_X1 U7589 ( .A1(n6065), .A2(n6127), .ZN(n6051) );
  XNOR2_X1 U7590 ( .A(n6051), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U7591 ( .A1(n7110), .A2(n9752), .ZN(n6052) );
  OAI211_X1 U7592 ( .C1(n6850), .C2(n6054), .A(n6053), .B(n6052), .ZN(n7719)
         );
  OR2_X1 U7593 ( .A1(n9320), .A2(n9861), .ZN(n6418) );
  NAND2_X1 U7594 ( .A1(n9320), .A2(n9861), .ZN(n6415) );
  NAND2_X1 U7595 ( .A1(n6418), .A2(n6415), .ZN(n7584) );
  NAND2_X1 U7596 ( .A1(n9321), .A2(n7521), .ZN(n6422) );
  NAND3_X1 U7597 ( .A1(n6055), .A2(n7583), .A3(n6422), .ZN(n6070) );
  NAND2_X1 U7598 ( .A1(n6358), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7599 ( .A1(n6355), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6060) );
  OR2_X1 U7600 ( .A1(n6056), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6057) );
  AND2_X1 U7601 ( .A1(n6074), .A2(n6057), .ZN(n7726) );
  NAND2_X1 U7602 ( .A1(n6020), .A2(n7726), .ZN(n6059) );
  NAND2_X1 U7603 ( .A1(n6347), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6058) );
  NAND4_X1 U7604 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n9319)
         );
  NAND2_X1 U7605 ( .A1(n6855), .A2(n6342), .ZN(n6069) );
  INV_X1 U7606 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U7607 ( .A1(n6065), .A2(n6064), .ZN(n6080) );
  NAND2_X1 U7608 ( .A1(n6080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6066) );
  XNOR2_X1 U7609 ( .A(n6066), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9756) );
  INV_X1 U7610 ( .A(n9756), .ZN(n6856) );
  OAI22_X1 U7611 ( .A1(n6062), .A2(n6857), .B1(n7106), .B2(n6856), .ZN(n6067)
         );
  INV_X1 U7612 ( .A(n6067), .ZN(n6068) );
  NAND2_X1 U7613 ( .A1(n6069), .A2(n6068), .ZN(n7817) );
  NAND3_X1 U7614 ( .A1(n6070), .A2(n6418), .A3(n7867), .ZN(n6071) );
  NAND2_X1 U7615 ( .A1(n9319), .A2(n9867), .ZN(n6487) );
  NAND2_X1 U7616 ( .A1(n6071), .A2(n6487), .ZN(n6090) );
  INV_X1 U7617 ( .A(n6397), .ZN(n6420) );
  INV_X1 U7618 ( .A(n6422), .ZN(n7571) );
  OAI211_X1 U7619 ( .C1(n7711), .C2(n7571), .A(n7583), .B(n6419), .ZN(n6073)
         );
  AND2_X1 U7620 ( .A1(n6487), .A2(n6415), .ZN(n6424) );
  NAND2_X1 U7621 ( .A1(n6073), .A2(n6424), .ZN(n6088) );
  NAND2_X1 U7622 ( .A1(n6355), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7623 ( .A1(n6356), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7624 ( .A1(n6074), .A2(n10095), .ZN(n6075) );
  AND2_X1 U7625 ( .A1(n6101), .A2(n6075), .ZN(n7879) );
  NAND2_X1 U7626 ( .A1(n6020), .A2(n7879), .ZN(n6077) );
  NAND2_X1 U7627 ( .A1(n6358), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6076) );
  NAND4_X1 U7628 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n9318)
         );
  INV_X1 U7629 ( .A(n9318), .ZN(n7983) );
  NAND2_X1 U7630 ( .A1(n6863), .A2(n6342), .ZN(n6087) );
  NAND2_X1 U7631 ( .A1(n6083), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6082) );
  MUX2_X1 U7632 ( .A(n6082), .B(P1_IR_REG_31__SCAN_IN), .S(n6081), .Z(n6084)
         );
  INV_X1 U7633 ( .A(n9769), .ZN(n7171) );
  OAI22_X1 U7634 ( .A1(n6062), .A2(n6866), .B1(n7106), .B2(n7171), .ZN(n6085)
         );
  INV_X1 U7635 ( .A(n6085), .ZN(n6086) );
  NAND2_X1 U7636 ( .A1(n7983), .A2(n9871), .ZN(n6401) );
  AND2_X1 U7637 ( .A1(n6401), .A2(n7867), .ZN(n7820) );
  NAND2_X1 U7638 ( .A1(n6088), .A2(n7820), .ZN(n6089) );
  NAND2_X1 U7639 ( .A1(n6872), .A2(n6342), .ZN(n6099) );
  NAND2_X1 U7640 ( .A1(n6091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6092) );
  MUX2_X1 U7641 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6092), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6096) );
  INV_X1 U7642 ( .A(n6094), .ZN(n6095) );
  NAND2_X1 U7643 ( .A1(n6096), .A2(n6095), .ZN(n7179) );
  OAI22_X1 U7644 ( .A1(n6062), .A2(n6873), .B1(n7106), .B2(n7179), .ZN(n6097)
         );
  INV_X1 U7645 ( .A(n6097), .ZN(n6098) );
  NAND2_X1 U7646 ( .A1(n6099), .A2(n6098), .ZN(n7987) );
  AND2_X1 U7647 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  NOR2_X1 U7648 ( .A1(n6113), .A2(n6102), .ZN(n7980) );
  NAND2_X1 U7649 ( .A1(n6020), .A2(n7980), .ZN(n6106) );
  NAND2_X1 U7650 ( .A1(n6355), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7651 ( .A1(n6347), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7652 ( .A1(n6358), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6103) );
  NAND4_X1 U7653 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n7995)
         );
  INV_X1 U7654 ( .A(n7995), .ZN(n8070) );
  OR2_X1 U7655 ( .A1(n7987), .A2(n8070), .ZN(n6400) );
  OR2_X1 U7656 ( .A1(n7983), .A2(n9871), .ZN(n7821) );
  AND2_X1 U7657 ( .A1(n6400), .A2(n7821), .ZN(n7991) );
  NAND2_X1 U7658 ( .A1(n6875), .A2(n6342), .ZN(n6112) );
  NOR2_X1 U7659 ( .A1(n6094), .A2(n6127), .ZN(n6107) );
  MUX2_X1 U7660 ( .A(n6127), .B(n6107), .S(P1_IR_REG_10__SCAN_IN), .Z(n6109)
         );
  OR2_X1 U7661 ( .A1(n6109), .A2(n6108), .ZN(n7169) );
  OAI22_X1 U7662 ( .A1(n6062), .A2(n6879), .B1(n7106), .B2(n7169), .ZN(n6110)
         );
  INV_X1 U7663 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7664 ( .A1(n6112), .A2(n6111), .ZN(n8005) );
  NAND2_X1 U7665 ( .A1(n6355), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7666 ( .A1(n6358), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6117) );
  NOR2_X1 U7667 ( .A1(n6113), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7668 ( .A1(n6020), .A2(n4966), .ZN(n6116) );
  NAND2_X1 U7669 ( .A1(n6356), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6115) );
  NAND4_X1 U7670 ( .A1(n6118), .A2(n6117), .A3(n6116), .A4(n6115), .ZN(n8004)
         );
  OR2_X1 U7671 ( .A1(n8005), .A2(n8199), .ZN(n6434) );
  NAND3_X1 U7672 ( .A1(n6121), .A2(n7991), .A3(n6434), .ZN(n6119) );
  NAND2_X1 U7673 ( .A1(n8005), .A2(n8199), .ZN(n8011) );
  NAND2_X1 U7674 ( .A1(n7987), .A2(n8070), .ZN(n7993) );
  NAND2_X1 U7675 ( .A1(n8011), .A2(n7993), .ZN(n6435) );
  NAND2_X1 U7676 ( .A1(n6435), .A2(n6434), .ZN(n6427) );
  NAND2_X1 U7677 ( .A1(n6119), .A2(n6427), .ZN(n6125) );
  INV_X1 U7678 ( .A(n7821), .ZN(n6120) );
  AND2_X1 U7679 ( .A1(n6434), .A2(n6400), .ZN(n6122) );
  AOI21_X1 U7680 ( .B1(n6123), .B2(n6122), .A(n4742), .ZN(n6124) );
  NAND2_X1 U7681 ( .A1(n6880), .A2(n6342), .ZN(n6132) );
  NOR2_X1 U7682 ( .A1(n6108), .A2(n6127), .ZN(n6126) );
  MUX2_X1 U7683 ( .A(n6127), .B(n6126), .S(P1_IR_REG_11__SCAN_IN), .Z(n6129)
         );
  OR2_X1 U7684 ( .A1(n6129), .A2(n6128), .ZN(n7250) );
  OAI22_X1 U7685 ( .A1(n6062), .A2(n10244), .B1(n7106), .B2(n7250), .ZN(n6130)
         );
  INV_X1 U7686 ( .A(n6130), .ZN(n6131) );
  NAND2_X1 U7687 ( .A1(n6355), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7688 ( .A1(n6356), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7689 ( .A1(n6133), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6134) );
  AND2_X1 U7690 ( .A1(n6148), .A2(n6134), .ZN(n8196) );
  NAND2_X1 U7691 ( .A1(n6020), .A2(n8196), .ZN(n6136) );
  NAND2_X1 U7692 ( .A1(n6358), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6135) );
  NAND4_X1 U7693 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n9317)
         );
  XNOR2_X1 U7694 ( .A(n8207), .B(n9317), .ZN(n8013) );
  NAND2_X1 U7695 ( .A1(n6139), .A2(n8013), .ZN(n6180) );
  NAND2_X1 U7696 ( .A1(n6884), .A2(n6342), .ZN(n6147) );
  NAND2_X1 U7697 ( .A1(n6140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6141) );
  MUX2_X1 U7698 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6141), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6144) );
  AND2_X1 U7699 ( .A1(n6144), .A2(n6143), .ZN(n7399) );
  INV_X1 U7700 ( .A(n7399), .ZN(n6885) );
  OAI22_X1 U7701 ( .A1(n6062), .A2(n6886), .B1(n7106), .B2(n6885), .ZN(n6145)
         );
  INV_X1 U7702 ( .A(n6145), .ZN(n6146) );
  NAND2_X1 U7703 ( .A1(n6355), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7704 ( .A1(n6358), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7705 ( .A1(n6148), .A2(n10166), .ZN(n6149) );
  AND2_X1 U7706 ( .A1(n6170), .A2(n6149), .ZN(n8121) );
  NAND2_X1 U7707 ( .A1(n6020), .A2(n8121), .ZN(n6151) );
  NAND2_X1 U7708 ( .A1(n6347), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6150) );
  NAND4_X1 U7709 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n9316)
         );
  INV_X1 U7710 ( .A(n9316), .ZN(n8141) );
  OR2_X1 U7711 ( .A1(n8158), .A2(n8141), .ZN(n6403) );
  INV_X1 U7712 ( .A(n9317), .ZN(n8119) );
  OR2_X1 U7713 ( .A1(n8207), .A2(n8119), .ZN(n8054) );
  AND2_X1 U7714 ( .A1(n6403), .A2(n8054), .ZN(n8147) );
  NAND2_X1 U7715 ( .A1(n6180), .A2(n8147), .ZN(n6178) );
  NAND2_X1 U7716 ( .A1(n8158), .A2(n8141), .ZN(n8149) );
  NAND2_X1 U7717 ( .A1(n7004), .A2(n6342), .ZN(n6160) );
  OR2_X1 U7718 ( .A1(n6143), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7719 ( .A1(n6154), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6156) );
  INV_X1 U7720 ( .A(n6156), .ZN(n6155) );
  NAND2_X1 U7721 ( .A1(n6155), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6157) );
  INV_X1 U7722 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U7723 ( .A1(n6156), .A2(n10195), .ZN(n6186) );
  AND2_X1 U7724 ( .A1(n6157), .A2(n6186), .ZN(n9807) );
  INV_X1 U7725 ( .A(n9807), .ZN(n7921) );
  OAI22_X1 U7726 ( .A1(n6062), .A2(n10315), .B1(n7106), .B2(n7921), .ZN(n6158)
         );
  INV_X1 U7727 ( .A(n6158), .ZN(n6159) );
  NAND2_X2 U7728 ( .A1(n6160), .A2(n6159), .ZN(n9179) );
  NAND2_X1 U7729 ( .A1(n6358), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7730 ( .A1(n6355), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6164) );
  AND2_X1 U7731 ( .A1(n6172), .A2(n9173), .ZN(n6161) );
  NOR2_X1 U7732 ( .A1(n6192), .A2(n6161), .ZN(n9174) );
  NAND2_X1 U7733 ( .A1(n6020), .A2(n9174), .ZN(n6163) );
  NAND2_X1 U7734 ( .A1(n6347), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6162) );
  NAND4_X1 U7735 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n9314)
         );
  INV_X1 U7736 ( .A(n9314), .ZN(n8288) );
  OR2_X2 U7737 ( .A1(n9179), .A2(n8288), .ZN(n8283) );
  NAND2_X1 U7738 ( .A1(n6964), .A2(n6342), .ZN(n6168) );
  NAND2_X1 U7739 ( .A1(n6143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  XNOR2_X1 U7740 ( .A(n6166), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7923) );
  AOI22_X1 U7741 ( .A1(n6344), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7110), .B2(
        n7923), .ZN(n6167) );
  NAND2_X1 U7742 ( .A1(n6358), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7743 ( .A1(n6355), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7744 ( .A1(n6170), .A2(n6169), .ZN(n6171) );
  AND2_X1 U7745 ( .A1(n6172), .A2(n6171), .ZN(n8182) );
  NAND2_X1 U7746 ( .A1(n6020), .A2(n8182), .ZN(n6174) );
  NAND2_X1 U7747 ( .A1(n6356), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6173) );
  NAND4_X1 U7748 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n9315)
         );
  INV_X1 U7749 ( .A(n9315), .ZN(n9177) );
  OR2_X1 U7750 ( .A1(n8183), .A2(n9177), .ZN(n6395) );
  AND2_X1 U7751 ( .A1(n8283), .A2(n6395), .ZN(n6439) );
  INV_X1 U7752 ( .A(n6439), .ZN(n6177) );
  AOI21_X1 U7753 ( .B1(n6178), .B2(n8149), .A(n6177), .ZN(n6185) );
  AND2_X1 U7754 ( .A1(n8207), .A2(n8119), .ZN(n8053) );
  INV_X1 U7755 ( .A(n8053), .ZN(n6179) );
  AND2_X1 U7756 ( .A1(n8149), .A2(n6179), .ZN(n6437) );
  NAND2_X1 U7757 ( .A1(n6180), .A2(n6437), .ZN(n6181) );
  NAND2_X1 U7758 ( .A1(n6181), .A2(n6403), .ZN(n6182) );
  NAND2_X1 U7759 ( .A1(n6182), .A2(n8151), .ZN(n6183) );
  NAND2_X1 U7760 ( .A1(n9179), .A2(n8288), .ZN(n6433) );
  INV_X1 U7761 ( .A(n6433), .ZN(n6429) );
  AOI21_X1 U7762 ( .B1(n6183), .B2(n6439), .A(n6429), .ZN(n6184) );
  NAND2_X1 U7763 ( .A1(n7186), .A2(n6342), .ZN(n6191) );
  NAND2_X1 U7764 ( .A1(n6186), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6188) );
  XNOR2_X1 U7765 ( .A(n6188), .B(n6187), .ZN(n8099) );
  OAI22_X1 U7766 ( .A1(n6062), .A2(n7189), .B1(n7106), .B2(n8099), .ZN(n6189)
         );
  INV_X1 U7767 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7768 ( .A1(n6358), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7769 ( .A1(n6355), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6196) );
  OR2_X1 U7770 ( .A1(n6192), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6193) );
  AND2_X1 U7771 ( .A1(n6193), .A2(n6207), .ZN(n9307) );
  NAND2_X1 U7772 ( .A1(n6020), .A2(n9307), .ZN(n6195) );
  NAND2_X1 U7773 ( .A1(n6356), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6194) );
  NAND4_X1 U7774 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n9313)
         );
  XNOR2_X1 U7775 ( .A(n8303), .B(n9313), .ZN(n8285) );
  NAND2_X1 U7776 ( .A1(n6433), .A2(n8151), .ZN(n6198) );
  NAND3_X1 U7777 ( .A1(n6198), .A2(n7007), .A3(n8283), .ZN(n6199) );
  NAND2_X1 U7778 ( .A1(n8285), .A2(n6199), .ZN(n6216) );
  NAND2_X1 U7779 ( .A1(n7271), .A2(n6342), .ZN(n6205) );
  INV_X1 U7780 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7781 ( .A1(n6201), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6202) );
  XNOR2_X1 U7782 ( .A(n6202), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8352) );
  INV_X1 U7783 ( .A(n8352), .ZN(n8106) );
  OAI22_X1 U7784 ( .A1(n6062), .A2(n7285), .B1(n7106), .B2(n8106), .ZN(n6203)
         );
  INV_X1 U7785 ( .A(n6203), .ZN(n6204) );
  NAND2_X2 U7786 ( .A1(n6205), .A2(n6204), .ZN(n9617) );
  NAND2_X1 U7787 ( .A1(n6358), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7788 ( .A1(n6355), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7789 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  AND2_X1 U7790 ( .A1(n6226), .A2(n6208), .ZN(n9213) );
  NAND2_X1 U7791 ( .A1(n6020), .A2(n9213), .ZN(n6210) );
  NAND2_X1 U7792 ( .A1(n6356), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6209) );
  NAND4_X1 U7793 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(n9538)
         );
  INV_X1 U7794 ( .A(n9538), .ZN(n9302) );
  NAND2_X1 U7795 ( .A1(n9617), .A2(n9302), .ZN(n8503) );
  NAND2_X2 U7796 ( .A1(n6445), .A2(n8503), .ZN(n8500) );
  INV_X1 U7797 ( .A(n9313), .ZN(n8309) );
  NOR2_X1 U7798 ( .A1(n8303), .A2(n8309), .ZN(n8306) );
  NAND2_X1 U7799 ( .A1(n8303), .A2(n8309), .ZN(n8305) );
  INV_X1 U7800 ( .A(n8305), .ZN(n6213) );
  MUX2_X1 U7801 ( .A(n8306), .B(n6213), .S(n6371), .Z(n6214) );
  NOR2_X1 U7802 ( .A1(n8500), .A2(n6214), .ZN(n6215) );
  NAND2_X1 U7803 ( .A1(n7309), .A2(n6342), .ZN(n6224) );
  NAND2_X1 U7804 ( .A1(n6218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7805 ( .A1(n6220), .A2(n6219), .ZN(n6234) );
  OR2_X1 U7806 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  NAND2_X1 U7807 ( .A1(n6234), .A2(n6221), .ZN(n9338) );
  OAI22_X1 U7808 ( .A1(n6062), .A2(n7343), .B1(n7106), .B2(n9338), .ZN(n6222)
         );
  INV_X1 U7809 ( .A(n6222), .ZN(n6223) );
  AND2_X1 U7810 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  NOR2_X1 U7811 ( .A1(n6240), .A2(n6227), .ZN(n9531) );
  NAND2_X1 U7812 ( .A1(n9531), .A2(n6020), .ZN(n6231) );
  NAND2_X1 U7813 ( .A1(n6355), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7814 ( .A1(n6358), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7815 ( .A1(n6356), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6228) );
  NAND4_X1 U7816 ( .A1(n6231), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(n9522)
         );
  INV_X1 U7817 ( .A(n9522), .ZN(n9216) );
  OR2_X1 U7818 ( .A1(n9610), .A2(n9216), .ZN(n9517) );
  NAND2_X1 U7819 ( .A1(n9610), .A2(n9216), .ZN(n6246) );
  MUX2_X1 U7820 ( .A(n6445), .B(n8503), .S(n7007), .Z(n6232) );
  NAND3_X1 U7821 ( .A1(n6233), .A2(n9535), .A3(n6232), .ZN(n6249) );
  NAND2_X1 U7822 ( .A1(n7473), .A2(n6342), .ZN(n6239) );
  INV_X1 U7823 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U7824 ( .A1(n6234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6236) );
  XNOR2_X1 U7825 ( .A(n6236), .B(n6235), .ZN(n9829) );
  OAI22_X1 U7826 ( .A1(n6062), .A2(n7475), .B1(n7106), .B2(n9829), .ZN(n6237)
         );
  INV_X1 U7827 ( .A(n6237), .ZN(n6238) );
  NAND2_X2 U7828 ( .A1(n6239), .A2(n6238), .ZN(n9605) );
  NOR2_X1 U7829 ( .A1(n6240), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6241) );
  OR2_X1 U7830 ( .A1(n6253), .A2(n6241), .ZN(n9513) );
  INV_X1 U7831 ( .A(n6020), .ZN(n6301) );
  NAND2_X1 U7832 ( .A1(n6355), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7833 ( .A1(n6356), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6242) );
  AND2_X1 U7834 ( .A1(n6243), .A2(n6242), .ZN(n6245) );
  NAND2_X1 U7835 ( .A1(n6358), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6244) );
  OAI211_X1 U7836 ( .C1(n9513), .C2(n6301), .A(n6245), .B(n6244), .ZN(n9540)
         );
  INV_X1 U7837 ( .A(n9540), .ZN(n9224) );
  NAND2_X1 U7838 ( .A1(n9605), .A2(n9224), .ZN(n6449) );
  NAND2_X1 U7839 ( .A1(n6449), .A2(n6246), .ZN(n8505) );
  OR2_X1 U7840 ( .A1(n9605), .A2(n9224), .ZN(n6394) );
  NAND2_X1 U7841 ( .A1(n6394), .A2(n9517), .ZN(n6450) );
  MUX2_X1 U7842 ( .A(n8505), .B(n6450), .S(n7007), .Z(n6247) );
  INV_X1 U7843 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U7844 ( .A1(n7588), .A2(n6342), .ZN(n6252) );
  OAI22_X1 U7845 ( .A1(n6062), .A2(n7589), .B1(n6482), .B2(n7106), .ZN(n6250)
         );
  INV_X1 U7846 ( .A(n6250), .ZN(n6251) );
  NOR2_X1 U7847 ( .A1(n6253), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6254) );
  OR2_X1 U7848 ( .A1(n6259), .A2(n6254), .ZN(n9497) );
  AOI22_X1 U7849 ( .A1(n6355), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n6347), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7850 ( .A1(n6358), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6255) );
  OAI211_X1 U7851 ( .C1(n9497), .C2(n6301), .A(n6256), .B(n6255), .ZN(n9521)
         );
  INV_X1 U7852 ( .A(n9521), .ZN(n9278) );
  OR2_X1 U7853 ( .A1(n9600), .A2(n9278), .ZN(n6393) );
  NAND2_X1 U7854 ( .A1(n7732), .A2(n6342), .ZN(n6258) );
  NAND2_X1 U7855 ( .A1(n6344), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6257) );
  NOR2_X1 U7856 ( .A1(n6259), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6260) );
  OR2_X1 U7857 ( .A1(n6269), .A2(n6260), .ZN(n9490) );
  AOI22_X1 U7858 ( .A1(n6355), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n6347), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7859 ( .A1(n6358), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6261) );
  OAI211_X1 U7860 ( .C1(n9490), .C2(n6301), .A(n6262), .B(n6261), .ZN(n9504)
         );
  INV_X1 U7861 ( .A(n9504), .ZN(n9194) );
  NAND2_X1 U7862 ( .A1(n9595), .A2(n9194), .ZN(n6392) );
  OR2_X1 U7863 ( .A1(n9595), .A2(n9194), .ZN(n8511) );
  AND2_X1 U7864 ( .A1(n8511), .A2(n6393), .ZN(n6451) );
  NAND2_X1 U7865 ( .A1(n7802), .A2(n6342), .ZN(n6268) );
  NAND2_X1 U7866 ( .A1(n6344), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6267) );
  OR2_X1 U7867 ( .A1(n6269), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6270) );
  AND2_X1 U7868 ( .A1(n6270), .A2(n6280), .ZN(n9468) );
  NAND2_X1 U7869 ( .A1(n9468), .A2(n6020), .ZN(n6276) );
  INV_X1 U7870 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U7871 ( .A1(n6355), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7872 ( .A1(n6356), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6271) );
  OAI211_X1 U7873 ( .C1(n6273), .C2(n10258), .A(n6272), .B(n6271), .ZN(n6274)
         );
  INV_X1 U7874 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U7875 ( .A1(n6276), .A2(n6275), .ZN(n9488) );
  INV_X1 U7876 ( .A(n9488), .ZN(n6286) );
  NAND2_X1 U7877 ( .A1(n9592), .A2(n6286), .ZN(n6391) );
  INV_X1 U7878 ( .A(n6391), .ZN(n6277) );
  AOI21_X1 U7879 ( .B1(n6309), .B2(n8511), .A(n6277), .ZN(n6288) );
  NAND2_X1 U7880 ( .A1(n8342), .A2(n6342), .ZN(n6279) );
  NAND2_X1 U7881 ( .A1(n6344), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7882 ( .A1(n6358), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7883 ( .A1(n6355), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6284) );
  INV_X1 U7884 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6281) );
  AOI21_X1 U7885 ( .B1(n6281), .B2(n6280), .A(n6300), .ZN(n9446) );
  NAND2_X1 U7886 ( .A1(n6020), .A2(n9446), .ZN(n6283) );
  NAND2_X1 U7887 ( .A1(n6356), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6282) );
  NAND4_X1 U7888 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n9462)
         );
  INV_X1 U7889 ( .A(n9462), .ZN(n9432) );
  OR2_X1 U7890 ( .A1(n9586), .A2(n9432), .ZN(n6455) );
  NAND2_X1 U7891 ( .A1(n6455), .A2(n8512), .ZN(n6287) );
  NAND2_X1 U7892 ( .A1(n9586), .A2(n9432), .ZN(n8513) );
  OAI21_X1 U7893 ( .B1(n6288), .B2(n6287), .A(n8513), .ZN(n6307) );
  NAND2_X1 U7894 ( .A1(n8001), .A2(n6342), .ZN(n6290) );
  NAND2_X1 U7895 ( .A1(n6344), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7896 ( .A1(n6358), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7897 ( .A1(n6355), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6295) );
  INV_X1 U7898 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U7899 ( .A1(n6299), .A2(n9232), .ZN(n6291) );
  AND2_X1 U7900 ( .A1(n6292), .A2(n6291), .ZN(n9418) );
  NAND2_X1 U7901 ( .A1(n6020), .A2(n9418), .ZN(n6294) );
  NAND2_X1 U7902 ( .A1(n6356), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6293) );
  NAND4_X1 U7903 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n9439)
         );
  OR2_X1 U7904 ( .A1(n9406), .A2(n8490), .ZN(n6316) );
  NAND2_X1 U7905 ( .A1(n7929), .A2(n6342), .ZN(n6298) );
  NAND2_X1 U7906 ( .A1(n6344), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6297) );
  OAI21_X1 U7907 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6300), .A(n6299), .ZN(
        n9427) );
  OR2_X1 U7908 ( .A1(n6301), .A2(n9427), .ZN(n6305) );
  NAND2_X1 U7909 ( .A1(n6355), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7910 ( .A1(n6356), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7911 ( .A1(n6358), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6302) );
  NAND4_X1 U7912 ( .A1(n6305), .A2(n6304), .A3(n6303), .A4(n6302), .ZN(n9452)
         );
  INV_X1 U7913 ( .A(n6316), .ZN(n6306) );
  NAND2_X1 U7914 ( .A1(n9581), .A2(n9256), .ZN(n6461) );
  NOR2_X1 U7915 ( .A1(n6306), .A2(n6461), .ZN(n6484) );
  NAND2_X1 U7916 ( .A1(n8517), .A2(n4746), .ZN(n6462) );
  INV_X1 U7917 ( .A(n8512), .ZN(n6308) );
  INV_X1 U7918 ( .A(n6392), .ZN(n6310) );
  NAND2_X1 U7919 ( .A1(n8512), .A2(n6310), .ZN(n6311) );
  AND2_X1 U7920 ( .A1(n6311), .A2(n6391), .ZN(n6312) );
  NAND2_X1 U7921 ( .A1(n8513), .A2(n6312), .ZN(n6448) );
  OAI21_X1 U7922 ( .B1(n6313), .B2(n6448), .A(n6455), .ZN(n6315) );
  INV_X1 U7923 ( .A(n9410), .ZN(n6314) );
  AOI21_X1 U7924 ( .B1(n6321), .B2(n6320), .A(n6319), .ZN(n6322) );
  NAND2_X1 U7925 ( .A1(n8330), .A2(n6342), .ZN(n6325) );
  NAND2_X1 U7926 ( .A1(n6344), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7927 ( .A1(n6355), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7928 ( .A1(n6358), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6334) );
  INV_X1 U7929 ( .A(n6330), .ZN(n6327) );
  AND2_X1 U7930 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6326) );
  NAND2_X1 U7931 ( .A1(n6327), .A2(n6326), .ZN(n6357) );
  INV_X1 U7932 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6329) );
  INV_X1 U7933 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6328) );
  OAI21_X1 U7934 ( .B1(n6330), .B2(n6329), .A(n6328), .ZN(n6331) );
  NAND2_X1 U7935 ( .A1(n6020), .A2(n9348), .ZN(n6333) );
  NAND2_X1 U7936 ( .A1(n6356), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6332) );
  MUX2_X1 U7937 ( .A(n8521), .B(n6464), .S(n7007), .Z(n6336) );
  NAND2_X1 U7938 ( .A1(n9352), .A2(n6336), .ZN(n6353) );
  NAND2_X1 U7939 ( .A1(n9160), .A2(n6342), .ZN(n6338) );
  NAND2_X1 U7940 ( .A1(n6344), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7941 ( .A1(n6356), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U7942 ( .A1(n6355), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7943 ( .A1(n6358), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6339) );
  NAND3_X1 U7944 ( .A1(n6341), .A2(n6340), .A3(n6339), .ZN(n9312) );
  NAND2_X1 U7945 ( .A1(n6343), .A2(n6342), .ZN(n6346) );
  NAND2_X1 U7946 ( .A1(n6344), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U7947 ( .A1(n6358), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7948 ( .A1(n6355), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7949 ( .A1(n6356), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6348) );
  NAND3_X1 U7950 ( .A1(n6350), .A2(n6349), .A3(n6348), .ZN(n9311) );
  INV_X1 U7951 ( .A(n9311), .ZN(n6384) );
  NAND2_X1 U7952 ( .A1(n9339), .A2(n6384), .ZN(n6471) );
  INV_X1 U7953 ( .A(n9312), .ZN(n6351) );
  NAND2_X1 U7954 ( .A1(n9339), .A2(n6351), .ZN(n6390) );
  NAND2_X1 U7955 ( .A1(n6471), .A2(n6390), .ZN(n6372) );
  MUX2_X1 U7956 ( .A(n8522), .B(n6469), .S(n7007), .Z(n6352) );
  NAND2_X1 U7957 ( .A1(n6355), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U7958 ( .A1(n6356), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6361) );
  INV_X1 U7959 ( .A(n6357), .ZN(n8497) );
  NAND2_X1 U7960 ( .A1(n6020), .A2(n8497), .ZN(n6360) );
  NAND2_X1 U7961 ( .A1(n6358), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6359) );
  INV_X1 U7962 ( .A(n6825), .ZN(n9354) );
  OAI21_X1 U7963 ( .B1(n9354), .B2(n9551), .A(n6363), .ZN(n6364) );
  NAND2_X1 U7964 ( .A1(n6367), .A2(n6364), .ZN(n6369) );
  OAI21_X1 U7965 ( .B1(n6367), .B2(n6825), .A(n4818), .ZN(n6365) );
  AOI21_X1 U7966 ( .B1(n8499), .B2(n6369), .A(n6365), .ZN(n6366) );
  NAND2_X1 U7967 ( .A1(n6366), .A2(n6371), .ZN(n6378) );
  INV_X1 U7968 ( .A(n6367), .ZN(n6368) );
  NAND2_X1 U7969 ( .A1(n6369), .A2(n6825), .ZN(n6375) );
  INV_X1 U7970 ( .A(n6370), .ZN(n6373) );
  NAND3_X1 U7971 ( .A1(n6376), .A2(n6375), .A3(n6374), .ZN(n6377) );
  NAND2_X1 U7972 ( .A1(n6378), .A2(n6377), .ZN(n6388) );
  NAND2_X1 U7973 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  NAND2_X1 U7974 ( .A1(n6382), .A2(n6381), .ZN(n6540) );
  NOR2_X1 U7975 ( .A1(n6544), .A2(n6383), .ZN(n6387) );
  OAI21_X1 U7976 ( .B1(n6482), .B2(n7296), .A(n6388), .ZN(n6386) );
  INV_X1 U7977 ( .A(n9550), .ZN(n6385) );
  NAND2_X1 U7978 ( .A1(n9551), .A2(n6825), .ZN(n8494) );
  NAND2_X1 U7979 ( .A1(n6390), .A2(n8494), .ZN(n6470) );
  INV_X1 U7980 ( .A(n9363), .ZN(n6412) );
  NAND2_X1 U7981 ( .A1(n9565), .A2(n9361), .ZN(n6463) );
  XNOR2_X1 U7982 ( .A(n9406), .B(n8490), .ZN(n9411) );
  NAND2_X1 U7983 ( .A1(n9410), .A2(n6461), .ZN(n9436) );
  INV_X1 U7984 ( .A(n9436), .ZN(n9425) );
  NAND2_X1 U7985 ( .A1(n8512), .A2(n6391), .ZN(n9457) );
  INV_X1 U7986 ( .A(n9457), .ZN(n9460) );
  NAND2_X1 U7987 ( .A1(n8511), .A2(n6392), .ZN(n9485) );
  INV_X1 U7988 ( .A(n9503), .ZN(n6408) );
  INV_X1 U7989 ( .A(n8172), .ZN(n8174) );
  NAND2_X1 U7990 ( .A1(n6396), .A2(n6490), .ZN(n7286) );
  NAND2_X1 U7991 ( .A1(n9325), .A2(n7022), .ZN(n6489) );
  NOR4_X1 U7992 ( .A1(n7543), .A2(n7292), .A3(n7286), .A4(n7018), .ZN(n6399)
         );
  NAND2_X1 U7993 ( .A1(n6419), .A2(n6422), .ZN(n7502) );
  NAND2_X1 U7994 ( .A1(n6397), .A2(n6423), .ZN(n7424) );
  INV_X1 U7995 ( .A(n7424), .ZN(n6398) );
  NAND4_X1 U7996 ( .A1(n6399), .A2(n7583), .A3(n7572), .A4(n6398), .ZN(n6402)
         );
  NAND2_X1 U7997 ( .A1(n6400), .A2(n7993), .ZN(n7822) );
  NAND2_X1 U7998 ( .A1(n7867), .A2(n6487), .ZN(n7722) );
  NOR4_X1 U7999 ( .A1(n6402), .A2(n7822), .A3(n7869), .A4(n7722), .ZN(n6404)
         );
  NAND2_X1 U8000 ( .A1(n6403), .A2(n8149), .ZN(n8168) );
  INV_X1 U8001 ( .A(n8168), .ZN(n8055) );
  NAND2_X1 U8002 ( .A1(n6434), .A2(n8011), .ZN(n8007) );
  INV_X1 U8003 ( .A(n8007), .ZN(n8009) );
  NAND4_X1 U8004 ( .A1(n6404), .A2(n8055), .A3(n8009), .A4(n8013), .ZN(n6405)
         );
  NOR4_X1 U8005 ( .A1(n8500), .A2(n8280), .A3(n8174), .A4(n6405), .ZN(n6406)
         );
  NAND3_X1 U8006 ( .A1(n6406), .A2(n9535), .A3(n8285), .ZN(n6407) );
  NOR4_X1 U8007 ( .A1(n9485), .A2(n6408), .A3(n9519), .A4(n6407), .ZN(n6409)
         );
  NAND4_X1 U8008 ( .A1(n9425), .A2(n9451), .A3(n9460), .A4(n6409), .ZN(n6410)
         );
  NOR4_X1 U8009 ( .A1(n9384), .A2(n9411), .A3(n9397), .A4(n6410), .ZN(n6411)
         );
  NAND2_X1 U8010 ( .A1(n8499), .A2(n9354), .ZN(n8495) );
  NAND4_X1 U8011 ( .A1(n9352), .A2(n6412), .A3(n6411), .A4(n8495), .ZN(n6413)
         );
  NOR3_X1 U8012 ( .A1(n6516), .A2(n6470), .A3(n6413), .ZN(n6414) );
  AOI21_X1 U8013 ( .B1(n6518), .B2(n6414), .A(n7412), .ZN(n6475) );
  INV_X1 U8014 ( .A(n6475), .ZN(n6477) );
  NAND2_X1 U8015 ( .A1(n6422), .A2(n6415), .ZN(n6416) );
  NAND2_X1 U8016 ( .A1(n6416), .A2(n6418), .ZN(n7712) );
  AND4_X1 U8017 ( .A1(n7712), .A2(n6487), .A3(n6423), .A4(n6417), .ZN(n6485)
         );
  NAND2_X1 U8018 ( .A1(n6419), .A2(n6418), .ZN(n7709) );
  NOR2_X1 U8019 ( .A1(n7709), .A2(n6420), .ZN(n6486) );
  AND2_X1 U8020 ( .A1(n6486), .A2(n6421), .ZN(n6493) );
  AOI21_X1 U8021 ( .B1(n6423), .B2(n6422), .A(n7709), .ZN(n6426) );
  INV_X1 U8022 ( .A(n6424), .ZN(n6425) );
  NOR3_X1 U8023 ( .A1(n6493), .A2(n6426), .A3(n6425), .ZN(n6432) );
  INV_X1 U8024 ( .A(n8505), .ZN(n6431) );
  NAND4_X1 U8025 ( .A1(n8151), .A2(n7820), .A3(n6437), .A4(n6427), .ZN(n6428)
         );
  NOR2_X1 U8026 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  NAND4_X1 U8027 ( .A1(n6431), .A2(n6430), .A3(n8305), .A4(n8503), .ZN(n6502)
         );
  AOI211_X1 U8028 ( .C1(n6485), .C2(n7538), .A(n6432), .B(n6502), .ZN(n6447)
         );
  AND2_X1 U8029 ( .A1(n8305), .A2(n6433), .ZN(n6443) );
  INV_X1 U8030 ( .A(n8147), .ZN(n6438) );
  OAI21_X1 U8031 ( .B1(n6435), .B2(n7991), .A(n6434), .ZN(n6436) );
  AOI22_X1 U8032 ( .A1(n6438), .A2(n8149), .B1(n6437), .B2(n6436), .ZN(n6441)
         );
  INV_X1 U8033 ( .A(n8151), .ZN(n6440) );
  OAI21_X1 U8034 ( .B1(n6441), .B2(n6440), .A(n6439), .ZN(n6442) );
  AOI21_X1 U8035 ( .B1(n6443), .B2(n6442), .A(n8306), .ZN(n6446) );
  INV_X1 U8036 ( .A(n8503), .ZN(n6444) );
  AOI211_X1 U8037 ( .C1(n6446), .C2(n6445), .A(n6444), .B(n8505), .ZN(n6504)
         );
  NOR2_X1 U8038 ( .A1(n6447), .A2(n6504), .ZN(n6457) );
  INV_X1 U8039 ( .A(n6448), .ZN(n6454) );
  NAND2_X1 U8040 ( .A1(n6454), .A2(n8509), .ZN(n6506) );
  INV_X1 U8041 ( .A(n8509), .ZN(n6452) );
  NAND2_X1 U8042 ( .A1(n6450), .A2(n6449), .ZN(n8506) );
  OAI211_X1 U8043 ( .C1(n6452), .C2(n8506), .A(n8512), .B(n6451), .ZN(n6453)
         );
  NAND2_X1 U8044 ( .A1(n6454), .A2(n6453), .ZN(n6456) );
  AND2_X1 U8045 ( .A1(n6456), .A2(n6455), .ZN(n6505) );
  OAI21_X1 U8046 ( .B1(n6457), .B2(n6506), .A(n6505), .ZN(n6460) );
  INV_X1 U8047 ( .A(n8515), .ZN(n6459) );
  AND2_X1 U8048 ( .A1(n8519), .A2(n8516), .ZN(n6458) );
  NAND2_X1 U8049 ( .A1(n8521), .A2(n6458), .ZN(n6508) );
  AOI211_X1 U8050 ( .C1(n6461), .C2(n6460), .A(n6459), .B(n6508), .ZN(n6468)
         );
  INV_X1 U8051 ( .A(n6462), .ZN(n6467) );
  NAND2_X1 U8052 ( .A1(n6464), .A2(n6463), .ZN(n6465) );
  NAND2_X1 U8053 ( .A1(n6465), .A2(n8521), .ZN(n6466) );
  OAI211_X1 U8054 ( .C1(n6508), .C2(n6467), .A(n8522), .B(n6466), .ZN(n6512)
         );
  NOR2_X1 U8055 ( .A1(n6468), .A2(n6512), .ZN(n6472) );
  NAND2_X1 U8056 ( .A1(n8495), .A2(n6469), .ZN(n6514) );
  INV_X1 U8057 ( .A(n6470), .ZN(n6513) );
  OAI211_X1 U8058 ( .C1(n6472), .C2(n6514), .A(n6513), .B(n6471), .ZN(n6473)
         );
  AOI211_X1 U8059 ( .C1(n4818), .C2(n6473), .A(n6383), .B(n6516), .ZN(n6474)
         );
  OR2_X1 U8060 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  MUX2_X1 U8061 ( .A(n6477), .B(n6476), .S(n6482), .Z(n6481) );
  NOR2_X1 U8062 ( .A1(n6483), .A2(n6482), .ZN(n6520) );
  INV_X1 U8063 ( .A(n6484), .ZN(n6510) );
  INV_X1 U8064 ( .A(n6485), .ZN(n6500) );
  INV_X1 U8065 ( .A(n6486), .ZN(n6488) );
  NAND3_X1 U8066 ( .A1(n6488), .A2(n6487), .A3(n7712), .ZN(n6499) );
  NAND3_X1 U8067 ( .A1(n6490), .A2(n6489), .A3(n7412), .ZN(n6491) );
  NAND2_X1 U8068 ( .A1(n7293), .A2(n6491), .ZN(n6496) );
  INV_X1 U8069 ( .A(n6492), .ZN(n6495) );
  INV_X1 U8070 ( .A(n6493), .ZN(n6494) );
  AOI211_X1 U8071 ( .C1(n6497), .C2(n6496), .A(n6495), .B(n6494), .ZN(n6498)
         );
  AOI21_X1 U8072 ( .B1(n6500), .B2(n6499), .A(n6498), .ZN(n6501) );
  NOR2_X1 U8073 ( .A1(n6502), .A2(n6501), .ZN(n6503) );
  NOR2_X1 U8074 ( .A1(n6504), .A2(n6503), .ZN(n6507) );
  OAI211_X1 U8075 ( .C1(n6507), .C2(n6506), .A(n8515), .B(n6505), .ZN(n6509)
         );
  AOI21_X1 U8076 ( .B1(n6510), .B2(n6509), .A(n6508), .ZN(n6511) );
  NOR2_X1 U8077 ( .A1(n6512), .A2(n6511), .ZN(n6515) );
  OAI21_X1 U8078 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(n6517) );
  AOI21_X1 U8079 ( .B1(n6518), .B2(n6517), .A(n6516), .ZN(n6519) );
  MUX2_X1 U8080 ( .A(n6552), .B(n6520), .S(n6519), .Z(n6524) );
  NAND2_X1 U8081 ( .A1(n6522), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6523) );
  XNOR2_X1 U8082 ( .A(n6523), .B(n4754), .ZN(n7114) );
  NOR2_X1 U8083 ( .A1(n7114), .A2(P1_U3084), .ZN(n7931) );
  INV_X1 U8084 ( .A(n6552), .ZN(n6525) );
  INV_X1 U8085 ( .A(n6526), .ZN(n9710) );
  INV_X1 U8086 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U8087 ( .A1(n6529), .A2(n6528), .ZN(n6531) );
  NAND2_X1 U8088 ( .A1(n6531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6527) );
  XNOR2_X1 U8089 ( .A(n6527), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6793) );
  OR2_X1 U8090 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  NAND2_X1 U8091 ( .A1(n6531), .A2(n6530), .ZN(n8190) );
  NAND2_X1 U8092 ( .A1(n4453), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6533) );
  XNOR2_X1 U8093 ( .A(n6533), .B(n6532), .ZN(n8003) );
  NOR2_X1 U8094 ( .A1(n8190), .A2(n8003), .ZN(n6534) );
  AND2_X1 U8095 ( .A1(n7114), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6862) );
  INV_X1 U8096 ( .A(n6860), .ZN(n7411) );
  NOR4_X1 U8097 ( .A1(n7509), .A2(n8348), .A3(n7411), .A4(n6535), .ZN(n6538)
         );
  INV_X1 U8098 ( .A(n7931), .ZN(n6536) );
  OAI21_X1 U8099 ( .B1(n6544), .B2(n6536), .A(P1_B_REG_SCAN_IN), .ZN(n6537) );
  OR2_X1 U8100 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  INV_X1 U8101 ( .A(n6540), .ZN(n6541) );
  NAND2_X2 U8102 ( .A1(n6541), .A2(n4794), .ZN(n6545) );
  CLKBUF_X3 U8103 ( .A(n6554), .Z(n6761) );
  NAND2_X1 U8104 ( .A1(n8303), .A2(n6784), .ZN(n6543) );
  NOR2_X2 U8105 ( .A1(n6545), .A2(n6548), .ZN(n6572) );
  NAND2_X1 U8106 ( .A1(n9313), .A2(n6693), .ZN(n6542) );
  NAND2_X1 U8107 ( .A1(n6543), .A2(n6542), .ZN(n6547) );
  NAND2_X1 U8108 ( .A1(n6544), .A2(n6482), .ZN(n6546) );
  XNOR2_X1 U8109 ( .A(n6547), .B(n7510), .ZN(n6690) );
  NAND2_X1 U8110 ( .A1(n9325), .A2(n6572), .ZN(n6550) );
  AOI22_X1 U8111 ( .A1(n6554), .A2(n7457), .B1(n6548), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8112 ( .A1(n6550), .A2(n6549), .ZN(n7153) );
  INV_X1 U8113 ( .A(n7153), .ZN(n6551) );
  NAND2_X1 U8114 ( .A1(n6551), .A2(n6562), .ZN(n6559) );
  NOR2_X1 U8115 ( .A1(n7116), .A2(n5986), .ZN(n6555) );
  AOI21_X1 U8116 ( .B1(n6572), .B2(n7457), .A(n6555), .ZN(n6556) );
  INV_X1 U8117 ( .A(n6556), .ZN(n6557) );
  NAND2_X1 U8118 ( .A1(n6564), .A2(n6572), .ZN(n6561) );
  NAND2_X1 U8119 ( .A1(n6761), .A2(n7456), .ZN(n6560) );
  NAND2_X1 U8120 ( .A1(n6561), .A2(n6560), .ZN(n6563) );
  XNOR2_X1 U8121 ( .A(n6563), .B(n6562), .ZN(n6568) );
  NAND2_X1 U8122 ( .A1(n4423), .A2(n6564), .ZN(n6566) );
  INV_X1 U8123 ( .A(n6786), .ZN(n6585) );
  NAND2_X1 U8124 ( .A1(n6585), .A2(n7456), .ZN(n6565) );
  AND2_X1 U8125 ( .A1(n6566), .A2(n6565), .ZN(n7264) );
  NAND2_X1 U8126 ( .A1(n7262), .A2(n7264), .ZN(n6571) );
  INV_X1 U8127 ( .A(n6567), .ZN(n6570) );
  INV_X1 U8128 ( .A(n6568), .ZN(n6569) );
  NAND2_X1 U8129 ( .A1(n6570), .A2(n6569), .ZN(n7263) );
  NAND2_X1 U8130 ( .A1(n6571), .A2(n7263), .ZN(n9260) );
  NAND2_X1 U8131 ( .A1(n6761), .A2(n4530), .ZN(n6575) );
  NAND2_X1 U8132 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  NAND2_X1 U8133 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  NAND2_X1 U8134 ( .A1(n4424), .A2(n6573), .ZN(n6578) );
  NAND2_X1 U8135 ( .A1(n6572), .A2(n4530), .ZN(n6577) );
  AND2_X1 U8136 ( .A1(n6578), .A2(n6577), .ZN(n6580) );
  NAND2_X1 U8137 ( .A1(n6579), .A2(n6580), .ZN(n6584) );
  NAND2_X1 U8138 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  NAND2_X1 U8139 ( .A1(n9261), .A2(n6584), .ZN(n7218) );
  NAND2_X1 U8140 ( .A1(n9323), .A2(n6585), .ZN(n6587) );
  NAND2_X1 U8141 ( .A1(n6761), .A2(n4422), .ZN(n6586) );
  NAND2_X1 U8142 ( .A1(n6587), .A2(n6586), .ZN(n6589) );
  XNOR2_X1 U8143 ( .A(n6589), .B(n6782), .ZN(n6597) );
  NAND2_X1 U8144 ( .A1(n4423), .A2(n9323), .ZN(n6591) );
  NAND2_X1 U8145 ( .A1(n6693), .A2(n4422), .ZN(n6590) );
  NAND2_X1 U8146 ( .A1(n6591), .A2(n6590), .ZN(n6595) );
  XNOR2_X1 U8147 ( .A(n6597), .B(n6595), .ZN(n7219) );
  NAND2_X1 U8148 ( .A1(n6761), .A2(n7504), .ZN(n6592) );
  NAND2_X1 U8149 ( .A1(n4424), .A2(n9322), .ZN(n6594) );
  NAND2_X1 U8150 ( .A1(n6693), .A2(n7504), .ZN(n6593) );
  NAND2_X1 U8151 ( .A1(n6594), .A2(n6593), .ZN(n6600) );
  XNOR2_X1 U8152 ( .A(n6599), .B(n6600), .ZN(n7276) );
  INV_X1 U8153 ( .A(n6595), .ZN(n6596) );
  NAND2_X1 U8154 ( .A1(n6597), .A2(n6596), .ZN(n7273) );
  NAND2_X1 U8155 ( .A1(n7274), .A2(n6598), .ZN(n7275) );
  INV_X1 U8156 ( .A(n6599), .ZN(n6601) );
  NAND2_X1 U8157 ( .A1(n6601), .A2(n6600), .ZN(n6602) );
  NAND2_X1 U8158 ( .A1(n7275), .A2(n6602), .ZN(n6607) );
  NAND2_X1 U8159 ( .A1(n9321), .A2(n6693), .ZN(n6604) );
  NAND2_X1 U8160 ( .A1(n6784), .A2(n7580), .ZN(n6603) );
  NAND2_X1 U8161 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  XNOR2_X1 U8162 ( .A(n6605), .B(n7510), .ZN(n6606) );
  OR2_X1 U8163 ( .A1(n6607), .A2(n6606), .ZN(n6612) );
  NAND2_X1 U8164 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  NAND2_X1 U8165 ( .A1(n4423), .A2(n9321), .ZN(n6610) );
  NAND2_X1 U8166 ( .A1(n6693), .A2(n7580), .ZN(n6609) );
  NAND2_X1 U8167 ( .A1(n6610), .A2(n6609), .ZN(n7520) );
  INV_X1 U8168 ( .A(n7520), .ZN(n6611) );
  NAND2_X1 U8169 ( .A1(n9320), .A2(n6693), .ZN(n6614) );
  NAND2_X1 U8170 ( .A1(n6784), .A2(n7719), .ZN(n6613) );
  NAND2_X1 U8171 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  XNOR2_X1 U8172 ( .A(n6615), .B(n6782), .ZN(n7529) );
  NAND2_X1 U8173 ( .A1(n4423), .A2(n9320), .ZN(n6617) );
  NAND2_X1 U8174 ( .A1(n6693), .A2(n7719), .ZN(n6616) );
  AND2_X1 U8175 ( .A1(n7529), .A2(n7528), .ZN(n6619) );
  NAND2_X1 U8176 ( .A1(n9319), .A2(n6693), .ZN(n6621) );
  NAND2_X1 U8177 ( .A1(n7817), .A2(n6761), .ZN(n6620) );
  NAND2_X1 U8178 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  XNOR2_X1 U8179 ( .A(n6622), .B(n6782), .ZN(n6625) );
  NAND2_X1 U8180 ( .A1(n4423), .A2(n9319), .ZN(n6624) );
  NAND2_X1 U8181 ( .A1(n6693), .A2(n7817), .ZN(n6623) );
  NAND2_X1 U8182 ( .A1(n6624), .A2(n6623), .ZN(n6626) );
  XNOR2_X1 U8183 ( .A(n6625), .B(n6626), .ZN(n7702) );
  INV_X1 U8184 ( .A(n6625), .ZN(n6627) );
  NAND2_X1 U8185 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  NAND2_X1 U8186 ( .A1(n9871), .A2(n6784), .ZN(n6631) );
  NAND2_X1 U8187 ( .A1(n9318), .A2(n6693), .ZN(n6630) );
  NAND2_X1 U8188 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  XNOR2_X1 U8189 ( .A(n6632), .B(n7510), .ZN(n7793) );
  NAND2_X1 U8190 ( .A1(n9871), .A2(n6778), .ZN(n6634) );
  NAND2_X1 U8191 ( .A1(n4423), .A2(n9318), .ZN(n6633) );
  NAND2_X1 U8192 ( .A1(n6634), .A2(n6633), .ZN(n7794) );
  NAND2_X1 U8193 ( .A1(n7987), .A2(n6784), .ZN(n6636) );
  NAND2_X1 U8194 ( .A1(n7995), .A2(n6693), .ZN(n6635) );
  NAND2_X1 U8195 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  XNOR2_X1 U8196 ( .A(n6637), .B(n6782), .ZN(n6639) );
  AND2_X1 U8197 ( .A1(n4424), .A2(n7995), .ZN(n6638) );
  AOI21_X1 U8198 ( .B1(n4621), .B2(n6693), .A(n6638), .ZN(n6640) );
  NAND2_X1 U8199 ( .A1(n6639), .A2(n6640), .ZN(n6644) );
  INV_X1 U8200 ( .A(n6639), .ZN(n6642) );
  INV_X1 U8201 ( .A(n6640), .ZN(n6641) );
  NAND2_X1 U8202 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  NAND2_X1 U8203 ( .A1(n6644), .A2(n6643), .ZN(n7979) );
  NAND2_X1 U8204 ( .A1(n7977), .A2(n6644), .ZN(n8064) );
  NAND2_X1 U8205 ( .A1(n8005), .A2(n6784), .ZN(n6646) );
  NAND2_X1 U8206 ( .A1(n8004), .A2(n6693), .ZN(n6645) );
  NAND2_X1 U8207 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XNOR2_X1 U8208 ( .A(n6647), .B(n7510), .ZN(n6653) );
  AND2_X1 U8209 ( .A1(n4424), .A2(n8004), .ZN(n6648) );
  AOI21_X1 U8210 ( .B1(n8005), .B2(n6693), .A(n6648), .ZN(n6654) );
  XNOR2_X1 U8211 ( .A(n6653), .B(n6654), .ZN(n8065) );
  NAND2_X1 U8212 ( .A1(n8064), .A2(n8065), .ZN(n8063) );
  NAND2_X1 U8213 ( .A1(n8207), .A2(n6761), .ZN(n6650) );
  NAND2_X1 U8214 ( .A1(n9317), .A2(n6693), .ZN(n6649) );
  NAND2_X1 U8215 ( .A1(n6650), .A2(n6649), .ZN(n6651) );
  XNOR2_X1 U8216 ( .A(n6651), .B(n7510), .ZN(n6663) );
  AND2_X1 U8217 ( .A1(n4424), .A2(n9317), .ZN(n6652) );
  AOI21_X1 U8218 ( .B1(n8207), .B2(n6778), .A(n6652), .ZN(n6661) );
  XNOR2_X1 U8219 ( .A(n6663), .B(n6661), .ZN(n8201) );
  INV_X1 U8220 ( .A(n6653), .ZN(n6655) );
  NAND2_X1 U8221 ( .A1(n6655), .A2(n6654), .ZN(n8202) );
  AND2_X1 U8222 ( .A1(n8201), .A2(n8202), .ZN(n6656) );
  NAND2_X1 U8223 ( .A1(n8063), .A2(n6656), .ZN(n8111) );
  NAND2_X1 U8224 ( .A1(n8158), .A2(n6761), .ZN(n6658) );
  NAND2_X1 U8225 ( .A1(n9316), .A2(n6693), .ZN(n6657) );
  NAND2_X1 U8226 ( .A1(n6658), .A2(n6657), .ZN(n6659) );
  XNOR2_X1 U8227 ( .A(n6659), .B(n7510), .ZN(n6665) );
  AND2_X1 U8228 ( .A1(n4424), .A2(n9316), .ZN(n6660) );
  AOI21_X1 U8229 ( .B1(n8158), .B2(n6778), .A(n6660), .ZN(n6666) );
  XNOR2_X1 U8230 ( .A(n6665), .B(n6666), .ZN(n8112) );
  INV_X1 U8231 ( .A(n6661), .ZN(n6662) );
  NAND2_X1 U8232 ( .A1(n6663), .A2(n6662), .ZN(n8113) );
  AND2_X1 U8233 ( .A1(n8112), .A2(n8113), .ZN(n6664) );
  INV_X1 U8234 ( .A(n6665), .ZN(n6667) );
  NAND2_X1 U8235 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  NAND2_X1 U8236 ( .A1(n8183), .A2(n6784), .ZN(n6670) );
  NAND2_X1 U8237 ( .A1(n9315), .A2(n6693), .ZN(n6669) );
  NAND2_X1 U8238 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  XNOR2_X1 U8239 ( .A(n6671), .B(n6782), .ZN(n6673) );
  AND2_X1 U8240 ( .A1(n4424), .A2(n9315), .ZN(n6672) );
  AOI21_X1 U8241 ( .B1(n8183), .B2(n6778), .A(n6672), .ZN(n6674) );
  AND2_X1 U8242 ( .A1(n6673), .A2(n6674), .ZN(n8133) );
  INV_X1 U8243 ( .A(n6673), .ZN(n6676) );
  INV_X1 U8244 ( .A(n6674), .ZN(n6675) );
  NAND2_X1 U8245 ( .A1(n6676), .A2(n6675), .ZN(n8134) );
  NAND2_X1 U8246 ( .A1(n9179), .A2(n6761), .ZN(n6678) );
  NAND2_X1 U8247 ( .A1(n9314), .A2(n6693), .ZN(n6677) );
  NAND2_X1 U8248 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  XNOR2_X1 U8249 ( .A(n6679), .B(n7510), .ZN(n6681) );
  NAND2_X1 U8250 ( .A1(n6682), .A2(n6681), .ZN(n6688) );
  INV_X1 U8251 ( .A(n6688), .ZN(n6680) );
  NOR2_X1 U8252 ( .A1(n6690), .A2(n6680), .ZN(n6685) );
  NAND2_X1 U8253 ( .A1(n9179), .A2(n6778), .ZN(n6684) );
  NAND2_X1 U8254 ( .A1(n4423), .A2(n9314), .ZN(n6683) );
  NAND2_X1 U8255 ( .A1(n6684), .A2(n6683), .ZN(n9172) );
  NAND2_X1 U8256 ( .A1(n6685), .A2(n6689), .ZN(n9295) );
  NAND2_X1 U8257 ( .A1(n8303), .A2(n6778), .ZN(n6687) );
  NAND2_X1 U8258 ( .A1(n4423), .A2(n9313), .ZN(n6686) );
  NAND2_X1 U8259 ( .A1(n6687), .A2(n6686), .ZN(n9297) );
  NAND2_X1 U8260 ( .A1(n9295), .A2(n9297), .ZN(n6692) );
  NAND2_X1 U8261 ( .A1(n6689), .A2(n6688), .ZN(n6691) );
  NAND2_X1 U8262 ( .A1(n6691), .A2(n6690), .ZN(n9294) );
  NAND2_X1 U8263 ( .A1(n9617), .A2(n6784), .ZN(n6695) );
  NAND2_X1 U8264 ( .A1(n9538), .A2(n6693), .ZN(n6694) );
  NAND2_X1 U8265 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  XNOR2_X1 U8266 ( .A(n6696), .B(n7510), .ZN(n6699) );
  NAND2_X1 U8267 ( .A1(n9617), .A2(n6778), .ZN(n6698) );
  NAND2_X1 U8268 ( .A1(n4423), .A2(n9538), .ZN(n6697) );
  NAND2_X1 U8269 ( .A1(n6698), .A2(n6697), .ZN(n6700) );
  INV_X1 U8270 ( .A(n6699), .ZN(n6702) );
  INV_X1 U8271 ( .A(n6700), .ZN(n6701) );
  NAND2_X1 U8272 ( .A1(n6702), .A2(n6701), .ZN(n9209) );
  NAND2_X1 U8273 ( .A1(n9610), .A2(n6784), .ZN(n6704) );
  NAND2_X1 U8274 ( .A1(n9522), .A2(n6778), .ZN(n6703) );
  NAND2_X1 U8275 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  XNOR2_X1 U8276 ( .A(n6705), .B(n6782), .ZN(n6710) );
  INV_X1 U8277 ( .A(n6710), .ZN(n6708) );
  AND2_X1 U8278 ( .A1(n4424), .A2(n9522), .ZN(n6706) );
  AOI21_X1 U8279 ( .B1(n9610), .B2(n6778), .A(n6706), .ZN(n6709) );
  INV_X1 U8280 ( .A(n6709), .ZN(n6707) );
  NAND2_X1 U8281 ( .A1(n6708), .A2(n6707), .ZN(n9220) );
  NAND2_X1 U8282 ( .A1(n9605), .A2(n6784), .ZN(n6712) );
  NAND2_X1 U8283 ( .A1(n9540), .A2(n6778), .ZN(n6711) );
  NAND2_X1 U8284 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  AND2_X1 U8285 ( .A1(n9540), .A2(n4424), .ZN(n6714) );
  NAND2_X1 U8286 ( .A1(n9274), .A2(n9276), .ZN(n6715) );
  NAND2_X1 U8287 ( .A1(n9600), .A2(n6784), .ZN(n6717) );
  NAND2_X1 U8288 ( .A1(n9521), .A2(n6778), .ZN(n6716) );
  NAND2_X1 U8289 ( .A1(n6717), .A2(n6716), .ZN(n6718) );
  XNOR2_X1 U8290 ( .A(n6718), .B(n7510), .ZN(n6720) );
  AND2_X1 U8291 ( .A1(n9521), .A2(n4424), .ZN(n6719) );
  AOI21_X1 U8292 ( .B1(n9600), .B2(n6778), .A(n6719), .ZN(n6721) );
  XNOR2_X1 U8293 ( .A(n6720), .B(n6721), .ZN(n9192) );
  INV_X1 U8294 ( .A(n6720), .ZN(n6722) );
  NAND2_X1 U8295 ( .A1(n6722), .A2(n6721), .ZN(n6723) );
  NAND2_X1 U8296 ( .A1(n9595), .A2(n6784), .ZN(n6725) );
  NAND2_X1 U8297 ( .A1(n9504), .A2(n6778), .ZN(n6724) );
  NAND2_X1 U8298 ( .A1(n6725), .A2(n6724), .ZN(n6726) );
  XNOR2_X1 U8299 ( .A(n6726), .B(n6782), .ZN(n9243) );
  AND2_X1 U8300 ( .A1(n9504), .A2(n4424), .ZN(n6727) );
  AOI21_X1 U8301 ( .B1(n9595), .B2(n6778), .A(n6727), .ZN(n9242) );
  AND2_X1 U8302 ( .A1(n9243), .A2(n9242), .ZN(n6731) );
  INV_X1 U8303 ( .A(n9243), .ZN(n6729) );
  INV_X1 U8304 ( .A(n9242), .ZN(n6728) );
  NAND2_X1 U8305 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  NAND2_X1 U8306 ( .A1(n9592), .A2(n6784), .ZN(n6733) );
  NAND2_X1 U8307 ( .A1(n9488), .A2(n6778), .ZN(n6732) );
  NAND2_X1 U8308 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  XNOR2_X1 U8309 ( .A(n6734), .B(n7510), .ZN(n6737) );
  NAND2_X1 U8310 ( .A1(n9592), .A2(n6778), .ZN(n6736) );
  NAND2_X1 U8311 ( .A1(n9488), .A2(n4423), .ZN(n6735) );
  NAND2_X1 U8312 ( .A1(n6736), .A2(n6735), .ZN(n6738) );
  INV_X1 U8313 ( .A(n6737), .ZN(n6740) );
  INV_X1 U8314 ( .A(n6738), .ZN(n6739) );
  NAND2_X1 U8315 ( .A1(n6740), .A2(n6739), .ZN(n8475) );
  NAND2_X1 U8316 ( .A1(n6741), .A2(n8475), .ZN(n6746) );
  AND2_X1 U8317 ( .A1(n4424), .A2(n9462), .ZN(n6742) );
  AOI21_X1 U8318 ( .B1(n9586), .B2(n6778), .A(n6742), .ZN(n6747) );
  NAND2_X1 U8319 ( .A1(n6746), .A2(n6747), .ZN(n9250) );
  NAND2_X1 U8320 ( .A1(n9586), .A2(n6761), .ZN(n6744) );
  NAND2_X1 U8321 ( .A1(n9462), .A2(n6778), .ZN(n6743) );
  NAND2_X1 U8322 ( .A1(n6744), .A2(n6743), .ZN(n6745) );
  INV_X1 U8323 ( .A(n6746), .ZN(n6749) );
  INV_X1 U8324 ( .A(n6747), .ZN(n6748) );
  NAND2_X1 U8325 ( .A1(n9581), .A2(n6761), .ZN(n6752) );
  NAND2_X1 U8326 ( .A1(n9452), .A2(n6778), .ZN(n6751) );
  NAND2_X1 U8327 ( .A1(n6752), .A2(n6751), .ZN(n6753) );
  XNOR2_X1 U8328 ( .A(n6753), .B(n7510), .ZN(n6754) );
  AOI22_X1 U8329 ( .A1(n9581), .A2(n6778), .B1(n4423), .B2(n9452), .ZN(n9183)
         );
  AOI22_X1 U8330 ( .A1(n9406), .A2(n6778), .B1(n4424), .B2(n9439), .ZN(n6759)
         );
  NAND2_X1 U8331 ( .A1(n9406), .A2(n6761), .ZN(n6756) );
  NAND2_X1 U8332 ( .A1(n9439), .A2(n6778), .ZN(n6755) );
  NAND2_X1 U8333 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  XNOR2_X1 U8334 ( .A(n6757), .B(n7510), .ZN(n6758) );
  XOR2_X1 U8335 ( .A(n6759), .B(n6758), .Z(n9231) );
  INV_X1 U8336 ( .A(n6758), .ZN(n6760) );
  NOR2_X2 U8337 ( .A1(n9229), .A2(n4978), .ZN(n9201) );
  AOI22_X1 U8338 ( .A1(n9570), .A2(n6778), .B1(n4423), .B2(n9414), .ZN(n6765)
         );
  NAND2_X1 U8339 ( .A1(n9570), .A2(n6761), .ZN(n6763) );
  NAND2_X1 U8340 ( .A1(n9414), .A2(n6778), .ZN(n6762) );
  NAND2_X1 U8341 ( .A1(n6763), .A2(n6762), .ZN(n6764) );
  XNOR2_X1 U8342 ( .A(n6764), .B(n7510), .ZN(n6767) );
  XOR2_X1 U8343 ( .A(n6765), .B(n6767), .Z(n9200) );
  INV_X1 U8344 ( .A(n6765), .ZN(n6766) );
  AOI22_X1 U8345 ( .A1(n9565), .A2(n6784), .B1(n6778), .B2(n9399), .ZN(n6768)
         );
  XOR2_X1 U8346 ( .A(n7510), .B(n6768), .Z(n6771) );
  INV_X1 U8347 ( .A(n9565), .ZN(n9379) );
  INV_X1 U8348 ( .A(n4424), .ZN(n6769) );
  OAI22_X1 U8349 ( .A1(n9379), .A2(n6786), .B1(n9361), .B2(n6769), .ZN(n6770)
         );
  NAND2_X1 U8350 ( .A1(n6771), .A2(n6770), .ZN(n9285) );
  NAND2_X1 U8351 ( .A1(n9561), .A2(n6784), .ZN(n6773) );
  NAND2_X1 U8352 ( .A1(n9353), .A2(n6778), .ZN(n6772) );
  NAND2_X1 U8353 ( .A1(n6773), .A2(n6772), .ZN(n6774) );
  XNOR2_X1 U8354 ( .A(n6774), .B(n6782), .ZN(n6777) );
  AND2_X1 U8355 ( .A1(n4424), .A2(n9353), .ZN(n6775) );
  AOI21_X1 U8356 ( .B1(n9561), .B2(n6778), .A(n6775), .ZN(n6776) );
  NAND2_X1 U8357 ( .A1(n6777), .A2(n6776), .ZN(n6826) );
  OAI21_X1 U8358 ( .B1(n6777), .B2(n6776), .A(n6826), .ZN(n8531) );
  NAND2_X1 U8359 ( .A1(n9555), .A2(n6778), .ZN(n6781) );
  INV_X1 U8360 ( .A(n8534), .ZN(n9367) );
  NAND2_X1 U8361 ( .A1(n9367), .A2(n4423), .ZN(n6780) );
  NAND2_X1 U8362 ( .A1(n6781), .A2(n6780), .ZN(n6783) );
  XNOR2_X1 U8363 ( .A(n6783), .B(n6782), .ZN(n6788) );
  NAND2_X1 U8364 ( .A1(n9555), .A2(n6784), .ZN(n6785) );
  OAI21_X1 U8365 ( .B1(n8534), .B2(n6786), .A(n6785), .ZN(n6787) );
  XNOR2_X1 U8366 ( .A(n6788), .B(n6787), .ZN(n6809) );
  INV_X1 U8367 ( .A(n6809), .ZN(n6827) );
  NAND3_X1 U8368 ( .A1(n8190), .A2(P1_B_REG_SCAN_IN), .A3(n8003), .ZN(n6791)
         );
  INV_X1 U8369 ( .A(n8003), .ZN(n6789) );
  INV_X1 U8370 ( .A(P1_B_REG_SCAN_IN), .ZN(n8347) );
  NAND2_X1 U8371 ( .A1(n6789), .A2(n8347), .ZN(n6790) );
  AND2_X1 U8372 ( .A1(n6791), .A2(n6790), .ZN(n6792) );
  NAND2_X1 U8373 ( .A1(n6793), .A2(n6792), .ZN(n7011) );
  OR2_X1 U8374 ( .A1(n7011), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6795) );
  INV_X1 U8375 ( .A(n6793), .ZN(n8194) );
  NAND2_X1 U8376 ( .A1(n8194), .A2(n8003), .ZN(n6794) );
  NOR4_X1 U8377 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6799) );
  NOR4_X1 U8378 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6798) );
  NOR4_X1 U8379 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6797) );
  NOR4_X1 U8380 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6796) );
  AND4_X1 U8381 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n6805)
         );
  NOR2_X1 U8382 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .ZN(
        n6803) );
  NOR4_X1 U8383 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6802) );
  NOR4_X1 U8384 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6801) );
  NOR4_X1 U8385 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6800) );
  AND4_X1 U8386 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6804)
         );
  NAND2_X1 U8387 ( .A1(n6805), .A2(n6804), .ZN(n7009) );
  INV_X1 U8388 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U8389 ( .A1(n7009), .A2(n10136), .ZN(n6806) );
  OR2_X1 U8390 ( .A1(n7011), .A2(n6806), .ZN(n6807) );
  NAND2_X1 U8391 ( .A1(n8194), .A2(n8190), .ZN(n7008) );
  AND2_X1 U8392 ( .A1(n6807), .A2(n7008), .ZN(n7409) );
  AND2_X1 U8393 ( .A1(n7052), .A2(n7409), .ZN(n6818) );
  NAND2_X1 U8394 ( .A1(n6818), .A2(n6860), .ZN(n6815) );
  NAND2_X1 U8395 ( .A1(n6553), .A2(n6383), .ZN(n7302) );
  NAND2_X1 U8396 ( .A1(n9881), .A2(n7296), .ZN(n6819) );
  NAND3_X1 U8397 ( .A1(n6827), .A2(n9264), .A3(n6826), .ZN(n6808) );
  AND2_X1 U8398 ( .A1(n6809), .A2(n9264), .ZN(n6810) );
  NAND2_X1 U8399 ( .A1(n8530), .A2(n6810), .ZN(n6831) );
  OR2_X1 U8400 ( .A1(n7302), .A2(n4794), .ZN(n7414) );
  NAND2_X1 U8401 ( .A1(n7509), .A2(n7414), .ZN(n6813) );
  INV_X1 U8402 ( .A(n6818), .ZN(n6811) );
  AND2_X1 U8403 ( .A1(n6811), .A2(n6860), .ZN(n6812) );
  NAND2_X1 U8404 ( .A1(n6813), .A2(n6812), .ZN(n6821) );
  OR2_X1 U8405 ( .A1(n7296), .A2(n6552), .ZN(n7017) );
  AND2_X1 U8406 ( .A1(n7116), .A2(n7114), .ZN(n6814) );
  AND2_X1 U8407 ( .A1(n7017), .A2(n6814), .ZN(n7054) );
  NAND3_X1 U8408 ( .A1(n6821), .A2(n7054), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n9237) );
  NOR2_X1 U8409 ( .A1(n7509), .A2(n6815), .ZN(n6817) );
  INV_X1 U8410 ( .A(n6817), .ZN(n6816) );
  AOI22_X1 U8411 ( .A1(n9298), .A2(n9353), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6824) );
  OR2_X1 U8412 ( .A1(n6819), .A2(n6818), .ZN(n7149) );
  NAND2_X1 U8413 ( .A1(n7149), .A2(n7054), .ZN(n6820) );
  NAND2_X1 U8414 ( .A1(n6820), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6822) );
  NAND2_X1 U8415 ( .A1(n9306), .A2(n9348), .ZN(n6823) );
  OAI211_X1 U8416 ( .C1(n6825), .C2(n9301), .A(n6824), .B(n6823), .ZN(n6829)
         );
  NOR3_X1 U8417 ( .A1(n6827), .A2(n6826), .A3(n9309), .ZN(n6828) );
  AOI211_X1 U8418 ( .C1(n9291), .C2(n9555), .A(n6829), .B(n6828), .ZN(n6830)
         );
  NAND3_X1 U8419 ( .A1(n6832), .A2(n6831), .A3(n6830), .ZN(P1_U3218) );
  INV_X1 U8420 ( .A(n6862), .ZN(n6833) );
  OR2_X2 U8421 ( .A1(n7116), .A2(n6833), .ZN(n9324) );
  NOR2_X1 U8422 ( .A1(n4538), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9649) );
  INV_X1 U8423 ( .A(n9649), .ZN(n8540) );
  INV_X1 U8424 ( .A(n7123), .ZN(n7338) );
  OAI222_X1 U8425 ( .A1(n8540), .A2(n6835), .B1(n9651), .B2(n6846), .C1(
        P1_U3084), .C2(n7338), .ZN(P1_U3351) );
  AOI22_X1 U8426 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n9649), .B1(n9718), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6836) );
  OAI21_X1 U8427 ( .B1(n6851), .B2(n9651), .A(n6836), .ZN(P1_U3349) );
  AND2_X1 U8428 ( .A1(n4538), .A2(n4420), .ZN(n9165) );
  AOI22_X1 U8429 ( .A1(n9165), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n8709), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8430 ( .B1(n6841), .B2(n9163), .A(n6838), .ZN(P2_U3357) );
  INV_X1 U8431 ( .A(n7177), .ZN(n9729) );
  OAI222_X1 U8432 ( .A1(n8540), .A2(n6839), .B1(n9651), .B2(n6844), .C1(
        P1_U3084), .C2(n9729), .ZN(P1_U3348) );
  AOI22_X1 U8433 ( .A1(n9752), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9649), .ZN(n6840) );
  OAI21_X1 U8434 ( .B1(n6850), .B2(n9651), .A(n6840), .ZN(P1_U3347) );
  INV_X1 U8435 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6842) );
  INV_X1 U8436 ( .A(n7121), .ZN(n7147) );
  OAI222_X1 U8437 ( .A1(n8540), .A2(n6842), .B1(n9651), .B2(n6841), .C1(
        P1_U3084), .C2(n7147), .ZN(P1_U3352) );
  INV_X1 U8438 ( .A(n7175), .ZN(n7129) );
  OAI222_X1 U8439 ( .A1(n8540), .A2(n6843), .B1(n9651), .B2(n6848), .C1(
        P1_U3084), .C2(n7129), .ZN(P1_U3350) );
  INV_X1 U8440 ( .A(n9165), .ZN(n8345) );
  INV_X1 U8441 ( .A(n8724), .ZN(n6949) );
  OAI222_X1 U8442 ( .A1(n8345), .A2(n6845), .B1(n9163), .B2(n6844), .C1(
        P2_U3152), .C2(n6949), .ZN(P2_U3353) );
  INV_X1 U8443 ( .A(n6907), .ZN(n9657) );
  OAI222_X1 U8444 ( .A1(n8345), .A2(n6847), .B1(n9163), .B2(n6846), .C1(
        P2_U3152), .C2(n9657), .ZN(P2_U3356) );
  INV_X1 U8445 ( .A(n6906), .ZN(n6933) );
  OAI222_X1 U8446 ( .A1(n8345), .A2(n6849), .B1(n9163), .B2(n6848), .C1(
        P2_U3152), .C2(n6933), .ZN(P2_U3355) );
  INV_X1 U8447 ( .A(n7032), .ZN(n6955) );
  OAI222_X1 U8448 ( .A1(n8345), .A2(n10292), .B1(n9163), .B2(n6850), .C1(
        P2_U3152), .C2(n6955), .ZN(P2_U3352) );
  INV_X1 U8449 ( .A(n6950), .ZN(n6920) );
  OAI222_X1 U8450 ( .A1(n8345), .A2(n6852), .B1(n9163), .B2(n6851), .C1(
        P2_U3152), .C2(n6920), .ZN(P2_U3354) );
  INV_X1 U8451 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U8452 ( .A1(n7052), .A2(n6860), .ZN(n6853) );
  OAI21_X1 U8453 ( .B1(n6860), .B2(n6854), .A(n6853), .ZN(P1_U3440) );
  INV_X1 U8454 ( .A(n6855), .ZN(n6858) );
  OAI222_X1 U8455 ( .A1(n8540), .A2(n6857), .B1(n9651), .B2(n6858), .C1(
        P1_U3084), .C2(n6856), .ZN(P1_U3346) );
  INV_X1 U8456 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6859) );
  INV_X1 U8457 ( .A(n8737), .ZN(n6948) );
  OAI222_X1 U8458 ( .A1(n8345), .A2(n6859), .B1(n9163), .B2(n6858), .C1(
        P2_U3152), .C2(n6948), .ZN(P2_U3351) );
  NAND2_X1 U8459 ( .A1(n6860), .A2(n7011), .ZN(n9840) );
  INV_X1 U8460 ( .A(n7008), .ZN(n6861) );
  AOI22_X1 U8461 ( .A1(n9840), .A2(n10136), .B1(n6862), .B2(n6861), .ZN(
        P1_U3441) );
  INV_X1 U8462 ( .A(n6863), .ZN(n6865) );
  INV_X1 U8463 ( .A(n7070), .ZN(n6957) );
  OAI222_X1 U8464 ( .A1(n8345), .A2(n6864), .B1(n9163), .B2(n6865), .C1(
        P2_U3152), .C2(n6957), .ZN(P2_U3350) );
  OAI222_X1 U8465 ( .A1(n8540), .A2(n6866), .B1(n9651), .B2(n6865), .C1(
        P1_U3084), .C2(n7171), .ZN(P1_U3345) );
  NAND2_X1 U8466 ( .A1(n5810), .A2(P2_U3966), .ZN(n6867) );
  OAI21_X1 U8467 ( .B1(n5028), .B2(P2_U3966), .A(n6867), .ZN(P2_U3552) );
  INV_X1 U8468 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U8469 ( .A1(n8779), .A2(P2_U3966), .ZN(n6868) );
  OAI21_X1 U8470 ( .B1(n6869), .B2(P2_U3966), .A(n6868), .ZN(P2_U3583) );
  OAI21_X1 U8471 ( .B1(n9945), .B2(n7085), .A(n6893), .ZN(n6871) );
  NAND2_X1 U8472 ( .A1(n9945), .A2(n6889), .ZN(n6870) );
  NAND2_X1 U8473 ( .A1(n6871), .A2(n6870), .ZN(n9658) );
  INV_X1 U8474 ( .A(n9658), .ZN(n9917) );
  NOR2_X1 U8475 ( .A1(n9917), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8476 ( .A(n6872), .ZN(n6874) );
  OAI222_X1 U8477 ( .A1(n9651), .A2(n6874), .B1(n7179), .B2(P1_U3084), .C1(
        n6873), .C2(n8540), .ZN(P1_U3344) );
  INV_X1 U8478 ( .A(n7045), .ZN(n6959) );
  OAI222_X1 U8479 ( .A1(P2_U3152), .A2(n6959), .B1(n8345), .B2(n5196), .C1(
        n6874), .C2(n9163), .ZN(P2_U3349) );
  INV_X1 U8480 ( .A(n6972), .ZN(n6967) );
  INV_X1 U8481 ( .A(n6875), .ZN(n6878) );
  OAI222_X1 U8482 ( .A1(P2_U3152), .A2(n6967), .B1(n8345), .B2(n5210), .C1(
        n6878), .C2(n9163), .ZN(P2_U3348) );
  NAND2_X1 U8483 ( .A1(n7995), .A2(P1_U4006), .ZN(n6876) );
  OAI21_X1 U8484 ( .B1(P1_U4006), .B2(n5196), .A(n6876), .ZN(P1_U3564) );
  NAND2_X1 U8485 ( .A1(n8004), .A2(P1_U4006), .ZN(n6877) );
  OAI21_X1 U8486 ( .B1(n5210), .B2(P1_U4006), .A(n6877), .ZN(P1_U3565) );
  OAI222_X1 U8487 ( .A1(n8540), .A2(n6879), .B1(n7169), .B2(P1_U3084), .C1(
        n9651), .C2(n6878), .ZN(P1_U3343) );
  INV_X1 U8488 ( .A(n6880), .ZN(n6882) );
  INV_X1 U8489 ( .A(n6976), .ZN(n6992) );
  OAI222_X1 U8490 ( .A1(n8345), .A2(n6881), .B1(n9163), .B2(n6882), .C1(n6992), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  OAI222_X1 U8491 ( .A1(n8540), .A2(n10244), .B1(n7250), .B2(P1_U3084), .C1(
        n9651), .C2(n6882), .ZN(P1_U3342) );
  NAND2_X1 U8492 ( .A1(n9488), .A2(P1_U4006), .ZN(n6883) );
  OAI21_X1 U8493 ( .B1(n5432), .B2(P1_U4006), .A(n6883), .ZN(P1_U3576) );
  INV_X1 U8494 ( .A(n6884), .ZN(n6887) );
  OAI222_X1 U8495 ( .A1(n8540), .A2(n6886), .B1(n9651), .B2(n6887), .C1(
        P1_U3084), .C2(n6885), .ZN(P1_U3341) );
  OAI222_X1 U8496 ( .A1(n8345), .A2(n6888), .B1(n9163), .B2(n6887), .C1(
        P2_U3152), .C2(n6986), .ZN(P2_U3346) );
  INV_X1 U8497 ( .A(n7085), .ZN(n6892) );
  NOR2_X1 U8498 ( .A1(n6913), .A2(n4420), .ZN(n8331) );
  AOI21_X1 U8499 ( .B1(n6890), .B2(n8331), .A(n5793), .ZN(n6891) );
  OAI21_X1 U8500 ( .B1(n9945), .B2(n6892), .A(n6891), .ZN(n6894) );
  NAND2_X1 U8501 ( .A1(n6894), .A2(n6893), .ZN(n6900) );
  INV_X2 U8502 ( .A(P2_U3966), .ZN(n8706) );
  NAND2_X1 U8503 ( .A1(n6900), .A2(n8706), .ZN(n6915) );
  NAND2_X1 U8504 ( .A1(n6915), .A2(n6913), .ZN(n9905) );
  NAND2_X1 U8505 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(n4420), .ZN(n10339) );
  INV_X1 U8506 ( .A(n10339), .ZN(n6905) );
  XNOR2_X1 U8507 ( .A(n8709), .B(n6895), .ZN(n8716) );
  AND2_X1 U8508 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8715) );
  NAND2_X1 U8509 ( .A1(n8716), .A2(n8715), .ZN(n8714) );
  NAND2_X1 U8510 ( .A1(n8709), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8511 ( .A1(n8714), .A2(n6896), .ZN(n9655) );
  XNOR2_X1 U8512 ( .A(n6907), .B(n9989), .ZN(n9656) );
  NAND2_X1 U8513 ( .A1(n9655), .A2(n9656), .ZN(n9654) );
  NAND2_X1 U8514 ( .A1(n6907), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6897) );
  AND2_X1 U8515 ( .A1(n9654), .A2(n6897), .ZN(n6923) );
  OR2_X1 U8516 ( .A1(n6906), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8517 ( .A1(P2_REG1_REG_3__SCAN_IN), .A2(n6906), .ZN(n6898) );
  NAND2_X1 U8518 ( .A1(n6899), .A2(n6898), .ZN(n6922) );
  NOR2_X1 U8519 ( .A1(n6923), .A2(n6922), .ZN(n6921) );
  AOI21_X1 U8520 ( .B1(n6906), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6921), .ZN(
        n6903) );
  XNOR2_X1 U8521 ( .A(n6950), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6902) );
  OR2_X1 U8522 ( .A1(n6902), .A2(n6903), .ZN(n6936) );
  INV_X1 U8523 ( .A(n6936), .ZN(n6901) );
  OR2_X1 U8524 ( .A1(n6900), .A2(n8277), .ZN(n9906) );
  AOI211_X1 U8525 ( .C1(n6903), .C2(n6902), .A(n6901), .B(n9906), .ZN(n6904)
         );
  AOI211_X1 U8526 ( .C1(n9917), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6905), .B(
        n6904), .ZN(n6919) );
  NAND2_X1 U8527 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n6906), .ZN(n6910) );
  AOI22_X1 U8528 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n6906), .B1(n6933), .B2(
        n5076), .ZN(n6930) );
  AOI22_X1 U8529 ( .A1(n6907), .A2(P2_REG2_REG_2__SCAN_IN), .B1(n5050), .B2(
        n9657), .ZN(n9666) );
  INV_X1 U8530 ( .A(n8709), .ZN(n6909) );
  OAI21_X1 U8531 ( .B1(n5050), .B2(n9657), .A(n9664), .ZN(n6929) );
  NAND2_X1 U8532 ( .A1(n6930), .A2(n6929), .ZN(n6928) );
  NAND2_X1 U8533 ( .A1(n6910), .A2(n6928), .ZN(n6917) );
  MUX2_X1 U8534 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6911), .S(n6950), .Z(n6916)
         );
  NOR2_X1 U8535 ( .A1(n6913), .A2(n6912), .ZN(n6914) );
  NAND2_X1 U8536 ( .A1(n6916), .A2(n6917), .ZN(n6951) );
  OAI211_X1 U8537 ( .C1(n6917), .C2(n6916), .A(n9904), .B(n6951), .ZN(n6918)
         );
  OAI211_X1 U8538 ( .C1(n9905), .C2(n6920), .A(n6919), .B(n6918), .ZN(P2_U3249) );
  INV_X1 U8539 ( .A(n9906), .ZN(n9922) );
  AOI21_X1 U8540 ( .B1(n6923), .B2(n6922), .A(n6921), .ZN(n6927) );
  INV_X1 U8541 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6925) );
  INV_X1 U8542 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7226) );
  OR2_X1 U8543 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7226), .ZN(n6924) );
  OAI21_X1 U8544 ( .B1(n9658), .B2(n6925), .A(n6924), .ZN(n6926) );
  AOI21_X1 U8545 ( .B1(n9922), .B2(n6927), .A(n6926), .ZN(n6932) );
  OAI211_X1 U8546 ( .C1(n6930), .C2(n6929), .A(n9904), .B(n6928), .ZN(n6931)
         );
  OAI211_X1 U8547 ( .C1(n9905), .C2(n6933), .A(n6932), .B(n6931), .ZN(P2_U3248) );
  NAND2_X1 U8548 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(n4420), .ZN(n7952) );
  INV_X1 U8549 ( .A(n7952), .ZN(n6947) );
  MUX2_X1 U8550 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n5218), .S(n6972), .Z(n6944)
         );
  NAND2_X1 U8551 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n8724), .ZN(n6937) );
  OAI21_X1 U8552 ( .B1(n8724), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6937), .ZN(
        n6934) );
  INV_X1 U8553 ( .A(n6934), .ZN(n8728) );
  NAND2_X1 U8554 ( .A1(n6950), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U8555 ( .A1(n6936), .A2(n6935), .ZN(n8727) );
  NAND2_X1 U8556 ( .A1(n8728), .A2(n8727), .ZN(n8726) );
  NAND2_X1 U8557 ( .A1(n8726), .A2(n6937), .ZN(n7026) );
  MUX2_X1 U8558 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n5126), .S(n7032), .Z(n7027)
         );
  NAND2_X1 U8559 ( .A1(n7026), .A2(n7027), .ZN(n7025) );
  NAND2_X1 U8560 ( .A1(n7032), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8561 ( .A1(n7025), .A2(n6938), .ZN(n8740) );
  NAND2_X1 U8562 ( .A1(n8737), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6940) );
  OAI21_X1 U8563 ( .B1(n8737), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6940), .ZN(
        n6939) );
  INV_X1 U8564 ( .A(n6939), .ZN(n8741) );
  NAND2_X1 U8565 ( .A1(n8740), .A2(n8741), .ZN(n8739) );
  NAND2_X1 U8566 ( .A1(n8739), .A2(n6940), .ZN(n7060) );
  MUX2_X1 U8567 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n5187), .S(n7070), .Z(n7061)
         );
  NAND2_X1 U8568 ( .A1(n7060), .A2(n7061), .ZN(n7059) );
  NAND2_X1 U8569 ( .A1(n7070), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8570 ( .A1(n7059), .A2(n6941), .ZN(n7039) );
  MUX2_X1 U8571 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n5203), .S(n7045), .Z(n7040)
         );
  NAND2_X1 U8572 ( .A1(n7039), .A2(n7040), .ZN(n7038) );
  NAND2_X1 U8573 ( .A1(n7045), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8574 ( .A1(n7038), .A2(n6942), .ZN(n6943) );
  NAND2_X1 U8575 ( .A1(n6943), .A2(n6944), .ZN(n6974) );
  OAI211_X1 U8576 ( .C1(n6944), .C2(n6943), .A(n9922), .B(n6974), .ZN(n6945)
         );
  INV_X1 U8577 ( .A(n6945), .ZN(n6946) );
  AOI211_X1 U8578 ( .C1(n9917), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6947), .B(
        n6946), .ZN(n6963) );
  NAND2_X1 U8579 ( .A1(n8737), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6956) );
  AOI22_X1 U8580 ( .A1(n8737), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n5158), .B2(
        n6948), .ZN(n8736) );
  NAND2_X1 U8581 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n8724), .ZN(n6953) );
  AOI22_X1 U8582 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n8724), .B1(n6949), .B2(
        n7760), .ZN(n8723) );
  NAND2_X1 U8583 ( .A1(n6950), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8584 ( .A1(n6952), .A2(n6951), .ZN(n8722) );
  NAND2_X1 U8585 ( .A1(n8723), .A2(n8722), .ZN(n8721) );
  NAND2_X1 U8586 ( .A1(n6953), .A2(n8721), .ZN(n7035) );
  MUX2_X1 U8587 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6954), .S(n7032), .Z(n7034)
         );
  NAND2_X1 U8588 ( .A1(n7035), .A2(n7034), .ZN(n7033) );
  OAI21_X1 U8589 ( .B1(n6954), .B2(n6955), .A(n7033), .ZN(n8735) );
  NAND2_X1 U8590 ( .A1(n8736), .A2(n8735), .ZN(n8734) );
  AND2_X1 U8591 ( .A1(n6956), .A2(n8734), .ZN(n7067) );
  MUX2_X1 U8592 ( .A(n5186), .B(P2_REG2_REG_8__SCAN_IN), .S(n7070), .Z(n7066)
         );
  NOR2_X1 U8593 ( .A1(n6957), .A2(n5186), .ZN(n7047) );
  MUX2_X1 U8594 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6958), .S(n7045), .Z(n7046)
         );
  AOI22_X1 U8595 ( .A1(n6972), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7945), .B2(
        n6967), .ZN(n6960) );
  OAI211_X1 U8596 ( .C1(n6961), .C2(n6960), .A(n9904), .B(n6966), .ZN(n6962)
         );
  OAI211_X1 U8597 ( .C1(n9905), .C2(n6967), .A(n6963), .B(n6962), .ZN(P2_U3255) );
  INV_X1 U8598 ( .A(n6964), .ZN(n7002) );
  AOI22_X1 U8599 ( .A1(n7923), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9649), .ZN(n6965) );
  OAI21_X1 U8600 ( .B1(n7002), .B2(n9651), .A(n6965), .ZN(P1_U3340) );
  NOR2_X1 U8601 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n6976), .ZN(n6968) );
  OAI21_X1 U8602 ( .B1(n7945), .B2(n6967), .A(n6966), .ZN(n6989) );
  AOI22_X1 U8603 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n6992), .B1(n6976), .B2(
        n8039), .ZN(n6988) );
  NOR2_X1 U8604 ( .A1(n6989), .A2(n6988), .ZN(n6987) );
  NOR2_X1 U8605 ( .A1(n6968), .A2(n6987), .ZN(n6971) );
  MUX2_X1 U8606 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n5266), .S(n6986), .Z(n6969)
         );
  INV_X1 U8607 ( .A(n6969), .ZN(n6970) );
  NAND2_X1 U8608 ( .A1(n6970), .A2(n6971), .ZN(n7201) );
  OAI211_X1 U8609 ( .C1(n6971), .C2(n6970), .A(n9904), .B(n7201), .ZN(n6985)
         );
  NAND2_X1 U8610 ( .A1(n6972), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6973) );
  AND2_X1 U8611 ( .A1(n6974), .A2(n6973), .ZN(n6996) );
  INV_X1 U8612 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6975) );
  MUX2_X1 U8613 ( .A(n6975), .B(P2_REG1_REG_11__SCAN_IN), .S(n6976), .Z(n6995)
         );
  NOR2_X1 U8614 ( .A1(n6996), .A2(n6995), .ZN(n6994) );
  AOI21_X1 U8615 ( .B1(n6976), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6994), .ZN(
        n6979) );
  MUX2_X1 U8616 ( .A(n6977), .B(P2_REG1_REG_12__SCAN_IN), .S(n6986), .Z(n6978)
         );
  NAND2_X1 U8617 ( .A1(n6978), .A2(n6979), .ZN(n7208) );
  OAI21_X1 U8618 ( .B1(n6979), .B2(n6978), .A(n7208), .ZN(n6983) );
  NAND2_X1 U8619 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(n4420), .ZN(n8030) );
  INV_X1 U8620 ( .A(n8030), .ZN(n6982) );
  INV_X1 U8621 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U8622 ( .A1(n9658), .A2(n6980), .ZN(n6981) );
  AOI211_X1 U8623 ( .C1(n9922), .C2(n6983), .A(n6982), .B(n6981), .ZN(n6984)
         );
  OAI211_X1 U8624 ( .C1(n9905), .C2(n6986), .A(n6985), .B(n6984), .ZN(P2_U3257) );
  AOI21_X1 U8625 ( .B1(n6989), .B2(n6988), .A(n6987), .ZN(n7001) );
  INV_X1 U8626 ( .A(n9904), .ZN(n9927) );
  NOR2_X1 U8627 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7858), .ZN(n6990) );
  AOI21_X1 U8628 ( .B1(n9917), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6990), .ZN(
        n6991) );
  OAI21_X1 U8629 ( .B1(n9905), .B2(n6992), .A(n6991), .ZN(n6993) );
  INV_X1 U8630 ( .A(n6993), .ZN(n7000) );
  INV_X1 U8631 ( .A(n6994), .ZN(n6998) );
  NAND2_X1 U8632 ( .A1(n6996), .A2(n6995), .ZN(n6997) );
  NAND3_X1 U8633 ( .A1(n9922), .A2(n6998), .A3(n6997), .ZN(n6999) );
  OAI211_X1 U8634 ( .C1(n7001), .C2(n9927), .A(n7000), .B(n6999), .ZN(P2_U3256) );
  INV_X1 U8635 ( .A(n9923), .ZN(n7207) );
  OAI222_X1 U8636 ( .A1(n8345), .A2(n7003), .B1(n9163), .B2(n7002), .C1(n7207), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8637 ( .A(n7004), .ZN(n7005) );
  OAI222_X1 U8638 ( .A1(n9651), .A2(n7005), .B1(n7921), .B2(P1_U3084), .C1(
        n10315), .C2(n8540), .ZN(P1_U3339) );
  INV_X1 U8639 ( .A(n7660), .ZN(n7212) );
  OAI222_X1 U8640 ( .A1(n8345), .A2(n7006), .B1(n9163), .B2(n7005), .C1(n7212), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OR2_X1 U8641 ( .A1(n9876), .A2(n7412), .ZN(n7015) );
  OAI21_X1 U8642 ( .B1(n7011), .B2(P1_D_REG_1__SCAN_IN), .A(n7008), .ZN(n7013)
         );
  INV_X1 U8643 ( .A(n7009), .ZN(n7010) );
  OR2_X1 U8644 ( .A1(n7011), .A2(n7010), .ZN(n7012) );
  AND2_X1 U8645 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  NOR2_X1 U8646 ( .A1(n7411), .A2(n7052), .ZN(n7016) );
  INV_X1 U8647 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7024) );
  NAND3_X1 U8648 ( .A1(n7018), .A2(n7509), .A3(n7302), .ZN(n7020) );
  NAND2_X1 U8649 ( .A1(n9539), .A2(n6564), .ZN(n7019) );
  NAND2_X1 U8650 ( .A1(n7020), .A2(n7019), .ZN(n7416) );
  INV_X1 U8651 ( .A(n7416), .ZN(n7021) );
  OAI21_X1 U8652 ( .B1(n7022), .B2(n7302), .A(n7021), .ZN(n7057) );
  NAND2_X1 U8653 ( .A1(n7057), .A2(n9891), .ZN(n7023) );
  OAI21_X1 U8654 ( .B1(n9891), .B2(n7024), .A(n7023), .ZN(P1_U3454) );
  INV_X1 U8655 ( .A(n9905), .ZN(n9924) );
  OAI21_X1 U8656 ( .B1(n7027), .B2(n7026), .A(n7025), .ZN(n7030) );
  NOR2_X1 U8657 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7370), .ZN(n7028) );
  AOI21_X1 U8658 ( .B1(n9917), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7028), .ZN(
        n7029) );
  OAI21_X1 U8659 ( .B1(n9906), .B2(n7030), .A(n7029), .ZN(n7031) );
  AOI21_X1 U8660 ( .B1(n7032), .B2(n9924), .A(n7031), .ZN(n7037) );
  OAI211_X1 U8661 ( .C1(n7035), .C2(n7034), .A(n9904), .B(n7033), .ZN(n7036)
         );
  NAND2_X1 U8662 ( .A1(n7037), .A2(n7036), .ZN(P2_U3251) );
  OAI21_X1 U8663 ( .B1(n7040), .B2(n7039), .A(n7038), .ZN(n7043) );
  AND2_X1 U8664 ( .A1(n4420), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7041) );
  AOI21_X1 U8665 ( .B1(n9917), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7041), .ZN(
        n7042) );
  OAI21_X1 U8666 ( .B1(n9906), .B2(n7043), .A(n7042), .ZN(n7044) );
  AOI21_X1 U8667 ( .B1(n7045), .B2(n9924), .A(n7044), .ZN(n7051) );
  OR3_X1 U8668 ( .A1(n7065), .A2(n7047), .A3(n7046), .ZN(n7048) );
  NAND3_X1 U8669 ( .A1(n7049), .A2(n9904), .A3(n7048), .ZN(n7050) );
  NAND2_X1 U8670 ( .A1(n7051), .A2(n7050), .ZN(P2_U3254) );
  AND2_X1 U8671 ( .A1(n7052), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7053) );
  INV_X1 U8672 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U8673 ( .A1(n7057), .A2(n9903), .ZN(n7058) );
  OAI21_X1 U8674 ( .B1(n9903), .B2(n10227), .A(n7058), .ZN(P1_U3523) );
  OAI21_X1 U8675 ( .B1(n7061), .B2(n7060), .A(n7059), .ZN(n7064) );
  NOR2_X1 U8676 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10175), .ZN(n7062) );
  AOI21_X1 U8677 ( .B1(n9917), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7062), .ZN(
        n7063) );
  OAI21_X1 U8678 ( .B1(n9906), .B2(n7064), .A(n7063), .ZN(n7069) );
  AOI211_X1 U8679 ( .C1(n7067), .C2(n7066), .A(n7065), .B(n9927), .ZN(n7068)
         );
  AOI211_X1 U8680 ( .C1(n9924), .C2(n7070), .A(n7069), .B(n7068), .ZN(n7071)
         );
  INV_X1 U8681 ( .A(n7071), .ZN(P2_U3253) );
  NAND2_X1 U8682 ( .A1(n7073), .A2(n7072), .ZN(n7074) );
  OR2_X1 U8683 ( .A1(n7075), .A2(n7074), .ZN(n7081) );
  OAI21_X1 U8684 ( .B1(n7076), .B2(n9979), .A(n7081), .ZN(n7079) );
  INV_X1 U8685 ( .A(n7077), .ZN(n7078) );
  NAND2_X1 U8686 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  NAND2_X1 U8687 ( .A1(n7080), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10341) );
  INV_X1 U8688 ( .A(n10341), .ZN(n8674) );
  NOR2_X1 U8689 ( .A1(n8674), .A2(n4420), .ZN(n8641) );
  NOR2_X1 U8690 ( .A1(n7081), .A2(n9945), .ZN(n7098) );
  NAND2_X1 U8691 ( .A1(n7098), .A2(n7082), .ZN(n8637) );
  INV_X1 U8692 ( .A(n8637), .ZN(n7482) );
  NAND2_X1 U8693 ( .A1(n8705), .A2(n8945), .ZN(n7084) );
  INV_X1 U8694 ( .A(n8977), .ZN(n8943) );
  NAND2_X1 U8695 ( .A1(n5810), .A2(n8943), .ZN(n7083) );
  NAND2_X1 U8696 ( .A1(n7084), .A2(n7083), .ZN(n7197) );
  AND2_X1 U8697 ( .A1(n9979), .A2(n7085), .ZN(n7086) );
  INV_X2 U8698 ( .A(n8432), .ZN(n8455) );
  OR2_X1 U8699 ( .A1(n7191), .A2(n8455), .ZN(n7131) );
  NAND2_X4 U8700 ( .A1(n7090), .A2(n7089), .ZN(n8453) );
  NAND2_X1 U8701 ( .A1(n8448), .A2(n7192), .ZN(n7091) );
  AND2_X1 U8702 ( .A1(n8707), .A2(n8432), .ZN(n7231) );
  OAI21_X1 U8703 ( .B1(n7094), .B2(n7093), .A(n8646), .ZN(n7095) );
  AOI22_X1 U8704 ( .A1(n7482), .A2(n7197), .B1(n8629), .B2(n7095), .ZN(n7101)
         );
  INV_X1 U8705 ( .A(n7096), .ZN(n7097) );
  NAND2_X1 U8706 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  NAND2_X1 U8707 ( .A1(n7099), .A2(n8989), .ZN(n8668) );
  NAND2_X1 U8708 ( .A1(n8668), .A2(n5046), .ZN(n7100) );
  OAI211_X1 U8709 ( .C1(n8641), .C2(n7594), .A(n7101), .B(n7100), .ZN(P2_U3224) );
  INV_X1 U8710 ( .A(n8982), .ZN(n8954) );
  OAI22_X1 U8711 ( .A1(n7759), .A2(n8954), .B1(n5047), .B2(n8979), .ZN(n7755)
         );
  INV_X1 U8712 ( .A(n9985), .ZN(n9090) );
  OAI22_X1 U8713 ( .A1(n7759), .A2(n9090), .B1(n7102), .B2(n7192), .ZN(n7103)
         );
  OR2_X1 U8714 ( .A1(n7755), .A2(n7103), .ZN(n7344) );
  NAND2_X1 U8715 ( .A1(n9996), .A2(n7344), .ZN(n7104) );
  OAI21_X1 U8716 ( .B1(n9996), .B2(n5041), .A(n7104), .ZN(P2_U3520) );
  NAND2_X1 U8717 ( .A1(n7296), .A2(n7116), .ZN(n7105) );
  NAND2_X1 U8718 ( .A1(n7105), .A2(n7114), .ZN(n7108) );
  NAND2_X1 U8719 ( .A1(n7108), .A2(n7106), .ZN(n7107) );
  NAND2_X1 U8720 ( .A1(n7107), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U8721 ( .A1(n7108), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7111) );
  OR2_X1 U8722 ( .A1(n7111), .A2(n8348), .ZN(n8371) );
  INV_X1 U8723 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7109) );
  MUX2_X1 U8724 ( .A(n7109), .B(P1_REG1_REG_1__SCAN_IN), .S(n7121), .Z(n7138)
         );
  NOR3_X1 U8725 ( .A1(n7138), .A2(n10227), .A3(n5986), .ZN(n7137) );
  AOI21_X1 U8726 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n7121), .A(n7137), .ZN(
        n7333) );
  XNOR2_X1 U8727 ( .A(n7123), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7332) );
  NOR2_X1 U8728 ( .A1(n7333), .A2(n7332), .ZN(n7331) );
  AOI21_X1 U8729 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n7123), .A(n7331), .ZN(
        n7113) );
  XNOR2_X1 U8730 ( .A(n7175), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n7112) );
  NOR2_X1 U8731 ( .A1(n7113), .A2(n7112), .ZN(n7174) );
  OR2_X1 U8732 ( .A1(n7111), .A2(n7110), .ZN(n9713) );
  AOI211_X1 U8733 ( .C1(n7113), .C2(n7112), .A(n7174), .B(n9833), .ZN(n7120)
         );
  NOR2_X1 U8734 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10165), .ZN(n7221) );
  INV_X1 U8735 ( .A(n7114), .ZN(n7115) );
  NOR2_X1 U8736 ( .A1(n7116), .A2(n7115), .ZN(n7117) );
  OR2_X1 U8737 ( .A1(P1_U3083), .A2(n7117), .ZN(n9821) );
  INV_X1 U8738 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7118) );
  NOR2_X1 U8739 ( .A1(n9821), .A2(n7118), .ZN(n7119) );
  NOR3_X1 U8740 ( .A1(n7120), .A2(n7221), .A3(n7119), .ZN(n7128) );
  OR2_X1 U8741 ( .A1(n8371), .A2(n6535), .ZN(n9782) );
  XOR2_X1 U8742 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7123), .Z(n7336) );
  INV_X1 U8743 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7122) );
  MUX2_X1 U8744 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7122), .S(n7121), .Z(n7144)
         );
  INV_X1 U8745 ( .A(n7325), .ZN(n7143) );
  NAND2_X1 U8746 ( .A1(n7144), .A2(n7143), .ZN(n7142) );
  NAND2_X1 U8747 ( .A1(n7175), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7159) );
  OAI21_X1 U8748 ( .B1(n7175), .B2(P1_REG2_REG_3__SCAN_IN), .A(n7159), .ZN(
        n7124) );
  OR2_X1 U8749 ( .A1(n7125), .A2(n7124), .ZN(n7160) );
  NAND2_X1 U8750 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  NAND3_X1 U8751 ( .A1(n9823), .A2(n7160), .A3(n7126), .ZN(n7127) );
  OAI211_X1 U8752 ( .C1(n9828), .C2(n7129), .A(n7128), .B(n7127), .ZN(P1_U3244) );
  AND2_X1 U8753 ( .A1(n8629), .A2(n8432), .ZN(n8627) );
  INV_X1 U8754 ( .A(n5810), .ZN(n7130) );
  OAI22_X1 U8755 ( .A1(n8456), .A2(n7130), .B1(n7192), .B2(n10351), .ZN(n7132)
         );
  NAND2_X1 U8756 ( .A1(n7132), .A2(n7131), .ZN(n7134) );
  AOI22_X1 U8757 ( .A1(n8675), .A2(n8707), .B1(n7754), .B2(n8668), .ZN(n7133)
         );
  OAI211_X1 U8758 ( .C1(n8641), .C2(n7135), .A(n7134), .B(n7133), .ZN(P2_U3234) );
  INV_X1 U8759 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7136) );
  NOR2_X1 U8760 ( .A1(n9821), .A2(n7136), .ZN(n7141) );
  AOI211_X1 U8761 ( .C1(n7139), .C2(n7138), .A(n7137), .B(n9833), .ZN(n7140)
         );
  AOI211_X1 U8762 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n7141), .B(
        n7140), .ZN(n7146) );
  OAI211_X1 U8763 ( .C1(n7144), .C2(n7143), .A(n9823), .B(n7142), .ZN(n7145)
         );
  OAI211_X1 U8764 ( .C1(n9828), .C2(n7147), .A(n7146), .B(n7145), .ZN(P1_U3242) );
  NAND2_X1 U8765 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8706), .ZN(n7148) );
  OAI21_X1 U8766 ( .B1(n8460), .B2(n8706), .A(n7148), .ZN(P2_U3581) );
  INV_X1 U8767 ( .A(n7149), .ZN(n7150) );
  OR2_X1 U8768 ( .A1(n7150), .A2(n9237), .ZN(n9269) );
  AOI22_X1 U8769 ( .A1(n9291), .A2(n7457), .B1(n9269), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7155) );
  OAI21_X1 U8770 ( .B1(n7151), .B2(n7153), .A(n7152), .ZN(n7326) );
  AOI22_X1 U8771 ( .A1(n7326), .A2(n9264), .B1(n9266), .B2(n6564), .ZN(n7154)
         );
  NAND2_X1 U8772 ( .A1(n7155), .A2(n7154), .ZN(P1_U3230) );
  INV_X1 U8773 ( .A(n9828), .ZN(n9808) );
  INV_X1 U8774 ( .A(n7169), .ZN(n7252) );
  INV_X1 U8775 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U8776 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8066) );
  OAI21_X1 U8777 ( .B1(n9821), .B2(n7156), .A(n8066), .ZN(n7168) );
  INV_X1 U8778 ( .A(n7179), .ZN(n9787) );
  NOR2_X1 U8779 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9769), .ZN(n7157) );
  AOI21_X1 U8780 ( .B1(n9769), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7157), .ZN(
        n9775) );
  NOR2_X1 U8781 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9756), .ZN(n7158) );
  AOI21_X1 U8782 ( .B1(n9756), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7158), .ZN(
        n9761) );
  NOR2_X1 U8783 ( .A1(n7177), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7162) );
  AOI21_X1 U8784 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7177), .A(n7162), .ZN(
        n9733) );
  NOR2_X1 U8785 ( .A1(n9718), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7161) );
  AOI21_X1 U8786 ( .B1(n9718), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7161), .ZN(
        n9721) );
  NAND2_X1 U8787 ( .A1(n9733), .A2(n9732), .ZN(n9731) );
  INV_X1 U8788 ( .A(n7162), .ZN(n7163) );
  NAND2_X1 U8789 ( .A1(n9731), .A2(n7163), .ZN(n9748) );
  XNOR2_X1 U8790 ( .A(n9752), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9749) );
  NOR2_X1 U8791 ( .A1(n9748), .A2(n9749), .ZN(n9747) );
  OAI21_X1 U8792 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9769), .A(n9773), .ZN(
        n9783) );
  XNOR2_X1 U8793 ( .A(n9787), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n9784) );
  NOR2_X1 U8794 ( .A1(n9783), .A2(n9784), .ZN(n9781) );
  NAND2_X1 U8795 ( .A1(n7252), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7164) );
  OAI21_X1 U8796 ( .B1(n7252), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7164), .ZN(
        n7165) );
  AOI211_X1 U8797 ( .C1(n7166), .C2(n7165), .A(n9782), .B(n7251), .ZN(n7167)
         );
  AOI211_X1 U8798 ( .C1(n9808), .C2(n7252), .A(n7168), .B(n7167), .ZN(n7185)
         );
  INV_X1 U8799 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7170) );
  MUX2_X1 U8800 ( .A(n7170), .B(P1_REG1_REG_10__SCAN_IN), .S(n7169), .Z(n7182)
         );
  INV_X1 U8801 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U8802 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n9769), .B1(n7171), .B2(
        n9899), .ZN(n9772) );
  NOR2_X1 U8803 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9756), .ZN(n7172) );
  AOI21_X1 U8804 ( .B1(n9756), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7172), .ZN(
        n9759) );
  XNOR2_X1 U8805 ( .A(n9752), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U8806 ( .A1(n7177), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7173) );
  OAI21_X1 U8807 ( .B1(n7177), .B2(P1_REG1_REG_5__SCAN_IN), .A(n7173), .ZN(
        n9735) );
  AOI21_X1 U8808 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n7175), .A(n7174), .ZN(
        n9716) );
  NOR2_X1 U8809 ( .A1(n9718), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7176) );
  AOI21_X1 U8810 ( .B1(n9718), .B2(P1_REG1_REG_4__SCAN_IN), .A(n7176), .ZN(
        n9717) );
  NAND2_X1 U8811 ( .A1(n9716), .A2(n9717), .ZN(n9715) );
  OAI21_X1 U8812 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9718), .A(n9715), .ZN(
        n9736) );
  NOR2_X1 U8813 ( .A1(n9735), .A2(n9736), .ZN(n9734) );
  AOI21_X1 U8814 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n7177), .A(n9734), .ZN(
        n9742) );
  INV_X1 U8815 ( .A(n9742), .ZN(n7178) );
  OAI22_X1 U8816 ( .A1(n9743), .A2(n7178), .B1(n9752), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U8817 ( .A1(n9759), .A2(n9758), .ZN(n9757) );
  OAI21_X1 U8818 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n9756), .A(n9757), .ZN(
        n9771) );
  NAND2_X1 U8819 ( .A1(n9772), .A2(n9771), .ZN(n9770) );
  OAI21_X1 U8820 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9769), .A(n9770), .ZN(
        n9790) );
  INV_X1 U8821 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7180) );
  MUX2_X1 U8822 ( .A(n7180), .B(P1_REG1_REG_9__SCAN_IN), .S(n7179), .Z(n9789)
         );
  NAND2_X1 U8823 ( .A1(n9790), .A2(n9789), .ZN(n9788) );
  OAI21_X1 U8824 ( .B1(n9787), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9788), .ZN(
        n7181) );
  NAND2_X1 U8825 ( .A1(n7181), .A2(n7182), .ZN(n7244) );
  OAI21_X1 U8826 ( .B1(n7182), .B2(n7181), .A(n7244), .ZN(n7183) );
  NAND2_X1 U8827 ( .A1(n7183), .A2(n9816), .ZN(n7184) );
  NAND2_X1 U8828 ( .A1(n7185), .A2(n7184), .ZN(P1_U3251) );
  INV_X1 U8829 ( .A(n7186), .ZN(n7188) );
  INV_X1 U8830 ( .A(n7679), .ZN(n7668) );
  OAI222_X1 U8831 ( .A1(n8345), .A2(n7187), .B1(n9163), .B2(n7188), .C1(
        P2_U3152), .C2(n7668), .ZN(P2_U3343) );
  OAI222_X1 U8832 ( .A1(n8540), .A2(n7189), .B1(n9651), .B2(n7188), .C1(
        P1_U3084), .C2(n8099), .ZN(P1_U3338) );
  OAI21_X1 U8833 ( .B1(n5811), .B2(n7191), .A(n7190), .ZN(n7592) );
  OAI21_X1 U8834 ( .B1(n7408), .B2(n7192), .A(n9959), .ZN(n7193) );
  NOR2_X1 U8835 ( .A1(n7193), .A2(n7622), .ZN(n7596) );
  INV_X1 U8836 ( .A(n7194), .ZN(n7195) );
  XNOR2_X1 U8837 ( .A(n7196), .B(n7195), .ZN(n7198) );
  AOI21_X1 U8838 ( .B1(n7198), .B2(n8982), .A(n7197), .ZN(n7593) );
  INV_X1 U8839 ( .A(n7593), .ZN(n7199) );
  AOI211_X1 U8840 ( .C1(n9985), .C2(n7592), .A(n7596), .B(n7199), .ZN(n7406)
         );
  MUX2_X1 U8841 ( .A(n6895), .B(n7406), .S(n9996), .Z(n7200) );
  OAI21_X1 U8842 ( .B1(n7408), .B2(n9071), .A(n7200), .ZN(P2_U3521) );
  NOR2_X1 U8843 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n9923), .ZN(n7203) );
  NAND2_X1 U8844 ( .A1(n7209), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U8845 ( .A1(n7202), .A2(n7201), .ZN(n9914) );
  AOI22_X1 U8846 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n7207), .B1(n9923), .B2(
        n8243), .ZN(n9913) );
  NOR2_X1 U8847 ( .A1(n9914), .A2(n9913), .ZN(n9912) );
  AOI22_X1 U8848 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7212), .B1(n7660), .B2(
        n5309), .ZN(n7204) );
  AOI21_X1 U8849 ( .B1(n7205), .B2(n7204), .A(n7655), .ZN(n7217) );
  AOI22_X1 U8850 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7660), .B1(n7212), .B2(
        n7206), .ZN(n7211) );
  AOI22_X1 U8851 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9923), .B1(n7207), .B2(
        n5285), .ZN(n9919) );
  OAI21_X1 U8852 ( .B1(n7209), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7208), .ZN(
        n9920) );
  NAND2_X1 U8853 ( .A1(n9919), .A2(n9920), .ZN(n9918) );
  OAI21_X1 U8854 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9923), .A(n9918), .ZN(
        n7210) );
  NAND2_X1 U8855 ( .A1(n7211), .A2(n7210), .ZN(n7659) );
  OAI21_X1 U8856 ( .B1(n7211), .B2(n7210), .A(n7659), .ZN(n7215) );
  NOR2_X1 U8857 ( .A1(n9905), .A2(n7212), .ZN(n7214) );
  INV_X1 U8858 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U8859 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(n4420), .ZN(n8223) );
  OAI21_X1 U8860 ( .B1(n9658), .B2(n10300), .A(n8223), .ZN(n7213) );
  AOI211_X1 U8861 ( .C1(n7215), .C2(n9922), .A(n7214), .B(n7213), .ZN(n7216)
         );
  OAI21_X1 U8862 ( .B1(n7217), .B2(n9927), .A(n7216), .ZN(P2_U3259) );
  INV_X1 U8863 ( .A(n9306), .ZN(n9281) );
  OAI21_X1 U8864 ( .B1(n7219), .B2(n7218), .A(n7274), .ZN(n7220) );
  NAND2_X1 U8865 ( .A1(n7220), .A2(n9264), .ZN(n7225) );
  INV_X1 U8866 ( .A(n9322), .ZN(n7541) );
  AOI21_X1 U8867 ( .B1(n9298), .B2(n6573), .A(n7221), .ZN(n7222) );
  OAI21_X1 U8868 ( .B1(n7541), .B2(n9301), .A(n7222), .ZN(n7223) );
  AOI21_X1 U8869 ( .B1(n9291), .B2(n4422), .A(n7223), .ZN(n7224) );
  OAI211_X1 U8870 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9281), .A(n7225), .B(
        n7224), .ZN(P1_U3216) );
  OAI22_X1 U8871 ( .A1(n10341), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n7226), .ZN(n7229) );
  OAI22_X1 U8872 ( .A1(n10345), .A2(n7436), .B1(n10343), .B2(n7227), .ZN(n7228) );
  AOI211_X1 U8873 ( .C1(n10349), .C2(n8705), .A(n7229), .B(n7228), .ZN(n7243)
         );
  XNOR2_X1 U8874 ( .A(n7436), .B(n8453), .ZN(n7352) );
  NAND2_X1 U8875 ( .A1(n10348), .A2(n8432), .ZN(n7353) );
  XNOR2_X1 U8876 ( .A(n7352), .B(n7353), .ZN(n7239) );
  INV_X1 U8877 ( .A(n7231), .ZN(n7232) );
  NAND2_X1 U8878 ( .A1(n7230), .A2(n7232), .ZN(n7233) );
  XNOR2_X1 U8879 ( .A(n9962), .B(n8453), .ZN(n7236) );
  AND2_X1 U8880 ( .A1(n8705), .A2(n8432), .ZN(n7234) );
  XNOR2_X1 U8881 ( .A(n7236), .B(n7234), .ZN(n8645) );
  INV_X1 U8882 ( .A(n7234), .ZN(n7235) );
  NAND2_X1 U8883 ( .A1(n7236), .A2(n7235), .ZN(n7237) );
  AOI21_X1 U8884 ( .B1(n7239), .B2(n7238), .A(n10351), .ZN(n7241) );
  NAND2_X1 U8885 ( .A1(n7241), .A2(n7357), .ZN(n7242) );
  NAND2_X1 U8886 ( .A1(n7243), .A2(n7242), .ZN(P2_U3220) );
  INV_X1 U8887 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10241) );
  MUX2_X1 U8888 ( .A(n10241), .B(P1_REG1_REG_12__SCAN_IN), .S(n7399), .Z(n7248) );
  INV_X1 U8889 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7246) );
  MUX2_X1 U8890 ( .A(n7246), .B(P1_REG1_REG_11__SCAN_IN), .S(n7250), .Z(n9797)
         );
  OAI21_X1 U8891 ( .B1(n7252), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7244), .ZN(
        n9798) );
  NAND2_X1 U8892 ( .A1(n9797), .A2(n9798), .ZN(n9796) );
  INV_X1 U8893 ( .A(n9796), .ZN(n7245) );
  AOI21_X1 U8894 ( .B1(n7246), .B2(n7250), .A(n7245), .ZN(n7247) );
  NOR2_X1 U8895 ( .A1(n7247), .A2(n7248), .ZN(n7390) );
  AOI21_X1 U8896 ( .B1(n7248), .B2(n7247), .A(n7390), .ZN(n7261) );
  NAND2_X1 U8897 ( .A1(n7399), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7249) );
  OAI21_X1 U8898 ( .B1(n7399), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7249), .ZN(
        n7255) );
  INV_X1 U8899 ( .A(n7250), .ZN(n9795) );
  XNOR2_X1 U8900 ( .A(n7250), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n9800) );
  OAI21_X1 U8901 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9795), .A(n7253), .ZN(
        n7254) );
  NOR2_X1 U8902 ( .A1(n7254), .A2(n7255), .ZN(n7398) );
  AOI211_X1 U8903 ( .C1(n7255), .C2(n7254), .A(n7398), .B(n9782), .ZN(n7256)
         );
  AOI21_X1 U8904 ( .B1(n9808), .B2(n7399), .A(n7256), .ZN(n7260) );
  INV_X1 U8905 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U8906 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8116) );
  OAI21_X1 U8907 ( .B1(n9821), .B2(n7257), .A(n8116), .ZN(n7258) );
  INV_X1 U8908 ( .A(n7258), .ZN(n7259) );
  OAI211_X1 U8909 ( .C1(n7261), .C2(n9833), .A(n7260), .B(n7259), .ZN(P1_U3253) );
  NAND2_X1 U8910 ( .A1(n7262), .A2(n7263), .ZN(n7265) );
  XNOR2_X1 U8911 ( .A(n7265), .B(n7264), .ZN(n7270) );
  AOI22_X1 U8912 ( .A1(n9266), .A2(n6573), .B1(n9298), .B2(n9325), .ZN(n7267)
         );
  OAI21_X1 U8913 ( .B1(n7266), .B2(n9303), .A(n7267), .ZN(n7268) );
  AOI21_X1 U8914 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n9269), .A(n7268), .ZN(
        n7269) );
  OAI21_X1 U8915 ( .B1(n7270), .B2(n9309), .A(n7269), .ZN(P1_U3220) );
  INV_X1 U8916 ( .A(n7271), .ZN(n7284) );
  INV_X1 U8917 ( .A(n7781), .ZN(n7682) );
  OAI222_X1 U8918 ( .A1(n8345), .A2(n7272), .B1(n9163), .B2(n7284), .C1(n7682), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8919 ( .A(n7555), .ZN(n7283) );
  AND2_X1 U8920 ( .A1(n7274), .A2(n7273), .ZN(n7277) );
  OAI211_X1 U8921 ( .C1(n7277), .C2(n7276), .A(n9264), .B(n7275), .ZN(n7282)
         );
  INV_X1 U8922 ( .A(n9323), .ZN(n7279) );
  INV_X1 U8923 ( .A(n9298), .ZN(n9234) );
  INV_X1 U8924 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10286) );
  NOR2_X1 U8925 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10286), .ZN(n9723) );
  AOI21_X1 U8926 ( .B1(n9266), .B2(n9321), .A(n9723), .ZN(n7278) );
  OAI21_X1 U8927 ( .B1(n7279), .B2(n9234), .A(n7278), .ZN(n7280) );
  AOI21_X1 U8928 ( .B1(n9291), .B2(n7504), .A(n7280), .ZN(n7281) );
  OAI211_X1 U8929 ( .C1(n9281), .C2(n7283), .A(n7282), .B(n7281), .ZN(P1_U3228) );
  OAI222_X1 U8930 ( .A1(n8540), .A2(n7285), .B1(n8106), .B2(P1_U3084), .C1(
        n9651), .C2(n7284), .ZN(P1_U3337) );
  INV_X1 U8931 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U8932 ( .A1(n9325), .A2(n7457), .ZN(n7287) );
  INV_X1 U8933 ( .A(n7287), .ZN(n7463) );
  OAI21_X1 U8934 ( .B1(n7289), .B2(n7292), .A(n7421), .ZN(n7568) );
  INV_X1 U8935 ( .A(n7568), .ZN(n7304) );
  NAND2_X1 U8936 ( .A1(n6553), .A2(n6483), .ZN(n7290) );
  AND3_X1 U8937 ( .A1(n7302), .A2(n6482), .A3(n7290), .ZN(n7291) );
  NAND2_X1 U8938 ( .A1(n7291), .A2(n7509), .ZN(n9672) );
  INV_X1 U8939 ( .A(n9672), .ZN(n8282) );
  XOR2_X1 U8940 ( .A(n7293), .B(n7292), .Z(n7298) );
  OR2_X1 U8941 ( .A1(n6553), .A2(n6482), .ZN(n7295) );
  OR2_X1 U8942 ( .A1(n6383), .A2(n4794), .ZN(n7294) );
  NAND2_X1 U8943 ( .A1(n7295), .A2(n7294), .ZN(n9542) );
  AOI22_X1 U8944 ( .A1(n9537), .A2(n6564), .B1(n9539), .B2(n9323), .ZN(n7297)
         );
  OAI21_X1 U8945 ( .B1(n7298), .B2(n9484), .A(n7297), .ZN(n7299) );
  AOI21_X1 U8946 ( .B1(n8282), .B2(n7568), .A(n7299), .ZN(n7570) );
  NOR2_X1 U8947 ( .A1(n7456), .A2(n7457), .ZN(n7300) );
  INV_X1 U8948 ( .A(n7300), .ZN(n7459) );
  INV_X1 U8949 ( .A(n7545), .ZN(n7301) );
  AOI21_X1 U8950 ( .B1(n4530), .B2(n7459), .A(n7301), .ZN(n7563) );
  NOR2_X1 U8951 ( .A1(n9881), .A2(n7566), .ZN(n9267) );
  AOI21_X1 U8952 ( .B1(n7563), .B2(n9873), .A(n9267), .ZN(n7303) );
  OAI211_X1 U8953 ( .C1(n7304), .C2(n9876), .A(n7570), .B(n7303), .ZN(n7306)
         );
  NAND2_X1 U8954 ( .A1(n7306), .A2(n9891), .ZN(n7305) );
  OAI21_X1 U8955 ( .B1(n9891), .B2(n10155), .A(n7305), .ZN(P1_U3460) );
  INV_X1 U8956 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7308) );
  NAND2_X1 U8957 ( .A1(n7306), .A2(n9903), .ZN(n7307) );
  OAI21_X1 U8958 ( .B1(n9903), .B2(n7308), .A(n7307), .ZN(P1_U3525) );
  INV_X1 U8959 ( .A(n7309), .ZN(n7342) );
  OAI222_X1 U8960 ( .A1(n8345), .A2(n7310), .B1(n9163), .B2(n7342), .C1(n7791), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8961 ( .A(n9096), .ZN(n9978) );
  OAI21_X1 U8962 ( .B1(n7313), .B2(n7312), .A(n7311), .ZN(n9003) );
  NAND2_X1 U8963 ( .A1(n9958), .A2(n4823), .ZN(n7314) );
  NAND2_X1 U8964 ( .A1(n7314), .A2(n9959), .ZN(n7315) );
  NOR2_X1 U8965 ( .A1(n4507), .A2(n7315), .ZN(n9005) );
  INV_X1 U8966 ( .A(n9003), .ZN(n7321) );
  AOI22_X1 U8967 ( .A1(n8943), .A2(n8705), .B1(n8704), .B2(n8945), .ZN(n7320)
         );
  OAI21_X1 U8968 ( .B1(n7317), .B2(n4516), .A(n7316), .ZN(n7318) );
  NAND2_X1 U8969 ( .A1(n7318), .A2(n8982), .ZN(n7319) );
  OAI211_X1 U8970 ( .C1(n7321), .C2(n8972), .A(n7320), .B(n7319), .ZN(n9000)
         );
  AOI211_X1 U8971 ( .C1(n9978), .C2(n9003), .A(n9005), .B(n9000), .ZN(n7439)
         );
  OAI22_X1 U8972 ( .A1(n9071), .A2(n7436), .B1(n9996), .B2(n5077), .ZN(n7322)
         );
  INV_X1 U8973 ( .A(n7322), .ZN(n7323) );
  OAI21_X1 U8974 ( .B1(n7439), .B2(n9994), .A(n7323), .ZN(P2_U3523) );
  INV_X1 U8975 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7324) );
  AOI21_X1 U8976 ( .B1(n9710), .B2(n7324), .A(n6535), .ZN(n9709) );
  INV_X1 U8977 ( .A(n9709), .ZN(n7330) );
  NOR2_X1 U8978 ( .A1(n6535), .A2(n7325), .ZN(n7328) );
  NOR2_X1 U8979 ( .A1(n7326), .A2(n6535), .ZN(n7327) );
  MUX2_X1 U8980 ( .A(n7328), .B(n7327), .S(n8348), .Z(n7329) );
  AOI211_X1 U8981 ( .C1(n5986), .C2(n7330), .A(n9324), .B(n7329), .ZN(n9722)
         );
  AOI211_X1 U8982 ( .C1(n7333), .C2(n7332), .A(n7331), .B(n9833), .ZN(n7341)
         );
  OAI211_X1 U8983 ( .C1(n7336), .C2(n7335), .A(n9823), .B(n7334), .ZN(n7337)
         );
  OAI21_X1 U8984 ( .B1(n9828), .B2(n7338), .A(n7337), .ZN(n7340) );
  INV_X1 U8985 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7890) );
  INV_X1 U8986 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10271) );
  OAI22_X1 U8987 ( .A1(n9821), .A2(n7890), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10271), .ZN(n7339) );
  OR4_X1 U8988 ( .A1(n9722), .A2(n7341), .A3(n7340), .A4(n7339), .ZN(P1_U3243)
         );
  OAI222_X1 U8989 ( .A1(n8540), .A2(n7343), .B1(n9338), .B2(P1_U3084), .C1(
        n9651), .C2(n7342), .ZN(P1_U3336) );
  INV_X1 U8990 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U8991 ( .A1(n9155), .A2(n7344), .ZN(n7345) );
  OAI21_X1 U8992 ( .B1(n9155), .B2(n7346), .A(n7345), .ZN(P2_U3451) );
  NOR2_X1 U8993 ( .A1(n7493), .A2(n8455), .ZN(n7348) );
  XNOR2_X1 U8994 ( .A(n7451), .B(n8453), .ZN(n7347) );
  NAND2_X1 U8995 ( .A1(n7348), .A2(n7347), .ZN(n7351) );
  INV_X1 U8996 ( .A(n7347), .ZN(n7350) );
  INV_X1 U8997 ( .A(n7348), .ZN(n7349) );
  NAND2_X1 U8998 ( .A1(n7350), .A2(n7349), .ZN(n7375) );
  AND2_X1 U8999 ( .A1(n7351), .A2(n7375), .ZN(n7369) );
  INV_X1 U9000 ( .A(n7352), .ZN(n7355) );
  INV_X1 U9001 ( .A(n7353), .ZN(n7354) );
  NAND2_X1 U9002 ( .A1(n7355), .A2(n7354), .ZN(n7356) );
  XNOR2_X1 U9003 ( .A(n8448), .B(n10344), .ZN(n7361) );
  INV_X1 U9004 ( .A(n7361), .ZN(n7359) );
  AND2_X1 U9005 ( .A1(n8704), .A2(n8432), .ZN(n7360) );
  INV_X1 U9006 ( .A(n7360), .ZN(n7358) );
  AND2_X1 U9007 ( .A1(n7361), .A2(n7360), .ZN(n10336) );
  NOR2_X1 U9008 ( .A1(n10342), .A2(n8455), .ZN(n7362) );
  XNOR2_X1 U9009 ( .A(n8594), .B(n8453), .ZN(n7363) );
  NAND2_X1 U9010 ( .A1(n7362), .A2(n7363), .ZN(n7366) );
  INV_X1 U9011 ( .A(n7362), .ZN(n7365) );
  INV_X1 U9012 ( .A(n7363), .ZN(n7364) );
  NAND2_X1 U9013 ( .A1(n7365), .A2(n7364), .ZN(n7367) );
  AND2_X1 U9014 ( .A1(n7366), .A2(n7367), .ZN(n8596) );
  NAND2_X1 U9015 ( .A1(n7368), .A2(n7369), .ZN(n7376) );
  OAI21_X1 U9016 ( .B1(n7369), .B2(n7368), .A(n7376), .ZN(n7373) );
  AOI22_X1 U9017 ( .A1(n8943), .A2(n8703), .B1(n8701), .B2(n8945), .ZN(n7447)
         );
  OAI22_X1 U9018 ( .A1(n8637), .A2(n7447), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7370), .ZN(n7372) );
  OAI22_X1 U9019 ( .A1(n10345), .A2(n7695), .B1(n10341), .B2(n7691), .ZN(n7371) );
  AOI211_X1 U9020 ( .C1(n8629), .C2(n7373), .A(n7372), .B(n7371), .ZN(n7374)
         );
  INV_X1 U9021 ( .A(n7374), .ZN(P2_U3241) );
  XNOR2_X1 U9022 ( .A(n7632), .B(n8453), .ZN(n7477) );
  NOR2_X1 U9023 ( .A1(n7377), .A2(n8455), .ZN(n7476) );
  XNOR2_X1 U9024 ( .A(n7477), .B(n7476), .ZN(n7479) );
  XNOR2_X1 U9025 ( .A(n7480), .B(n7479), .ZN(n7381) );
  AOI22_X1 U9026 ( .A1(n8675), .A2(n8700), .B1(n7632), .B2(n8668), .ZN(n7380)
         );
  AND2_X1 U9027 ( .A1(n4420), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8738) );
  NOR2_X1 U9028 ( .A1(n10341), .A2(n7629), .ZN(n7378) );
  AOI211_X1 U9029 ( .C1(n10349), .C2(n8702), .A(n8738), .B(n7378), .ZN(n7379)
         );
  OAI211_X1 U9030 ( .C1(n7381), .C2(n10351), .A(n7380), .B(n7379), .ZN(
        P2_U3215) );
  XNOR2_X1 U9031 ( .A(n7382), .B(n7384), .ZN(n7766) );
  INV_X1 U9032 ( .A(n7766), .ZN(n7388) );
  INV_X1 U9033 ( .A(n7450), .ZN(n7383) );
  AOI211_X1 U9034 ( .C1(n8594), .C2(n7601), .A(n9981), .B(n7383), .ZN(n7762)
         );
  OAI211_X1 U9035 ( .C1(n7385), .C2(n7384), .A(n7445), .B(n8982), .ZN(n7387)
         );
  AOI22_X1 U9036 ( .A1(n8702), .A2(n8945), .B1(n8943), .B2(n8704), .ZN(n7386)
         );
  NAND2_X1 U9037 ( .A1(n7387), .A2(n7386), .ZN(n7763) );
  AOI211_X1 U9038 ( .C1(n9985), .C2(n7388), .A(n7762), .B(n7763), .ZN(n7443)
         );
  AOI22_X1 U9039 ( .A1(n9081), .A2(n8594), .B1(n9994), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7389) );
  OAI21_X1 U9040 ( .B1(n7443), .B2(n9994), .A(n7389), .ZN(P2_U3525) );
  INV_X1 U9041 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7397) );
  INV_X1 U9042 ( .A(n7390), .ZN(n7391) );
  OAI21_X1 U9043 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7399), .A(n7391), .ZN(
        n7394) );
  INV_X1 U9044 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7392) );
  MUX2_X1 U9045 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7392), .S(n7923), .Z(n7393)
         );
  NAND2_X1 U9046 ( .A1(n7393), .A2(n7394), .ZN(n7922) );
  OAI21_X1 U9047 ( .B1(n7394), .B2(n7393), .A(n7922), .ZN(n7395) );
  NAND2_X1 U9048 ( .A1(n9816), .A2(n7395), .ZN(n7396) );
  NAND2_X1 U9049 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8137) );
  OAI211_X1 U9050 ( .C1(n9821), .C2(n7397), .A(n7396), .B(n8137), .ZN(n7404)
         );
  INV_X1 U9051 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7400) );
  MUX2_X1 U9052 ( .A(n7400), .B(P1_REG2_REG_13__SCAN_IN), .S(n7923), .Z(n7401)
         );
  AOI211_X1 U9053 ( .C1(n7402), .C2(n7401), .A(n7916), .B(n9782), .ZN(n7403)
         );
  AOI211_X1 U9054 ( .C1(n9808), .C2(n7923), .A(n7404), .B(n7403), .ZN(n7405)
         );
  INV_X1 U9055 ( .A(n7405), .ZN(P1_U3254) );
  INV_X1 U9056 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10152) );
  MUX2_X1 U9057 ( .A(n10152), .B(n7406), .S(n9155), .Z(n7407) );
  OAI21_X1 U9058 ( .B1(n9152), .B2(n7408), .A(n7407), .ZN(P2_U3454) );
  NAND2_X1 U9059 ( .A1(n7410), .A2(n7409), .ZN(n7413) );
  NOR2_X1 U9060 ( .A1(n7413), .A2(n9420), .ZN(n9467) );
  INV_X1 U9061 ( .A(n7414), .ZN(n7415) );
  INV_X1 U9062 ( .A(n9533), .ZN(n9405) );
  OAI21_X1 U9063 ( .B1(n9545), .B2(n9405), .A(n7457), .ZN(n7418) );
  AOI22_X1 U9064 ( .A1(n9477), .A2(n7416), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9530), .ZN(n7417) );
  OAI211_X1 U9065 ( .C1(n9477), .C2(n7324), .A(n7418), .B(n7417), .ZN(P1_U3291) );
  INV_X1 U9066 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7431) );
  OR2_X1 U9067 ( .A1(n6573), .A2(n4530), .ZN(n7420) );
  OR2_X1 U9068 ( .A1(n9323), .A2(n4422), .ZN(n7422) );
  OAI21_X1 U9069 ( .B1(n7423), .B2(n7424), .A(n7506), .ZN(n7560) );
  INV_X1 U9070 ( .A(n7560), .ZN(n7429) );
  XNOR2_X1 U9071 ( .A(n6072), .B(n7424), .ZN(n7426) );
  AOI22_X1 U9072 ( .A1(n9539), .A2(n9321), .B1(n9537), .B2(n9323), .ZN(n7425)
         );
  OAI21_X1 U9073 ( .B1(n7426), .B2(n9484), .A(n7425), .ZN(n7427) );
  AOI21_X1 U9074 ( .B1(n7560), .B2(n8282), .A(n7427), .ZN(n7562) );
  AOI21_X1 U9075 ( .B1(n7504), .B2(n7547), .A(n7513), .ZN(n7554) );
  AOI22_X1 U9076 ( .A1(n7554), .A2(n9873), .B1(n9872), .B2(n7504), .ZN(n7428)
         );
  OAI211_X1 U9077 ( .C1(n7429), .C2(n9876), .A(n7562), .B(n7428), .ZN(n7432)
         );
  NAND2_X1 U9078 ( .A1(n7432), .A2(n9891), .ZN(n7430) );
  OAI21_X1 U9079 ( .B1(n9891), .B2(n7431), .A(n7430), .ZN(P1_U3466) );
  INV_X1 U9080 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U9081 ( .A1(n7432), .A2(n9903), .ZN(n7433) );
  OAI21_X1 U9082 ( .B1(n9903), .B2(n7434), .A(n7433), .ZN(P1_U3527) );
  INV_X1 U9083 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7435) );
  OAI22_X1 U9084 ( .A1(n9152), .A2(n7436), .B1(n9155), .B2(n7435), .ZN(n7437)
         );
  INV_X1 U9085 ( .A(n7437), .ZN(n7438) );
  OAI21_X1 U9086 ( .B1(n7439), .B2(n9987), .A(n7438), .ZN(P2_U3460) );
  OAI22_X1 U9087 ( .A1(n9152), .A2(n7440), .B1(n9155), .B2(n5105), .ZN(n7441)
         );
  INV_X1 U9088 ( .A(n7441), .ZN(n7442) );
  OAI21_X1 U9089 ( .B1(n7443), .B2(n9987), .A(n7442), .ZN(P2_U3466) );
  NAND2_X1 U9090 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  XNOR2_X1 U9091 ( .A(n7446), .B(n7452), .ZN(n7448) );
  OAI21_X1 U9092 ( .B1(n7448), .B2(n8954), .A(n7447), .ZN(n7696) );
  INV_X1 U9093 ( .A(n7488), .ZN(n7449) );
  AOI211_X1 U9094 ( .C1(n7451), .C2(n7450), .A(n9981), .B(n7449), .ZN(n7693)
         );
  NOR2_X1 U9095 ( .A1(n7696), .A2(n7693), .ZN(n7690) );
  XNOR2_X1 U9096 ( .A(n7453), .B(n7452), .ZN(n7699) );
  INV_X1 U9097 ( .A(n9060), .ZN(n9082) );
  OAI22_X1 U9098 ( .A1(n9071), .A2(n7695), .B1(n9996), .B2(n5126), .ZN(n7454)
         );
  AOI21_X1 U9099 ( .B1(n7699), .B2(n9082), .A(n7454), .ZN(n7455) );
  OAI21_X1 U9100 ( .B1(n7690), .B2(n9994), .A(n7455), .ZN(P2_U3526) );
  NAND2_X1 U9101 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  AND3_X1 U9102 ( .A1(n7459), .A2(n9873), .A3(n7458), .ZN(n9845) );
  INV_X1 U9103 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U9104 ( .A1(n9537), .A2(n9325), .ZN(n9843) );
  OAI21_X1 U9105 ( .B1(n9489), .B2(n10169), .A(n9843), .ZN(n7465) );
  INV_X1 U9106 ( .A(n6573), .ZN(n7540) );
  INV_X1 U9107 ( .A(n7286), .ZN(n7462) );
  INV_X1 U9108 ( .A(n7460), .ZN(n7461) );
  AOI21_X1 U9109 ( .B1(n7463), .B2(n7462), .A(n7461), .ZN(n9842) );
  OAI222_X1 U9110 ( .A1(n9380), .A2(n7540), .B1(n9672), .B2(n9842), .C1(n7464), 
        .C2(n9484), .ZN(n9847) );
  AOI211_X1 U9111 ( .C1(n9845), .C2(n6482), .A(n7465), .B(n9847), .ZN(n7472)
         );
  INV_X1 U9112 ( .A(n6545), .ZN(n7467) );
  NAND2_X1 U9113 ( .A1(n7467), .A2(n9420), .ZN(n7468) );
  NOR2_X1 U9114 ( .A1(n4421), .A2(n7468), .ZN(n8298) );
  INV_X1 U9115 ( .A(n9842), .ZN(n7470) );
  OAI22_X1 U9116 ( .A1(n9477), .A2(n7122), .B1(n9533), .B2(n7266), .ZN(n7469)
         );
  AOI21_X1 U9117 ( .B1(n8298), .B2(n7470), .A(n7469), .ZN(n7471) );
  OAI21_X1 U9118 ( .B1(n7472), .B2(n4421), .A(n7471), .ZN(P1_U3290) );
  INV_X1 U9119 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10184) );
  INV_X1 U9120 ( .A(n7473), .ZN(n7474) );
  INV_X1 U9121 ( .A(n8752), .ZN(n8764) );
  OAI222_X1 U9122 ( .A1(n8345), .A2(n10184), .B1(n9163), .B2(n7474), .C1(
        P2_U3152), .C2(n8764), .ZN(P2_U3340) );
  OAI222_X1 U9123 ( .A1(n8540), .A2(n7475), .B1(n9651), .B2(n7474), .C1(
        P1_U3084), .C2(n9829), .ZN(P1_U3335) );
  NAND2_X1 U9124 ( .A1(n7477), .A2(n7476), .ZN(n7478) );
  XNOR2_X1 U9125 ( .A(n7771), .B(n8448), .ZN(n7641) );
  NOR2_X1 U9126 ( .A1(n7646), .A2(n8455), .ZN(n7642) );
  XNOR2_X1 U9127 ( .A(n7641), .B(n7642), .ZN(n7639) );
  XNOR2_X1 U9128 ( .A(n7640), .B(n7639), .ZN(n7486) );
  AOI22_X1 U9129 ( .A1(n8943), .A2(n8701), .B1(n8699), .B2(n8945), .ZN(n7742)
         );
  INV_X1 U9130 ( .A(n7742), .ZN(n7481) );
  AOI22_X1 U9131 ( .A1(n7482), .A2(n7481), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n7485) );
  INV_X1 U9132 ( .A(n7483), .ZN(n7744) );
  AOI22_X1 U9133 ( .A1(n7771), .A2(n8668), .B1(n8674), .B2(n7744), .ZN(n7484)
         );
  OAI211_X1 U9134 ( .C1(n7486), .C2(n10351), .A(n7485), .B(n7484), .ZN(
        P2_U3223) );
  XNOR2_X1 U9135 ( .A(n7487), .B(n5163), .ZN(n7637) );
  INV_X1 U9136 ( .A(n7746), .ZN(n7490) );
  NAND2_X1 U9137 ( .A1(n7488), .A2(n7632), .ZN(n7489) );
  NAND2_X1 U9138 ( .A1(n7490), .A2(n7489), .ZN(n7627) );
  AOI21_X1 U9139 ( .B1(n7492), .B2(n7491), .A(n8954), .ZN(n7496) );
  OAI22_X1 U9140 ( .A1(n7493), .A2(n8977), .B1(n7646), .B2(n8979), .ZN(n7494)
         );
  AOI21_X1 U9141 ( .B1(n7496), .B2(n7495), .A(n7494), .ZN(n7635) );
  OAI21_X1 U9142 ( .B1(n9981), .B2(n7627), .A(n7635), .ZN(n7497) );
  AOI21_X1 U9143 ( .B1(n7637), .B2(n9985), .A(n7497), .ZN(n7501) );
  AOI22_X1 U9144 ( .A1(n9081), .A2(n7632), .B1(n9994), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7498) );
  OAI21_X1 U9145 ( .B1(n7501), .B2(n9994), .A(n7498), .ZN(P2_U3527) );
  NOR2_X1 U9146 ( .A1(n9155), .A2(n5153), .ZN(n7499) );
  AOI21_X1 U9147 ( .B1(n9142), .B2(n7632), .A(n7499), .ZN(n7500) );
  OAI21_X1 U9148 ( .B1(n7501), .B2(n9987), .A(n7500), .ZN(P2_U3472) );
  XNOR2_X1 U9149 ( .A(n7711), .B(n7502), .ZN(n7503) );
  AOI222_X1 U9150 ( .A1(n9542), .A2(n7503), .B1(n9322), .B2(n9537), .C1(n9320), 
        .C2(n9539), .ZN(n9856) );
  OR2_X1 U9151 ( .A1(n9322), .A2(n7504), .ZN(n7505) );
  INV_X1 U9152 ( .A(n7582), .ZN(n7507) );
  AOI21_X1 U9153 ( .B1(n7572), .B2(n7508), .A(n7507), .ZN(n9858) );
  AND2_X1 U9154 ( .A1(n7510), .A2(n7509), .ZN(n7511) );
  INV_X1 U9155 ( .A(n9547), .ZN(n8162) );
  INV_X1 U9156 ( .A(n7575), .ZN(n7512) );
  OAI211_X1 U9157 ( .C1(n7521), .C2(n7513), .A(n7512), .B(n9873), .ZN(n9854)
         );
  INV_X1 U9158 ( .A(n9467), .ZN(n7516) );
  AOI22_X1 U9159 ( .A1(n4421), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7525), .B2(
        n9530), .ZN(n7515) );
  NAND2_X1 U9160 ( .A1(n9405), .A2(n7580), .ZN(n7514) );
  OAI211_X1 U9161 ( .C1(n9854), .C2(n7516), .A(n7515), .B(n7514), .ZN(n7517)
         );
  AOI21_X1 U9162 ( .B1(n9858), .B2(n8162), .A(n7517), .ZN(n7518) );
  OAI21_X1 U9163 ( .B1(n7466), .B2(n9856), .A(n7518), .ZN(P1_U3286) );
  AOI21_X1 U9164 ( .B1(n7520), .B2(n7519), .A(n4510), .ZN(n7527) );
  OR2_X1 U9165 ( .A1(n9881), .A2(n7521), .ZN(n9855) );
  INV_X1 U9166 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U9167 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10171), .ZN(n9738) );
  AOI21_X1 U9168 ( .B1(n9266), .B2(n9320), .A(n9738), .ZN(n7523) );
  NAND2_X1 U9169 ( .A1(n9298), .A2(n9322), .ZN(n7522) );
  OAI211_X1 U9170 ( .C1(n9855), .C2(n9269), .A(n7523), .B(n7522), .ZN(n7524)
         );
  AOI21_X1 U9171 ( .B1(n7525), .B2(n9306), .A(n7524), .ZN(n7526) );
  OAI21_X1 U9172 ( .B1(n7527), .B2(n9309), .A(n7526), .ZN(P1_U3225) );
  XNOR2_X1 U9173 ( .A(n7529), .B(n7528), .ZN(n7530) );
  XNOR2_X1 U9174 ( .A(n7531), .B(n7530), .ZN(n7537) );
  NOR2_X1 U9175 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7532), .ZN(n9751) );
  AOI21_X1 U9176 ( .B1(n9266), .B2(n9319), .A(n9751), .ZN(n7534) );
  NAND2_X1 U9177 ( .A1(n9298), .A2(n9321), .ZN(n7533) );
  OAI211_X1 U9178 ( .C1(n9861), .C2(n9303), .A(n7534), .B(n7533), .ZN(n7535)
         );
  AOI21_X1 U9179 ( .B1(n7576), .B2(n9306), .A(n7535), .ZN(n7536) );
  OAI21_X1 U9180 ( .B1(n7537), .B2(n9309), .A(n7536), .ZN(P1_U3237) );
  XNOR2_X1 U9181 ( .A(n7543), .B(n7538), .ZN(n7539) );
  OAI222_X1 U9182 ( .A1(n9380), .A2(n7541), .B1(n9431), .B2(n7540), .C1(n7539), 
        .C2(n9484), .ZN(n9850) );
  INV_X1 U9183 ( .A(n9850), .ZN(n7553) );
  OAI21_X1 U9184 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n9852) );
  INV_X1 U9185 ( .A(n9545), .ZN(n8296) );
  NAND2_X1 U9186 ( .A1(n7545), .A2(n4422), .ZN(n7546) );
  NAND2_X1 U9187 ( .A1(n7547), .A2(n7546), .ZN(n9849) );
  AOI22_X1 U9188 ( .A1(n7466), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9530), .B2(
        n10165), .ZN(n7550) );
  NAND2_X1 U9189 ( .A1(n9405), .A2(n4422), .ZN(n7549) );
  OAI211_X1 U9190 ( .C1(n8296), .C2(n9849), .A(n7550), .B(n7549), .ZN(n7551)
         );
  AOI21_X1 U9191 ( .B1(n8162), .B2(n9852), .A(n7551), .ZN(n7552) );
  OAI21_X1 U9192 ( .B1(n7553), .B2(n4421), .A(n7552), .ZN(P1_U3288) );
  NAND2_X1 U9193 ( .A1(n7554), .A2(n9545), .ZN(n7557) );
  AOI22_X1 U9194 ( .A1(n4421), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7555), .B2(
        n9530), .ZN(n7556) );
  OAI211_X1 U9195 ( .C1(n7558), .C2(n9533), .A(n7557), .B(n7556), .ZN(n7559)
         );
  AOI21_X1 U9196 ( .B1(n7560), .B2(n8298), .A(n7559), .ZN(n7561) );
  OAI21_X1 U9197 ( .B1(n7562), .B2(n4421), .A(n7561), .ZN(P1_U3287) );
  NAND2_X1 U9198 ( .A1(n9545), .A2(n7563), .ZN(n7565) );
  INV_X1 U9199 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U9200 ( .A1(n4421), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9530), .ZN(n7564) );
  OAI211_X1 U9201 ( .C1(n7566), .C2(n9533), .A(n7565), .B(n7564), .ZN(n7567)
         );
  AOI21_X1 U9202 ( .B1(n8298), .B2(n7568), .A(n7567), .ZN(n7569) );
  OAI21_X1 U9203 ( .B1(n7570), .B2(n4421), .A(n7569), .ZN(P1_U3289) );
  AOI21_X1 U9204 ( .B1(n7711), .B2(n7572), .A(n7571), .ZN(n7573) );
  XNOR2_X1 U9205 ( .A(n7573), .B(n7583), .ZN(n7574) );
  AOI222_X1 U9206 ( .A1(n9542), .A2(n7574), .B1(n9319), .B2(n9539), .C1(n9321), 
        .C2(n9537), .ZN(n9860) );
  OAI211_X1 U9207 ( .C1(n7575), .C2(n9861), .A(n9873), .B(n7724), .ZN(n9859)
         );
  INV_X1 U9208 ( .A(n9859), .ZN(n7579) );
  AOI22_X1 U9209 ( .A1(n4421), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7576), .B2(
        n9530), .ZN(n7577) );
  OAI21_X1 U9210 ( .B1(n9861), .B2(n9533), .A(n7577), .ZN(n7578) );
  AOI21_X1 U9211 ( .B1(n7579), .B2(n9467), .A(n7578), .ZN(n7587) );
  NAND2_X1 U9212 ( .A1(n9321), .A2(n7580), .ZN(n7581) );
  OAI21_X1 U9213 ( .B1(n7585), .B2(n7584), .A(n7721), .ZN(n9863) );
  NAND2_X1 U9214 ( .A1(n9863), .A2(n8162), .ZN(n7586) );
  OAI211_X1 U9215 ( .C1(n9860), .C2(n7466), .A(n7587), .B(n7586), .ZN(P1_U3285) );
  INV_X1 U9216 ( .A(n7588), .ZN(n7590) );
  OAI222_X1 U9217 ( .A1(n8540), .A2(n7589), .B1(n9651), .B2(n7590), .C1(n6482), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U9218 ( .A1(n8345), .A2(n7591), .B1(n9163), .B2(n7590), .C1(
        P2_U3152), .C2(n8929), .ZN(P2_U3339) );
  AOI22_X1 U9219 ( .A1(n9940), .A2(n7592), .B1(n9002), .B2(n5046), .ZN(n7598)
         );
  INV_X1 U9220 ( .A(n8995), .ZN(n9930) );
  OAI21_X1 U9221 ( .B1(n7594), .B2(n8989), .A(n7593), .ZN(n7595) );
  AOI22_X1 U9222 ( .A1(n7596), .A2(n9930), .B1(n9001), .B2(n7595), .ZN(n7597)
         );
  OAI211_X1 U9223 ( .C1(n8710), .C2(n9001), .A(n7598), .B(n7597), .ZN(P2_U3295) );
  OAI21_X1 U9224 ( .B1(n7600), .B2(n7604), .A(n7599), .ZN(n9971) );
  INV_X1 U9225 ( .A(n9001), .ZN(n9944) );
  AND2_X1 U9226 ( .A1(n9944), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7603) );
  OAI211_X1 U9227 ( .C1(n4507), .C2(n10344), .A(n9959), .B(n7601), .ZN(n9968)
         );
  OAI22_X1 U9228 ( .A1(n8995), .A2(n9968), .B1(n10340), .B2(n8989), .ZN(n7602)
         );
  AOI211_X1 U9229 ( .C1(n9940), .C2(n9971), .A(n7603), .B(n7602), .ZN(n7611)
         );
  INV_X1 U9230 ( .A(n7604), .ZN(n7605) );
  XNOR2_X1 U9231 ( .A(n7606), .B(n7605), .ZN(n7607) );
  NAND2_X1 U9232 ( .A1(n7607), .A2(n8982), .ZN(n7609) );
  AOI22_X1 U9233 ( .A1(n8703), .A2(n8945), .B1(n8943), .B2(n10348), .ZN(n7608)
         );
  NAND2_X1 U9234 ( .A1(n7609), .A2(n7608), .ZN(n9969) );
  NAND2_X1 U9235 ( .A1(n9001), .A2(n9969), .ZN(n7610) );
  OAI211_X1 U9236 ( .C1(n10344), .C2(n9937), .A(n7611), .B(n7610), .ZN(
        P2_U3292) );
  OAI21_X1 U9237 ( .B1(n7614), .B2(n7613), .A(n7612), .ZN(n9964) );
  AND2_X1 U9238 ( .A1(n9944), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7621) );
  XNOR2_X1 U9239 ( .A(n7616), .B(n7615), .ZN(n7617) );
  NAND2_X1 U9240 ( .A1(n7617), .A2(n8982), .ZN(n7619) );
  AOI22_X1 U9241 ( .A1(n8943), .A2(n8707), .B1(n10348), .B2(n8945), .ZN(n7618)
         );
  AND2_X1 U9242 ( .A1(n7619), .A2(n7618), .ZN(n9965) );
  OAI22_X1 U9243 ( .A1(n9944), .A2(n9965), .B1(n5049), .B2(n8989), .ZN(n7620)
         );
  AOI211_X1 U9244 ( .C1(n9940), .C2(n9964), .A(n7621), .B(n7620), .ZN(n7626)
         );
  NOR2_X1 U9245 ( .A1(n8995), .A2(n9981), .ZN(n8950) );
  INV_X1 U9246 ( .A(n7622), .ZN(n7624) );
  NAND2_X1 U9247 ( .A1(n7624), .A2(n7623), .ZN(n9960) );
  NAND3_X1 U9248 ( .A1(n8950), .A2(n9958), .A3(n9960), .ZN(n7625) );
  OAI211_X1 U9249 ( .C1(n9962), .C2(n9937), .A(n7626), .B(n7625), .ZN(P2_U3294) );
  INV_X1 U9250 ( .A(n7627), .ZN(n7631) );
  NAND2_X1 U9251 ( .A1(n9944), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7628) );
  OAI21_X1 U9252 ( .B1(n8989), .B2(n7629), .A(n7628), .ZN(n7630) );
  AOI21_X1 U9253 ( .B1(n8950), .B2(n7631), .A(n7630), .ZN(n7634) );
  NAND2_X1 U9254 ( .A1(n9002), .A2(n7632), .ZN(n7633) );
  OAI211_X1 U9255 ( .C1(n7635), .C2(n8998), .A(n7634), .B(n7633), .ZN(n7636)
         );
  AOI21_X1 U9256 ( .B1(n9940), .B2(n7637), .A(n7636), .ZN(n7638) );
  INV_X1 U9257 ( .A(n7638), .ZN(P2_U3289) );
  INV_X1 U9258 ( .A(n7641), .ZN(n7643) );
  NAND2_X1 U9259 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  XNOR2_X1 U9260 ( .A(n9929), .B(n8453), .ZN(n7838) );
  OR2_X1 U9261 ( .A1(n7941), .A2(n8455), .ZN(n7835) );
  XNOR2_X1 U9262 ( .A(n7838), .B(n7835), .ZN(n7645) );
  XNOR2_X1 U9263 ( .A(n7837), .B(n7645), .ZN(n7654) );
  NOR2_X1 U9264 ( .A1(n10341), .A2(n9932), .ZN(n7652) );
  OR2_X1 U9265 ( .A1(n7859), .A2(n8979), .ZN(n7648) );
  OR2_X1 U9266 ( .A1(n7646), .A2(n8977), .ZN(n7647) );
  NAND2_X1 U9267 ( .A1(n7648), .A2(n7647), .ZN(n7809) );
  INV_X1 U9268 ( .A(n7809), .ZN(n7650) );
  OAI22_X1 U9269 ( .A1(n8637), .A2(n7650), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7649), .ZN(n7651) );
  AOI211_X1 U9270 ( .C1(n9929), .C2(n8668), .A(n7652), .B(n7651), .ZN(n7653)
         );
  OAI21_X1 U9271 ( .B1(n7654), .B2(n10351), .A(n7653), .ZN(P2_U3233) );
  NOR2_X1 U9272 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7660), .ZN(n7656) );
  NOR2_X1 U9273 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7657), .ZN(n7680) );
  AOI21_X1 U9274 ( .B1(n7657), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7680), .ZN(
        n7658) );
  NOR2_X1 U9275 ( .A1(n7658), .A2(n9927), .ZN(n7666) );
  OAI21_X1 U9276 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7660), .A(n7659), .ZN(
        n7667) );
  XNOR2_X1 U9277 ( .A(n7667), .B(n7668), .ZN(n7661) );
  NOR2_X1 U9278 ( .A1(n9079), .A2(n7661), .ZN(n7669) );
  AOI211_X1 U9279 ( .C1(n7661), .C2(n9079), .A(n7669), .B(n9906), .ZN(n7665)
         );
  AND2_X1 U9280 ( .A1(n4420), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7662) );
  AOI21_X1 U9281 ( .B1(n9917), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7662), .ZN(
        n7663) );
  OAI21_X1 U9282 ( .B1(n9905), .B2(n7668), .A(n7663), .ZN(n7664) );
  OR3_X1 U9283 ( .A1(n7666), .A2(n7665), .A3(n7664), .ZN(P2_U3260) );
  NOR2_X1 U9284 ( .A1(n7668), .A2(n7667), .ZN(n7670) );
  NOR2_X1 U9285 ( .A1(n7670), .A2(n7669), .ZN(n7673) );
  XNOR2_X1 U9286 ( .A(n7781), .B(n7671), .ZN(n7672) );
  NAND2_X1 U9287 ( .A1(n7672), .A2(n7673), .ZN(n7780) );
  OAI21_X1 U9288 ( .B1(n7673), .B2(n7672), .A(n7780), .ZN(n7677) );
  NAND2_X1 U9289 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(n4420), .ZN(n8465) );
  INV_X1 U9290 ( .A(n8465), .ZN(n7674) );
  AOI21_X1 U9291 ( .B1(n9917), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7674), .ZN(
        n7675) );
  OAI21_X1 U9292 ( .B1(n9905), .B2(n7682), .A(n7675), .ZN(n7676) );
  AOI21_X1 U9293 ( .B1(n7677), .B2(n9922), .A(n7676), .ZN(n7686) );
  NOR2_X1 U9294 ( .A1(n7679), .A2(n7678), .ZN(n7681) );
  AOI22_X1 U9295 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7781), .B1(n7682), .B2(
        n8991), .ZN(n7683) );
  OAI211_X1 U9296 ( .C1(n7684), .C2(n7683), .A(n9904), .B(n7776), .ZN(n7685)
         );
  NAND2_X1 U9297 ( .A1(n7686), .A2(n7685), .ZN(P2_U3261) );
  INV_X1 U9298 ( .A(n9146), .ZN(n8339) );
  INV_X1 U9299 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7687) );
  OAI22_X1 U9300 ( .A1(n9152), .A2(n7695), .B1(n9155), .B2(n7687), .ZN(n7688)
         );
  AOI21_X1 U9301 ( .B1(n7699), .B2(n8339), .A(n7688), .ZN(n7689) );
  OAI21_X1 U9302 ( .B1(n7690), .B2(n9987), .A(n7689), .ZN(P2_U3469) );
  INV_X1 U9303 ( .A(n7691), .ZN(n7692) );
  INV_X1 U9304 ( .A(n8989), .ZN(n9933) );
  AOI22_X1 U9305 ( .A1(n9930), .A2(n7693), .B1(n7692), .B2(n9933), .ZN(n7694)
         );
  OAI21_X1 U9306 ( .B1(n9937), .B2(n7695), .A(n7694), .ZN(n7698) );
  MUX2_X1 U9307 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7696), .S(n9001), .Z(n7697)
         );
  AOI211_X1 U9308 ( .C1(n9940), .C2(n7699), .A(n7698), .B(n7697), .ZN(n7700)
         );
  INV_X1 U9309 ( .A(n7700), .ZN(P2_U3290) );
  XNOR2_X1 U9310 ( .A(n7701), .B(n7702), .ZN(n7708) );
  AND2_X1 U9311 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9755) );
  AOI21_X1 U9312 ( .B1(n9266), .B2(n9318), .A(n9755), .ZN(n7705) );
  NAND2_X1 U9313 ( .A1(n9306), .A2(n7726), .ZN(n7704) );
  NAND2_X1 U9314 ( .A1(n9298), .A2(n9320), .ZN(n7703) );
  AND3_X1 U9315 ( .A1(n7705), .A2(n7704), .A3(n7703), .ZN(n7707) );
  NAND2_X1 U9316 ( .A1(n9291), .A2(n7817), .ZN(n7706) );
  OAI211_X1 U9317 ( .C1(n7708), .C2(n9309), .A(n7707), .B(n7706), .ZN(P1_U3211) );
  INV_X1 U9318 ( .A(n7709), .ZN(n7710) );
  NAND2_X1 U9319 ( .A1(n7711), .A2(n7710), .ZN(n7713) );
  NAND2_X1 U9320 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  NAND2_X1 U9321 ( .A1(n7714), .A2(n7722), .ZN(n7715) );
  NAND2_X1 U9322 ( .A1(n7868), .A2(n7715), .ZN(n7718) );
  NAND2_X1 U9323 ( .A1(n9537), .A2(n9320), .ZN(n7716) );
  OAI21_X1 U9324 ( .B1(n7983), .B2(n9380), .A(n7716), .ZN(n7717) );
  AOI21_X1 U9325 ( .B1(n7718), .B2(n9542), .A(n7717), .ZN(n9866) );
  OR2_X1 U9326 ( .A1(n9320), .A2(n7719), .ZN(n7720) );
  NAND2_X1 U9327 ( .A1(n7721), .A2(n7720), .ZN(n7723) );
  OAI21_X1 U9328 ( .B1(n7723), .B2(n7722), .A(n7819), .ZN(n9869) );
  NAND2_X1 U9329 ( .A1(n9869), .A2(n8162), .ZN(n7731) );
  INV_X1 U9330 ( .A(n7724), .ZN(n7725) );
  OAI211_X1 U9331 ( .C1(n7725), .C2(n9867), .A(n9873), .B(n7878), .ZN(n9865)
         );
  INV_X1 U9332 ( .A(n9865), .ZN(n7729) );
  AOI22_X1 U9333 ( .A1(n4421), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7726), .B2(
        n9530), .ZN(n7727) );
  OAI21_X1 U9334 ( .B1(n9867), .B2(n9533), .A(n7727), .ZN(n7728) );
  AOI21_X1 U9335 ( .B1(n7729), .B2(n9467), .A(n7728), .ZN(n7730) );
  OAI211_X1 U9336 ( .C1(n7466), .C2(n9866), .A(n7731), .B(n7730), .ZN(P1_U3284) );
  INV_X1 U9337 ( .A(n7732), .ZN(n7775) );
  OAI222_X1 U9338 ( .A1(n8345), .A2(n7734), .B1(n9163), .B2(n7775), .C1(n7733), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U9339 ( .A(n7735), .ZN(n7736) );
  AOI21_X1 U9340 ( .B1(n5192), .B2(n7737), .A(n7736), .ZN(n7769) );
  INV_X1 U9341 ( .A(n7769), .ZN(n7753) );
  INV_X1 U9342 ( .A(n7738), .ZN(n7739) );
  AOI21_X1 U9343 ( .B1(n7741), .B2(n7740), .A(n7739), .ZN(n7743) );
  OAI21_X1 U9344 ( .B1(n7743), .B2(n8954), .A(n7742), .ZN(n7767) );
  NAND2_X1 U9345 ( .A1(n9002), .A2(n7771), .ZN(n7750) );
  AOI22_X1 U9346 ( .A1(n8998), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7744), .B2(
        n9933), .ZN(n7749) );
  OR2_X1 U9347 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  AND3_X1 U9348 ( .A1(n7807), .A2(n7747), .A3(n9959), .ZN(n7768) );
  NAND2_X1 U9349 ( .A1(n9930), .A2(n7768), .ZN(n7748) );
  NAND3_X1 U9350 ( .A1(n7750), .A2(n7749), .A3(n7748), .ZN(n7751) );
  AOI21_X1 U9351 ( .B1(n7767), .B2(n9001), .A(n7751), .ZN(n7752) );
  OAI21_X1 U9352 ( .B1(n7753), .B2(n5915), .A(n7752), .ZN(P2_U3288) );
  OAI21_X1 U9353 ( .B1(n8950), .B2(n9002), .A(n7754), .ZN(n7758) );
  AOI21_X1 U9354 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n9933), .A(n7755), .ZN(
        n7756) );
  MUX2_X1 U9355 ( .A(n7756), .B(n6908), .S(n9944), .Z(n7757) );
  OAI211_X1 U9356 ( .C1(n7759), .C2(n5915), .A(n7758), .B(n7757), .ZN(P2_U3296) );
  OAI22_X1 U9357 ( .A1(n9001), .A2(n7760), .B1(n8592), .B2(n8989), .ZN(n7761)
         );
  AOI21_X1 U9358 ( .B1(n9930), .B2(n7762), .A(n7761), .ZN(n7765) );
  AOI22_X1 U9359 ( .A1(n9002), .A2(n8594), .B1(n7763), .B2(n9001), .ZN(n7764)
         );
  OAI211_X1 U9360 ( .C1(n7766), .C2(n5915), .A(n7765), .B(n7764), .ZN(P2_U3291) );
  AOI211_X1 U9361 ( .C1(n7769), .C2(n9985), .A(n7768), .B(n7767), .ZN(n7773)
         );
  AOI22_X1 U9362 ( .A1(n9081), .A2(n7771), .B1(n9994), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n7770) );
  OAI21_X1 U9363 ( .B1(n7773), .B2(n9994), .A(n7770), .ZN(P2_U3528) );
  AOI22_X1 U9364 ( .A1(n9142), .A2(n7771), .B1(n9987), .B2(
        P2_REG0_REG_8__SCAN_IN), .ZN(n7772) );
  OAI21_X1 U9365 ( .B1(n7773), .B2(n9987), .A(n7772), .ZN(P2_U3475) );
  OAI222_X1 U9366 ( .A1(n9651), .A2(n7775), .B1(P1_U3084), .B2(n4794), .C1(
        n7774), .C2(n8540), .ZN(P1_U3333) );
  NAND2_X1 U9367 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7781), .ZN(n7777) );
  AOI22_X1 U9368 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n8754), .B1(n7791), .B2(
        n5375), .ZN(n7778) );
  OAI211_X1 U9369 ( .C1(n7779), .C2(n7778), .A(n9904), .B(n8747), .ZN(n7790)
         );
  XNOR2_X1 U9370 ( .A(n7791), .B(n9069), .ZN(n7783) );
  OAI21_X1 U9371 ( .B1(n7781), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7780), .ZN(
        n7782) );
  NOR2_X1 U9372 ( .A1(n7783), .A2(n7782), .ZN(n8753) );
  AOI21_X1 U9373 ( .B1(n7783), .B2(n7782), .A(n8753), .ZN(n7788) );
  INV_X1 U9374 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7786) );
  OR2_X1 U9375 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7784), .ZN(n7785) );
  OAI21_X1 U9376 ( .B1(n9658), .B2(n7786), .A(n7785), .ZN(n7787) );
  AOI21_X1 U9377 ( .B1(n9922), .B2(n7788), .A(n7787), .ZN(n7789) );
  OAI211_X1 U9378 ( .C1(n9905), .C2(n7791), .A(n7790), .B(n7789), .ZN(P2_U3262) );
  XOR2_X1 U9379 ( .A(n7794), .B(n7793), .Z(n7795) );
  XNOR2_X1 U9380 ( .A(n7792), .B(n7795), .ZN(n7801) );
  NOR2_X1 U9381 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10095), .ZN(n9768) );
  AOI21_X1 U9382 ( .B1(n9266), .B2(n7995), .A(n9768), .ZN(n7798) );
  NAND2_X1 U9383 ( .A1(n9306), .A2(n7879), .ZN(n7797) );
  NAND2_X1 U9384 ( .A1(n9298), .A2(n9319), .ZN(n7796) );
  AND3_X1 U9385 ( .A1(n7798), .A2(n7797), .A3(n7796), .ZN(n7800) );
  NAND2_X1 U9386 ( .A1(n9291), .A2(n9871), .ZN(n7799) );
  OAI211_X1 U9387 ( .C1(n7801), .C2(n9309), .A(n7800), .B(n7799), .ZN(P1_U3219) );
  INV_X1 U9388 ( .A(n7802), .ZN(n7834) );
  OAI222_X1 U9389 ( .A1(P2_U3152), .A2(n7803), .B1(n8345), .B2(n5432), .C1(
        n7834), .C2(n9163), .ZN(P2_U3337) );
  XNOR2_X1 U9390 ( .A(n7805), .B(n4704), .ZN(n9941) );
  INV_X1 U9391 ( .A(n7806), .ZN(n7947) );
  AOI211_X1 U9392 ( .C1(n9929), .C2(n7807), .A(n9981), .B(n7947), .ZN(n9931)
         );
  XNOR2_X1 U9393 ( .A(n7808), .B(n4704), .ZN(n7810) );
  AOI21_X1 U9394 ( .B1(n7810), .B2(n8982), .A(n7809), .ZN(n9943) );
  INV_X1 U9395 ( .A(n9943), .ZN(n7811) );
  AOI211_X1 U9396 ( .C1(n9941), .C2(n9985), .A(n9931), .B(n7811), .ZN(n7816)
         );
  AOI22_X1 U9397 ( .A1(n9081), .A2(n9929), .B1(n9994), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7812) );
  OAI21_X1 U9398 ( .B1(n7816), .B2(n9994), .A(n7812), .ZN(P2_U3529) );
  INV_X1 U9399 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7813) );
  NOR2_X1 U9400 ( .A1(n9155), .A2(n7813), .ZN(n7814) );
  AOI21_X1 U9401 ( .B1(n9142), .B2(n9929), .A(n7814), .ZN(n7815) );
  OAI21_X1 U9402 ( .B1(n7816), .B2(n9987), .A(n7815), .ZN(P2_U3478) );
  OR2_X1 U9403 ( .A1(n9319), .A2(n7817), .ZN(n7864) );
  XOR2_X1 U9404 ( .A(n7822), .B(n7988), .Z(n9888) );
  INV_X1 U9405 ( .A(n9888), .ZN(n7832) );
  NAND2_X1 U9406 ( .A1(n7992), .A2(n7821), .ZN(n7823) );
  XNOR2_X1 U9407 ( .A(n7823), .B(n7822), .ZN(n7824) );
  NAND2_X1 U9408 ( .A1(n7824), .A2(n9542), .ZN(n7826) );
  AOI22_X1 U9409 ( .A1(n9537), .A2(n9318), .B1(n9539), .B2(n8004), .ZN(n7825)
         );
  NAND2_X1 U9410 ( .A1(n7826), .A2(n7825), .ZN(n9886) );
  INV_X1 U9411 ( .A(n7987), .ZN(n9882) );
  INV_X1 U9412 ( .A(n7989), .ZN(n7827) );
  OAI21_X1 U9413 ( .B1(n9882), .B2(n7877), .A(n7827), .ZN(n9884) );
  AOI22_X1 U9414 ( .A1(n7466), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7980), .B2(
        n9530), .ZN(n7829) );
  NAND2_X1 U9415 ( .A1(n9405), .A2(n7987), .ZN(n7828) );
  OAI211_X1 U9416 ( .C1(n9884), .C2(n8296), .A(n7829), .B(n7828), .ZN(n7830)
         );
  AOI21_X1 U9417 ( .B1(n9886), .B2(n9477), .A(n7830), .ZN(n7831) );
  OAI21_X1 U9418 ( .B1(n7832), .B2(n9547), .A(n7831), .ZN(P1_U3282) );
  OAI222_X1 U9419 ( .A1(n9651), .A2(n7834), .B1(P1_U3084), .B2(n6383), .C1(
        n7833), .C2(n8540), .ZN(P1_U3332) );
  NAND2_X1 U9420 ( .A1(n7836), .A2(n7835), .ZN(n7841) );
  XNOR2_X1 U9421 ( .A(n7961), .B(n8453), .ZN(n7842) );
  NOR2_X1 U9422 ( .A1(n7859), .A2(n8455), .ZN(n7843) );
  NAND2_X1 U9423 ( .A1(n7842), .A2(n7843), .ZN(n7853) );
  INV_X1 U9424 ( .A(n7842), .ZN(n7852) );
  INV_X1 U9425 ( .A(n7843), .ZN(n7844) );
  NAND2_X1 U9426 ( .A1(n7852), .A2(n7844), .ZN(n7845) );
  NAND2_X1 U9427 ( .A1(n7853), .A2(n7845), .ZN(n7958) );
  XNOR2_X1 U9428 ( .A(n8043), .B(n8453), .ZN(n7847) );
  NOR2_X1 U9429 ( .A1(n8081), .A2(n8455), .ZN(n7848) );
  NAND2_X1 U9430 ( .A1(n7847), .A2(n7848), .ZN(n8027) );
  INV_X1 U9431 ( .A(n7847), .ZN(n8024) );
  INV_X1 U9432 ( .A(n7848), .ZN(n7849) );
  NAND2_X1 U9433 ( .A1(n8024), .A2(n7849), .ZN(n7850) );
  AND2_X1 U9434 ( .A1(n8027), .A2(n7850), .ZN(n7854) );
  INV_X1 U9435 ( .A(n7854), .ZN(n7851) );
  AOI21_X1 U9436 ( .B1(n7955), .B2(n7851), .A(n10351), .ZN(n7857) );
  NOR3_X1 U9437 ( .A1(n8456), .A2(n7852), .A3(n7859), .ZN(n7856) );
  NAND2_X1 U9438 ( .A1(n7855), .A2(n7854), .ZN(n8029) );
  OAI21_X1 U9439 ( .B1(n7857), .B2(n7856), .A(n8029), .ZN(n7863) );
  OAI22_X1 U9440 ( .A1(n10341), .A2(n8038), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7858), .ZN(n7861) );
  OAI22_X1 U9441 ( .A1(n7859), .A2(n8665), .B1(n10343), .B2(n8237), .ZN(n7860)
         );
  AOI211_X1 U9442 ( .C1(n8043), .C2(n8668), .A(n7861), .B(n7860), .ZN(n7862)
         );
  NAND2_X1 U9443 ( .A1(n7863), .A2(n7862), .ZN(P2_U3238) );
  AND2_X1 U9444 ( .A1(n7819), .A2(n7864), .ZN(n7866) );
  OAI21_X1 U9445 ( .B1(n7866), .B2(n7869), .A(n7865), .ZN(n9877) );
  INV_X1 U9446 ( .A(n8298), .ZN(n7884) );
  OR2_X1 U9447 ( .A1(n9877), .A2(n9672), .ZN(n7876) );
  NAND2_X1 U9448 ( .A1(n7868), .A2(n7867), .ZN(n7871) );
  INV_X1 U9449 ( .A(n7869), .ZN(n7870) );
  XNOR2_X1 U9450 ( .A(n7871), .B(n7870), .ZN(n7874) );
  NAND2_X1 U9451 ( .A1(n9537), .A2(n9319), .ZN(n7872) );
  OAI21_X1 U9452 ( .B1(n8070), .B2(n9380), .A(n7872), .ZN(n7873) );
  AOI21_X1 U9453 ( .B1(n7874), .B2(n9542), .A(n7873), .ZN(n7875) );
  NAND2_X1 U9454 ( .A1(n7876), .A2(n7875), .ZN(n9879) );
  NAND2_X1 U9455 ( .A1(n9879), .A2(n9477), .ZN(n7883) );
  AOI21_X1 U9456 ( .B1(n9871), .B2(n7878), .A(n7877), .ZN(n9874) );
  AOI22_X1 U9457 ( .A1(n4421), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7879), .B2(
        n9530), .ZN(n7880) );
  OAI21_X1 U9458 ( .B1(n4620), .B2(n9533), .A(n7880), .ZN(n7881) );
  AOI21_X1 U9459 ( .B1(n9874), .B2(n9545), .A(n7881), .ZN(n7882) );
  OAI211_X1 U9460 ( .C1(n9877), .C2(n7884), .A(n7883), .B(n7882), .ZN(P1_U3283) );
  INV_X1 U9461 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10361) );
  NOR2_X1 U9462 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n7885) );
  AOI21_X1 U9463 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n7885), .ZN(n10005) );
  NOR2_X1 U9464 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7886) );
  AOI21_X1 U9465 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7886), .ZN(n10008) );
  NOR2_X1 U9466 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7887) );
  AOI21_X1 U9467 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n7887), .ZN(n10011) );
  NOR2_X1 U9468 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7888) );
  AOI21_X1 U9469 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7888), .ZN(n10014) );
  NOR2_X1 U9470 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7889) );
  AOI21_X1 U9471 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7889), .ZN(n10017) );
  NOR2_X1 U9472 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7896) );
  INV_X1 U9473 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9727) );
  XOR2_X1 U9474 ( .A(n9727), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10374) );
  NAND2_X1 U9475 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7894) );
  XOR2_X1 U9476 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10372) );
  NAND2_X1 U9477 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7892) );
  XNOR2_X1 U9478 ( .A(n7890), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n10368) );
  AOI21_X1 U9479 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9997) );
  INV_X1 U9480 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10001) );
  NAND3_X1 U9481 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9999) );
  OAI21_X1 U9482 ( .B1(n9997), .B2(n10001), .A(n9999), .ZN(n10367) );
  NAND2_X1 U9483 ( .A1(n10368), .A2(n10367), .ZN(n7891) );
  NAND2_X1 U9484 ( .A1(n7892), .A2(n7891), .ZN(n10371) );
  NAND2_X1 U9485 ( .A1(n10372), .A2(n10371), .ZN(n7893) );
  NAND2_X1 U9486 ( .A1(n7894), .A2(n7893), .ZN(n10373) );
  NOR2_X1 U9487 ( .A1(n10374), .A2(n10373), .ZN(n7895) );
  NOR2_X1 U9488 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  NOR2_X1 U9489 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7897), .ZN(n10357) );
  AND2_X1 U9490 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7897), .ZN(n10356) );
  NOR2_X1 U9491 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10356), .ZN(n7898) );
  NOR2_X1 U9492 ( .A1(n10357), .A2(n7898), .ZN(n7899) );
  NAND2_X1 U9493 ( .A1(n7899), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7901) );
  XOR2_X1 U9494 ( .A(n7899), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10355) );
  NAND2_X1 U9495 ( .A1(n10355), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U9496 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  NAND2_X1 U9497 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7902), .ZN(n7904) );
  INV_X1 U9498 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9767) );
  XNOR2_X1 U9499 ( .A(n9767), .B(n7902), .ZN(n10370) );
  NAND2_X1 U9500 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10370), .ZN(n7903) );
  NAND2_X1 U9501 ( .A1(n7904), .A2(n7903), .ZN(n7905) );
  NAND2_X1 U9502 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7905), .ZN(n7907) );
  INV_X1 U9503 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9780) );
  XNOR2_X1 U9504 ( .A(n9780), .B(n7905), .ZN(n10369) );
  NAND2_X1 U9505 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10369), .ZN(n7906) );
  NAND2_X1 U9506 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  AND2_X1 U9507 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7908), .ZN(n7909) );
  INV_X1 U9508 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10366) );
  XNOR2_X1 U9509 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7908), .ZN(n10365) );
  NOR2_X1 U9510 ( .A1(n10366), .A2(n10365), .ZN(n10364) );
  NOR2_X1 U9511 ( .A1(n7909), .A2(n10364), .ZN(n10026) );
  NAND2_X1 U9512 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7910) );
  OAI21_X1 U9513 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7910), .ZN(n10025) );
  NOR2_X1 U9514 ( .A1(n10026), .A2(n10025), .ZN(n10024) );
  AOI21_X1 U9515 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10024), .ZN(n10023) );
  NAND2_X1 U9516 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7911) );
  OAI21_X1 U9517 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7911), .ZN(n10022) );
  NOR2_X1 U9518 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  AOI21_X1 U9519 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10021), .ZN(n10020) );
  NOR2_X1 U9520 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7912) );
  AOI21_X1 U9521 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7912), .ZN(n10019) );
  NAND2_X1 U9522 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  OAI21_X1 U9523 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10018), .ZN(n10016) );
  NAND2_X1 U9524 ( .A1(n10017), .A2(n10016), .ZN(n10015) );
  OAI21_X1 U9525 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10015), .ZN(n10013) );
  NAND2_X1 U9526 ( .A1(n10014), .A2(n10013), .ZN(n10012) );
  OAI21_X1 U9527 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10012), .ZN(n10010) );
  NAND2_X1 U9528 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  OAI21_X1 U9529 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10009), .ZN(n10007) );
  NAND2_X1 U9530 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  OAI21_X1 U9531 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10006), .ZN(n10004) );
  NAND2_X1 U9532 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  OAI21_X1 U9533 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10003), .ZN(n10360) );
  NOR2_X1 U9534 ( .A1(n10361), .A2(n10360), .ZN(n7913) );
  NAND2_X1 U9535 ( .A1(n10361), .A2(n10360), .ZN(n10359) );
  OAI21_X1 U9536 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7913), .A(n10359), .ZN(
        n7915) );
  XNOR2_X1 U9537 ( .A(n8376), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7914) );
  XNOR2_X1 U9538 ( .A(n7915), .B(n7914), .ZN(ADD_1071_U4) );
  NAND2_X1 U9539 ( .A1(n7917), .A2(n7921), .ZN(n7918) );
  INV_X1 U9540 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9810) );
  NAND2_X1 U9541 ( .A1(n9811), .A2(n9810), .ZN(n9809) );
  NAND2_X1 U9542 ( .A1(n7918), .A2(n9809), .ZN(n8093) );
  XNOR2_X1 U9543 ( .A(n8093), .B(n8099), .ZN(n7920) );
  INV_X1 U9544 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7919) );
  NOR2_X1 U9545 ( .A1(n7919), .A2(n7920), .ZN(n8094) );
  AOI211_X1 U9546 ( .C1(n7920), .C2(n7919), .A(n8094), .B(n9782), .ZN(n7928)
         );
  INV_X1 U9547 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9689) );
  AOI22_X1 U9548 ( .A1(n9807), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9689), .B2(
        n7921), .ZN(n9814) );
  OAI21_X1 U9549 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7923), .A(n7922), .ZN(
        n9813) );
  NAND2_X1 U9550 ( .A1(n9814), .A2(n9813), .ZN(n9812) );
  OAI21_X1 U9551 ( .B1(n9807), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9812), .ZN(
        n8098) );
  XNOR2_X1 U9552 ( .A(n8098), .B(n8099), .ZN(n7924) );
  INV_X1 U9553 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U9554 ( .A1(n10274), .A2(n7924), .ZN(n8100) );
  AOI211_X1 U9555 ( .C1(n7924), .C2(n10274), .A(n8100), .B(n9833), .ZN(n7927)
         );
  INV_X1 U9556 ( .A(n9821), .ZN(n9837) );
  NAND2_X1 U9557 ( .A1(n9837), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U9558 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9299) );
  OAI211_X1 U9559 ( .C1(n8099), .C2(n9828), .A(n7925), .B(n9299), .ZN(n7926)
         );
  OR3_X1 U9560 ( .A1(n7928), .A2(n7927), .A3(n7926), .ZN(P1_U3256) );
  INV_X1 U9561 ( .A(n7929), .ZN(n7933) );
  AOI21_X1 U9562 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9165), .A(n5793), .ZN(
        n7930) );
  OAI21_X1 U9563 ( .B1(n7933), .B2(n9163), .A(n7930), .ZN(P2_U3335) );
  AOI21_X1 U9564 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9649), .A(n7931), .ZN(
        n7932) );
  OAI21_X1 U9565 ( .B1(n7933), .B2(n9651), .A(n7932), .ZN(P1_U3330) );
  NAND2_X1 U9566 ( .A1(n7936), .A2(n7935), .ZN(n7937) );
  NAND2_X1 U9567 ( .A1(n7934), .A2(n7937), .ZN(n9972) );
  NOR2_X1 U9568 ( .A1(n8998), .A2(n7938), .ZN(n9004) );
  INV_X1 U9569 ( .A(n9004), .ZN(n8249) );
  XNOR2_X1 U9570 ( .A(n7940), .B(n7939), .ZN(n7943) );
  OAI22_X1 U9571 ( .A1(n8081), .A2(n8979), .B1(n7941), .B2(n8977), .ZN(n7942)
         );
  AOI21_X1 U9572 ( .B1(n7943), .B2(n8982), .A(n7942), .ZN(n7944) );
  OAI21_X1 U9573 ( .B1(n9972), .B2(n8972), .A(n7944), .ZN(n9975) );
  NAND2_X1 U9574 ( .A1(n9975), .A2(n9001), .ZN(n7951) );
  OAI22_X1 U9575 ( .A1(n9001), .A2(n7945), .B1(n7954), .B2(n8989), .ZN(n7949)
         );
  INV_X1 U9576 ( .A(n7961), .ZN(n9974) );
  INV_X1 U9577 ( .A(n7969), .ZN(n7946) );
  OAI211_X1 U9578 ( .C1(n9974), .C2(n7947), .A(n7946), .B(n9959), .ZN(n9973)
         );
  NOR2_X1 U9579 ( .A1(n9973), .A2(n8995), .ZN(n7948) );
  AOI211_X1 U9580 ( .C1(n9002), .C2(n7961), .A(n7949), .B(n7948), .ZN(n7950)
         );
  OAI211_X1 U9581 ( .C1(n9972), .C2(n8249), .A(n7951), .B(n7950), .ZN(P2_U3286) );
  AOI22_X1 U9582 ( .A1(n8675), .A2(n8697), .B1(n10349), .B2(n8699), .ZN(n7953)
         );
  OAI211_X1 U9583 ( .C1(n7954), .C2(n10341), .A(n7953), .B(n7952), .ZN(n7960)
         );
  INV_X1 U9584 ( .A(n7955), .ZN(n7956) );
  AOI211_X1 U9585 ( .C1(n7958), .C2(n7957), .A(n10351), .B(n7956), .ZN(n7959)
         );
  AOI211_X1 U9586 ( .C1(n7961), .C2(n8668), .A(n7960), .B(n7959), .ZN(n7962)
         );
  INV_X1 U9587 ( .A(n7962), .ZN(P2_U3219) );
  XNOR2_X1 U9588 ( .A(n7963), .B(n7964), .ZN(n8044) );
  INV_X1 U9589 ( .A(n7964), .ZN(n7966) );
  OAI21_X1 U9590 ( .B1(n7967), .B2(n7966), .A(n7965), .ZN(n7968) );
  AOI222_X1 U9591 ( .A1(n8982), .A2(n7968), .B1(n8696), .B2(n8945), .C1(n8698), 
        .C2(n8943), .ZN(n8048) );
  OAI21_X1 U9592 ( .B1(n7969), .B2(n7973), .A(n9959), .ZN(n7970) );
  OR2_X1 U9593 ( .A1(n8082), .A2(n7970), .ZN(n8040) );
  NAND2_X1 U9594 ( .A1(n8048), .A2(n8040), .ZN(n7975) );
  OAI22_X1 U9595 ( .A1(n9071), .A2(n7973), .B1(n9996), .B2(n6975), .ZN(n7971)
         );
  AOI21_X1 U9596 ( .B1(n7975), .B2(n9996), .A(n7971), .ZN(n7972) );
  OAI21_X1 U9597 ( .B1(n9060), .B2(n8044), .A(n7972), .ZN(P2_U3531) );
  OAI22_X1 U9598 ( .A1(n9152), .A2(n7973), .B1(n9155), .B2(n5236), .ZN(n7974)
         );
  AOI21_X1 U9599 ( .B1(n7975), .B2(n9155), .A(n7974), .ZN(n7976) );
  OAI21_X1 U9600 ( .B1(n9146), .B2(n8044), .A(n7976), .ZN(P2_U3484) );
  INV_X1 U9601 ( .A(n7977), .ZN(n7978) );
  AOI21_X1 U9602 ( .B1(n7979), .B2(n4929), .A(n7978), .ZN(n7986) );
  NAND2_X1 U9603 ( .A1(n9306), .A2(n7980), .ZN(n7982) );
  AND2_X1 U9604 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9786) );
  AOI21_X1 U9605 ( .B1(n9266), .B2(n8004), .A(n9786), .ZN(n7981) );
  OAI211_X1 U9606 ( .C1(n7983), .C2(n9234), .A(n7982), .B(n7981), .ZN(n7984)
         );
  AOI21_X1 U9607 ( .B1(n9291), .B2(n4621), .A(n7984), .ZN(n7985) );
  OAI21_X1 U9608 ( .B1(n7986), .B2(n9309), .A(n7985), .ZN(P1_U3229) );
  XNOR2_X1 U9609 ( .A(n8008), .B(n8009), .ZN(n9673) );
  INV_X1 U9610 ( .A(n8005), .ZN(n9671) );
  NAND2_X1 U9611 ( .A1(n7989), .A2(n9671), .ZN(n8015) );
  OAI211_X1 U9612 ( .C1(n7989), .C2(n9671), .A(n9873), .B(n8015), .ZN(n9669)
         );
  INV_X1 U9613 ( .A(n9669), .ZN(n7999) );
  AOI22_X1 U9614 ( .A1(n4421), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n4966), .B2(
        n9530), .ZN(n7990) );
  OAI21_X1 U9615 ( .B1(n9671), .B2(n9533), .A(n7990), .ZN(n7998) );
  XNOR2_X1 U9616 ( .A(n8010), .B(n8009), .ZN(n7996) );
  AOI222_X1 U9617 ( .A1(n9542), .A2(n7996), .B1(n9317), .B2(n9539), .C1(n7995), 
        .C2(n9537), .ZN(n9670) );
  NOR2_X1 U9618 ( .A1(n9670), .A2(n7466), .ZN(n7997) );
  AOI211_X1 U9619 ( .C1(n7999), .C2(n9467), .A(n7998), .B(n7997), .ZN(n8000)
         );
  OAI21_X1 U9620 ( .B1(n9547), .B2(n9673), .A(n8000), .ZN(P1_U3281) );
  INV_X1 U9621 ( .A(n8001), .ZN(n8022) );
  OAI222_X1 U9622 ( .A1(n9651), .A2(n8022), .B1(P1_U3084), .B2(n8003), .C1(
        n8002), .C2(n8540), .ZN(P1_U3329) );
  NOR2_X1 U9623 ( .A1(n8005), .A2(n8004), .ZN(n8006) );
  XNOR2_X1 U9624 ( .A(n8050), .B(n8013), .ZN(n9701) );
  INV_X1 U9625 ( .A(n9701), .ZN(n8021) );
  XOR2_X1 U9626 ( .A(n8052), .B(n8013), .Z(n8014) );
  OAI222_X1 U9627 ( .A1(n9380), .A2(n8141), .B1(n9431), .B2(n8199), .C1(n9484), 
        .C2(n8014), .ZN(n9700) );
  INV_X1 U9628 ( .A(n8015), .ZN(n8016) );
  INV_X1 U9629 ( .A(n8207), .ZN(n9697) );
  OAI21_X1 U9630 ( .B1(n8016), .B2(n9697), .A(n8058), .ZN(n9698) );
  AOI22_X1 U9631 ( .A1(n4421), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8196), .B2(
        n9530), .ZN(n8018) );
  NAND2_X1 U9632 ( .A1(n9405), .A2(n8207), .ZN(n8017) );
  OAI211_X1 U9633 ( .C1(n9698), .C2(n8296), .A(n8018), .B(n8017), .ZN(n8019)
         );
  AOI21_X1 U9634 ( .B1(n9700), .B2(n9477), .A(n8019), .ZN(n8020) );
  OAI21_X1 U9635 ( .B1(n8021), .B2(n9547), .A(n8020), .ZN(P1_U3280) );
  OAI222_X1 U9636 ( .A1(P2_U3152), .A2(n8023), .B1(n9163), .B2(n8022), .C1(
        n10187), .C2(n8345), .ZN(P2_U3334) );
  INV_X1 U9637 ( .A(n8029), .ZN(n8026) );
  NOR3_X1 U9638 ( .A1(n8456), .A2(n8024), .A3(n8081), .ZN(n8025) );
  AOI21_X1 U9639 ( .B1(n8026), .B2(n8629), .A(n8025), .ZN(n8037) );
  XNOR2_X1 U9640 ( .A(n8087), .B(n8448), .ZN(n8211) );
  NOR2_X1 U9641 ( .A1(n8237), .A2(n8455), .ZN(n8209) );
  XNOR2_X1 U9642 ( .A(n8211), .B(n8209), .ZN(n8036) );
  AND2_X1 U9643 ( .A1(n8036), .A2(n8027), .ZN(n8028) );
  NOR2_X1 U9644 ( .A1(n8213), .A2(n10351), .ZN(n8034) );
  AND2_X1 U9645 ( .A1(n8668), .A2(n8087), .ZN(n8033) );
  OAI21_X1 U9646 ( .B1(n10341), .B2(n8085), .A(n8030), .ZN(n8032) );
  OAI22_X1 U9647 ( .A1(n8269), .A2(n10343), .B1(n8665), .B2(n8081), .ZN(n8031)
         );
  NOR4_X1 U9648 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n8035)
         );
  OAI21_X1 U9649 ( .B1(n8037), .B2(n8036), .A(n8035), .ZN(P2_U3226) );
  OAI22_X1 U9650 ( .A1(n9001), .A2(n8039), .B1(n8038), .B2(n8989), .ZN(n8042)
         );
  NOR2_X1 U9651 ( .A1(n8040), .A2(n8995), .ZN(n8041) );
  AOI211_X1 U9652 ( .C1(n9002), .C2(n8043), .A(n8042), .B(n8041), .ZN(n8047)
         );
  INV_X1 U9653 ( .A(n8044), .ZN(n8045) );
  NAND2_X1 U9654 ( .A1(n8045), .A2(n9940), .ZN(n8046) );
  OAI211_X1 U9655 ( .C1(n8048), .C2(n8998), .A(n8047), .B(n8046), .ZN(P2_U3285) );
  OR2_X1 U9656 ( .A1(n8207), .A2(n9317), .ZN(n8049) );
  NAND2_X1 U9657 ( .A1(n8207), .A2(n9317), .ZN(n8051) );
  XNOR2_X1 U9658 ( .A(n8169), .B(n8168), .ZN(n8128) );
  NAND2_X1 U9659 ( .A1(n8148), .A2(n8054), .ZN(n8056) );
  XNOR2_X1 U9660 ( .A(n8056), .B(n8055), .ZN(n8057) );
  OAI222_X1 U9661 ( .A1(n9431), .A2(n8119), .B1(n9380), .B2(n9177), .C1(n9484), 
        .C2(n8057), .ZN(n8125) );
  INV_X1 U9662 ( .A(n8158), .ZN(n8124) );
  AOI211_X1 U9663 ( .C1(n8158), .C2(n8058), .A(n9883), .B(n8179), .ZN(n8126)
         );
  NAND2_X1 U9664 ( .A1(n8126), .A2(n9467), .ZN(n8060) );
  AOI22_X1 U9665 ( .A1(n4421), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8121), .B2(
        n9530), .ZN(n8059) );
  OAI211_X1 U9666 ( .C1(n8124), .C2(n9533), .A(n8060), .B(n8059), .ZN(n8061)
         );
  AOI21_X1 U9667 ( .B1(n8125), .B2(n9477), .A(n8061), .ZN(n8062) );
  OAI21_X1 U9668 ( .B1(n8128), .B2(n9547), .A(n8062), .ZN(P1_U3279) );
  OAI21_X1 U9669 ( .B1(n8065), .B2(n8064), .A(n8063), .ZN(n8073) );
  NOR2_X1 U9670 ( .A1(n9671), .A2(n9303), .ZN(n8072) );
  INV_X1 U9671 ( .A(n8066), .ZN(n8067) );
  AOI21_X1 U9672 ( .B1(n9266), .B2(n9317), .A(n8067), .ZN(n8069) );
  NAND2_X1 U9673 ( .A1(n9306), .A2(n4966), .ZN(n8068) );
  OAI211_X1 U9674 ( .C1(n8070), .C2(n9234), .A(n8069), .B(n8068), .ZN(n8071)
         );
  AOI211_X1 U9675 ( .C1(n8073), .C2(n9264), .A(n8072), .B(n8071), .ZN(n8074)
         );
  INV_X1 U9676 ( .A(n8074), .ZN(P1_U3215) );
  XNOR2_X1 U9677 ( .A(n8076), .B(n8075), .ZN(n9986) );
  INV_X1 U9678 ( .A(n9986), .ZN(n8092) );
  NAND2_X1 U9679 ( .A1(n7965), .A2(n8077), .ZN(n8079) );
  XNOR2_X1 U9680 ( .A(n8079), .B(n8078), .ZN(n8080) );
  OAI222_X1 U9681 ( .A1(n8977), .A2(n8081), .B1(n8979), .B2(n8269), .C1(n8080), 
        .C2(n8954), .ZN(n9983) );
  OR2_X1 U9682 ( .A1(n8082), .A2(n9980), .ZN(n8083) );
  NAND2_X1 U9683 ( .A1(n8241), .A2(n8083), .ZN(n9982) );
  INV_X1 U9684 ( .A(n8950), .ZN(n8089) );
  NAND2_X1 U9685 ( .A1(n9944), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8084) );
  OAI21_X1 U9686 ( .B1(n8989), .B2(n8085), .A(n8084), .ZN(n8086) );
  AOI21_X1 U9687 ( .B1(n9002), .B2(n8087), .A(n8086), .ZN(n8088) );
  OAI21_X1 U9688 ( .B1(n9982), .B2(n8089), .A(n8088), .ZN(n8090) );
  AOI21_X1 U9689 ( .B1(n9983), .B2(n9001), .A(n8090), .ZN(n8091) );
  OAI21_X1 U9690 ( .B1(n5915), .B2(n8092), .A(n8091), .ZN(P2_U3284) );
  NOR2_X1 U9691 ( .A1(n8099), .A2(n8093), .ZN(n8095) );
  NAND2_X1 U9692 ( .A1(n8352), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8365) );
  OAI21_X1 U9693 ( .B1(n8352), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8365), .ZN(
        n8096) );
  AOI211_X1 U9694 ( .C1(n8097), .C2(n8096), .A(n8364), .B(n9782), .ZN(n8109)
         );
  NOR2_X1 U9695 ( .A1(n8099), .A2(n8098), .ZN(n8101) );
  NOR2_X1 U9696 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  XNOR2_X1 U9697 ( .A(n8352), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8102) );
  NOR2_X1 U9698 ( .A1(n8103), .A2(n8102), .ZN(n8353) );
  AOI211_X1 U9699 ( .C1(n8103), .C2(n8102), .A(n8353), .B(n9833), .ZN(n8108)
         );
  NAND2_X1 U9700 ( .A1(n9837), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U9701 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n8104) );
  OAI211_X1 U9702 ( .C1(n9828), .C2(n8106), .A(n8105), .B(n8104), .ZN(n8107)
         );
  OR3_X1 U9703 ( .A1(n8109), .A2(n8108), .A3(n8107), .ZN(P1_U3257) );
  INV_X1 U9704 ( .A(n8110), .ZN(n8115) );
  AOI21_X1 U9705 ( .B1(n8200), .B2(n8113), .A(n8112), .ZN(n8114) );
  OAI21_X1 U9706 ( .B1(n8115), .B2(n8114), .A(n9264), .ZN(n8123) );
  INV_X1 U9707 ( .A(n8116), .ZN(n8117) );
  AOI21_X1 U9708 ( .B1(n9266), .B2(n9315), .A(n8117), .ZN(n8118) );
  OAI21_X1 U9709 ( .B1(n8119), .B2(n9234), .A(n8118), .ZN(n8120) );
  AOI21_X1 U9710 ( .B1(n8121), .B2(n9306), .A(n8120), .ZN(n8122) );
  OAI211_X1 U9711 ( .C1(n8124), .C2(n9303), .A(n8123), .B(n8122), .ZN(P1_U3222) );
  AOI211_X1 U9712 ( .C1(n9872), .C2(n8158), .A(n8126), .B(n8125), .ZN(n8127)
         );
  OAI21_X1 U9713 ( .B1(n8128), .B2(n9683), .A(n8127), .ZN(n8130) );
  NAND2_X1 U9714 ( .A1(n8130), .A2(n9903), .ZN(n8129) );
  OAI21_X1 U9715 ( .B1(n9903), .B2(n10241), .A(n8129), .ZN(P1_U3535) );
  INV_X1 U9716 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U9717 ( .A1(n8130), .A2(n9891), .ZN(n8131) );
  OAI21_X1 U9718 ( .B1(n9891), .B2(n10321), .A(n8131), .ZN(P1_U3490) );
  INV_X1 U9719 ( .A(n8133), .ZN(n8135) );
  NAND2_X1 U9720 ( .A1(n8135), .A2(n8134), .ZN(n8136) );
  XNOR2_X1 U9721 ( .A(n8132), .B(n8136), .ZN(n8144) );
  INV_X1 U9722 ( .A(n8137), .ZN(n8138) );
  AOI21_X1 U9723 ( .B1(n9266), .B2(n9314), .A(n8138), .ZN(n8140) );
  NAND2_X1 U9724 ( .A1(n9306), .A2(n8182), .ZN(n8139) );
  OAI211_X1 U9725 ( .C1(n8141), .C2(n9234), .A(n8140), .B(n8139), .ZN(n8142)
         );
  AOI21_X1 U9726 ( .B1(n8183), .B2(n9291), .A(n8142), .ZN(n8143) );
  OAI21_X1 U9727 ( .B1(n8144), .B2(n9309), .A(n8143), .ZN(P1_U3232) );
  INV_X1 U9728 ( .A(n8145), .ZN(n8195) );
  AOI22_X1 U9729 ( .A1(n9952), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9165), .ZN(n8146) );
  OAI21_X1 U9730 ( .B1(n8195), .B2(n9163), .A(n8146), .ZN(P2_U3332) );
  AOI21_X1 U9731 ( .B1(n8152), .B2(n8280), .A(n9484), .ZN(n8156) );
  INV_X1 U9732 ( .A(n8280), .ZN(n8153) );
  NAND2_X1 U9733 ( .A1(n9539), .A2(n9313), .ZN(n8154) );
  OAI21_X1 U9734 ( .B1(n9177), .B2(n9431), .A(n8154), .ZN(n8155) );
  AOI21_X1 U9735 ( .B1(n8156), .B2(n8284), .A(n8155), .ZN(n9685) );
  OR2_X1 U9736 ( .A1(n8183), .A2(n9315), .ZN(n8157) );
  AND2_X1 U9737 ( .A1(n8168), .A2(n8157), .ZN(n8161) );
  INV_X1 U9738 ( .A(n8157), .ZN(n8160) );
  NAND2_X1 U9739 ( .A1(n8158), .A2(n9316), .ZN(n8170) );
  AND2_X1 U9740 ( .A1(n4977), .A2(n8170), .ZN(n8159) );
  XNOR2_X1 U9741 ( .A(n8281), .B(n8280), .ZN(n9688) );
  NAND2_X1 U9742 ( .A1(n9688), .A2(n8162), .ZN(n8167) );
  INV_X1 U9743 ( .A(n8183), .ZN(n9690) );
  INV_X1 U9744 ( .A(n9179), .ZN(n9686) );
  OAI211_X1 U9745 ( .C1(n8181), .C2(n9686), .A(n9873), .B(n4509), .ZN(n9684)
         );
  INV_X1 U9746 ( .A(n9684), .ZN(n8165) );
  AOI22_X1 U9747 ( .A1(n4421), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9174), .B2(
        n9530), .ZN(n8163) );
  OAI21_X1 U9748 ( .B1(n9686), .B2(n9533), .A(n8163), .ZN(n8164) );
  AOI21_X1 U9749 ( .B1(n8165), .B2(n9467), .A(n8164), .ZN(n8166) );
  OAI211_X1 U9750 ( .C1(n7466), .C2(n9685), .A(n8167), .B(n8166), .ZN(P1_U3277) );
  NAND2_X1 U9751 ( .A1(n8169), .A2(n8168), .ZN(n8171) );
  NAND2_X1 U9752 ( .A1(n8171), .A2(n8170), .ZN(n8173) );
  XNOR2_X1 U9753 ( .A(n8173), .B(n8172), .ZN(n9694) );
  XNOR2_X1 U9754 ( .A(n8175), .B(n8174), .ZN(n8177) );
  AOI22_X1 U9755 ( .A1(n9539), .A2(n9314), .B1(n9537), .B2(n9316), .ZN(n8176)
         );
  OAI21_X1 U9756 ( .B1(n8177), .B2(n9484), .A(n8176), .ZN(n8178) );
  AOI21_X1 U9757 ( .B1(n9694), .B2(n8282), .A(n8178), .ZN(n9696) );
  NOR2_X1 U9758 ( .A1(n8179), .A2(n9690), .ZN(n8180) );
  OR2_X1 U9759 ( .A1(n8181), .A2(n8180), .ZN(n9691) );
  AOI22_X1 U9760 ( .A1(n4421), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8182), .B2(
        n9530), .ZN(n8185) );
  NAND2_X1 U9761 ( .A1(n8183), .A2(n9405), .ZN(n8184) );
  OAI211_X1 U9762 ( .C1(n9691), .C2(n8296), .A(n8185), .B(n8184), .ZN(n8186)
         );
  AOI21_X1 U9763 ( .B1(n9694), .B2(n8298), .A(n8186), .ZN(n8187) );
  OAI21_X1 U9764 ( .B1(n9696), .B2(n4421), .A(n8187), .ZN(P1_U3278) );
  INV_X1 U9765 ( .A(n8188), .ZN(n8191) );
  OAI222_X1 U9766 ( .A1(n8345), .A2(n10218), .B1(n9163), .B2(n8191), .C1(
        P2_U3152), .C2(n8189), .ZN(P2_U3333) );
  OAI222_X1 U9767 ( .A1(n8540), .A2(n8192), .B1(n9651), .B2(n8191), .C1(n8190), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9768 ( .A1(n9651), .A2(n8195), .B1(P1_U3084), .B2(n8194), .C1(
        n8193), .C2(n8540), .ZN(P1_U3327) );
  AND2_X1 U9769 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9794) );
  AOI21_X1 U9770 ( .B1(n9266), .B2(n9316), .A(n9794), .ZN(n8198) );
  NAND2_X1 U9771 ( .A1(n9306), .A2(n8196), .ZN(n8197) );
  OAI211_X1 U9772 ( .C1(n8199), .C2(n9234), .A(n8198), .B(n8197), .ZN(n8206)
         );
  INV_X1 U9773 ( .A(n8200), .ZN(n8204) );
  AOI21_X1 U9774 ( .B1(n8063), .B2(n8202), .A(n8201), .ZN(n8203) );
  NOR3_X1 U9775 ( .A1(n8204), .A2(n8203), .A3(n9309), .ZN(n8205) );
  AOI211_X1 U9776 ( .C1(n9291), .C2(n8207), .A(n8206), .B(n8205), .ZN(n8208)
         );
  INV_X1 U9777 ( .A(n8208), .ZN(P1_U3234) );
  INV_X1 U9778 ( .A(n8209), .ZN(n8210) );
  NAND2_X1 U9779 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  XNOR2_X1 U9780 ( .A(n9092), .B(n8453), .ZN(n8214) );
  NOR2_X1 U9781 ( .A1(n8269), .A2(n8455), .ZN(n8215) );
  NAND2_X1 U9782 ( .A1(n8214), .A2(n8215), .ZN(n8220) );
  INV_X1 U9783 ( .A(n8214), .ZN(n8218) );
  INV_X1 U9784 ( .A(n8215), .ZN(n8216) );
  NAND2_X1 U9785 ( .A1(n8218), .A2(n8216), .ZN(n8217) );
  NAND2_X1 U9786 ( .A1(n8220), .A2(n8217), .ZN(n8253) );
  INV_X1 U9787 ( .A(n8222), .ZN(n8252) );
  NOR3_X1 U9788 ( .A1(n8218), .A2(n8456), .A3(n8269), .ZN(n8219) );
  AOI21_X1 U9789 ( .B1(n8252), .B2(n8629), .A(n8219), .ZN(n8230) );
  XNOR2_X1 U9790 ( .A(n9087), .B(n8448), .ZN(n8389) );
  NOR2_X1 U9791 ( .A1(n8322), .A2(n8455), .ZN(n8387) );
  XNOR2_X1 U9792 ( .A(n8389), .B(n8387), .ZN(n8229) );
  AND2_X1 U9793 ( .A1(n8229), .A2(n8220), .ZN(n8221) );
  NOR2_X1 U9794 ( .A1(n8391), .A2(n10351), .ZN(n8227) );
  AND2_X1 U9795 ( .A1(n9087), .A2(n8668), .ZN(n8226) );
  OAI21_X1 U9796 ( .B1(n10341), .B2(n8261), .A(n8223), .ZN(n8225) );
  OAI22_X1 U9797 ( .A1(n8978), .A2(n10343), .B1(n8665), .B2(n8269), .ZN(n8224)
         );
  NOR4_X1 U9798 ( .A1(n8227), .A2(n8226), .A3(n8225), .A4(n8224), .ZN(n8228)
         );
  OAI21_X1 U9799 ( .B1(n8230), .B2(n8229), .A(n8228), .ZN(P2_U3217) );
  NAND2_X1 U9800 ( .A1(n8231), .A2(n5294), .ZN(n8232) );
  NAND2_X1 U9801 ( .A1(n8233), .A2(n8232), .ZN(n9097) );
  NAND2_X1 U9802 ( .A1(n8234), .A2(n8235), .ZN(n8236) );
  NAND2_X1 U9803 ( .A1(n8267), .A2(n8236), .ZN(n8239) );
  OAI22_X1 U9804 ( .A1(n8322), .A2(n8979), .B1(n8237), .B2(n8977), .ZN(n8238)
         );
  AOI21_X1 U9805 ( .B1(n8239), .B2(n8982), .A(n8238), .ZN(n8240) );
  OAI21_X1 U9806 ( .B1(n9097), .B2(n8972), .A(n8240), .ZN(n9099) );
  NAND2_X1 U9807 ( .A1(n9099), .A2(n9001), .ZN(n8248) );
  NAND2_X1 U9808 ( .A1(n8241), .A2(n9092), .ZN(n8242) );
  AND2_X1 U9809 ( .A1(n8260), .A2(n8242), .ZN(n9094) );
  OAI22_X1 U9810 ( .A1(n9001), .A2(n8243), .B1(n8251), .B2(n8989), .ZN(n8246)
         );
  INV_X1 U9811 ( .A(n9092), .ZN(n8244) );
  NOR2_X1 U9812 ( .A1(n9937), .A2(n8244), .ZN(n8245) );
  AOI211_X1 U9813 ( .C1(n9094), .C2(n8950), .A(n8246), .B(n8245), .ZN(n8247)
         );
  OAI211_X1 U9814 ( .C1(n9097), .C2(n8249), .A(n8248), .B(n8247), .ZN(P2_U3283) );
  AOI22_X1 U9815 ( .A1(n8675), .A2(n8694), .B1(n10349), .B2(n8696), .ZN(n8250)
         );
  NAND2_X1 U9816 ( .A1(n4420), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9915) );
  OAI211_X1 U9817 ( .C1(n10341), .C2(n8251), .A(n8250), .B(n9915), .ZN(n8256)
         );
  AOI211_X1 U9818 ( .C1(n8254), .C2(n8253), .A(n10351), .B(n8252), .ZN(n8255)
         );
  AOI211_X1 U9819 ( .C1(n9092), .C2(n8668), .A(n8256), .B(n8255), .ZN(n8257)
         );
  INV_X1 U9820 ( .A(n8257), .ZN(P2_U3236) );
  XNOR2_X1 U9821 ( .A(n8259), .B(n8258), .ZN(n9091) );
  AOI211_X1 U9822 ( .C1(n9087), .C2(n8260), .A(n9981), .B(n8323), .ZN(n9086)
         );
  INV_X1 U9823 ( .A(n9087), .ZN(n8264) );
  INV_X1 U9824 ( .A(n8261), .ZN(n8262) );
  AOI22_X1 U9825 ( .A1(n9944), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8262), .B2(
        n9933), .ZN(n8263) );
  OAI21_X1 U9826 ( .B1(n9937), .B2(n8264), .A(n8263), .ZN(n8274) );
  AOI21_X1 U9827 ( .B1(n8267), .B2(n8266), .A(n8265), .ZN(n8268) );
  NOR2_X1 U9828 ( .A1(n8268), .A2(n8954), .ZN(n8272) );
  OAI22_X1 U9829 ( .A1(n8978), .A2(n8979), .B1(n8269), .B2(n8977), .ZN(n8270)
         );
  AOI21_X1 U9830 ( .B1(n8272), .B2(n8271), .A(n8270), .ZN(n9089) );
  NOR2_X1 U9831 ( .A1(n9089), .A2(n8998), .ZN(n8273) );
  AOI211_X1 U9832 ( .C1(n9086), .C2(n9930), .A(n8274), .B(n8273), .ZN(n8275)
         );
  OAI21_X1 U9833 ( .B1(n5915), .B2(n9091), .A(n8275), .ZN(P2_U3282) );
  INV_X1 U9834 ( .A(n8276), .ZN(n8336) );
  AOI22_X1 U9835 ( .A1(n8277), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9165), .ZN(n8278) );
  OAI21_X1 U9836 ( .B1(n8336), .B2(n9163), .A(n8278), .ZN(P2_U3331) );
  NOR2_X1 U9837 ( .A1(n9179), .A2(n9314), .ZN(n8279) );
  XNOR2_X1 U9838 ( .A(n8302), .B(n8285), .ZN(n9620) );
  NAND2_X1 U9839 ( .A1(n9620), .A2(n8282), .ZN(n8292) );
  NAND2_X1 U9840 ( .A1(n8284), .A2(n8283), .ZN(n8307) );
  INV_X1 U9841 ( .A(n8285), .ZN(n8286) );
  XNOR2_X1 U9842 ( .A(n8307), .B(n8286), .ZN(n8290) );
  NAND2_X1 U9843 ( .A1(n9539), .A2(n9538), .ZN(n8287) );
  OAI21_X1 U9844 ( .B1(n8288), .B2(n9431), .A(n8287), .ZN(n8289) );
  AOI21_X1 U9845 ( .B1(n8290), .B2(n9542), .A(n8289), .ZN(n8291) );
  NAND2_X1 U9846 ( .A1(n8292), .A2(n8291), .ZN(n9625) );
  INV_X1 U9847 ( .A(n9625), .ZN(n8300) );
  NAND2_X1 U9848 ( .A1(n4509), .A2(n8303), .ZN(n8293) );
  NAND2_X1 U9849 ( .A1(n4447), .A2(n8293), .ZN(n9622) );
  AOI22_X1 U9850 ( .A1(n4421), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9307), .B2(
        n9530), .ZN(n8295) );
  NAND2_X1 U9851 ( .A1(n8303), .A2(n9405), .ZN(n8294) );
  OAI211_X1 U9852 ( .C1(n9622), .C2(n8296), .A(n8295), .B(n8294), .ZN(n8297)
         );
  AOI21_X1 U9853 ( .B1(n9620), .B2(n8298), .A(n8297), .ZN(n8299) );
  OAI21_X1 U9854 ( .B1(n8300), .B2(n4421), .A(n8299), .ZN(P1_U3276) );
  NAND2_X1 U9855 ( .A1(n8302), .A2(n8301), .ZN(n8304) );
  INV_X1 U9856 ( .A(n8303), .ZN(n9621) );
  NAND2_X1 U9857 ( .A1(n8304), .A2(n4970), .ZN(n8484) );
  XNOR2_X1 U9858 ( .A(n8484), .B(n8500), .ZN(n9619) );
  XNOR2_X1 U9859 ( .A(n8502), .B(n8500), .ZN(n8308) );
  OAI222_X1 U9860 ( .A1(n9380), .A2(n9216), .B1(n9431), .B2(n8309), .C1(n8308), 
        .C2(n9484), .ZN(n9615) );
  INV_X1 U9861 ( .A(n9617), .ZN(n8313) );
  INV_X1 U9862 ( .A(n9529), .ZN(n8310) );
  AOI211_X1 U9863 ( .C1(n9617), .C2(n4447), .A(n9883), .B(n8310), .ZN(n9616)
         );
  NAND2_X1 U9864 ( .A1(n9616), .A2(n9467), .ZN(n8312) );
  AOI22_X1 U9865 ( .A1(n4421), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9213), .B2(
        n9530), .ZN(n8311) );
  OAI211_X1 U9866 ( .C1(n8313), .C2(n9533), .A(n8312), .B(n8311), .ZN(n8314)
         );
  AOI21_X1 U9867 ( .B1(n9615), .B2(n9477), .A(n8314), .ZN(n8315) );
  OAI21_X1 U9868 ( .B1(n9619), .B2(n9547), .A(n8315), .ZN(P1_U3275) );
  OAI21_X1 U9869 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(n9083) );
  INV_X1 U9870 ( .A(n9083), .ZN(n8329) );
  XNOR2_X1 U9871 ( .A(n8320), .B(n8319), .ZN(n8321) );
  OAI222_X1 U9872 ( .A1(n8979), .A2(n8956), .B1(n8977), .B2(n8322), .C1(n8954), 
        .C2(n8321), .ZN(n8338) );
  AOI211_X1 U9873 ( .C1(n9080), .C2(n4614), .A(n9981), .B(n8988), .ZN(n8337)
         );
  NAND2_X1 U9874 ( .A1(n8337), .A2(n9930), .ZN(n8326) );
  INV_X1 U9875 ( .A(n8324), .ZN(n8673) );
  AOI22_X1 U9876 ( .A1(n9944), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8673), .B2(
        n9933), .ZN(n8325) );
  OAI211_X1 U9877 ( .C1(n8678), .C2(n9937), .A(n8326), .B(n8325), .ZN(n8327)
         );
  AOI21_X1 U9878 ( .B1(n8338), .B2(n9001), .A(n8327), .ZN(n8328) );
  OAI21_X1 U9879 ( .B1(n8329), .B2(n5915), .A(n8328), .ZN(P2_U3281) );
  INV_X1 U9880 ( .A(n8330), .ZN(n8334) );
  AOI21_X1 U9881 ( .B1(n9165), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8331), .ZN(
        n8332) );
  OAI21_X1 U9882 ( .B1(n8334), .B2(n9163), .A(n8332), .ZN(P2_U3330) );
  AOI22_X1 U9883 ( .A1(n4727), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9649), .ZN(n8333) );
  OAI21_X1 U9884 ( .B1(n8334), .B2(n9651), .A(n8333), .ZN(P1_U3325) );
  OAI222_X1 U9885 ( .A1(n9651), .A2(n8336), .B1(P1_U3084), .B2(n8348), .C1(
        n8335), .C2(n8540), .ZN(P1_U3326) );
  NOR2_X1 U9886 ( .A1(n8338), .A2(n8337), .ZN(n9078) );
  MUX2_X1 U9887 ( .A(n10314), .B(n9078), .S(n9155), .Z(n8341) );
  AOI22_X1 U9888 ( .A1(n9083), .A2(n8339), .B1(n9142), .B2(n9080), .ZN(n8340)
         );
  NAND2_X1 U9889 ( .A1(n8341), .A2(n8340), .ZN(P2_U3496) );
  INV_X1 U9890 ( .A(n8342), .ZN(n8538) );
  OAI222_X1 U9891 ( .A1(n8345), .A2(n8344), .B1(n9163), .B2(n8538), .C1(
        P2_U3152), .C2(n8343), .ZN(P2_U3336) );
  INV_X1 U9892 ( .A(n9605), .ZN(n9516) );
  NAND2_X1 U9893 ( .A1(n9528), .A2(n9516), .ZN(n9510) );
  INV_X1 U9894 ( .A(n9592), .ZN(n9471) );
  INV_X1 U9895 ( .A(n9586), .ZN(n9448) );
  INV_X1 U9896 ( .A(n9561), .ZN(n9360) );
  NAND2_X1 U9897 ( .A1(n9340), .A2(n9679), .ZN(n8346) );
  XNOR2_X1 U9898 ( .A(n9550), .B(n8346), .ZN(n9548) );
  NAND2_X1 U9899 ( .A1(n9548), .A2(n9545), .ZN(n8351) );
  NOR2_X1 U9900 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  NOR2_X1 U9901 ( .A1(n9380), .A2(n8349), .ZN(n8525) );
  NAND2_X1 U9902 ( .A1(n8525), .A2(n9311), .ZN(n9678) );
  NOR2_X1 U9903 ( .A1(n4421), .A2(n9678), .ZN(n9341) );
  AOI21_X1 U9904 ( .B1(n4421), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9341), .ZN(
        n8350) );
  OAI211_X1 U9905 ( .C1(n9550), .C2(n9533), .A(n8351), .B(n8350), .ZN(P1_U3261) );
  INV_X1 U9906 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8358) );
  XNOR2_X1 U9907 ( .A(n9829), .B(n8358), .ZN(n9832) );
  XNOR2_X1 U9908 ( .A(n9338), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U9909 ( .A1(n8352), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8355) );
  INV_X1 U9910 ( .A(n8353), .ZN(n8354) );
  NAND2_X1 U9911 ( .A1(n8355), .A2(n8354), .ZN(n9327) );
  NAND2_X1 U9912 ( .A1(n9328), .A2(n9327), .ZN(n9326) );
  INV_X1 U9913 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8356) );
  OR2_X1 U9914 ( .A1(n9338), .A2(n8356), .ZN(n8357) );
  NAND2_X1 U9915 ( .A1(n9326), .A2(n8357), .ZN(n9831) );
  NAND2_X1 U9916 ( .A1(n9829), .A2(n8358), .ZN(n8359) );
  NAND2_X1 U9917 ( .A1(n9835), .A2(n8359), .ZN(n8361) );
  INV_X1 U9918 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8360) );
  XNOR2_X1 U9919 ( .A(n8361), .B(n8360), .ZN(n8373) );
  INV_X1 U9920 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8362) );
  OR2_X1 U9921 ( .A1(n9829), .A2(n8362), .ZN(n8368) );
  NAND2_X1 U9922 ( .A1(n9829), .A2(n8362), .ZN(n8363) );
  AND2_X1 U9923 ( .A1(n8368), .A2(n8363), .ZN(n9825) );
  XNOR2_X1 U9924 ( .A(n9338), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U9925 ( .A1(n9335), .A2(n9334), .ZN(n9333) );
  INV_X1 U9926 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8366) );
  OR2_X1 U9927 ( .A1(n9338), .A2(n8366), .ZN(n8367) );
  NAND2_X1 U9928 ( .A1(n9333), .A2(n8367), .ZN(n9824) );
  NAND2_X1 U9929 ( .A1(n9825), .A2(n9824), .ZN(n9822) );
  NAND2_X1 U9930 ( .A1(n9822), .A2(n8368), .ZN(n8369) );
  XNOR2_X1 U9931 ( .A(n8369), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8372) );
  INV_X1 U9932 ( .A(n8372), .ZN(n8370) );
  OAI22_X1 U9933 ( .A1(n9833), .A2(n8373), .B1(n9782), .B2(n8372), .ZN(n8374)
         );
  NAND2_X1 U9934 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9193) );
  OAI211_X1 U9935 ( .C1(n8376), .C2(n9821), .A(n8375), .B(n9193), .ZN(P1_U3260) );
  OAI21_X1 U9936 ( .B1(n8386), .B2(n9146), .A(n8381), .ZN(P2_U3517) );
  OAI21_X1 U9937 ( .B1(n8386), .B2(n9060), .A(n8385), .ZN(P2_U3549) );
  INV_X1 U9938 ( .A(n8387), .ZN(n8388) );
  NAND2_X1 U9939 ( .A1(n8389), .A2(n8388), .ZN(n8390) );
  XNOR2_X1 U9940 ( .A(n9080), .B(n8448), .ZN(n8393) );
  NOR2_X1 U9941 ( .A1(n8978), .A2(n8455), .ZN(n8679) );
  NAND2_X1 U9942 ( .A1(n8671), .A2(n8679), .ZN(n8396) );
  INV_X1 U9943 ( .A(n8392), .ZN(n8395) );
  INV_X1 U9944 ( .A(n8393), .ZN(n8394) );
  XNOR2_X1 U9945 ( .A(n8993), .B(n8448), .ZN(n8399) );
  NOR2_X1 U9946 ( .A1(n8956), .A2(n8455), .ZN(n8397) );
  XNOR2_X1 U9947 ( .A(n8399), .B(n8397), .ZN(n8468) );
  INV_X1 U9948 ( .A(n8397), .ZN(n8398) );
  NAND2_X1 U9949 ( .A1(n8399), .A2(n8398), .ZN(n8400) );
  XNOR2_X1 U9950 ( .A(n8960), .B(n8453), .ZN(n8401) );
  NOR2_X1 U9951 ( .A1(n8980), .A2(n8455), .ZN(n8402) );
  NAND2_X1 U9952 ( .A1(n8401), .A2(n8402), .ZN(n8406) );
  INV_X1 U9953 ( .A(n8401), .ZN(n8655) );
  INV_X1 U9954 ( .A(n8402), .ZN(n8403) );
  NAND2_X1 U9955 ( .A1(n8655), .A2(n8403), .ZN(n8404) );
  NAND2_X1 U9956 ( .A1(n8406), .A2(n8404), .ZN(n8603) );
  XNOR2_X1 U9957 ( .A(n9061), .B(n8453), .ZN(n8407) );
  NOR2_X1 U9958 ( .A1(n8955), .A2(n8455), .ZN(n8408) );
  NAND2_X1 U9959 ( .A1(n8407), .A2(n8408), .ZN(n8411) );
  INV_X1 U9960 ( .A(n8407), .ZN(n8561) );
  INV_X1 U9961 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U9962 ( .A1(n8561), .A2(n8409), .ZN(n8410) );
  AND2_X1 U9963 ( .A1(n8411), .A2(n8410), .ZN(n8652) );
  XNOR2_X1 U9964 ( .A(n9143), .B(n8453), .ZN(n8413) );
  NAND2_X1 U9965 ( .A1(n8946), .A2(n8432), .ZN(n8414) );
  XNOR2_X1 U9966 ( .A(n8413), .B(n8414), .ZN(n8562) );
  AND2_X1 U9967 ( .A1(n8562), .A2(n8411), .ZN(n8412) );
  INV_X1 U9968 ( .A(n8413), .ZN(n8415) );
  NAND2_X1 U9969 ( .A1(n8415), .A2(n8414), .ZN(n8416) );
  XNOR2_X1 U9970 ( .A(n9049), .B(n8453), .ZN(n8417) );
  NOR2_X1 U9971 ( .A1(n8892), .A2(n8455), .ZN(n8418) );
  NAND2_X1 U9972 ( .A1(n8417), .A2(n8418), .ZN(n8421) );
  INV_X1 U9973 ( .A(n8417), .ZN(n8570) );
  INV_X1 U9974 ( .A(n8418), .ZN(n8419) );
  NAND2_X1 U9975 ( .A1(n8570), .A2(n8419), .ZN(n8420) );
  AND2_X1 U9976 ( .A1(n8421), .A2(n8420), .ZN(n8621) );
  XNOR2_X1 U9977 ( .A(n8904), .B(n8453), .ZN(n8425) );
  NAND2_X1 U9978 ( .A1(n8915), .A2(n8432), .ZN(n8423) );
  XNOR2_X1 U9979 ( .A(n8425), .B(n8423), .ZN(n8568) );
  NAND2_X1 U9980 ( .A1(n8422), .A2(n8568), .ZN(n8571) );
  INV_X1 U9981 ( .A(n8423), .ZN(n8424) );
  NAND2_X1 U9982 ( .A1(n8425), .A2(n8424), .ZN(n8426) );
  NAND2_X1 U9983 ( .A1(n8571), .A2(n8426), .ZN(n8429) );
  XNOR2_X1 U9984 ( .A(n9131), .B(n8448), .ZN(n8427) );
  XNOR2_X1 U9985 ( .A(n8429), .B(n8427), .ZN(n8630) );
  OR2_X1 U9986 ( .A1(n8893), .A2(n8455), .ZN(n8628) );
  NAND2_X1 U9987 ( .A1(n8630), .A2(n8628), .ZN(n8431) );
  INV_X1 U9988 ( .A(n8427), .ZN(n8428) );
  OR2_X1 U9989 ( .A1(n8429), .A2(n8428), .ZN(n8430) );
  XNOR2_X1 U9990 ( .A(n9036), .B(n8453), .ZN(n8434) );
  XNOR2_X1 U9991 ( .A(n8858), .B(n8448), .ZN(n8611) );
  INV_X1 U9992 ( .A(n8634), .ZN(n8691) );
  NAND2_X1 U9993 ( .A1(n8691), .A2(n8432), .ZN(n8549) );
  AOI21_X1 U9994 ( .B1(n8611), .B2(n8690), .A(n8549), .ZN(n8433) );
  NAND2_X1 U9995 ( .A1(n8550), .A2(n8433), .ZN(n8441) );
  NOR2_X1 U9996 ( .A1(n8690), .A2(n8455), .ZN(n8438) );
  INV_X1 U9997 ( .A(n8611), .ZN(n8437) );
  OAI21_X1 U9998 ( .B1(n8438), .B2(n8437), .A(n8609), .ZN(n8440) );
  INV_X1 U9999 ( .A(n8438), .ZN(n8614) );
  NAND3_X1 U10000 ( .A1(n8441), .A2(n8440), .A3(n8439), .ZN(n8583) );
  XNOR2_X1 U10001 ( .A(n9027), .B(n8453), .ZN(n8442) );
  NOR2_X1 U10002 ( .A1(n8822), .A2(n8455), .ZN(n8443) );
  AND2_X1 U10003 ( .A1(n8442), .A2(n8443), .ZN(n8579) );
  INV_X1 U10004 ( .A(n8442), .ZN(n8580) );
  INV_X1 U10005 ( .A(n8443), .ZN(n8444) );
  NAND2_X1 U10006 ( .A1(n8580), .A2(n8444), .ZN(n8578) );
  OAI21_X1 U10007 ( .B1(n8583), .B2(n8579), .A(n8578), .ZN(n8663) );
  XNOR2_X1 U10008 ( .A(n9115), .B(n8453), .ZN(n8446) );
  NOR2_X1 U10009 ( .A1(n8802), .A2(n8455), .ZN(n8445) );
  XNOR2_X1 U10010 ( .A(n8446), .B(n8445), .ZN(n8662) );
  NAND2_X1 U10011 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  XNOR2_X1 U10012 ( .A(n8814), .B(n8448), .ZN(n8449) );
  NOR2_X1 U10013 ( .A1(n8823), .A2(n8455), .ZN(n8450) );
  XNOR2_X1 U10014 ( .A(n8449), .B(n8450), .ZN(n8542) );
  NAND2_X1 U10015 ( .A1(n8541), .A2(n8542), .ZN(n8452) );
  INV_X1 U10016 ( .A(n8449), .ZN(n8451) );
  XNOR2_X1 U10017 ( .A(n8794), .B(n8453), .ZN(n8454) );
  OAI21_X1 U10018 ( .B1(n8803), .B2(n8455), .A(n8629), .ZN(n8464) );
  INV_X1 U10019 ( .A(n8803), .ZN(n8686) );
  INV_X1 U10020 ( .A(n8458), .ZN(n8789) );
  OAI22_X1 U10021 ( .A1(n8789), .A2(n10341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8459), .ZN(n8462) );
  OAI22_X1 U10022 ( .A1(n8460), .A2(n10343), .B1(n8665), .B2(n8823), .ZN(n8461) );
  AOI211_X1 U10023 ( .C1(n8794), .C2(n8668), .A(n8462), .B(n8461), .ZN(n8463)
         );
  AOI22_X1 U10024 ( .A1(n10349), .A2(n8693), .B1(n8675), .B2(n8944), .ZN(n8466) );
  OAI211_X1 U10025 ( .C1(n8990), .C2(n10341), .A(n8466), .B(n8465), .ZN(n8471)
         );
  INV_X1 U10026 ( .A(n8672), .ZN(n8467) );
  NOR2_X1 U10027 ( .A1(n8456), .A2(n8978), .ZN(n8683) );
  AOI22_X1 U10028 ( .A1(n8467), .A2(n8629), .B1(n8683), .B2(n8671), .ZN(n8469)
         );
  NOR2_X1 U10029 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  AOI211_X1 U10030 ( .C1(n8993), .C2(n8668), .A(n8471), .B(n8470), .ZN(n8472)
         );
  OAI21_X1 U10031 ( .B1(n8473), .B2(n10351), .A(n8472), .ZN(P2_U3228) );
  INV_X1 U10032 ( .A(n8475), .ZN(n8477) );
  NOR2_X1 U10033 ( .A1(n8477), .A2(n8476), .ZN(n8478) );
  XNOR2_X1 U10034 ( .A(n8474), .B(n8478), .ZN(n8483) );
  AOI22_X1 U10035 ( .A1(n9266), .A2(n9462), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8480) );
  NAND2_X1 U10036 ( .A1(n9306), .A2(n9468), .ZN(n8479) );
  OAI211_X1 U10037 ( .C1(n9194), .C2(n9234), .A(n8480), .B(n8479), .ZN(n8481)
         );
  AOI21_X1 U10038 ( .B1(n9592), .B2(n9291), .A(n8481), .ZN(n8482) );
  OAI21_X1 U10039 ( .B1(n8483), .B2(n9309), .A(n8482), .ZN(P1_U3221) );
  INV_X1 U10040 ( .A(n9406), .ZN(n8489) );
  INV_X1 U10041 ( .A(n9581), .ZN(n9430) );
  INV_X1 U10042 ( .A(n9610), .ZN(n9534) );
  INV_X1 U10043 ( .A(n9600), .ZN(n9500) );
  NAND2_X1 U10044 ( .A1(n9474), .A2(n8485), .ZN(n8486) );
  INV_X1 U10045 ( .A(n9595), .ZN(n9479) );
  NAND2_X1 U10046 ( .A1(n8486), .A2(n4971), .ZN(n9458) );
  NAND2_X1 U10047 ( .A1(n8489), .A2(n8490), .ZN(n8491) );
  NAND2_X1 U10048 ( .A1(n9346), .A2(n9345), .ZN(n9344) );
  NAND2_X1 U10049 ( .A1(n8495), .A2(n8494), .ZN(n8524) );
  AOI21_X1 U10050 ( .B1(n9551), .B2(n8496), .A(n9340), .ZN(n9552) );
  AOI22_X1 U10051 ( .A1(n4421), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8497), .B2(
        n9530), .ZN(n8498) );
  OAI21_X1 U10052 ( .B1(n8499), .B2(n9533), .A(n8498), .ZN(n8529) );
  INV_X1 U10053 ( .A(n8500), .ZN(n8501) );
  NAND2_X1 U10054 ( .A1(n8502), .A2(n8501), .ZN(n8504) );
  NAND2_X1 U10055 ( .A1(n8504), .A2(n8503), .ZN(n9536) );
  INV_X1 U10056 ( .A(n9536), .ZN(n8508) );
  INV_X1 U10057 ( .A(n8506), .ZN(n8507) );
  NAND2_X1 U10058 ( .A1(n9502), .A2(n9503), .ZN(n9501) );
  NAND2_X1 U10059 ( .A1(n9461), .A2(n9460), .ZN(n9459) );
  AND2_X2 U10060 ( .A1(n9459), .A2(n8512), .ZN(n9450) );
  INV_X1 U10061 ( .A(n8516), .ZN(n8518) );
  OAI21_X1 U10062 ( .B1(n9398), .B2(n8518), .A(n8517), .ZN(n9383) );
  INV_X1 U10063 ( .A(n8519), .ZN(n8520) );
  NAND2_X1 U10064 ( .A1(n9350), .A2(n8522), .ZN(n8523) );
  INV_X1 U10065 ( .A(n8525), .ZN(n8526) );
  OAI222_X1 U10066 ( .A1(n9484), .A2(n8527), .B1(n6351), .B2(n8526), .C1(n8534), .C2(n9431), .ZN(n8528) );
  AOI22_X1 U10067 ( .A1(n9298), .A2(n9399), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8533) );
  NAND2_X1 U10068 ( .A1(n9306), .A2(n9370), .ZN(n8532) );
  OAI211_X1 U10069 ( .C1(n8534), .C2(n9301), .A(n8533), .B(n8532), .ZN(n8535)
         );
  AOI21_X1 U10070 ( .B1(n9561), .B2(n9291), .A(n8535), .ZN(n8536) );
  OAI21_X1 U10071 ( .B1(n8537), .B2(n9309), .A(n8536), .ZN(P1_U3212) );
  OAI222_X1 U10072 ( .A1(n8540), .A2(n8539), .B1(n9651), .B2(n8538), .C1(n6553), .C2(P1_U3084), .ZN(P1_U3331) );
  XNOR2_X1 U10073 ( .A(n8541), .B(n8542), .ZN(n8548) );
  INV_X1 U10074 ( .A(n8543), .ZN(n8809) );
  OAI22_X1 U10075 ( .A1(n10341), .A2(n8809), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8544), .ZN(n8546) );
  OAI22_X1 U10076 ( .A1(n8803), .A2(n10343), .B1(n8665), .B2(n8802), .ZN(n8545) );
  AOI211_X1 U10077 ( .C1(n8814), .C2(n8668), .A(n8546), .B(n8545), .ZN(n8547)
         );
  OAI21_X1 U10078 ( .B1(n8548), .B2(n10351), .A(n8547), .ZN(P2_U3216) );
  AOI22_X1 U10079 ( .A1(n8550), .A2(n8629), .B1(n8627), .B2(n8691), .ZN(n8555)
         );
  OAI22_X1 U10080 ( .A1(n10341), .A2(n8869), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8551), .ZN(n8553) );
  OAI22_X1 U10081 ( .A1(n8690), .A2(n10343), .B1(n8665), .B2(n8893), .ZN(n8552) );
  AOI211_X1 U10082 ( .C1(n9036), .C2(n8668), .A(n8553), .B(n8552), .ZN(n8554)
         );
  OAI21_X1 U10083 ( .B1(n8610), .B2(n8555), .A(n8554), .ZN(P2_U3218) );
  OAI21_X1 U10084 ( .B1(n8562), .B2(n8556), .A(n8557), .ZN(n8558) );
  NAND2_X1 U10085 ( .A1(n8558), .A2(n8629), .ZN(n8566) );
  NOR2_X1 U10086 ( .A1(n10343), .A2(n8892), .ZN(n8560) );
  NAND2_X1 U10087 ( .A1(n4420), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8776) );
  OAI21_X1 U10088 ( .B1(n10341), .B2(n8931), .A(n8776), .ZN(n8559) );
  AOI211_X1 U10089 ( .C1(n9143), .C2(n8668), .A(n8560), .B(n8559), .ZN(n8565)
         );
  NOR3_X1 U10090 ( .A1(n8562), .A2(n8561), .A3(n8456), .ZN(n8563) );
  OAI21_X1 U10091 ( .B1(n8563), .B2(n10349), .A(n5830), .ZN(n8564) );
  NAND3_X1 U10092 ( .A1(n8566), .A2(n8565), .A3(n8564), .ZN(P2_U3221) );
  INV_X1 U10093 ( .A(n8568), .ZN(n8569) );
  AOI21_X1 U10094 ( .B1(n8567), .B2(n8569), .A(n10351), .ZN(n8573) );
  NOR3_X1 U10095 ( .A1(n8570), .A2(n8892), .A3(n8456), .ZN(n8572) );
  OAI21_X1 U10096 ( .B1(n8573), .B2(n8572), .A(n8571), .ZN(n8577) );
  NOR2_X1 U10097 ( .A1(n10341), .A2(n8899), .ZN(n8575) );
  OAI22_X1 U10098 ( .A1(n8892), .A2(n8665), .B1(n10343), .B2(n8893), .ZN(n8574) );
  AOI211_X1 U10099 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(n4420), .A(n8575), .B(
        n8574), .ZN(n8576) );
  OAI211_X1 U10100 ( .C1(n9134), .C2(n10345), .A(n8577), .B(n8576), .ZN(
        P2_U3225) );
  INV_X1 U10101 ( .A(n8578), .ZN(n8582) );
  OR3_X1 U10102 ( .A1(n8579), .A2(n8582), .A3(n10351), .ZN(n8585) );
  NOR3_X1 U10103 ( .A1(n8580), .A2(n8822), .A3(n8456), .ZN(n8581) );
  AOI21_X1 U10104 ( .B1(n8629), .B2(n8582), .A(n8581), .ZN(n8584) );
  MUX2_X1 U10105 ( .A(n8585), .B(n8584), .S(n8583), .Z(n8591) );
  INV_X1 U10106 ( .A(n8802), .ZN(n8688) );
  NOR2_X1 U10107 ( .A1(n8690), .A2(n8977), .ZN(n8586) );
  AOI21_X1 U10108 ( .B1(n8688), .B2(n8945), .A(n8586), .ZN(n8842) );
  OAI22_X1 U10109 ( .A1(n8842), .A2(n8637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8587), .ZN(n8588) );
  AOI21_X1 U10110 ( .B1(n8589), .B2(n8674), .A(n8588), .ZN(n8590) );
  OAI211_X1 U10111 ( .C1(n5868), .C2(n10345), .A(n8591), .B(n8590), .ZN(
        P2_U3227) );
  NOR2_X1 U10112 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5107), .ZN(n8725) );
  NOR2_X1 U10113 ( .A1(n10341), .A2(n8592), .ZN(n8593) );
  AOI211_X1 U10114 ( .C1(n10349), .C2(n8704), .A(n8725), .B(n8593), .ZN(n8601)
         );
  AOI22_X1 U10115 ( .A1(n8675), .A2(n8702), .B1(n8594), .B2(n8668), .ZN(n8600)
         );
  OAI21_X1 U10116 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n8598) );
  NAND2_X1 U10117 ( .A1(n8598), .A2(n8629), .ZN(n8599) );
  NAND3_X1 U10118 ( .A1(n8601), .A2(n8600), .A3(n8599), .ZN(P2_U3229) );
  INV_X1 U10119 ( .A(n8654), .ZN(n8602) );
  AOI211_X1 U10120 ( .C1(n8604), .C2(n8603), .A(n10351), .B(n8602), .ZN(n8608)
         );
  AOI22_X1 U10121 ( .A1(n8674), .A2(n8963), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        n4420), .ZN(n8606) );
  AOI22_X1 U10122 ( .A1(n8675), .A2(n5830), .B1(n10349), .B2(n8692), .ZN(n8605) );
  OAI211_X1 U10123 ( .C1(n5829), .C2(n10345), .A(n8606), .B(n8605), .ZN(n8607)
         );
  OR2_X1 U10124 ( .A1(n8608), .A2(n8607), .ZN(P2_U3230) );
  XNOR2_X1 U10125 ( .A(n8612), .B(n8611), .ZN(n8615) );
  OAI22_X1 U10126 ( .A1(n8615), .A2(n10351), .B1(n8690), .B2(n8456), .ZN(n8613) );
  OAI21_X1 U10127 ( .B1(n8615), .B2(n8614), .A(n8613), .ZN(n8619) );
  INV_X1 U10128 ( .A(n8856), .ZN(n8617) );
  AOI22_X1 U10129 ( .A1(n8689), .A2(n8945), .B1(n8943), .B2(n8691), .ZN(n8847)
         );
  OAI22_X1 U10130 ( .A1(n8847), .A2(n8637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10230), .ZN(n8616) );
  AOI21_X1 U10131 ( .B1(n8617), .B2(n8674), .A(n8616), .ZN(n8618) );
  OAI211_X1 U10132 ( .C1(n9123), .C2(n10345), .A(n8619), .B(n8618), .ZN(
        P2_U3231) );
  OAI211_X1 U10133 ( .C1(n8621), .C2(n8620), .A(n8567), .B(n8629), .ZN(n8626)
         );
  NOR2_X1 U10134 ( .A1(n8622), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8624) );
  OAI22_X1 U10135 ( .A1(n8633), .A2(n10343), .B1(n8665), .B2(n8658), .ZN(n8623) );
  AOI211_X1 U10136 ( .C1(n8674), .C2(n8909), .A(n8624), .B(n8623), .ZN(n8625)
         );
  OAI211_X1 U10137 ( .C1(n8911), .C2(n10345), .A(n8626), .B(n8625), .ZN(
        P2_U3235) );
  NAND2_X1 U10138 ( .A1(n8627), .A2(n4669), .ZN(n8632) );
  NAND2_X1 U10139 ( .A1(n8629), .A2(n8628), .ZN(n8631) );
  MUX2_X1 U10140 ( .A(n8632), .B(n8631), .S(n8630), .Z(n8640) );
  OAI22_X1 U10141 ( .A1(n8634), .A2(n8979), .B1(n8633), .B2(n8977), .ZN(n8880)
         );
  INV_X1 U10142 ( .A(n8880), .ZN(n8636) );
  OAI22_X1 U10143 ( .A1(n8637), .A2(n8636), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8635), .ZN(n8638) );
  AOI21_X1 U10144 ( .B1(n8885), .B2(n8674), .A(n8638), .ZN(n8639) );
  OAI211_X1 U10145 ( .C1(n4606), .C2(n10345), .A(n8640), .B(n8639), .ZN(
        P2_U3237) );
  INV_X1 U10146 ( .A(n8641), .ZN(n8644) );
  OAI22_X1 U10147 ( .A1(n9962), .A2(n10345), .B1(n10351), .B2(n8642), .ZN(
        n8643) );
  AOI21_X1 U10148 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n8644), .A(n8643), .ZN(
        n8651) );
  AOI22_X1 U10149 ( .A1(n10349), .A2(n8707), .B1(n8675), .B2(n10348), .ZN(
        n8650) );
  OAI22_X1 U10150 ( .A1(n8456), .A2(n5047), .B1(n7230), .B2(n10351), .ZN(n8648) );
  INV_X1 U10151 ( .A(n8645), .ZN(n8647) );
  NAND3_X1 U10152 ( .A1(n8648), .A2(n8647), .A3(n8646), .ZN(n8649) );
  NAND3_X1 U10153 ( .A1(n8651), .A2(n8650), .A3(n8649), .ZN(P2_U3239) );
  INV_X1 U10154 ( .A(n8652), .ZN(n8653) );
  AOI21_X1 U10155 ( .B1(n8654), .B2(n8653), .A(n10351), .ZN(n8657) );
  NOR3_X1 U10156 ( .A1(n8655), .A2(n8980), .A3(n8456), .ZN(n8656) );
  OAI21_X1 U10157 ( .B1(n8657), .B2(n8656), .A(n8556), .ZN(n8661) );
  AND2_X1 U10158 ( .A1(n4420), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8755) );
  OAI22_X1 U10159 ( .A1(n8980), .A2(n8665), .B1(n10343), .B2(n8658), .ZN(n8659) );
  AOI211_X1 U10160 ( .C1(n8674), .C2(n8937), .A(n8755), .B(n8659), .ZN(n8660)
         );
  OAI211_X1 U10161 ( .C1(n8939), .C2(n10345), .A(n8661), .B(n8660), .ZN(
        P2_U3240) );
  XNOR2_X1 U10162 ( .A(n8663), .B(n8662), .ZN(n8670) );
  OAI22_X1 U10163 ( .A1(n10341), .A2(n8828), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8664), .ZN(n8667) );
  OAI22_X1 U10164 ( .A1(n8822), .A2(n8665), .B1(n10343), .B2(n8823), .ZN(n8666) );
  AOI211_X1 U10165 ( .C1(n9115), .C2(n8668), .A(n8667), .B(n8666), .ZN(n8669)
         );
  OAI21_X1 U10166 ( .B1(n8670), .B2(n10351), .A(n8669), .ZN(P2_U3242) );
  NAND2_X1 U10167 ( .A1(n8672), .A2(n8671), .ZN(n8682) );
  AOI22_X1 U10168 ( .A1(n8674), .A2(n8673), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        n4420), .ZN(n8677) );
  AOI22_X1 U10169 ( .A1(n10349), .A2(n8694), .B1(n8675), .B2(n8692), .ZN(n8676) );
  OAI211_X1 U10170 ( .C1(n8678), .C2(n10345), .A(n8677), .B(n8676), .ZN(n8681)
         );
  NOR3_X1 U10171 ( .A1(n8682), .A2(n8679), .A3(n10351), .ZN(n8680) );
  AOI211_X1 U10172 ( .C1(n8683), .C2(n8682), .A(n8681), .B(n8680), .ZN(n8684)
         );
  INV_X1 U10173 ( .A(n8684), .ZN(P2_U3243) );
  MUX2_X1 U10174 ( .A(n8685), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8706), .Z(
        P2_U3582) );
  MUX2_X1 U10175 ( .A(n8686), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8706), .Z(
        P2_U3580) );
  MUX2_X1 U10176 ( .A(n8687), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8706), .Z(
        P2_U3579) );
  MUX2_X1 U10177 ( .A(n8688), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8706), .Z(
        P2_U3578) );
  MUX2_X1 U10178 ( .A(n8689), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8706), .Z(
        P2_U3577) );
  MUX2_X1 U10179 ( .A(n4691), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8706), .Z(
        P2_U3576) );
  MUX2_X1 U10180 ( .A(n8691), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8706), .Z(
        P2_U3575) );
  MUX2_X1 U10181 ( .A(n4669), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8706), .Z(
        P2_U3574) );
  MUX2_X1 U10182 ( .A(n8915), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8706), .Z(
        P2_U3573) );
  MUX2_X1 U10183 ( .A(n8924), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8706), .Z(
        P2_U3572) );
  MUX2_X1 U10184 ( .A(n8946), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8706), .Z(
        P2_U3571) );
  MUX2_X1 U10185 ( .A(n5830), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8706), .Z(
        P2_U3570) );
  MUX2_X1 U10186 ( .A(n8944), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8706), .Z(
        P2_U3569) );
  MUX2_X1 U10187 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8692), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10188 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8693), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10189 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8694), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10190 ( .A(n8695), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8706), .Z(
        P2_U3565) );
  MUX2_X1 U10191 ( .A(n8696), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8706), .Z(
        P2_U3564) );
  MUX2_X1 U10192 ( .A(n8697), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8706), .Z(
        P2_U3563) );
  MUX2_X1 U10193 ( .A(n8698), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8706), .Z(
        P2_U3562) );
  MUX2_X1 U10194 ( .A(n8699), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8706), .Z(
        P2_U3561) );
  MUX2_X1 U10195 ( .A(n8700), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8706), .Z(
        P2_U3560) );
  MUX2_X1 U10196 ( .A(n8701), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8706), .Z(
        P2_U3559) );
  MUX2_X1 U10197 ( .A(n8702), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8706), .Z(
        P2_U3558) );
  MUX2_X1 U10198 ( .A(n8703), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8706), .Z(
        P2_U3557) );
  MUX2_X1 U10199 ( .A(n8704), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8706), .Z(
        P2_U3556) );
  MUX2_X1 U10200 ( .A(n10348), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8706), .Z(
        P2_U3555) );
  MUX2_X1 U10201 ( .A(n8705), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8706), .Z(
        P2_U3554) );
  MUX2_X1 U10202 ( .A(n8707), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8706), .Z(
        P2_U3553) );
  NAND2_X1 U10203 ( .A1(n9924), .A2(n8709), .ZN(n8720) );
  NOR2_X1 U10204 ( .A1(n8708), .A2(n6908), .ZN(n8713) );
  MUX2_X1 U10205 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n8710), .S(n8709), .Z(n8712)
         );
  OAI211_X1 U10206 ( .C1(n8713), .C2(n8712), .A(n9904), .B(n8711), .ZN(n8719)
         );
  AOI22_X1 U10207 ( .A1(n9917), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n4420), .ZN(n8718) );
  OAI211_X1 U10208 ( .C1(n8716), .C2(n8715), .A(n9922), .B(n8714), .ZN(n8717)
         );
  NAND4_X1 U10209 ( .A1(n8720), .A2(n8719), .A3(n8718), .A4(n8717), .ZN(
        P2_U3246) );
  OAI211_X1 U10210 ( .C1(n8723), .C2(n8722), .A(n9904), .B(n8721), .ZN(n8733)
         );
  NAND2_X1 U10211 ( .A1(n9924), .A2(n8724), .ZN(n8732) );
  AOI21_X1 U10212 ( .B1(n9917), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8725), .ZN(
        n8731) );
  OAI21_X1 U10213 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8729) );
  OR2_X1 U10214 ( .A1(n9906), .A2(n8729), .ZN(n8730) );
  NAND4_X1 U10215 ( .A1(n8733), .A2(n8732), .A3(n8731), .A4(n8730), .ZN(
        P2_U3250) );
  OAI211_X1 U10216 ( .C1(n8736), .C2(n8735), .A(n9904), .B(n8734), .ZN(n8746)
         );
  NAND2_X1 U10217 ( .A1(n9924), .A2(n8737), .ZN(n8745) );
  AOI21_X1 U10218 ( .B1(n9917), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8738), .ZN(
        n8744) );
  OAI21_X1 U10219 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n8742) );
  OR2_X1 U10220 ( .A1(n9906), .A2(n8742), .ZN(n8743) );
  NAND4_X1 U10221 ( .A1(n8746), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(
        P2_U3252) );
  NAND2_X1 U10222 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n8754), .ZN(n8748) );
  NAND2_X1 U10223 ( .A1(n8748), .A2(n8747), .ZN(n8749) );
  AOI21_X1 U10224 ( .B1(n8750), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8768), .ZN(
        n8751) );
  OR2_X1 U10225 ( .A1(n8751), .A2(n9927), .ZN(n8760) );
  XNOR2_X1 U10226 ( .A(n8752), .B(n8763), .ZN(n8762) );
  AOI21_X1 U10227 ( .B1(n8754), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8753), .ZN(
        n8761) );
  XNOR2_X1 U10228 ( .A(n8762), .B(n8761), .ZN(n8758) );
  INV_X1 U10229 ( .A(n8755), .ZN(n8756) );
  OAI21_X1 U10230 ( .B1(n9658), .B2(n10361), .A(n8756), .ZN(n8757) );
  AOI21_X1 U10231 ( .B1(n9922), .B2(n8758), .A(n8757), .ZN(n8759) );
  OAI211_X1 U10232 ( .C1(n9905), .C2(n8764), .A(n8760), .B(n8759), .ZN(
        P2_U3263) );
  NAND2_X1 U10233 ( .A1(n8762), .A2(n8761), .ZN(n8766) );
  NAND2_X1 U10234 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  NAND2_X1 U10235 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  XNOR2_X1 U10236 ( .A(n8767), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8772) );
  INV_X1 U10237 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U10238 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  XOR2_X1 U10239 ( .A(n10273), .B(n8770), .Z(n8774) );
  NAND2_X1 U10240 ( .A1(n8774), .A2(n9904), .ZN(n8771) );
  INV_X1 U10241 ( .A(n8772), .ZN(n8773) );
  OAI22_X1 U10242 ( .A1(n8774), .A2(n9927), .B1(n8773), .B2(n9906), .ZN(n8775)
         );
  NAND2_X1 U10243 ( .A1(n9107), .A2(n8784), .ZN(n8783) );
  NAND2_X1 U10244 ( .A1(n9010), .A2(n8950), .ZN(n8782) );
  INV_X1 U10245 ( .A(n8778), .ZN(n8780) );
  AND2_X1 U10246 ( .A1(n8780), .A2(n8779), .ZN(n9009) );
  INV_X1 U10247 ( .A(n9009), .ZN(n9012) );
  NOR2_X1 U10248 ( .A1(n8998), .A2(n9012), .ZN(n8786) );
  AOI21_X1 U10249 ( .B1(n9944), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8786), .ZN(
        n8781) );
  OAI211_X1 U10250 ( .C1(n9103), .C2(n9937), .A(n8782), .B(n8781), .ZN(
        P2_U3265) );
  OAI211_X1 U10251 ( .C1(n9107), .C2(n8784), .A(n9959), .B(n8783), .ZN(n9013)
         );
  NOR2_X1 U10252 ( .A1(n9107), .A2(n9937), .ZN(n8785) );
  AOI211_X1 U10253 ( .C1(n9944), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8786), .B(
        n8785), .ZN(n8787) );
  OAI21_X1 U10254 ( .B1(n8995), .B2(n9013), .A(n8787), .ZN(P2_U3266) );
  OAI22_X1 U10255 ( .A1(n9001), .A2(n8790), .B1(n8789), .B2(n8989), .ZN(n8793)
         );
  NOR2_X1 U10256 ( .A1(n8791), .A2(n8995), .ZN(n8792) );
  AOI211_X1 U10257 ( .C1(n9002), .C2(n8794), .A(n8793), .B(n8792), .ZN(n8795)
         );
  OAI211_X1 U10258 ( .C1(n9944), .C2(n8797), .A(n8796), .B(n8795), .ZN(
        P2_U3268) );
  NAND2_X1 U10259 ( .A1(n8798), .A2(n8799), .ZN(n8801) );
  XNOR2_X1 U10260 ( .A(n8801), .B(n8800), .ZN(n8805) );
  OAI22_X1 U10261 ( .A1(n8803), .A2(n8979), .B1(n8802), .B2(n8977), .ZN(n8804)
         );
  XNOR2_X1 U10262 ( .A(n8807), .B(n8806), .ZN(n9109) );
  INV_X1 U10263 ( .A(n9109), .ZN(n8808) );
  NAND2_X1 U10264 ( .A1(n8808), .A2(n9940), .ZN(n8816) );
  OAI22_X1 U10265 ( .A1(n9001), .A2(n8810), .B1(n8809), .B2(n8989), .ZN(n8813)
         );
  OAI211_X1 U10266 ( .C1(n9108), .C2(n8826), .A(n9959), .B(n8811), .ZN(n9016)
         );
  NOR2_X1 U10267 ( .A1(n9016), .A2(n8995), .ZN(n8812) );
  AOI211_X1 U10268 ( .C1(n9002), .C2(n8814), .A(n8813), .B(n8812), .ZN(n8815)
         );
  OAI211_X1 U10269 ( .C1(n9944), .C2(n9017), .A(n8816), .B(n8815), .ZN(
        P2_U3269) );
  XOR2_X1 U10270 ( .A(n8820), .B(n8817), .Z(n9118) );
  AOI22_X1 U10271 ( .A1(n9115), .A2(n9002), .B1(n9944), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8831) );
  INV_X1 U10272 ( .A(n8798), .ZN(n8819) );
  AOI21_X1 U10273 ( .B1(n8820), .B2(n8818), .A(n8819), .ZN(n8821) );
  OAI222_X1 U10274 ( .A1(n8979), .A2(n8823), .B1(n8977), .B2(n8822), .C1(n8954), .C2(n8821), .ZN(n9021) );
  NAND2_X1 U10275 ( .A1(n9115), .A2(n8834), .ZN(n8824) );
  NAND2_X1 U10276 ( .A1(n8824), .A2(n9959), .ZN(n8825) );
  NOR2_X1 U10277 ( .A1(n8826), .A2(n8825), .ZN(n9020) );
  NAND2_X1 U10278 ( .A1(n9020), .A2(n8929), .ZN(n8827) );
  OAI21_X1 U10279 ( .B1(n8989), .B2(n8828), .A(n8827), .ZN(n8829) );
  OAI21_X1 U10280 ( .B1(n9021), .B2(n8829), .A(n9001), .ZN(n8830) );
  OAI211_X1 U10281 ( .C1(n9118), .C2(n5915), .A(n8831), .B(n8830), .ZN(
        P2_U3270) );
  XOR2_X1 U10282 ( .A(n8840), .B(n8832), .Z(n9122) );
  INV_X1 U10283 ( .A(n8834), .ZN(n8835) );
  AOI211_X1 U10284 ( .C1(n9027), .C2(n8853), .A(n9981), .B(n8835), .ZN(n9026)
         );
  NOR2_X1 U10285 ( .A1(n5868), .A2(n9937), .ZN(n8839) );
  OAI22_X1 U10286 ( .A1(n9001), .A2(n8837), .B1(n8836), .B2(n8989), .ZN(n8838)
         );
  AOI211_X1 U10287 ( .C1(n9026), .C2(n9930), .A(n8839), .B(n8838), .ZN(n8845)
         );
  XNOR2_X1 U10288 ( .A(n8841), .B(n8840), .ZN(n8843) );
  OAI21_X1 U10289 ( .B1(n8843), .B2(n8954), .A(n8842), .ZN(n9025) );
  NAND2_X1 U10290 ( .A1(n9025), .A2(n9001), .ZN(n8844) );
  OAI211_X1 U10291 ( .C1(n9122), .C2(n5915), .A(n8845), .B(n8844), .ZN(
        P2_U3271) );
  XNOR2_X1 U10292 ( .A(n8846), .B(n8852), .ZN(n8849) );
  INV_X1 U10293 ( .A(n8847), .ZN(n8848) );
  AOI21_X1 U10294 ( .B1(n8849), .B2(n8982), .A(n8848), .ZN(n9031) );
  AOI21_X1 U10295 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n9124) );
  INV_X1 U10296 ( .A(n9124), .ZN(n8861) );
  AOI21_X1 U10297 ( .B1(n8871), .B2(n8858), .A(n9981), .ZN(n8854) );
  NAND2_X1 U10298 ( .A1(n8854), .A2(n8853), .ZN(n9030) );
  NAND2_X1 U10299 ( .A1(n9944), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8855) );
  OAI21_X1 U10300 ( .B1(n8989), .B2(n8856), .A(n8855), .ZN(n8857) );
  AOI21_X1 U10301 ( .B1(n8858), .B2(n9002), .A(n8857), .ZN(n8859) );
  OAI21_X1 U10302 ( .B1(n9030), .B2(n8995), .A(n8859), .ZN(n8860) );
  AOI21_X1 U10303 ( .B1(n8861), .B2(n9940), .A(n8860), .ZN(n8862) );
  OAI21_X1 U10304 ( .B1(n9944), .B2(n9031), .A(n8862), .ZN(P2_U3272) );
  OAI21_X1 U10305 ( .B1(n8865), .B2(n8864), .A(n8863), .ZN(n8866) );
  AOI222_X1 U10306 ( .A1(n8982), .A2(n8866), .B1(n4669), .B2(n8943), .C1(n4691), .C2(n8945), .ZN(n9039) );
  OR2_X1 U10307 ( .A1(n8868), .A2(n8867), .ZN(n9035) );
  NAND3_X1 U10308 ( .A1(n9035), .A2(n9034), .A3(n9940), .ZN(n8876) );
  OAI22_X1 U10309 ( .A1(n9001), .A2(n8870), .B1(n8869), .B2(n8989), .ZN(n8874)
         );
  OAI211_X1 U10310 ( .C1(n8872), .C2(n8883), .A(n9959), .B(n8871), .ZN(n9038)
         );
  NOR2_X1 U10311 ( .A1(n9038), .A2(n8995), .ZN(n8873) );
  AOI211_X1 U10312 ( .C1(n9002), .C2(n9036), .A(n8874), .B(n8873), .ZN(n8875)
         );
  OAI211_X1 U10313 ( .C1(n9944), .C2(n9039), .A(n8876), .B(n8875), .ZN(
        P2_U3273) );
  XNOR2_X1 U10314 ( .A(n8878), .B(n8877), .ZN(n9133) );
  AOI21_X1 U10315 ( .B1(n4466), .B2(n8879), .A(n8954), .ZN(n8882) );
  AOI21_X1 U10316 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n9042) );
  INV_X1 U10317 ( .A(n9042), .ZN(n8889) );
  INV_X1 U10318 ( .A(n8901), .ZN(n8884) );
  OAI211_X1 U10319 ( .C1(n4606), .C2(n8884), .A(n4608), .B(n9959), .ZN(n9041)
         );
  AOI22_X1 U10320 ( .A1(n9944), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8885), .B2(
        n9933), .ZN(n8887) );
  NAND2_X1 U10321 ( .A1(n9131), .A2(n9002), .ZN(n8886) );
  OAI211_X1 U10322 ( .C1(n9041), .C2(n8995), .A(n8887), .B(n8886), .ZN(n8888)
         );
  AOI21_X1 U10323 ( .B1(n8889), .B2(n9001), .A(n8888), .ZN(n8890) );
  OAI21_X1 U10324 ( .B1(n9133), .B2(n5915), .A(n8890), .ZN(P2_U3274) );
  XNOR2_X1 U10325 ( .A(n8891), .B(n8896), .ZN(n8895) );
  OAI22_X1 U10326 ( .A1(n8893), .A2(n8979), .B1(n8892), .B2(n8977), .ZN(n8894)
         );
  AOI21_X1 U10327 ( .B1(n8895), .B2(n8982), .A(n8894), .ZN(n9046) );
  XOR2_X1 U10328 ( .A(n8897), .B(n8896), .Z(n9135) );
  INV_X1 U10329 ( .A(n9135), .ZN(n8898) );
  NAND2_X1 U10330 ( .A1(n8898), .A2(n9940), .ZN(n8906) );
  OAI22_X1 U10331 ( .A1(n9001), .A2(n8900), .B1(n8899), .B2(n8989), .ZN(n8903)
         );
  OAI211_X1 U10332 ( .C1(n4490), .C2(n9134), .A(n9959), .B(n8901), .ZN(n9045)
         );
  NOR2_X1 U10333 ( .A1(n9045), .A2(n8995), .ZN(n8902) );
  AOI211_X1 U10334 ( .C1(n9002), .C2(n8904), .A(n8903), .B(n8902), .ZN(n8905)
         );
  OAI211_X1 U10335 ( .C1(n9944), .C2(n9046), .A(n8906), .B(n8905), .ZN(
        P2_U3275) );
  XNOR2_X1 U10336 ( .A(n8907), .B(n8914), .ZN(n9053) );
  INV_X1 U10337 ( .A(n8927), .ZN(n8908) );
  AOI21_X1 U10338 ( .B1(n9049), .B2(n8908), .A(n4490), .ZN(n9050) );
  AOI22_X1 U10339 ( .A1(n9944), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8909), .B2(
        n9933), .ZN(n8910) );
  OAI21_X1 U10340 ( .B1(n8911), .B2(n9937), .A(n8910), .ZN(n8918) );
  NAND2_X1 U10341 ( .A1(n8921), .A2(n8912), .ZN(n8913) );
  XOR2_X1 U10342 ( .A(n8914), .B(n8913), .Z(n8916) );
  AOI222_X1 U10343 ( .A1(n8982), .A2(n8916), .B1(n8946), .B2(n8943), .C1(n8915), .C2(n8945), .ZN(n9052) );
  NOR2_X1 U10344 ( .A1(n9052), .A2(n8998), .ZN(n8917) );
  AOI211_X1 U10345 ( .C1(n9050), .C2(n8950), .A(n8918), .B(n8917), .ZN(n8919)
         );
  OAI21_X1 U10346 ( .B1(n5915), .B2(n9053), .A(n8919), .ZN(P2_U3276) );
  XOR2_X1 U10347 ( .A(n8920), .B(n8923), .Z(n9147) );
  AOI22_X1 U10348 ( .A1(n9143), .A2(n9002), .B1(n9944), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8934) );
  OAI21_X1 U10349 ( .B1(n8923), .B2(n8922), .A(n8921), .ZN(n8925) );
  AOI222_X1 U10350 ( .A1(n8982), .A2(n8925), .B1(n8924), .B2(n8945), .C1(n5830), .C2(n8943), .ZN(n9054) );
  OAI21_X1 U10351 ( .B1(n8936), .B2(n8926), .A(n9959), .ZN(n8928) );
  NOR2_X1 U10352 ( .A1(n8928), .A2(n8927), .ZN(n9055) );
  NAND2_X1 U10353 ( .A1(n9055), .A2(n8929), .ZN(n8930) );
  OAI211_X1 U10354 ( .C1(n8989), .C2(n8931), .A(n9054), .B(n8930), .ZN(n8932)
         );
  NAND2_X1 U10355 ( .A1(n8932), .A2(n9001), .ZN(n8933) );
  OAI211_X1 U10356 ( .C1(n9147), .C2(n5915), .A(n8934), .B(n8933), .ZN(
        P2_U3277) );
  XOR2_X1 U10357 ( .A(n8935), .B(n8940), .Z(n9065) );
  AOI21_X1 U10358 ( .B1(n9061), .B2(n8961), .A(n8936), .ZN(n9062) );
  AOI22_X1 U10359 ( .A1(n9944), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8937), .B2(
        n9933), .ZN(n8938) );
  OAI21_X1 U10360 ( .B1(n8939), .B2(n9937), .A(n8938), .ZN(n8949) );
  INV_X1 U10361 ( .A(n8940), .ZN(n8942) );
  OAI21_X1 U10362 ( .B1(n4494), .B2(n8942), .A(n8941), .ZN(n8947) );
  AOI222_X1 U10363 ( .A1(n8982), .A2(n8947), .B1(n8946), .B2(n8945), .C1(n8944), .C2(n8943), .ZN(n9064) );
  NOR2_X1 U10364 ( .A1(n9064), .A2(n8998), .ZN(n8948) );
  AOI211_X1 U10365 ( .C1(n9062), .C2(n8950), .A(n8949), .B(n8948), .ZN(n8951)
         );
  OAI21_X1 U10366 ( .B1(n9065), .B2(n5915), .A(n8951), .ZN(P2_U3278) );
  XNOR2_X1 U10367 ( .A(n8952), .B(n8958), .ZN(n8953) );
  OAI222_X1 U10368 ( .A1(n8977), .A2(n8956), .B1(n8979), .B2(n8955), .C1(n8954), .C2(n8953), .ZN(n9066) );
  INV_X1 U10369 ( .A(n9066), .ZN(n8968) );
  OAI21_X1 U10370 ( .B1(n8959), .B2(n8958), .A(n8957), .ZN(n9068) );
  AOI21_X1 U10371 ( .B1(n8987), .B2(n8960), .A(n9981), .ZN(n8962) );
  AND2_X1 U10372 ( .A1(n8962), .A2(n8961), .ZN(n9067) );
  NAND2_X1 U10373 ( .A1(n9067), .A2(n9930), .ZN(n8965) );
  AOI22_X1 U10374 ( .A1(n8998), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8963), .B2(
        n9933), .ZN(n8964) );
  OAI211_X1 U10375 ( .C1(n5829), .C2(n9937), .A(n8965), .B(n8964), .ZN(n8966)
         );
  AOI21_X1 U10376 ( .B1(n9068), .B2(n9940), .A(n8966), .ZN(n8967) );
  OAI21_X1 U10377 ( .B1(n9944), .B2(n8968), .A(n8967), .ZN(P2_U3279) );
  AND2_X1 U10378 ( .A1(n8969), .A2(n5360), .ZN(n8970) );
  OR2_X1 U10379 ( .A1(n8971), .A2(n8970), .ZN(n8986) );
  OR2_X1 U10380 ( .A1(n8986), .A2(n8972), .ZN(n8985) );
  NAND2_X1 U10381 ( .A1(n8973), .A2(n8974), .ZN(n8975) );
  NAND2_X1 U10382 ( .A1(n8976), .A2(n8975), .ZN(n8983) );
  OAI22_X1 U10383 ( .A1(n8980), .A2(n8979), .B1(n8978), .B2(n8977), .ZN(n8981)
         );
  AOI21_X1 U10384 ( .B1(n8983), .B2(n8982), .A(n8981), .ZN(n8984) );
  AND2_X1 U10385 ( .A1(n8985), .A2(n8984), .ZN(n9076) );
  INV_X1 U10386 ( .A(n8986), .ZN(n9075) );
  OAI211_X1 U10387 ( .C1(n8988), .C2(n9073), .A(n9959), .B(n8987), .ZN(n9072)
         );
  OAI22_X1 U10388 ( .A1(n9001), .A2(n8991), .B1(n8990), .B2(n8989), .ZN(n8992)
         );
  AOI21_X1 U10389 ( .B1(n8993), .B2(n9002), .A(n8992), .ZN(n8994) );
  OAI21_X1 U10390 ( .B1(n9072), .B2(n8995), .A(n8994), .ZN(n8996) );
  AOI21_X1 U10391 ( .B1(n9075), .B2(n9004), .A(n8996), .ZN(n8997) );
  OAI21_X1 U10392 ( .B1(n9076), .B2(n8998), .A(n8997), .ZN(P2_U3280) );
  NOR2_X1 U10393 ( .A1(n9001), .A2(n5076), .ZN(n8999) );
  AOI21_X1 U10394 ( .B1(n9001), .B2(n9000), .A(n8999), .ZN(n9008) );
  AOI22_X1 U10395 ( .A1(n9004), .A2(n9003), .B1(n9002), .B2(n4823), .ZN(n9007)
         );
  AOI22_X1 U10396 ( .A1(n9930), .A2(n9005), .B1(n9933), .B2(n7226), .ZN(n9006)
         );
  NAND3_X1 U10397 ( .A1(n9008), .A2(n9007), .A3(n9006), .ZN(P2_U3293) );
  INV_X1 U10398 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9011) );
  INV_X1 U10399 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9014) );
  AND2_X1 U10400 ( .A1(n9013), .A2(n9012), .ZN(n9104) );
  MUX2_X1 U10401 ( .A(n9014), .B(n9104), .S(n9996), .Z(n9015) );
  OAI21_X1 U10402 ( .B1(n9107), .B2(n9071), .A(n9015), .ZN(P2_U3550) );
  OAI22_X1 U10403 ( .A1(n9109), .A2(n9060), .B1(n9108), .B2(n9071), .ZN(n9019)
         );
  NAND2_X1 U10404 ( .A1(n9017), .A2(n9016), .ZN(n9110) );
  MUX2_X1 U10405 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9110), .S(n9996), .Z(n9018) );
  OR2_X1 U10406 ( .A1(n9019), .A2(n9018), .ZN(P2_U3547) );
  INV_X1 U10407 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9022) );
  NOR2_X1 U10408 ( .A1(n9021), .A2(n9020), .ZN(n9113) );
  MUX2_X1 U10409 ( .A(n9022), .B(n9113), .S(n9996), .Z(n9024) );
  NAND2_X1 U10410 ( .A1(n9115), .A2(n9081), .ZN(n9023) );
  OAI211_X1 U10411 ( .C1(n9118), .C2(n9060), .A(n9024), .B(n9023), .ZN(
        P2_U3546) );
  INV_X1 U10412 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9028) );
  AOI211_X1 U10413 ( .C1(n9093), .C2(n9027), .A(n9026), .B(n9025), .ZN(n9119)
         );
  MUX2_X1 U10414 ( .A(n9028), .B(n9119), .S(n9996), .Z(n9029) );
  OAI21_X1 U10415 ( .B1(n9122), .B2(n9060), .A(n9029), .ZN(P2_U3545) );
  OAI22_X1 U10416 ( .A1(n9124), .A2(n9060), .B1(n9123), .B2(n9071), .ZN(n9033)
         );
  NAND2_X1 U10417 ( .A1(n9031), .A2(n9030), .ZN(n9125) );
  MUX2_X1 U10418 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9125), .S(n9996), .Z(n9032) );
  OR2_X1 U10419 ( .A1(n9033), .A2(n9032), .ZN(P2_U3544) );
  NAND3_X1 U10420 ( .A1(n9035), .A2(n9034), .A3(n9985), .ZN(n9040) );
  NAND2_X1 U10421 ( .A1(n9036), .A2(n9093), .ZN(n9037) );
  NAND4_X1 U10422 ( .A1(n9040), .A2(n9039), .A3(n9038), .A4(n9037), .ZN(n9128)
         );
  MUX2_X1 U10423 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9128), .S(n9996), .Z(
        P2_U3543) );
  NAND2_X1 U10424 ( .A1(n9042), .A2(n9041), .ZN(n9129) );
  MUX2_X1 U10425 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9129), .S(n9996), .Z(n9043) );
  AOI21_X1 U10426 ( .B1(n9081), .B2(n9131), .A(n9043), .ZN(n9044) );
  OAI21_X1 U10427 ( .B1(n9133), .B2(n9060), .A(n9044), .ZN(P2_U3542) );
  OAI22_X1 U10428 ( .A1(n9135), .A2(n9060), .B1(n9134), .B2(n9071), .ZN(n9048)
         );
  NAND2_X1 U10429 ( .A1(n9046), .A2(n9045), .ZN(n9136) );
  MUX2_X1 U10430 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9136), .S(n9996), .Z(n9047) );
  OR2_X1 U10431 ( .A1(n9048), .A2(n9047), .ZN(P2_U3541) );
  AOI22_X1 U10432 ( .A1(n9050), .A2(n9959), .B1(n9093), .B2(n9049), .ZN(n9051)
         );
  OAI211_X1 U10433 ( .C1(n9053), .C2(n9090), .A(n9052), .B(n9051), .ZN(n9139)
         );
  MUX2_X1 U10434 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9139), .S(n9996), .Z(
        P2_U3540) );
  INV_X1 U10435 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9057) );
  INV_X1 U10436 ( .A(n9054), .ZN(n9056) );
  NOR2_X1 U10437 ( .A1(n9056), .A2(n9055), .ZN(n9140) );
  MUX2_X1 U10438 ( .A(n9057), .B(n9140), .S(n9996), .Z(n9059) );
  NAND2_X1 U10439 ( .A1(n9143), .A2(n9081), .ZN(n9058) );
  OAI211_X1 U10440 ( .C1(n9147), .C2(n9060), .A(n9059), .B(n9058), .ZN(
        P2_U3539) );
  AOI22_X1 U10441 ( .A1(n9062), .A2(n9959), .B1(n9093), .B2(n9061), .ZN(n9063)
         );
  OAI211_X1 U10442 ( .C1(n9065), .C2(n9090), .A(n9064), .B(n9063), .ZN(n9148)
         );
  MUX2_X1 U10443 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9148), .S(n9996), .Z(
        P2_U3538) );
  AOI211_X1 U10444 ( .C1(n9068), .C2(n9985), .A(n9067), .B(n9066), .ZN(n9149)
         );
  MUX2_X1 U10445 ( .A(n9069), .B(n9149), .S(n9996), .Z(n9070) );
  OAI21_X1 U10446 ( .B1(n5829), .B2(n9071), .A(n9070), .ZN(P2_U3537) );
  OAI21_X1 U10447 ( .B1(n9073), .B2(n9979), .A(n9072), .ZN(n9074) );
  AOI21_X1 U10448 ( .B1(n9075), .B2(n9978), .A(n9074), .ZN(n9077) );
  NAND2_X1 U10449 ( .A1(n9077), .A2(n9076), .ZN(n9153) );
  MUX2_X1 U10450 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9153), .S(n9996), .Z(
        P2_U3536) );
  MUX2_X1 U10451 ( .A(n9079), .B(n9078), .S(n9996), .Z(n9085) );
  AOI22_X1 U10452 ( .A1(n9083), .A2(n9082), .B1(n9081), .B2(n9080), .ZN(n9084)
         );
  NAND2_X1 U10453 ( .A1(n9085), .A2(n9084), .ZN(P2_U3535) );
  AOI21_X1 U10454 ( .B1(n9093), .B2(n9087), .A(n9086), .ZN(n9088) );
  OAI211_X1 U10455 ( .C1(n9091), .C2(n9090), .A(n9089), .B(n9088), .ZN(n9154)
         );
  MUX2_X1 U10456 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9154), .S(n9996), .Z(
        P2_U3534) );
  AOI22_X1 U10457 ( .A1(n9094), .A2(n9959), .B1(n9093), .B2(n9092), .ZN(n9095)
         );
  OAI21_X1 U10458 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9098) );
  OR2_X1 U10459 ( .A1(n9099), .A2(n9098), .ZN(n9156) );
  MUX2_X1 U10460 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9156), .S(n9996), .Z(
        P2_U3533) );
  INV_X1 U10461 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U10462 ( .A(n9101), .B(n9100), .S(n9155), .Z(n9102) );
  OAI21_X1 U10463 ( .B1(n9103), .B2(n9152), .A(n9102), .ZN(P2_U3519) );
  INV_X1 U10464 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9105) );
  MUX2_X1 U10465 ( .A(n9105), .B(n9104), .S(n9155), .Z(n9106) );
  OAI21_X1 U10466 ( .B1(n9107), .B2(n9152), .A(n9106), .ZN(P2_U3518) );
  OAI22_X1 U10467 ( .A1(n9109), .A2(n9146), .B1(n9108), .B2(n9152), .ZN(n9112)
         );
  MUX2_X1 U10468 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9110), .S(n9155), .Z(n9111) );
  OR2_X1 U10469 ( .A1(n9112), .A2(n9111), .ZN(P2_U3515) );
  INV_X1 U10470 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9114) );
  MUX2_X1 U10471 ( .A(n9114), .B(n9113), .S(n9155), .Z(n9117) );
  NAND2_X1 U10472 ( .A1(n9115), .A2(n9142), .ZN(n9116) );
  OAI211_X1 U10473 ( .C1(n9118), .C2(n9146), .A(n9117), .B(n9116), .ZN(
        P2_U3514) );
  INV_X1 U10474 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9120) );
  MUX2_X1 U10475 ( .A(n9120), .B(n9119), .S(n9155), .Z(n9121) );
  OAI21_X1 U10476 ( .B1(n9122), .B2(n9146), .A(n9121), .ZN(P2_U3513) );
  OAI22_X1 U10477 ( .A1(n9124), .A2(n9146), .B1(n9123), .B2(n9152), .ZN(n9127)
         );
  MUX2_X1 U10478 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9125), .S(n9155), .Z(n9126) );
  OR2_X1 U10479 ( .A1(n9127), .A2(n9126), .ZN(P2_U3512) );
  MUX2_X1 U10480 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9128), .S(n9155), .Z(
        P2_U3511) );
  MUX2_X1 U10481 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9129), .S(n9155), .Z(n9130) );
  AOI21_X1 U10482 ( .B1(n9142), .B2(n9131), .A(n9130), .ZN(n9132) );
  OAI21_X1 U10483 ( .B1(n9133), .B2(n9146), .A(n9132), .ZN(P2_U3510) );
  OAI22_X1 U10484 ( .A1(n9135), .A2(n9146), .B1(n9134), .B2(n9152), .ZN(n9138)
         );
  MUX2_X1 U10485 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9136), .S(n9155), .Z(n9137) );
  OR2_X1 U10486 ( .A1(n9138), .A2(n9137), .ZN(P2_U3509) );
  MUX2_X1 U10487 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9139), .S(n9155), .Z(
        P2_U3508) );
  INV_X1 U10488 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U10489 ( .A(n9141), .B(n9140), .S(n9155), .Z(n9145) );
  NAND2_X1 U10490 ( .A1(n9143), .A2(n9142), .ZN(n9144) );
  OAI211_X1 U10491 ( .C1(n9147), .C2(n9146), .A(n9145), .B(n9144), .ZN(
        P2_U3507) );
  MUX2_X1 U10492 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9148), .S(n9155), .Z(
        P2_U3505) );
  INV_X1 U10493 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9150) );
  MUX2_X1 U10494 ( .A(n9150), .B(n9149), .S(n9155), .Z(n9151) );
  OAI21_X1 U10495 ( .B1(n5829), .B2(n9152), .A(n9151), .ZN(P2_U3502) );
  MUX2_X1 U10496 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9153), .S(n9155), .Z(
        P2_U3499) );
  MUX2_X1 U10497 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9154), .S(n9155), .Z(
        P2_U3493) );
  MUX2_X1 U10498 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9156), .S(n9155), .Z(
        P2_U3490) );
  INV_X1 U10499 ( .A(n6343), .ZN(n9645) );
  NOR4_X1 U10500 ( .A1(n5013), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9157), .A4(
        n4420), .ZN(n9158) );
  AOI21_X1 U10501 ( .B1(n9165), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9158), .ZN(
        n9159) );
  OAI21_X1 U10502 ( .B1(n9645), .B2(n9163), .A(n9159), .ZN(P2_U3327) );
  INV_X1 U10503 ( .A(n9160), .ZN(n9648) );
  AOI22_X1 U10504 ( .A1(n9161), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9165), .ZN(n9162) );
  OAI21_X1 U10505 ( .B1(n9648), .B2(n9163), .A(n9162), .ZN(P2_U3328) );
  INV_X1 U10506 ( .A(n9164), .ZN(n9652) );
  AOI22_X1 U10507 ( .A1(n9166), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9165), .ZN(n9167) );
  OAI21_X1 U10508 ( .B1(n9652), .B2(n9163), .A(n9167), .ZN(P2_U3329) );
  INV_X1 U10509 ( .A(n9168), .ZN(n9169) );
  MUX2_X1 U10510 ( .A(n9169), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10511 ( .A1(n9170), .A2(n6688), .ZN(n9171) );
  XOR2_X1 U10512 ( .A(n9172), .B(n9171), .Z(n9181) );
  NOR2_X1 U10513 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9173), .ZN(n9806) );
  AOI21_X1 U10514 ( .B1(n9266), .B2(n9313), .A(n9806), .ZN(n9176) );
  NAND2_X1 U10515 ( .A1(n9306), .A2(n9174), .ZN(n9175) );
  OAI211_X1 U10516 ( .C1(n9177), .C2(n9234), .A(n9176), .B(n9175), .ZN(n9178)
         );
  AOI21_X1 U10517 ( .B1(n9179), .B2(n9291), .A(n9178), .ZN(n9180) );
  OAI21_X1 U10518 ( .B1(n9181), .B2(n9309), .A(n9180), .ZN(P1_U3213) );
  NAND2_X1 U10519 ( .A1(n4470), .A2(n9182), .ZN(n9184) );
  XNOR2_X1 U10520 ( .A(n9184), .B(n9183), .ZN(n9190) );
  INV_X1 U10521 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9185) );
  OAI22_X1 U10522 ( .A1(n9301), .A2(n8490), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9185), .ZN(n9186) );
  AOI21_X1 U10523 ( .B1(n9298), .B2(n9462), .A(n9186), .ZN(n9187) );
  OAI21_X1 U10524 ( .B1(n9281), .B2(n9427), .A(n9187), .ZN(n9188) );
  AOI21_X1 U10525 ( .B1(n9581), .B2(n9291), .A(n9188), .ZN(n9189) );
  OAI21_X1 U10526 ( .B1(n9190), .B2(n9309), .A(n9189), .ZN(P1_U3214) );
  XOR2_X1 U10527 ( .A(n9191), .B(n9192), .Z(n9199) );
  OAI21_X1 U10528 ( .B1(n9194), .B2(n9301), .A(n9193), .ZN(n9195) );
  AOI21_X1 U10529 ( .B1(n9298), .B2(n9540), .A(n9195), .ZN(n9196) );
  OAI21_X1 U10530 ( .B1(n9281), .B2(n9497), .A(n9196), .ZN(n9197) );
  AOI21_X1 U10531 ( .B1(n9600), .B2(n9291), .A(n9197), .ZN(n9198) );
  OAI21_X1 U10532 ( .B1(n9199), .B2(n9309), .A(n9198), .ZN(P1_U3217) );
  XNOR2_X1 U10533 ( .A(n9201), .B(n9200), .ZN(n9202) );
  NAND2_X1 U10534 ( .A1(n9202), .A2(n9264), .ZN(n9207) );
  OAI22_X1 U10535 ( .A1(n9301), .A2(n9361), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9203), .ZN(n9205) );
  NOR2_X1 U10536 ( .A1(n9234), .A2(n8490), .ZN(n9204) );
  AOI211_X1 U10537 ( .C1(n9394), .C2(n9306), .A(n9205), .B(n9204), .ZN(n9206)
         );
  OAI211_X1 U10538 ( .C1(n9396), .C2(n9303), .A(n9207), .B(n9206), .ZN(
        P1_U3223) );
  INV_X1 U10539 ( .A(n9209), .ZN(n9211) );
  NOR2_X1 U10540 ( .A1(n9211), .A2(n9210), .ZN(n9212) );
  XNOR2_X1 U10541 ( .A(n9208), .B(n9212), .ZN(n9219) );
  AOI22_X1 U10542 ( .A1(n9298), .A2(n9313), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n9215) );
  NAND2_X1 U10543 ( .A1(n9306), .A2(n9213), .ZN(n9214) );
  OAI211_X1 U10544 ( .C1(n9216), .C2(n9301), .A(n9215), .B(n9214), .ZN(n9217)
         );
  AOI21_X1 U10545 ( .B1(n9617), .B2(n9291), .A(n9217), .ZN(n9218) );
  OAI21_X1 U10546 ( .B1(n9219), .B2(n9309), .A(n9218), .ZN(P1_U3224) );
  NAND2_X1 U10547 ( .A1(n4512), .A2(n9220), .ZN(n9221) );
  XNOR2_X1 U10548 ( .A(n9222), .B(n9221), .ZN(n9228) );
  NAND2_X1 U10549 ( .A1(n9298), .A2(n9538), .ZN(n9223) );
  NAND2_X1 U10550 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9329) );
  OAI211_X1 U10551 ( .C1(n9224), .C2(n9301), .A(n9223), .B(n9329), .ZN(n9226)
         );
  NOR2_X1 U10552 ( .A1(n9534), .A2(n9303), .ZN(n9225) );
  AOI211_X1 U10553 ( .C1(n9531), .C2(n9306), .A(n9226), .B(n9225), .ZN(n9227)
         );
  OAI21_X1 U10554 ( .B1(n9228), .B2(n9309), .A(n9227), .ZN(P1_U3226) );
  AOI21_X1 U10555 ( .B1(n9231), .B2(n9230), .A(n9229), .ZN(n9240) );
  OAI22_X1 U10556 ( .A1(n9301), .A2(n9233), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9232), .ZN(n9236) );
  NOR2_X1 U10557 ( .A1(n9234), .A2(n9256), .ZN(n9235) );
  AOI211_X1 U10558 ( .C1(n9418), .C2(n9306), .A(n9236), .B(n9235), .ZN(n9239)
         );
  NAND2_X1 U10559 ( .A1(n9406), .A2(n9872), .ZN(n9576) );
  OR2_X1 U10560 ( .A1(n9576), .A2(n9237), .ZN(n9238) );
  OAI211_X1 U10561 ( .C1(n9240), .C2(n9309), .A(n9239), .B(n9238), .ZN(
        P1_U3227) );
  XNOR2_X1 U10562 ( .A(n9243), .B(n9242), .ZN(n9244) );
  XNOR2_X1 U10563 ( .A(n9241), .B(n9244), .ZN(n9249) );
  AOI22_X1 U10564 ( .A1(n9488), .A2(n9266), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9246) );
  NAND2_X1 U10565 ( .A1(n9298), .A2(n9521), .ZN(n9245) );
  OAI211_X1 U10566 ( .C1(n9281), .C2(n9490), .A(n9246), .B(n9245), .ZN(n9247)
         );
  AOI21_X1 U10567 ( .B1(n9595), .B2(n9291), .A(n9247), .ZN(n9248) );
  OAI21_X1 U10568 ( .B1(n9249), .B2(n9309), .A(n9248), .ZN(P1_U3231) );
  NAND2_X1 U10569 ( .A1(n9251), .A2(n9250), .ZN(n9252) );
  XOR2_X1 U10570 ( .A(n9253), .B(n9252), .Z(n9259) );
  AOI22_X1 U10571 ( .A1(n9488), .A2(n9298), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9255) );
  NAND2_X1 U10572 ( .A1(n9306), .A2(n9446), .ZN(n9254) );
  OAI211_X1 U10573 ( .C1(n9256), .C2(n9301), .A(n9255), .B(n9254), .ZN(n9257)
         );
  AOI21_X1 U10574 ( .B1(n9586), .B2(n9291), .A(n9257), .ZN(n9258) );
  OAI21_X1 U10575 ( .B1(n9259), .B2(n9309), .A(n9258), .ZN(P1_U3233) );
  OAI21_X1 U10576 ( .B1(n9263), .B2(n9260), .A(n9261), .ZN(n9265) );
  NAND2_X1 U10577 ( .A1(n9265), .A2(n9264), .ZN(n9273) );
  AOI22_X1 U10578 ( .A1(n9266), .A2(n9323), .B1(n9298), .B2(n6564), .ZN(n9272)
         );
  INV_X1 U10579 ( .A(n9269), .ZN(n9268) );
  NAND2_X1 U10580 ( .A1(n9268), .A2(n9267), .ZN(n9271) );
  NAND2_X1 U10581 ( .A1(n9269), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9270) );
  NAND4_X1 U10582 ( .A1(n9273), .A2(n9272), .A3(n9271), .A4(n9270), .ZN(
        P1_U3235) );
  NAND2_X1 U10583 ( .A1(n9274), .A2(n9275), .ZN(n9277) );
  XNOR2_X1 U10584 ( .A(n9277), .B(n9276), .ZN(n9284) );
  NAND2_X1 U10585 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9826) );
  OAI21_X1 U10586 ( .B1(n9278), .B2(n9301), .A(n9826), .ZN(n9279) );
  AOI21_X1 U10587 ( .B1(n9298), .B2(n9522), .A(n9279), .ZN(n9280) );
  OAI21_X1 U10588 ( .B1(n9281), .B2(n9513), .A(n9280), .ZN(n9282) );
  AOI21_X1 U10589 ( .B1(n9605), .B2(n9291), .A(n9282), .ZN(n9283) );
  OAI21_X1 U10590 ( .B1(n9284), .B2(n9309), .A(n9283), .ZN(P1_U3236) );
  NAND2_X1 U10591 ( .A1(n4493), .A2(n9285), .ZN(n9286) );
  XNOR2_X1 U10592 ( .A(n9287), .B(n9286), .ZN(n9293) );
  AOI22_X1 U10593 ( .A1(n9298), .A2(n9414), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9289) );
  NAND2_X1 U10594 ( .A1(n9306), .A2(n9377), .ZN(n9288) );
  OAI211_X1 U10595 ( .C1(n9381), .C2(n9301), .A(n9289), .B(n9288), .ZN(n9290)
         );
  AOI21_X1 U10596 ( .B1(n9565), .B2(n9291), .A(n9290), .ZN(n9292) );
  OAI21_X1 U10597 ( .B1(n9293), .B2(n9309), .A(n9292), .ZN(P1_U3238) );
  NAND2_X1 U10598 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  XOR2_X1 U10599 ( .A(n9297), .B(n9296), .Z(n9310) );
  NAND2_X1 U10600 ( .A1(n9298), .A2(n9314), .ZN(n9300) );
  OAI211_X1 U10601 ( .C1(n9302), .C2(n9301), .A(n9300), .B(n9299), .ZN(n9305)
         );
  NOR2_X1 U10602 ( .A1(n9621), .A2(n9303), .ZN(n9304) );
  AOI211_X1 U10603 ( .C1(n9307), .C2(n9306), .A(n9305), .B(n9304), .ZN(n9308)
         );
  OAI21_X1 U10604 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(P1_U3239) );
  MUX2_X1 U10605 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9311), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10606 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9312), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9354), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10608 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9367), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10609 ( .A(n9353), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9324), .Z(
        P1_U3582) );
  MUX2_X1 U10610 ( .A(n9399), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9324), .Z(
        P1_U3581) );
  MUX2_X1 U10611 ( .A(n9414), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9324), .Z(
        P1_U3580) );
  MUX2_X1 U10612 ( .A(n9439), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9324), .Z(
        P1_U3579) );
  MUX2_X1 U10613 ( .A(n9452), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9324), .Z(
        P1_U3578) );
  MUX2_X1 U10614 ( .A(n9462), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9324), .Z(
        P1_U3577) );
  MUX2_X1 U10615 ( .A(n9504), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9324), .Z(
        P1_U3575) );
  MUX2_X1 U10616 ( .A(n9521), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9324), .Z(
        P1_U3574) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9540), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10618 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9522), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10619 ( .A(n9538), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9324), .Z(
        P1_U3571) );
  MUX2_X1 U10620 ( .A(n9313), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9324), .Z(
        P1_U3570) );
  MUX2_X1 U10621 ( .A(n9314), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9324), .Z(
        P1_U3569) );
  MUX2_X1 U10622 ( .A(n9315), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9324), .Z(
        P1_U3568) );
  MUX2_X1 U10623 ( .A(n9316), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9324), .Z(
        P1_U3567) );
  MUX2_X1 U10624 ( .A(n9317), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9324), .Z(
        P1_U3566) );
  MUX2_X1 U10625 ( .A(n9318), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9324), .Z(
        P1_U3563) );
  MUX2_X1 U10626 ( .A(n9319), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9324), .Z(
        P1_U3562) );
  MUX2_X1 U10627 ( .A(n9320), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9324), .Z(
        P1_U3561) );
  MUX2_X1 U10628 ( .A(n9321), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9324), .Z(
        P1_U3560) );
  MUX2_X1 U10629 ( .A(n9322), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9324), .Z(
        P1_U3559) );
  MUX2_X1 U10630 ( .A(n9323), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9324), .Z(
        P1_U3558) );
  MUX2_X1 U10631 ( .A(n6573), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9324), .Z(
        P1_U3557) );
  MUX2_X1 U10632 ( .A(n6564), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9324), .Z(
        P1_U3556) );
  MUX2_X1 U10633 ( .A(n9325), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9324), .Z(
        P1_U3555) );
  INV_X1 U10634 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9331) );
  OAI211_X1 U10635 ( .C1(n9328), .C2(n9327), .A(n9816), .B(n9326), .ZN(n9330)
         );
  OAI211_X1 U10636 ( .C1(n9821), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9332)
         );
  INV_X1 U10637 ( .A(n9332), .ZN(n9337) );
  OAI211_X1 U10638 ( .C1(n9335), .C2(n9334), .A(n9823), .B(n9333), .ZN(n9336)
         );
  OAI211_X1 U10639 ( .C1(n9828), .C2(n9338), .A(n9337), .B(n9336), .ZN(
        P1_U3258) );
  XNOR2_X1 U10640 ( .A(n9340), .B(n9339), .ZN(n9681) );
  NAND2_X1 U10641 ( .A1(n9681), .A2(n9545), .ZN(n9343) );
  AOI21_X1 U10642 ( .B1(n4421), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9341), .ZN(
        n9342) );
  OAI211_X1 U10643 ( .C1(n9679), .C2(n9533), .A(n9343), .B(n9342), .ZN(
        P1_U3262) );
  OAI21_X1 U10644 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(n9559) );
  AOI21_X1 U10645 ( .B1(n9555), .B2(n9368), .A(n9347), .ZN(n9556) );
  AOI22_X1 U10646 ( .A1(n4421), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9348), .B2(
        n9530), .ZN(n9349) );
  OAI21_X1 U10647 ( .B1(n4615), .B2(n9533), .A(n9349), .ZN(n9357) );
  OAI21_X1 U10648 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9355) );
  AOI222_X1 U10649 ( .A1(n9542), .A2(n9355), .B1(n9354), .B2(n9539), .C1(n9353), .C2(n9537), .ZN(n9558) );
  NOR2_X1 U10650 ( .A1(n9558), .A2(n7466), .ZN(n9356) );
  AOI211_X1 U10651 ( .C1(n9556), .C2(n9545), .A(n9357), .B(n9356), .ZN(n9358)
         );
  OAI21_X1 U10652 ( .B1(n9559), .B2(n9547), .A(n9358), .ZN(P1_U3263) );
  XOR2_X1 U10653 ( .A(n9363), .B(n9359), .Z(n9564) );
  NOR2_X1 U10654 ( .A1(n9360), .A2(n9533), .ZN(n9373) );
  NOR2_X1 U10655 ( .A1(n9361), .A2(n9431), .ZN(n9366) );
  AOI211_X1 U10656 ( .C1(n9364), .C2(n9363), .A(n9484), .B(n9362), .ZN(n9365)
         );
  INV_X1 U10657 ( .A(n9368), .ZN(n9369) );
  AOI211_X1 U10658 ( .C1(n9561), .C2(n4619), .A(n9883), .B(n9369), .ZN(n9560)
         );
  AOI22_X1 U10659 ( .A1(n9560), .A2(n6482), .B1(n9530), .B2(n9370), .ZN(n9371)
         );
  AOI21_X1 U10660 ( .B1(n9563), .B2(n9371), .A(n4421), .ZN(n9372) );
  AOI211_X1 U10661 ( .C1(n7466), .C2(P1_REG2_REG_27__SCAN_IN), .A(n9373), .B(
        n9372), .ZN(n9374) );
  OAI21_X1 U10662 ( .B1(n9564), .B2(n9547), .A(n9374), .ZN(P1_U3264) );
  XNOR2_X1 U10663 ( .A(n9375), .B(n9384), .ZN(n9569) );
  AOI21_X1 U10664 ( .B1(n9565), .B2(n9391), .A(n9376), .ZN(n9566) );
  AOI22_X1 U10665 ( .A1(n4421), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9377), .B2(
        n9530), .ZN(n9378) );
  OAI21_X1 U10666 ( .B1(n9379), .B2(n9533), .A(n9378), .ZN(n9388) );
  NOR2_X1 U10667 ( .A1(n9381), .A2(n9380), .ZN(n9386) );
  AOI211_X1 U10668 ( .C1(n9384), .C2(n9383), .A(n9484), .B(n9382), .ZN(n9385)
         );
  AOI211_X1 U10669 ( .C1(n9537), .C2(n9414), .A(n9386), .B(n9385), .ZN(n9568)
         );
  NOR2_X1 U10670 ( .A1(n9568), .A2(n4421), .ZN(n9387) );
  AOI211_X1 U10671 ( .C1(n9566), .C2(n9545), .A(n9388), .B(n9387), .ZN(n9389)
         );
  OAI21_X1 U10672 ( .B1(n9569), .B2(n9547), .A(n9389), .ZN(P1_U3265) );
  XOR2_X1 U10673 ( .A(n9397), .B(n9390), .Z(n9574) );
  INV_X1 U10674 ( .A(n9409), .ZN(n9393) );
  INV_X1 U10675 ( .A(n9391), .ZN(n9392) );
  AOI21_X1 U10676 ( .B1(n9570), .B2(n9393), .A(n9392), .ZN(n9571) );
  AOI22_X1 U10677 ( .A1(n4421), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9394), .B2(
        n9530), .ZN(n9395) );
  OAI21_X1 U10678 ( .B1(n9396), .B2(n9533), .A(n9395), .ZN(n9402) );
  XNOR2_X1 U10679 ( .A(n9398), .B(n9397), .ZN(n9400) );
  AOI222_X1 U10680 ( .A1(n9542), .A2(n9400), .B1(n9399), .B2(n9539), .C1(n9439), .C2(n9537), .ZN(n9573) );
  NOR2_X1 U10681 ( .A1(n9573), .A2(n7466), .ZN(n9401) );
  AOI211_X1 U10682 ( .C1(n9571), .C2(n9545), .A(n9402), .B(n9401), .ZN(n9403)
         );
  OAI21_X1 U10683 ( .B1(n9574), .B2(n9547), .A(n9403), .ZN(P1_U3266) );
  XOR2_X1 U10684 ( .A(n9411), .B(n9404), .Z(n9579) );
  AOI22_X1 U10685 ( .A1(n9406), .A2(n9405), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4421), .ZN(n9423) );
  NAND2_X1 U10686 ( .A1(n9426), .A2(n9406), .ZN(n9407) );
  NAND2_X1 U10687 ( .A1(n9407), .A2(n9873), .ZN(n9408) );
  OR2_X1 U10688 ( .A1(n9409), .A2(n9408), .ZN(n9575) );
  NAND2_X1 U10689 ( .A1(n9433), .A2(n9410), .ZN(n9412) );
  XNOR2_X1 U10690 ( .A(n9412), .B(n9411), .ZN(n9413) );
  NAND2_X1 U10691 ( .A1(n9413), .A2(n9542), .ZN(n9578) );
  NAND2_X1 U10692 ( .A1(n9537), .A2(n9452), .ZN(n9416) );
  NAND2_X1 U10693 ( .A1(n9539), .A2(n9414), .ZN(n9415) );
  AND2_X1 U10694 ( .A1(n9416), .A2(n9415), .ZN(n9577) );
  INV_X1 U10695 ( .A(n9577), .ZN(n9417) );
  AOI21_X1 U10696 ( .B1(n9418), .B2(n9530), .A(n9417), .ZN(n9419) );
  OAI211_X1 U10697 ( .C1(n9420), .C2(n9575), .A(n9578), .B(n9419), .ZN(n9421)
         );
  NAND2_X1 U10698 ( .A1(n9421), .A2(n9477), .ZN(n9422) );
  OAI211_X1 U10699 ( .C1(n9579), .C2(n9547), .A(n9423), .B(n9422), .ZN(
        P1_U3267) );
  XNOR2_X1 U10700 ( .A(n9424), .B(n9425), .ZN(n9584) );
  AOI211_X1 U10701 ( .C1(n9581), .C2(n9444), .A(n9883), .B(n4629), .ZN(n9580)
         );
  INV_X1 U10702 ( .A(n9427), .ZN(n9428) );
  AOI22_X1 U10703 ( .A1(n4421), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9428), .B2(
        n9530), .ZN(n9429) );
  OAI21_X1 U10704 ( .B1(n9430), .B2(n9533), .A(n9429), .ZN(n9441) );
  NOR2_X1 U10705 ( .A1(n9432), .A2(n9431), .ZN(n9438) );
  INV_X1 U10706 ( .A(n9433), .ZN(n9434) );
  AOI211_X1 U10707 ( .C1(n9436), .C2(n9435), .A(n9484), .B(n9434), .ZN(n9437)
         );
  AOI211_X1 U10708 ( .C1(n9539), .C2(n9439), .A(n9438), .B(n9437), .ZN(n9583)
         );
  NOR2_X1 U10709 ( .A1(n9583), .A2(n4421), .ZN(n9440) );
  AOI211_X1 U10710 ( .C1(n9580), .C2(n9467), .A(n9441), .B(n9440), .ZN(n9442)
         );
  OAI21_X1 U10711 ( .B1(n9584), .B2(n9547), .A(n9442), .ZN(P1_U3268) );
  XNOR2_X1 U10712 ( .A(n9443), .B(n9451), .ZN(n9589) );
  INV_X1 U10713 ( .A(n9465), .ZN(n9445) );
  AOI211_X1 U10714 ( .C1(n9586), .C2(n9445), .A(n9883), .B(n4630), .ZN(n9585)
         );
  AOI22_X1 U10715 ( .A1(n4421), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9446), .B2(
        n9530), .ZN(n9447) );
  OAI21_X1 U10716 ( .B1(n9448), .B2(n9533), .A(n9447), .ZN(n9455) );
  OAI21_X1 U10717 ( .B1(n9451), .B2(n9450), .A(n9449), .ZN(n9453) );
  AOI222_X1 U10718 ( .A1(n9542), .A2(n9453), .B1(n9452), .B2(n9539), .C1(n9488), .C2(n9537), .ZN(n9588) );
  NOR2_X1 U10719 ( .A1(n9588), .A2(n7466), .ZN(n9454) );
  AOI211_X1 U10720 ( .C1(n9585), .C2(n9467), .A(n9455), .B(n9454), .ZN(n9456)
         );
  OAI21_X1 U10721 ( .B1(n9589), .B2(n9547), .A(n9456), .ZN(P1_U3269) );
  XNOR2_X1 U10722 ( .A(n9458), .B(n9457), .ZN(n9594) );
  OAI211_X1 U10723 ( .C1(n9461), .C2(n9460), .A(n9459), .B(n9542), .ZN(n9464)
         );
  AOI22_X1 U10724 ( .A1(n9504), .A2(n9537), .B1(n9539), .B2(n9462), .ZN(n9463)
         );
  NAND2_X1 U10725 ( .A1(n9464), .A2(n9463), .ZN(n9590) );
  INV_X1 U10726 ( .A(n9476), .ZN(n9466) );
  AOI211_X1 U10727 ( .C1(n9592), .C2(n9466), .A(n9883), .B(n9465), .ZN(n9591)
         );
  NAND2_X1 U10728 ( .A1(n9591), .A2(n9467), .ZN(n9470) );
  AOI22_X1 U10729 ( .A1(n4421), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9468), .B2(
        n9530), .ZN(n9469) );
  OAI211_X1 U10730 ( .C1(n9471), .C2(n9533), .A(n9470), .B(n9469), .ZN(n9472)
         );
  AOI21_X1 U10731 ( .B1(n9477), .B2(n9590), .A(n9472), .ZN(n9473) );
  OAI21_X1 U10732 ( .B1(n9594), .B2(n9547), .A(n9473), .ZN(P1_U3270) );
  XNOR2_X1 U10733 ( .A(n9474), .B(n9485), .ZN(n9599) );
  AND2_X1 U10734 ( .A1(n9495), .A2(n9595), .ZN(n9475) );
  NOR2_X1 U10735 ( .A1(n9476), .A2(n9475), .ZN(n9596) );
  INV_X1 U10736 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9478) );
  OAI22_X1 U10737 ( .A1(n9479), .A2(n9533), .B1(n9478), .B2(n9477), .ZN(n9480)
         );
  AOI21_X1 U10738 ( .B1(n9596), .B2(n9545), .A(n9480), .ZN(n9493) );
  AND2_X1 U10739 ( .A1(n9521), .A2(n9537), .ZN(n9487) );
  INV_X1 U10740 ( .A(n9482), .ZN(n9483) );
  AOI211_X1 U10741 ( .C1(n9485), .C2(n9481), .A(n9484), .B(n9483), .ZN(n9486)
         );
  AOI211_X1 U10742 ( .C1(n9539), .C2(n9488), .A(n9487), .B(n9486), .ZN(n9598)
         );
  OAI21_X1 U10743 ( .B1(n9490), .B2(n9489), .A(n9598), .ZN(n9491) );
  NAND2_X1 U10744 ( .A1(n9491), .A2(n9477), .ZN(n9492) );
  OAI211_X1 U10745 ( .C1(n9599), .C2(n9547), .A(n9493), .B(n9492), .ZN(
        P1_U3271) );
  XNOR2_X1 U10746 ( .A(n9494), .B(n9503), .ZN(n9604) );
  INV_X1 U10747 ( .A(n9495), .ZN(n9496) );
  AOI21_X1 U10748 ( .B1(n9600), .B2(n9510), .A(n9496), .ZN(n9601) );
  INV_X1 U10749 ( .A(n9497), .ZN(n9498) );
  AOI22_X1 U10750 ( .A1(n4421), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9498), .B2(
        n9530), .ZN(n9499) );
  OAI21_X1 U10751 ( .B1(n9500), .B2(n9533), .A(n9499), .ZN(n9507) );
  OAI21_X1 U10752 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9505) );
  AOI222_X1 U10753 ( .A1(n9542), .A2(n9505), .B1(n9540), .B2(n9537), .C1(n9504), .C2(n9539), .ZN(n9603) );
  NOR2_X1 U10754 ( .A1(n9603), .A2(n7466), .ZN(n9506) );
  AOI211_X1 U10755 ( .C1(n9601), .C2(n9545), .A(n9507), .B(n9506), .ZN(n9508)
         );
  OAI21_X1 U10756 ( .B1(n9604), .B2(n9547), .A(n9508), .ZN(P1_U3272) );
  XNOR2_X1 U10757 ( .A(n9509), .B(n9519), .ZN(n9609) );
  INV_X1 U10758 ( .A(n9528), .ZN(n9512) );
  INV_X1 U10759 ( .A(n9510), .ZN(n9511) );
  AOI21_X1 U10760 ( .B1(n9605), .B2(n9512), .A(n9511), .ZN(n9606) );
  INV_X1 U10761 ( .A(n9513), .ZN(n9514) );
  AOI22_X1 U10762 ( .A1(n4421), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9514), .B2(
        n9530), .ZN(n9515) );
  OAI21_X1 U10763 ( .B1(n9516), .B2(n9533), .A(n9515), .ZN(n9525) );
  INV_X1 U10764 ( .A(n9535), .ZN(n9518) );
  OAI21_X1 U10765 ( .B1(n9536), .B2(n9518), .A(n9517), .ZN(n9520) );
  XNOR2_X1 U10766 ( .A(n9520), .B(n9519), .ZN(n9523) );
  AOI222_X1 U10767 ( .A1(n9542), .A2(n9523), .B1(n9522), .B2(n9537), .C1(n9521), .C2(n9539), .ZN(n9608) );
  NOR2_X1 U10768 ( .A1(n9608), .A2(n7466), .ZN(n9524) );
  AOI211_X1 U10769 ( .C1(n9606), .C2(n9545), .A(n9525), .B(n9524), .ZN(n9526)
         );
  OAI21_X1 U10770 ( .B1(n9609), .B2(n9547), .A(n9526), .ZN(P1_U3273) );
  XNOR2_X1 U10771 ( .A(n9527), .B(n9535), .ZN(n9614) );
  AOI21_X1 U10772 ( .B1(n9610), .B2(n9529), .A(n9528), .ZN(n9611) );
  AOI22_X1 U10773 ( .A1(n4421), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9531), .B2(
        n9530), .ZN(n9532) );
  OAI21_X1 U10774 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9544) );
  XNOR2_X1 U10775 ( .A(n9536), .B(n9535), .ZN(n9541) );
  AOI222_X1 U10776 ( .A1(n9542), .A2(n9541), .B1(n9540), .B2(n9539), .C1(n9538), .C2(n9537), .ZN(n9613) );
  NOR2_X1 U10777 ( .A1(n9613), .A2(n7466), .ZN(n9543) );
  AOI211_X1 U10778 ( .C1(n9611), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9546)
         );
  OAI21_X1 U10779 ( .B1(n9614), .B2(n9547), .A(n9546), .ZN(P1_U3274) );
  NAND2_X1 U10780 ( .A1(n9548), .A2(n9873), .ZN(n9549) );
  OAI211_X1 U10781 ( .C1(n9550), .C2(n9881), .A(n9549), .B(n9678), .ZN(n9626)
         );
  MUX2_X1 U10782 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9626), .S(n9903), .Z(
        P1_U3554) );
  AOI22_X1 U10783 ( .A1(n9556), .A2(n9873), .B1(n9872), .B2(n9555), .ZN(n9557)
         );
  OAI211_X1 U10784 ( .C1(n9559), .C2(n9683), .A(n9558), .B(n9557), .ZN(n9627)
         );
  MUX2_X1 U10785 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9627), .S(n9903), .Z(
        P1_U3551) );
  AOI21_X1 U10786 ( .B1(n9872), .B2(n9561), .A(n9560), .ZN(n9562) );
  OAI211_X1 U10787 ( .C1(n9564), .C2(n9683), .A(n9563), .B(n9562), .ZN(n9628)
         );
  MUX2_X1 U10788 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9628), .S(n9903), .Z(
        P1_U3550) );
  AOI22_X1 U10789 ( .A1(n9566), .A2(n9873), .B1(n9872), .B2(n9565), .ZN(n9567)
         );
  OAI211_X1 U10790 ( .C1(n9569), .C2(n9683), .A(n9568), .B(n9567), .ZN(n9629)
         );
  MUX2_X1 U10791 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9629), .S(n9903), .Z(
        P1_U3549) );
  AOI22_X1 U10792 ( .A1(n9571), .A2(n9873), .B1(n9872), .B2(n9570), .ZN(n9572)
         );
  OAI211_X1 U10793 ( .C1(n9574), .C2(n9683), .A(n9573), .B(n9572), .ZN(n9630)
         );
  MUX2_X1 U10794 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9630), .S(n9903), .Z(
        P1_U3548) );
  OAI21_X1 U10795 ( .B1(n9579), .B2(n9683), .A(n4979), .ZN(n9631) );
  MUX2_X1 U10796 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9631), .S(n9903), .Z(
        P1_U3547) );
  AOI21_X1 U10797 ( .B1(n9872), .B2(n9581), .A(n9580), .ZN(n9582) );
  OAI211_X1 U10798 ( .C1(n9584), .C2(n9683), .A(n9583), .B(n9582), .ZN(n9632)
         );
  MUX2_X1 U10799 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9632), .S(n9903), .Z(
        P1_U3546) );
  AOI21_X1 U10800 ( .B1(n9872), .B2(n9586), .A(n9585), .ZN(n9587) );
  OAI211_X1 U10801 ( .C1(n9589), .C2(n9683), .A(n9588), .B(n9587), .ZN(n9633)
         );
  MUX2_X1 U10802 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9633), .S(n9903), .Z(
        P1_U3545) );
  AOI211_X1 U10803 ( .C1(n9872), .C2(n9592), .A(n9591), .B(n9590), .ZN(n9593)
         );
  OAI21_X1 U10804 ( .B1(n9594), .B2(n9683), .A(n9593), .ZN(n9634) );
  MUX2_X1 U10805 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9634), .S(n9903), .Z(
        P1_U3544) );
  AOI22_X1 U10806 ( .A1(n9596), .A2(n9873), .B1(n9872), .B2(n9595), .ZN(n9597)
         );
  OAI211_X1 U10807 ( .C1(n9599), .C2(n9683), .A(n9598), .B(n9597), .ZN(n9635)
         );
  MUX2_X1 U10808 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9635), .S(n9903), .Z(
        P1_U3543) );
  AOI22_X1 U10809 ( .A1(n9601), .A2(n9873), .B1(n9872), .B2(n9600), .ZN(n9602)
         );
  OAI211_X1 U10810 ( .C1(n9604), .C2(n9683), .A(n9603), .B(n9602), .ZN(n9636)
         );
  MUX2_X1 U10811 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9636), .S(n9903), .Z(
        P1_U3542) );
  AOI22_X1 U10812 ( .A1(n9606), .A2(n9873), .B1(n9872), .B2(n9605), .ZN(n9607)
         );
  OAI211_X1 U10813 ( .C1(n9609), .C2(n9683), .A(n9608), .B(n9607), .ZN(n9637)
         );
  MUX2_X1 U10814 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9637), .S(n9903), .Z(
        P1_U3541) );
  AOI22_X1 U10815 ( .A1(n9611), .A2(n9873), .B1(n9872), .B2(n9610), .ZN(n9612)
         );
  OAI211_X1 U10816 ( .C1(n9614), .C2(n9683), .A(n9613), .B(n9612), .ZN(n9638)
         );
  MUX2_X1 U10817 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9638), .S(n9903), .Z(
        P1_U3540) );
  AOI211_X1 U10818 ( .C1(n9872), .C2(n9617), .A(n9616), .B(n9615), .ZN(n9618)
         );
  OAI21_X1 U10819 ( .B1(n9619), .B2(n9683), .A(n9618), .ZN(n9639) );
  MUX2_X1 U10820 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9639), .S(n9903), .Z(
        P1_U3539) );
  INV_X1 U10821 ( .A(n9876), .ZN(n9693) );
  AND2_X1 U10822 ( .A1(n9620), .A2(n9693), .ZN(n9624) );
  OAI22_X1 U10823 ( .A1(n9622), .A2(n9883), .B1(n9621), .B2(n9881), .ZN(n9623)
         );
  MUX2_X1 U10824 ( .A(n9640), .B(P1_REG1_REG_15__SCAN_IN), .S(n9901), .Z(
        P1_U3538) );
  MUX2_X1 U10825 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9626), .S(n9891), .Z(
        P1_U3522) );
  MUX2_X1 U10826 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9627), .S(n9891), .Z(
        P1_U3519) );
  MUX2_X1 U10827 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9628), .S(n9891), .Z(
        P1_U3518) );
  MUX2_X1 U10828 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9629), .S(n9891), .Z(
        P1_U3517) );
  MUX2_X1 U10829 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9630), .S(n9891), .Z(
        P1_U3516) );
  MUX2_X1 U10830 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9631), .S(n9891), .Z(
        P1_U3515) );
  MUX2_X1 U10831 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9632), .S(n9891), .Z(
        P1_U3514) );
  MUX2_X1 U10832 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9633), .S(n9891), .Z(
        P1_U3513) );
  MUX2_X1 U10833 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9634), .S(n9891), .Z(
        P1_U3512) );
  MUX2_X1 U10834 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9635), .S(n9891), .Z(
        P1_U3511) );
  MUX2_X1 U10835 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9636), .S(n9891), .Z(
        P1_U3510) );
  MUX2_X1 U10836 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9637), .S(n9891), .Z(
        P1_U3508) );
  MUX2_X1 U10837 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9638), .S(n9891), .Z(
        P1_U3505) );
  MUX2_X1 U10838 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9639), .S(n9891), .Z(
        P1_U3502) );
  MUX2_X1 U10839 ( .A(n9640), .B(P1_REG0_REG_15__SCAN_IN), .S(n9889), .Z(
        P1_U3499) );
  INV_X1 U10840 ( .A(n9641), .ZN(n9642) );
  NOR4_X1 U10841 ( .A1(n9642), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n6127), .ZN(n9643) );
  AOI21_X1 U10842 ( .B1(n9649), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9643), .ZN(
        n9644) );
  OAI21_X1 U10843 ( .B1(n9645), .B2(n9651), .A(n9644), .ZN(P1_U3322) );
  AOI22_X1 U10844 ( .A1(n9646), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9649), .ZN(n9647) );
  OAI21_X1 U10845 ( .B1(n9648), .B2(n9651), .A(n9647), .ZN(P1_U3323) );
  AOI22_X1 U10846 ( .A1(n5941), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9649), .ZN(n9650) );
  OAI21_X1 U10847 ( .B1(n9652), .B2(n9651), .A(n9650), .ZN(P1_U3324) );
  OAI21_X1 U10848 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n9662) );
  OR2_X1 U10849 ( .A1(n9905), .A2(n9657), .ZN(n9661) );
  INV_X1 U10850 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10150) );
  OAI22_X1 U10851 ( .A1(n9658), .A2(n10150), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5049), .ZN(n9659) );
  INV_X1 U10852 ( .A(n9659), .ZN(n9660) );
  OAI211_X1 U10853 ( .C1(n9906), .C2(n9662), .A(n9661), .B(n9660), .ZN(n9663)
         );
  INV_X1 U10854 ( .A(n9663), .ZN(n9668) );
  OAI211_X1 U10855 ( .C1(n9666), .C2(n9665), .A(n9904), .B(n9664), .ZN(n9667)
         );
  NAND2_X1 U10856 ( .A1(n9668), .A2(n9667), .ZN(P2_U3247) );
  INV_X1 U10857 ( .A(n9673), .ZN(n9676) );
  OAI211_X1 U10858 ( .C1(n9671), .C2(n9881), .A(n9670), .B(n9669), .ZN(n9675)
         );
  NOR2_X1 U10859 ( .A1(n9673), .A2(n9672), .ZN(n9674) );
  AOI211_X1 U10860 ( .C1(n9693), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9677)
         );
  INV_X1 U10861 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U10862 ( .A1(n9891), .A2(n9677), .B1(n10093), .B2(n9889), .ZN(
        P1_U3484) );
  AOI22_X1 U10863 ( .A1(n9903), .A2(n9677), .B1(n7170), .B2(n9901), .ZN(
        P1_U3533) );
  OAI21_X1 U10864 ( .B1(n9679), .B2(n9881), .A(n9678), .ZN(n9680) );
  AOI21_X1 U10865 ( .B1(n9681), .B2(n9873), .A(n9680), .ZN(n9703) );
  INV_X1 U10866 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9682) );
  AOI22_X1 U10867 ( .A1(n9903), .A2(n9703), .B1(n9682), .B2(n9901), .ZN(
        P1_U3553) );
  OAI211_X1 U10868 ( .C1(n9686), .C2(n9881), .A(n9685), .B(n9684), .ZN(n9687)
         );
  AOI21_X1 U10869 ( .B1(n9688), .B2(n9887), .A(n9687), .ZN(n9705) );
  AOI22_X1 U10870 ( .A1(n9903), .A2(n9705), .B1(n9689), .B2(n9901), .ZN(
        P1_U3537) );
  OAI22_X1 U10871 ( .A1(n9691), .A2(n9883), .B1(n9690), .B2(n9881), .ZN(n9692)
         );
  AOI21_X1 U10872 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9695) );
  AND2_X1 U10873 ( .A1(n9696), .A2(n9695), .ZN(n9706) );
  AOI22_X1 U10874 ( .A1(n9903), .A2(n9706), .B1(n7392), .B2(n9901), .ZN(
        P1_U3536) );
  OAI22_X1 U10875 ( .A1(n9698), .A2(n9883), .B1(n9697), .B2(n9881), .ZN(n9699)
         );
  AOI211_X1 U10876 ( .C1(n9701), .C2(n9887), .A(n9700), .B(n9699), .ZN(n9708)
         );
  AOI22_X1 U10877 ( .A1(n9903), .A2(n9708), .B1(n7246), .B2(n9901), .ZN(
        P1_U3534) );
  INV_X1 U10878 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10879 ( .A1(n9891), .A2(n9703), .B1(n9702), .B2(n9889), .ZN(
        P1_U3521) );
  INV_X1 U10880 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9704) );
  AOI22_X1 U10881 ( .A1(n9891), .A2(n9705), .B1(n9704), .B2(n9889), .ZN(
        P1_U3496) );
  INV_X1 U10882 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U10883 ( .A1(n9891), .A2(n9706), .B1(n10153), .B2(n9889), .ZN(
        P1_U3493) );
  INV_X1 U10884 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U10885 ( .A1(n9891), .A2(n9708), .B1(n9707), .B2(n9889), .ZN(
        P1_U3487) );
  XNOR2_X1 U10886 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10887 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10888 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9710), .A(n9709), .ZN(
        n9711) );
  XNOR2_X1 U10889 ( .A(n9711), .B(n5986), .ZN(n9714) );
  AOI22_X1 U10890 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9837), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n9712) );
  OAI21_X1 U10891 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(P1_U3241) );
  OAI21_X1 U10892 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n9719) );
  AOI22_X1 U10893 ( .A1(n9816), .A2(n9719), .B1(n9808), .B2(n9718), .ZN(n9726)
         );
  XOR2_X1 U10894 ( .A(n9721), .B(n9720), .Z(n9724) );
  AOI211_X1 U10895 ( .C1(n9823), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9725)
         );
  OAI211_X1 U10896 ( .C1(n9821), .C2(n9727), .A(n9726), .B(n9725), .ZN(
        P1_U3245) );
  INV_X1 U10897 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9728) );
  OAI22_X1 U10898 ( .A1(n9828), .A2(n9729), .B1(n9821), .B2(n9728), .ZN(n9730)
         );
  INV_X1 U10899 ( .A(n9730), .ZN(n9741) );
  OAI21_X1 U10900 ( .B1(n9733), .B2(n9732), .A(n9731), .ZN(n9739) );
  AOI211_X1 U10901 ( .C1(n9736), .C2(n9735), .A(n9734), .B(n9833), .ZN(n9737)
         );
  AOI211_X1 U10902 ( .C1(n9823), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9740)
         );
  NAND2_X1 U10903 ( .A1(n9741), .A2(n9740), .ZN(P1_U3246) );
  XNOR2_X1 U10904 ( .A(n9743), .B(n9742), .ZN(n9745) );
  INV_X1 U10905 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9744) );
  OAI22_X1 U10906 ( .A1(n9833), .A2(n9745), .B1(n9821), .B2(n9744), .ZN(n9746)
         );
  INV_X1 U10907 ( .A(n9746), .ZN(n9754) );
  AOI211_X1 U10908 ( .C1(n9749), .C2(n9748), .A(n9747), .B(n9782), .ZN(n9750)
         );
  AOI211_X1 U10909 ( .C1(n9808), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9753)
         );
  NAND2_X1 U10910 ( .A1(n9754), .A2(n9753), .ZN(P1_U3247) );
  AOI21_X1 U10911 ( .B1(n9808), .B2(n9756), .A(n9755), .ZN(n9766) );
  OAI21_X1 U10912 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(n9764) );
  OAI21_X1 U10913 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(n9763) );
  AOI22_X1 U10914 ( .A1(n9816), .A2(n9764), .B1(n9823), .B2(n9763), .ZN(n9765)
         );
  OAI211_X1 U10915 ( .C1(n9821), .C2(n9767), .A(n9766), .B(n9765), .ZN(
        P1_U3248) );
  AOI21_X1 U10916 ( .B1(n9808), .B2(n9769), .A(n9768), .ZN(n9779) );
  OAI21_X1 U10917 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9777) );
  OAI21_X1 U10918 ( .B1(n9775), .B2(n9774), .A(n9773), .ZN(n9776) );
  AOI22_X1 U10919 ( .A1(n9816), .A2(n9777), .B1(n9823), .B2(n9776), .ZN(n9778)
         );
  OAI211_X1 U10920 ( .C1(n9821), .C2(n9780), .A(n9779), .B(n9778), .ZN(
        P1_U3249) );
  AOI211_X1 U10921 ( .C1(n9784), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9785)
         );
  AOI211_X1 U10922 ( .C1(n9808), .C2(n9787), .A(n9786), .B(n9785), .ZN(n9793)
         );
  OAI21_X1 U10923 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9791) );
  NAND2_X1 U10924 ( .A1(n9791), .A2(n9816), .ZN(n9792) );
  OAI211_X1 U10925 ( .C1(n10366), .C2(n9821), .A(n9793), .B(n9792), .ZN(
        P1_U3250) );
  INV_X1 U10926 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9805) );
  AOI21_X1 U10927 ( .B1(n9808), .B2(n9795), .A(n9794), .ZN(n9804) );
  OAI21_X1 U10928 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(n9802) );
  XNOR2_X1 U10929 ( .A(n9800), .B(n9799), .ZN(n9801) );
  AOI22_X1 U10930 ( .A1(n9816), .A2(n9802), .B1(n9823), .B2(n9801), .ZN(n9803)
         );
  OAI211_X1 U10931 ( .C1(n9821), .C2(n9805), .A(n9804), .B(n9803), .ZN(
        P1_U3252) );
  INV_X1 U10932 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9820) );
  AOI21_X1 U10933 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9819) );
  OAI21_X1 U10934 ( .B1(n9811), .B2(n9810), .A(n9809), .ZN(n9817) );
  OAI21_X1 U10935 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9815) );
  AOI22_X1 U10936 ( .A1(n9817), .A2(n9823), .B1(n9816), .B2(n9815), .ZN(n9818)
         );
  OAI211_X1 U10937 ( .C1(n9821), .C2(n9820), .A(n9819), .B(n9818), .ZN(
        P1_U3255) );
  OAI211_X1 U10938 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9827)
         );
  OAI211_X1 U10939 ( .C1(n9829), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9830)
         );
  INV_X1 U10940 ( .A(n9830), .ZN(n9839) );
  NAND2_X1 U10941 ( .A1(n9832), .A2(n9831), .ZN(n9834) );
  AOI21_X1 U10942 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  AOI21_X1 U10943 ( .B1(n9837), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9836), .ZN(
        n9838) );
  NAND2_X1 U10944 ( .A1(n9839), .A2(n9838), .ZN(P1_U3259) );
  AND2_X1 U10945 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9840), .ZN(P1_U3292) );
  AND2_X1 U10946 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9840), .ZN(P1_U3293) );
  AND2_X1 U10947 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9840), .ZN(P1_U3294) );
  INV_X1 U10948 ( .A(n9840), .ZN(n9841) );
  INV_X1 U10949 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U10950 ( .A1(n9841), .A2(n10217), .ZN(P1_U3295) );
  AND2_X1 U10951 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9840), .ZN(P1_U3296) );
  AND2_X1 U10952 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9840), .ZN(P1_U3297) );
  AND2_X1 U10953 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9840), .ZN(P1_U3298) );
  INV_X1 U10954 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10287) );
  NOR2_X1 U10955 ( .A1(n9841), .A2(n10287), .ZN(P1_U3299) );
  AND2_X1 U10956 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9840), .ZN(P1_U3300) );
  AND2_X1 U10957 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9840), .ZN(P1_U3301) );
  AND2_X1 U10958 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9840), .ZN(P1_U3302) );
  AND2_X1 U10959 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9840), .ZN(P1_U3303) );
  INV_X1 U10960 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U10961 ( .A1(n9841), .A2(n10196), .ZN(P1_U3304) );
  AND2_X1 U10962 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9840), .ZN(P1_U3305) );
  AND2_X1 U10963 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9840), .ZN(P1_U3306) );
  INV_X1 U10964 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U10965 ( .A1(n9841), .A2(n10122), .ZN(P1_U3307) );
  AND2_X1 U10966 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9840), .ZN(P1_U3308) );
  AND2_X1 U10967 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9840), .ZN(P1_U3309) );
  INV_X1 U10968 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U10969 ( .A1(n9841), .A2(n10198), .ZN(P1_U3310) );
  AND2_X1 U10970 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9840), .ZN(P1_U3311) );
  INV_X1 U10971 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U10972 ( .A1(n9841), .A2(n10228), .ZN(P1_U3312) );
  AND2_X1 U10973 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9840), .ZN(P1_U3313) );
  INV_X1 U10974 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10233) );
  NOR2_X1 U10975 ( .A1(n9841), .A2(n10233), .ZN(P1_U3314) );
  AND2_X1 U10976 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9840), .ZN(P1_U3315) );
  AND2_X1 U10977 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9840), .ZN(P1_U3316) );
  INV_X1 U10978 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10109) );
  NOR2_X1 U10979 ( .A1(n9841), .A2(n10109), .ZN(P1_U3317) );
  AND2_X1 U10980 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9840), .ZN(P1_U3318) );
  AND2_X1 U10981 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9840), .ZN(P1_U3319) );
  AND2_X1 U10982 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9840), .ZN(P1_U3320) );
  INV_X1 U10983 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U10984 ( .A1(n9841), .A2(n10133), .ZN(P1_U3321) );
  NOR2_X1 U10985 ( .A1(n9842), .A2(n9876), .ZN(n9846) );
  OAI21_X1 U10986 ( .B1(n7266), .B2(n9881), .A(n9843), .ZN(n9844) );
  NOR4_X1 U10987 ( .A1(n9847), .A2(n9846), .A3(n9845), .A4(n9844), .ZN(n9892)
         );
  INV_X1 U10988 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U10989 ( .A1(n9891), .A2(n9892), .B1(n10183), .B2(n9889), .ZN(
        P1_U3457) );
  OAI22_X1 U10990 ( .A1(n9849), .A2(n9883), .B1(n9848), .B2(n9881), .ZN(n9851)
         );
  AOI211_X1 U10991 ( .C1(n9887), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9893)
         );
  INV_X1 U10992 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U10993 ( .A1(n9891), .A2(n9893), .B1(n9853), .B2(n9889), .ZN(
        P1_U3463) );
  NAND3_X1 U10994 ( .A1(n9856), .A2(n9855), .A3(n9854), .ZN(n9857) );
  AOI21_X1 U10995 ( .B1(n9858), .B2(n9887), .A(n9857), .ZN(n9895) );
  INV_X1 U10996 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10119) );
  AOI22_X1 U10997 ( .A1(n9891), .A2(n9895), .B1(n10119), .B2(n9889), .ZN(
        P1_U3469) );
  OAI211_X1 U10998 ( .C1(n9861), .C2(n9881), .A(n9860), .B(n9859), .ZN(n9862)
         );
  AOI21_X1 U10999 ( .B1(n9887), .B2(n9863), .A(n9862), .ZN(n9897) );
  INV_X1 U11000 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9864) );
  AOI22_X1 U11001 ( .A1(n9891), .A2(n9897), .B1(n9864), .B2(n9889), .ZN(
        P1_U3472) );
  OAI211_X1 U11002 ( .C1(n9867), .C2(n9881), .A(n9866), .B(n9865), .ZN(n9868)
         );
  AOI21_X1 U11003 ( .B1(n9869), .B2(n9887), .A(n9868), .ZN(n9898) );
  INV_X1 U11004 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U11005 ( .A1(n9891), .A2(n9898), .B1(n9870), .B2(n9889), .ZN(
        P1_U3475) );
  AOI22_X1 U11006 ( .A1(n9874), .A2(n9873), .B1(n9872), .B2(n9871), .ZN(n9875)
         );
  OAI21_X1 U11007 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  NOR2_X1 U11008 ( .A1(n9879), .A2(n9878), .ZN(n9900) );
  INV_X1 U11009 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U11010 ( .A1(n9891), .A2(n9900), .B1(n9880), .B2(n9889), .ZN(
        P1_U3478) );
  OAI22_X1 U11011 ( .A1(n9884), .A2(n9883), .B1(n9882), .B2(n9881), .ZN(n9885)
         );
  AOI211_X1 U11012 ( .C1(n9888), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9902)
         );
  INV_X1 U11013 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9890) );
  AOI22_X1 U11014 ( .A1(n9891), .A2(n9902), .B1(n9890), .B2(n9889), .ZN(
        P1_U3481) );
  AOI22_X1 U11015 ( .A1(n9903), .A2(n9892), .B1(n7109), .B2(n9901), .ZN(
        P1_U3524) );
  INV_X1 U11016 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U11017 ( .A1(n9903), .A2(n9893), .B1(n10255), .B2(n9901), .ZN(
        P1_U3526) );
  INV_X1 U11018 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9894) );
  AOI22_X1 U11019 ( .A1(n9903), .A2(n9895), .B1(n9894), .B2(n9901), .ZN(
        P1_U3528) );
  INV_X1 U11020 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U11021 ( .A1(n9903), .A2(n9897), .B1(n9896), .B2(n9901), .ZN(
        P1_U3529) );
  INV_X1 U11022 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U11023 ( .A1(n9903), .A2(n9898), .B1(n10214), .B2(n9901), .ZN(
        P1_U3530) );
  AOI22_X1 U11024 ( .A1(n9903), .A2(n9900), .B1(n9899), .B2(n9901), .ZN(
        P1_U3531) );
  AOI22_X1 U11025 ( .A1(n9903), .A2(n9902), .B1(n7180), .B2(n9901), .ZN(
        P1_U3532) );
  AOI22_X1 U11026 ( .A1(n9904), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9922), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U11027 ( .A1(n9917), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9910) );
  NOR2_X1 U11028 ( .A1(n9927), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9908) );
  OAI21_X1 U11029 ( .B1(n9906), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9905), .ZN(
        n9907) );
  OAI21_X1 U11030 ( .B1(n9908), .B2(n9907), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9909) );
  OAI211_X1 U11031 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9911), .A(n9910), .B(
        n9909), .ZN(P2_U3245) );
  AOI21_X1 U11032 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n9928) );
  INV_X1 U11033 ( .A(n9915), .ZN(n9916) );
  AOI21_X1 U11034 ( .B1(n9917), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n9916), .ZN(
        n9926) );
  OAI21_X1 U11035 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9921) );
  AOI22_X1 U11036 ( .A1(n9924), .A2(n9923), .B1(n9922), .B2(n9921), .ZN(n9925)
         );
  OAI211_X1 U11037 ( .C1(n9928), .C2(n9927), .A(n9926), .B(n9925), .ZN(
        P2_U3258) );
  INV_X1 U11038 ( .A(n9929), .ZN(n9938) );
  NAND2_X1 U11039 ( .A1(n9931), .A2(n9930), .ZN(n9936) );
  INV_X1 U11040 ( .A(n9932), .ZN(n9934) );
  AOI22_X1 U11041 ( .A1(n8998), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9934), .B2(
        n9933), .ZN(n9935) );
  OAI211_X1 U11042 ( .C1(n9938), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9939)
         );
  AOI21_X1 U11043 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9942) );
  OAI21_X1 U11044 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(P2_U3287) );
  INV_X1 U11045 ( .A(n9945), .ZN(n9947) );
  NAND2_X1 U11046 ( .A1(n9947), .A2(n9946), .ZN(n9954) );
  AND2_X1 U11047 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9954), .ZN(P2_U3297) );
  AND2_X1 U11048 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9954), .ZN(P2_U3298) );
  AND2_X1 U11049 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9954), .ZN(P2_U3299) );
  AND2_X1 U11050 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9954), .ZN(P2_U3300) );
  INV_X1 U11051 ( .A(n9954), .ZN(n9948) );
  NOR2_X1 U11052 ( .A1(n9948), .A2(n10289), .ZN(P2_U3301) );
  INV_X1 U11053 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10318) );
  NOR2_X1 U11054 ( .A1(n9948), .A2(n10318), .ZN(P2_U3302) );
  AND2_X1 U11055 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9954), .ZN(P2_U3303) );
  NOR2_X1 U11056 ( .A1(n9948), .A2(n10140), .ZN(P2_U3304) );
  NOR2_X1 U11057 ( .A1(n9948), .A2(n10105), .ZN(P2_U3305) );
  INV_X1 U11058 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10277) );
  NOR2_X1 U11059 ( .A1(n9948), .A2(n10277), .ZN(P2_U3306) );
  AND2_X1 U11060 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9954), .ZN(P2_U3307) );
  AND2_X1 U11061 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9954), .ZN(P2_U3308) );
  NOR2_X1 U11062 ( .A1(n9948), .A2(n10181), .ZN(P2_U3309) );
  AND2_X1 U11063 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9954), .ZN(P2_U3310) );
  AND2_X1 U11064 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9954), .ZN(P2_U3311) );
  AND2_X1 U11065 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9954), .ZN(P2_U3312) );
  INV_X1 U11066 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10253) );
  NOR2_X1 U11067 ( .A1(n9948), .A2(n10253), .ZN(P2_U3313) );
  INV_X1 U11068 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10168) );
  NOR2_X1 U11069 ( .A1(n9948), .A2(n10168), .ZN(P2_U3314) );
  AND2_X1 U11070 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9954), .ZN(P2_U3315) );
  AND2_X1 U11071 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9954), .ZN(P2_U3316) );
  AND2_X1 U11072 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9954), .ZN(P2_U3317) );
  AND2_X1 U11073 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9954), .ZN(P2_U3318) );
  INV_X1 U11074 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U11075 ( .A1(n9948), .A2(n10126), .ZN(P2_U3319) );
  AND2_X1 U11076 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9954), .ZN(P2_U3320) );
  AND2_X1 U11077 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9954), .ZN(P2_U3321) );
  AND2_X1 U11078 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9954), .ZN(P2_U3322) );
  INV_X1 U11079 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10291) );
  NOR2_X1 U11080 ( .A1(n9948), .A2(n10291), .ZN(P2_U3323) );
  AND2_X1 U11081 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9954), .ZN(P2_U3324) );
  AND2_X1 U11082 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9954), .ZN(P2_U3325) );
  AND2_X1 U11083 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9954), .ZN(P2_U3326) );
  NOR2_X1 U11084 ( .A1(n9949), .A2(n9952), .ZN(n9951) );
  INV_X1 U11085 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U11086 ( .A1(n9957), .A2(n9951), .B1(n9950), .B2(n9954), .ZN(
        P2_U3437) );
  NOR2_X1 U11087 ( .A1(n9953), .A2(n9952), .ZN(n9956) );
  INV_X1 U11088 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11089 ( .A1(n9957), .A2(n9956), .B1(n9955), .B2(n9954), .ZN(
        P2_U3438) );
  NAND3_X1 U11090 ( .A1(n9960), .A2(n9959), .A3(n9958), .ZN(n9961) );
  OAI21_X1 U11091 ( .B1(n9962), .B2(n9979), .A(n9961), .ZN(n9963) );
  AOI21_X1 U11092 ( .B1(n9964), .B2(n9985), .A(n9963), .ZN(n9966) );
  AND2_X1 U11093 ( .A1(n9966), .A2(n9965), .ZN(n9990) );
  INV_X1 U11094 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U11095 ( .A1(n9155), .A2(n9990), .B1(n9967), .B2(n9987), .ZN(
        P2_U3457) );
  OAI21_X1 U11096 ( .B1(n10344), .B2(n9979), .A(n9968), .ZN(n9970) );
  AOI211_X1 U11097 ( .C1(n9985), .C2(n9971), .A(n9970), .B(n9969), .ZN(n9992)
         );
  AOI22_X1 U11098 ( .A1(n9155), .A2(n9992), .B1(n5082), .B2(n9987), .ZN(
        P2_U3463) );
  INV_X1 U11099 ( .A(n9972), .ZN(n9977) );
  OAI21_X1 U11100 ( .B1(n9974), .B2(n9979), .A(n9973), .ZN(n9976) );
  AOI211_X1 U11101 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9993)
         );
  INV_X1 U11102 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U11103 ( .A1(n9155), .A2(n9993), .B1(n10132), .B2(n9987), .ZN(
        P2_U3481) );
  OAI22_X1 U11104 ( .A1(n9982), .A2(n9981), .B1(n9980), .B2(n9979), .ZN(n9984)
         );
  AOI211_X1 U11105 ( .C1(n9986), .C2(n9985), .A(n9984), .B(n9983), .ZN(n9995)
         );
  INV_X1 U11106 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11107 ( .A1(n9155), .A2(n9995), .B1(n9988), .B2(n9987), .ZN(
        P2_U3487) );
  AOI22_X1 U11108 ( .A1(n9996), .A2(n9990), .B1(n9989), .B2(n9994), .ZN(
        P2_U3522) );
  INV_X1 U11109 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11110 ( .A1(n9996), .A2(n9992), .B1(n9991), .B2(n9994), .ZN(
        P2_U3524) );
  AOI22_X1 U11111 ( .A1(n9996), .A2(n9993), .B1(n5218), .B2(n9994), .ZN(
        P2_U3530) );
  AOI22_X1 U11112 ( .A1(n9996), .A2(n9995), .B1(n6977), .B2(n9994), .ZN(
        P2_U3532) );
  INV_X1 U11113 ( .A(n9997), .ZN(n9998) );
  NAND2_X1 U11114 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  XOR2_X1 U11115 ( .A(n10001), .B(n10000), .Z(ADD_1071_U5) );
  INV_X1 U11116 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10215) );
  INV_X1 U11117 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U11118 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .B1(n10215), .B2(n10002), .ZN(ADD_1071_U46) );
  OAI21_X1 U11119 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(ADD_1071_U56) );
  OAI21_X1 U11120 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(ADD_1071_U57) );
  OAI21_X1 U11121 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(ADD_1071_U58) );
  OAI21_X1 U11122 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(ADD_1071_U59) );
  OAI21_X1 U11123 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(ADD_1071_U60) );
  OAI21_X1 U11124 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(ADD_1071_U61) );
  AOI21_X1 U11125 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(ADD_1071_U62) );
  AOI21_X1 U11126 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(ADD_1071_U63) );
  NAND2_X1 U11127 ( .A1(keyinput25), .A2(keyinput101), .ZN(n10027) );
  NOR3_X1 U11128 ( .A1(keyinput113), .A2(keyinput29), .A3(n10027), .ZN(n10028)
         );
  NAND3_X1 U11129 ( .A1(keyinput93), .A2(keyinput80), .A3(n10028), .ZN(n10041)
         );
  NOR2_X1 U11130 ( .A1(keyinput102), .A2(keyinput73), .ZN(n10029) );
  NAND3_X1 U11131 ( .A1(keyinput71), .A2(keyinput28), .A3(n10029), .ZN(n10030)
         );
  NOR3_X1 U11132 ( .A1(keyinput60), .A2(keyinput65), .A3(n10030), .ZN(n10039)
         );
  NOR2_X1 U11133 ( .A1(keyinput43), .A2(keyinput72), .ZN(n10031) );
  NAND3_X1 U11134 ( .A1(keyinput51), .A2(keyinput96), .A3(n10031), .ZN(n10037)
         );
  OR4_X1 U11135 ( .A1(keyinput1), .A2(keyinput63), .A3(keyinput126), .A4(
        keyinput45), .ZN(n10036) );
  INV_X1 U11136 ( .A(keyinput114), .ZN(n10032) );
  NAND4_X1 U11137 ( .A1(keyinput44), .A2(keyinput116), .A3(keyinput20), .A4(
        n10032), .ZN(n10035) );
  NOR2_X1 U11138 ( .A1(keyinput47), .A2(keyinput17), .ZN(n10033) );
  NAND3_X1 U11139 ( .A1(keyinput16), .A2(keyinput119), .A3(n10033), .ZN(n10034) );
  NOR4_X1 U11140 ( .A1(n10037), .A2(n10036), .A3(n10035), .A4(n10034), .ZN(
        n10038) );
  NAND4_X1 U11141 ( .A1(keyinput42), .A2(keyinput23), .A3(n10039), .A4(n10038), 
        .ZN(n10040) );
  NOR4_X1 U11142 ( .A1(keyinput125), .A2(keyinput57), .A3(n10041), .A4(n10040), 
        .ZN(n10089) );
  INV_X1 U11143 ( .A(keyinput66), .ZN(n10042) );
  NAND4_X1 U11144 ( .A1(keyinput91), .A2(keyinput95), .A3(keyinput33), .A4(
        n10042), .ZN(n10043) );
  NOR4_X1 U11145 ( .A1(keyinput87), .A2(keyinput100), .A3(keyinput5), .A4(
        n10043), .ZN(n10055) );
  NOR4_X1 U11146 ( .A1(keyinput11), .A2(keyinput61), .A3(keyinput83), .A4(
        keyinput76), .ZN(n10054) );
  NAND2_X1 U11147 ( .A1(keyinput55), .A2(keyinput26), .ZN(n10044) );
  NOR3_X1 U11148 ( .A1(keyinput67), .A2(keyinput122), .A3(n10044), .ZN(n10053)
         );
  OR4_X1 U11149 ( .A1(keyinput12), .A2(keyinput88), .A3(keyinput52), .A4(
        keyinput90), .ZN(n10051) );
  INV_X1 U11150 ( .A(keyinput103), .ZN(n10045) );
  NAND4_X1 U11151 ( .A1(keyinput15), .A2(keyinput111), .A3(keyinput68), .A4(
        n10045), .ZN(n10050) );
  NOR2_X1 U11152 ( .A1(keyinput106), .A2(keyinput27), .ZN(n10046) );
  NAND3_X1 U11153 ( .A1(keyinput98), .A2(keyinput70), .A3(n10046), .ZN(n10049)
         );
  NOR2_X1 U11154 ( .A1(keyinput64), .A2(keyinput54), .ZN(n10047) );
  NAND3_X1 U11155 ( .A1(keyinput123), .A2(keyinput115), .A3(n10047), .ZN(
        n10048) );
  NOR4_X1 U11156 ( .A1(n10051), .A2(n10050), .A3(n10049), .A4(n10048), .ZN(
        n10052) );
  NAND4_X1 U11157 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        n10087) );
  NAND2_X1 U11158 ( .A1(keyinput84), .A2(keyinput105), .ZN(n10056) );
  NOR3_X1 U11159 ( .A1(keyinput99), .A2(keyinput48), .A3(n10056), .ZN(n10057)
         );
  NAND3_X1 U11160 ( .A1(keyinput24), .A2(keyinput9), .A3(n10057), .ZN(n10058)
         );
  NOR3_X1 U11161 ( .A1(keyinput112), .A2(keyinput41), .A3(n10058), .ZN(n10070)
         );
  NOR4_X1 U11162 ( .A1(keyinput35), .A2(keyinput22), .A3(keyinput18), .A4(
        keyinput32), .ZN(n10069) );
  NAND2_X1 U11163 ( .A1(keyinput36), .A2(keyinput14), .ZN(n10059) );
  NOR3_X1 U11164 ( .A1(keyinput19), .A2(keyinput97), .A3(n10059), .ZN(n10068)
         );
  NAND4_X1 U11165 ( .A1(keyinput107), .A2(keyinput118), .A3(keyinput37), .A4(
        keyinput124), .ZN(n10066) );
  NOR2_X1 U11166 ( .A1(keyinput108), .A2(keyinput110), .ZN(n10060) );
  NAND3_X1 U11167 ( .A1(keyinput3), .A2(keyinput79), .A3(n10060), .ZN(n10065)
         );
  NOR2_X1 U11168 ( .A1(keyinput34), .A2(keyinput21), .ZN(n10061) );
  NAND3_X1 U11169 ( .A1(keyinput127), .A2(keyinput117), .A3(n10061), .ZN(
        n10064) );
  INV_X1 U11170 ( .A(keyinput8), .ZN(n10062) );
  NAND4_X1 U11171 ( .A1(keyinput6), .A2(keyinput59), .A3(keyinput81), .A4(
        n10062), .ZN(n10063) );
  NOR4_X1 U11172 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10067) );
  NAND4_X1 U11173 ( .A1(n10070), .A2(n10069), .A3(n10068), .A4(n10067), .ZN(
        n10086) );
  NAND2_X1 U11174 ( .A1(keyinput120), .A2(keyinput82), .ZN(n10071) );
  NOR3_X1 U11175 ( .A1(keyinput77), .A2(keyinput69), .A3(n10071), .ZN(n10077)
         );
  NOR4_X1 U11176 ( .A1(keyinput121), .A2(keyinput40), .A3(keyinput46), .A4(
        keyinput74), .ZN(n10076) );
  INV_X1 U11177 ( .A(keyinput50), .ZN(n10072) );
  NOR4_X1 U11178 ( .A1(keyinput109), .A2(keyinput30), .A3(keyinput13), .A4(
        n10072), .ZN(n10075) );
  NAND2_X1 U11179 ( .A1(keyinput2), .A2(keyinput92), .ZN(n10073) );
  NOR3_X1 U11180 ( .A1(keyinput53), .A2(keyinput38), .A3(n10073), .ZN(n10074)
         );
  NAND4_X1 U11181 ( .A1(n10077), .A2(n10076), .A3(n10075), .A4(n10074), .ZN(
        n10085) );
  NOR4_X1 U11182 ( .A1(keyinput75), .A2(keyinput58), .A3(keyinput4), .A4(
        keyinput49), .ZN(n10083) );
  INV_X1 U11183 ( .A(keyinput31), .ZN(n10078) );
  NOR4_X1 U11184 ( .A1(keyinput94), .A2(keyinput104), .A3(keyinput39), .A4(
        n10078), .ZN(n10082) );
  AND4_X1 U11185 ( .A1(keyinput85), .A2(keyinput0), .A3(keyinput89), .A4(
        keyinput86), .ZN(n10081) );
  INV_X1 U11186 ( .A(keyinput78), .ZN(n10079) );
  NOR4_X1 U11187 ( .A1(keyinput56), .A2(keyinput10), .A3(keyinput62), .A4(
        n10079), .ZN(n10080) );
  NAND4_X1 U11188 ( .A1(n10083), .A2(n10082), .A3(n10081), .A4(n10080), .ZN(
        n10084) );
  NOR4_X1 U11189 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10088) );
  AOI21_X1 U11190 ( .B1(n10089), .B2(n10088), .A(keyinput7), .ZN(n10335) );
  INV_X1 U11191 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U11192 ( .A1(n5526), .A2(keyinput63), .B1(keyinput43), .B2(n10091), 
        .ZN(n10090) );
  OAI221_X1 U11193 ( .B1(n5526), .B2(keyinput63), .C1(n10091), .C2(keyinput43), 
        .A(n10090), .ZN(n10103) );
  AOI22_X1 U11194 ( .A1(n10093), .A2(keyinput51), .B1(keyinput126), .B2(n9331), 
        .ZN(n10092) );
  OAI221_X1 U11195 ( .B1(n10093), .B2(keyinput51), .C1(n9331), .C2(keyinput126), .A(n10092), .ZN(n10102) );
  INV_X1 U11196 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U11197 ( .A1(n10096), .A2(keyinput45), .B1(n10095), .B2(keyinput96), 
        .ZN(n10094) );
  OAI221_X1 U11198 ( .B1(n10096), .B2(keyinput45), .C1(n10095), .C2(keyinput96), .A(n10094), .ZN(n10101) );
  INV_X1 U11199 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10099) );
  INV_X1 U11200 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U11201 ( .A1(n10099), .A2(keyinput72), .B1(n10098), .B2(keyinput42), 
        .ZN(n10097) );
  OAI221_X1 U11202 ( .B1(n10099), .B2(keyinput72), .C1(n10098), .C2(keyinput42), .A(n10097), .ZN(n10100) );
  NOR4_X1 U11203 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10148) );
  INV_X1 U11204 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11205 ( .A1(n10106), .A2(keyinput73), .B1(keyinput60), .B2(n10105), 
        .ZN(n10104) );
  OAI221_X1 U11206 ( .B1(n10106), .B2(keyinput73), .C1(n10105), .C2(keyinput60), .A(n10104), .ZN(n10116) );
  AOI22_X1 U11207 ( .A1(n5490), .A2(keyinput23), .B1(keyinput71), .B2(n6895), 
        .ZN(n10107) );
  OAI221_X1 U11208 ( .B1(n5490), .B2(keyinput23), .C1(n6895), .C2(keyinput71), 
        .A(n10107), .ZN(n10115) );
  AOI22_X1 U11209 ( .A1(n5210), .A2(keyinput65), .B1(n10109), .B2(keyinput102), 
        .ZN(n10108) );
  OAI221_X1 U11210 ( .B1(n5210), .B2(keyinput65), .C1(n10109), .C2(keyinput102), .A(n10108), .ZN(n10114) );
  INV_X1 U11211 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10110) );
  XOR2_X1 U11212 ( .A(n10110), .B(keyinput125), .Z(n10112) );
  XNOR2_X1 U11213 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput28), .ZN(n10111) );
  NAND2_X1 U11214 ( .A1(n10112), .A2(n10111), .ZN(n10113) );
  NOR4_X1 U11215 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10147) );
  AOI22_X1 U11216 ( .A1(n10119), .A2(keyinput57), .B1(n10118), .B2(keyinput101), .ZN(n10117) );
  OAI221_X1 U11217 ( .B1(n10119), .B2(keyinput57), .C1(n10118), .C2(
        keyinput101), .A(n10117), .ZN(n10130) );
  AOI22_X1 U11218 ( .A1(n4993), .A2(keyinput113), .B1(keyinput93), .B2(n5236), 
        .ZN(n10120) );
  OAI221_X1 U11219 ( .B1(n4993), .B2(keyinput113), .C1(n5236), .C2(keyinput93), 
        .A(n10120), .ZN(n10129) );
  AOI22_X1 U11220 ( .A1(n10123), .A2(keyinput80), .B1(n10122), .B2(keyinput25), 
        .ZN(n10121) );
  OAI221_X1 U11221 ( .B1(n10123), .B2(keyinput80), .C1(n10122), .C2(keyinput25), .A(n10121), .ZN(n10128) );
  INV_X1 U11222 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U11223 ( .A1(n10126), .A2(keyinput29), .B1(n10125), .B2(keyinput47), 
        .ZN(n10124) );
  OAI221_X1 U11224 ( .B1(n10126), .B2(keyinput29), .C1(n10125), .C2(keyinput47), .A(n10124), .ZN(n10127) );
  NOR4_X1 U11225 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10146) );
  AOI22_X1 U11226 ( .A1(n10133), .A2(keyinput17), .B1(keyinput114), .B2(n10132), .ZN(n10131) );
  OAI221_X1 U11227 ( .B1(n10133), .B2(keyinput17), .C1(n10132), .C2(
        keyinput114), .A(n10131), .ZN(n10144) );
  INV_X1 U11228 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U11229 ( .A1(n10136), .A2(keyinput44), .B1(keyinput116), .B2(n10135), .ZN(n10134) );
  OAI221_X1 U11230 ( .B1(n10136), .B2(keyinput44), .C1(n10135), .C2(
        keyinput116), .A(n10134), .ZN(n10143) );
  XNOR2_X1 U11231 ( .A(P2_REG0_REG_20__SCAN_IN), .B(keyinput20), .ZN(n10139)
         );
  XNOR2_X1 U11232 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput119), .ZN(n10138) );
  XNOR2_X1 U11233 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput94), .ZN(n10137) );
  NAND3_X1 U11234 ( .A1(n10139), .A2(n10138), .A3(n10137), .ZN(n10142) );
  XNOR2_X1 U11235 ( .A(n10140), .B(keyinput16), .ZN(n10141) );
  NOR4_X1 U11236 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10145) );
  NAND4_X1 U11237 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(
        n10333) );
  AOI22_X1 U11238 ( .A1(n6908), .A2(keyinput49), .B1(keyinput56), .B2(n10150), 
        .ZN(n10149) );
  OAI221_X1 U11239 ( .B1(n6908), .B2(keyinput49), .C1(n10150), .C2(keyinput56), 
        .A(n10149), .ZN(n10163) );
  AOI22_X1 U11240 ( .A1(n10153), .A2(keyinput58), .B1(keyinput4), .B2(n10152), 
        .ZN(n10151) );
  OAI221_X1 U11241 ( .B1(n10153), .B2(keyinput58), .C1(n10152), .C2(keyinput4), 
        .A(n10151), .ZN(n10162) );
  AOI22_X1 U11242 ( .A1(n10156), .A2(keyinput31), .B1(n10155), .B2(keyinput75), 
        .ZN(n10154) );
  OAI221_X1 U11243 ( .B1(n10156), .B2(keyinput31), .C1(n10155), .C2(keyinput75), .A(n10154), .ZN(n10161) );
  INV_X1 U11244 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10157) );
  XOR2_X1 U11245 ( .A(n10157), .B(keyinput104), .Z(n10159) );
  XNOR2_X1 U11246 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput39), .ZN(n10158) );
  NAND2_X1 U11247 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  NOR4_X1 U11248 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10212) );
  AOI22_X1 U11249 ( .A1(n10166), .A2(keyinput10), .B1(keyinput62), .B2(n10165), 
        .ZN(n10164) );
  OAI221_X1 U11250 ( .B1(n10166), .B2(keyinput10), .C1(n10165), .C2(keyinput62), .A(n10164), .ZN(n10179) );
  AOI22_X1 U11251 ( .A1(n10169), .A2(keyinput78), .B1(keyinput85), .B2(n10168), 
        .ZN(n10167) );
  OAI221_X1 U11252 ( .B1(n10169), .B2(keyinput78), .C1(n10168), .C2(keyinput85), .A(n10167), .ZN(n10178) );
  INV_X1 U11253 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U11254 ( .A1(n10172), .A2(keyinput0), .B1(n10171), .B2(keyinput89), 
        .ZN(n10170) );
  OAI221_X1 U11255 ( .B1(n10172), .B2(keyinput0), .C1(n10171), .C2(keyinput89), 
        .A(n10170), .ZN(n10177) );
  INV_X1 U11256 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11257 ( .A1(n10175), .A2(keyinput86), .B1(keyinput121), .B2(n10174), .ZN(n10173) );
  OAI221_X1 U11258 ( .B1(n10175), .B2(keyinput86), .C1(n10174), .C2(
        keyinput121), .A(n10173), .ZN(n10176) );
  NOR4_X1 U11259 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10211) );
  AOI22_X1 U11260 ( .A1(n10181), .A2(keyinput40), .B1(keyinput46), .B2(n10361), 
        .ZN(n10180) );
  OAI221_X1 U11261 ( .B1(n10181), .B2(keyinput40), .C1(n10361), .C2(keyinput46), .A(n10180), .ZN(n10193) );
  AOI22_X1 U11262 ( .A1(n10184), .A2(keyinput69), .B1(keyinput92), .B2(n10183), 
        .ZN(n10182) );
  OAI221_X1 U11263 ( .B1(n10184), .B2(keyinput69), .C1(n10183), .C2(keyinput92), .A(n10182), .ZN(n10192) );
  INV_X1 U11264 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U11265 ( .A1(n10187), .A2(keyinput77), .B1(keyinput120), .B2(n10186), .ZN(n10185) );
  OAI221_X1 U11266 ( .B1(n10187), .B2(keyinput77), .C1(n10186), .C2(
        keyinput120), .A(n10185), .ZN(n10191) );
  XNOR2_X1 U11267 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput82), .ZN(n10189) );
  XNOR2_X1 U11268 ( .A(keyinput74), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n10188)
         );
  NAND2_X1 U11269 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  NOR4_X1 U11270 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10210) );
  AOI22_X1 U11271 ( .A1(n10196), .A2(keyinput87), .B1(n10195), .B2(keyinput13), 
        .ZN(n10194) );
  OAI221_X1 U11272 ( .B1(n10196), .B2(keyinput87), .C1(n10195), .C2(keyinput13), .A(n10194), .ZN(n10208) );
  AOI22_X1 U11273 ( .A1(n10199), .A2(keyinput50), .B1(n10198), .B2(keyinput30), 
        .ZN(n10197) );
  OAI221_X1 U11274 ( .B1(n10199), .B2(keyinput50), .C1(n10198), .C2(keyinput30), .A(n10197), .ZN(n10207) );
  INV_X1 U11275 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10202) );
  INV_X1 U11276 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U11277 ( .A1(n10202), .A2(keyinput38), .B1(n10201), .B2(keyinput53), 
        .ZN(n10200) );
  OAI221_X1 U11278 ( .B1(n10202), .B2(keyinput38), .C1(n10201), .C2(keyinput53), .A(n10200), .ZN(n10206) );
  XNOR2_X1 U11279 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput2), .ZN(n10204) );
  XNOR2_X1 U11280 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput109), .ZN(n10203) );
  NAND2_X1 U11281 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  NOR4_X1 U11282 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10209) );
  NAND4_X1 U11283 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n10332) );
  AOI22_X1 U11284 ( .A1(n10215), .A2(keyinput97), .B1(n10214), .B2(keyinput18), 
        .ZN(n10213) );
  OAI221_X1 U11285 ( .B1(n10215), .B2(keyinput97), .C1(n10214), .C2(keyinput18), .A(n10213), .ZN(n10225) );
  AOI22_X1 U11286 ( .A1(n10218), .A2(keyinput32), .B1(n10217), .B2(keyinput3), 
        .ZN(n10216) );
  OAI221_X1 U11287 ( .B1(n10218), .B2(keyinput32), .C1(n10217), .C2(keyinput3), 
        .A(n10216), .ZN(n10224) );
  XNOR2_X1 U11288 ( .A(P1_REG1_REG_21__SCAN_IN), .B(keyinput36), .ZN(n10222)
         );
  XNOR2_X1 U11289 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput22), .ZN(n10221) );
  XNOR2_X1 U11290 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput35), .ZN(n10220) );
  XNOR2_X1 U11291 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput14), .ZN(n10219)
         );
  NAND4_X1 U11292 ( .A1(n10222), .A2(n10221), .A3(n10220), .A4(n10219), .ZN(
        n10223) );
  NOR3_X1 U11293 ( .A1(n10225), .A2(n10224), .A3(n10223), .ZN(n10269) );
  AOI22_X1 U11294 ( .A1(n10228), .A2(keyinput99), .B1(keyinput84), .B2(n10227), 
        .ZN(n10226) );
  OAI221_X1 U11295 ( .B1(n10228), .B2(keyinput99), .C1(n10227), .C2(keyinput84), .A(n10226), .ZN(n10239) );
  AOI22_X1 U11296 ( .A1(n6954), .A2(keyinput41), .B1(n10230), .B2(keyinput19), 
        .ZN(n10229) );
  OAI221_X1 U11297 ( .B1(n6954), .B2(keyinput41), .C1(n10230), .C2(keyinput19), 
        .A(n10229), .ZN(n10238) );
  AOI22_X1 U11298 ( .A1(n10233), .A2(keyinput48), .B1(keyinput112), .B2(n10232), .ZN(n10231) );
  OAI221_X1 U11299 ( .B1(n10233), .B2(keyinput48), .C1(n10232), .C2(
        keyinput112), .A(n10231), .ZN(n10237) );
  XNOR2_X1 U11300 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput9), .ZN(n10235) );
  XNOR2_X1 U11301 ( .A(SI_10_), .B(keyinput105), .ZN(n10234) );
  NAND2_X1 U11302 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  NOR4_X1 U11303 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10268) );
  AOI22_X1 U11304 ( .A1(n4420), .A2(keyinput81), .B1(n10241), .B2(keyinput34), 
        .ZN(n10240) );
  OAI221_X1 U11305 ( .B1(n4420), .B2(keyinput81), .C1(n10241), .C2(keyinput34), 
        .A(n10240), .ZN(n10251) );
  AOI22_X1 U11306 ( .A1(n10244), .A2(keyinput127), .B1(keyinput117), .B2(n8551), .ZN(n10243) );
  OAI221_X1 U11307 ( .B1(n10244), .B2(keyinput127), .C1(n8551), .C2(
        keyinput117), .A(n10243), .ZN(n10250) );
  XNOR2_X1 U11308 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput59), .ZN(n10248) );
  XNOR2_X1 U11309 ( .A(P1_REG2_REG_15__SCAN_IN), .B(keyinput8), .ZN(n10247) );
  XNOR2_X1 U11310 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput21), .ZN(n10246)
         );
  XNOR2_X1 U11311 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput1), .ZN(n10245) );
  NAND4_X1 U11312 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10249) );
  NOR3_X1 U11313 ( .A1(n10251), .A2(n10250), .A3(n10249), .ZN(n10267) );
  AOI22_X1 U11314 ( .A1(n10253), .A2(keyinput79), .B1(n7122), .B2(keyinput37), 
        .ZN(n10252) );
  OAI221_X1 U11315 ( .B1(n10253), .B2(keyinput79), .C1(n7122), .C2(keyinput37), 
        .A(n10252), .ZN(n10265) );
  INV_X1 U11316 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U11317 ( .A1(n10256), .A2(keyinput118), .B1(keyinput108), .B2(
        n10255), .ZN(n10254) );
  OAI221_X1 U11318 ( .B1(n10256), .B2(keyinput118), .C1(n10255), .C2(
        keyinput108), .A(n10254), .ZN(n10264) );
  INV_X1 U11319 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U11320 ( .A1(n10259), .A2(keyinput124), .B1(n10258), .B2(keyinput6), 
        .ZN(n10257) );
  OAI221_X1 U11321 ( .B1(n10259), .B2(keyinput124), .C1(n10258), .C2(keyinput6), .A(n10257), .ZN(n10263) );
  XNOR2_X1 U11322 ( .A(P2_REG2_REG_20__SCAN_IN), .B(keyinput107), .ZN(n10261)
         );
  XNOR2_X1 U11323 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput110), .ZN(n10260) );
  NAND2_X1 U11324 ( .A1(n10261), .A2(n10260), .ZN(n10262) );
  NOR4_X1 U11325 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n10266) );
  NAND4_X1 U11326 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10331) );
  INV_X1 U11327 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U11328 ( .A1(n10362), .A2(keyinput88), .B1(n10271), .B2(keyinput52), 
        .ZN(n10270) );
  OAI221_X1 U11329 ( .B1(n10362), .B2(keyinput88), .C1(n10271), .C2(keyinput52), .A(n10270), .ZN(n10284) );
  AOI22_X1 U11330 ( .A1(n10274), .A2(keyinput68), .B1(keyinput12), .B2(n10273), 
        .ZN(n10272) );
  OAI221_X1 U11331 ( .B1(n10274), .B2(keyinput68), .C1(n10273), .C2(keyinput12), .A(n10272), .ZN(n10283) );
  INV_X1 U11332 ( .A(SI_21_), .ZN(n10276) );
  AOI22_X1 U11333 ( .A1(n10277), .A2(keyinput90), .B1(n10276), .B2(keyinput26), 
        .ZN(n10275) );
  OAI221_X1 U11334 ( .B1(n10277), .B2(keyinput90), .C1(n10276), .C2(keyinput26), .A(n10275), .ZN(n10282) );
  INV_X1 U11335 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n10278) );
  XOR2_X1 U11336 ( .A(n10278), .B(keyinput111), .Z(n10280) );
  XNOR2_X1 U11337 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput15), .ZN(n10279) );
  NAND2_X1 U11338 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  NOR4_X1 U11339 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(
        n10329) );
  NAND2_X1 U11340 ( .A1(n10286), .A2(keyinput91), .ZN(n10285) );
  OAI221_X1 U11341 ( .B1(n10287), .B2(keyinput7), .C1(n10286), .C2(keyinput91), 
        .A(n10285), .ZN(n10298) );
  AOI22_X1 U11342 ( .A1(n5986), .A2(keyinput100), .B1(keyinput5), .B2(n10289), 
        .ZN(n10288) );
  OAI221_X1 U11343 ( .B1(n5986), .B2(keyinput100), .C1(n10289), .C2(keyinput5), 
        .A(n10288), .ZN(n10297) );
  AOI22_X1 U11344 ( .A1(n10292), .A2(keyinput33), .B1(keyinput103), .B2(n10291), .ZN(n10290) );
  OAI221_X1 U11345 ( .B1(n10292), .B2(keyinput33), .C1(n10291), .C2(
        keyinput103), .A(n10290), .ZN(n10296) );
  AOI22_X1 U11346 ( .A1(n10294), .A2(keyinput66), .B1(n7180), .B2(keyinput95), 
        .ZN(n10293) );
  OAI221_X1 U11347 ( .B1(n10294), .B2(keyinput66), .C1(n7180), .C2(keyinput95), 
        .A(n10293), .ZN(n10295) );
  NOR4_X1 U11348 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10328) );
  AOI22_X1 U11349 ( .A1(n10300), .A2(keyinput54), .B1(n5107), .B2(keyinput64), 
        .ZN(n10299) );
  OAI221_X1 U11350 ( .B1(n10300), .B2(keyinput54), .C1(n5107), .C2(keyinput64), 
        .A(n10299), .ZN(n10310) );
  INV_X1 U11351 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10303) );
  INV_X1 U11352 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U11353 ( .A1(n10303), .A2(keyinput70), .B1(n10302), .B2(keyinput24), 
        .ZN(n10301) );
  OAI221_X1 U11354 ( .B1(n10303), .B2(keyinput70), .C1(n10302), .C2(keyinput24), .A(n10301), .ZN(n10309) );
  XNOR2_X1 U11355 ( .A(SI_26_), .B(keyinput115), .ZN(n10307) );
  XNOR2_X1 U11356 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput98), .ZN(n10306) );
  XNOR2_X1 U11357 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(keyinput106), .ZN(n10305)
         );
  XNOR2_X1 U11358 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput27), .ZN(n10304) );
  NAND4_X1 U11359 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10308) );
  NOR3_X1 U11360 ( .A1(n10310), .A2(n10309), .A3(n10308), .ZN(n10327) );
  INV_X1 U11361 ( .A(keyinput61), .ZN(n10312) );
  AOI22_X1 U11362 ( .A1(n7400), .A2(keyinput83), .B1(SI_31_), .B2(n10312), 
        .ZN(n10311) );
  OAI221_X1 U11363 ( .B1(n7400), .B2(keyinput83), .C1(n10312), .C2(SI_31_), 
        .A(n10311), .ZN(n10325) );
  AOI22_X1 U11364 ( .A1(n10315), .A2(keyinput67), .B1(keyinput11), .B2(n10314), 
        .ZN(n10313) );
  OAI221_X1 U11365 ( .B1(n10315), .B2(keyinput67), .C1(n10314), .C2(keyinput11), .A(n10313), .ZN(n10324) );
  AOI22_X1 U11366 ( .A1(n10318), .A2(keyinput122), .B1(n10317), .B2(
        keyinput123), .ZN(n10316) );
  OAI221_X1 U11367 ( .B1(n10318), .B2(keyinput122), .C1(n10317), .C2(
        keyinput123), .A(n10316), .ZN(n10323) );
  AOI22_X1 U11368 ( .A1(n10321), .A2(keyinput76), .B1(n10320), .B2(keyinput55), 
        .ZN(n10319) );
  OAI221_X1 U11369 ( .B1(n10321), .B2(keyinput76), .C1(n10320), .C2(keyinput55), .A(n10319), .ZN(n10322) );
  NOR4_X1 U11370 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  NAND4_X1 U11371 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n10330) );
  NOR4_X1 U11372 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10334) );
  OAI21_X1 U11373 ( .B1(P1_D_REG_24__SCAN_IN), .B2(n10335), .A(n10334), .ZN(
        n10354) );
  NOR2_X1 U11374 ( .A1(n4515), .A2(n10336), .ZN(n10337) );
  XNOR2_X1 U11375 ( .A(n10338), .B(n10337), .ZN(n10352) );
  OAI21_X1 U11376 ( .B1(n10341), .B2(n10340), .A(n10339), .ZN(n10347) );
  OAI22_X1 U11377 ( .A1(n10345), .A2(n10344), .B1(n10343), .B2(n10342), .ZN(
        n10346) );
  AOI211_X1 U11378 ( .C1(n10349), .C2(n10348), .A(n10347), .B(n10346), .ZN(
        n10350) );
  OAI21_X1 U11379 ( .B1(n10352), .B2(n10351), .A(n10350), .ZN(n10353) );
  XNOR2_X1 U11380 ( .A(n10354), .B(n10353), .ZN(P2_U3232) );
  XOR2_X1 U11381 ( .A(n10355), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11382 ( .A1(n10357), .A2(n10356), .ZN(n10358) );
  XOR2_X1 U11383 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10358), .Z(ADD_1071_U51) );
  OAI21_X1 U11384 ( .B1(n10361), .B2(n10360), .A(n10359), .ZN(n10363) );
  XOR2_X1 U11385 ( .A(n10363), .B(n10362), .Z(ADD_1071_U55) );
  AOI21_X1 U11386 ( .B1(n10366), .B2(n10365), .A(n10364), .ZN(ADD_1071_U47) );
  XOR2_X1 U11387 ( .A(n10368), .B(n10367), .Z(ADD_1071_U54) );
  XOR2_X1 U11388 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10369), .Z(ADD_1071_U48) );
  XOR2_X1 U11389 ( .A(n10370), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11390 ( .A(n10372), .B(n10371), .Z(ADD_1071_U53) );
  XNOR2_X1 U11391 ( .A(n10374), .B(n10373), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4933 ( .A(n6761), .Z(n6784) );
  CLKBUF_X1 U4936 ( .A(n6562), .Z(n7510) );
  CLKBUF_X1 U4943 ( .A(n6478), .Z(n6480) );
endmodule

