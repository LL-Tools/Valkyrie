

module b20_C_gen_AntiSAT_k_256_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4507, n4508, n4509, n4510, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479;

  OR2_X1 U5013 ( .A1(n8585), .A2(n9380), .ZN(n9414) );
  BUF_X2 U5014 ( .A(n6704), .Z(n4508) );
  INV_X1 U5015 ( .A(n5984), .ZN(n9858) );
  INV_X1 U5016 ( .A(n6699), .ZN(n6675) );
  INV_X1 U5017 ( .A(n7413), .ZN(n10166) );
  INV_X1 U5019 ( .A(n5218), .ZN(n7420) );
  CLKBUF_X2 U5020 ( .A(n5206), .Z(n5539) );
  NAND2_X1 U5021 ( .A1(n5760), .A2(n8243), .ZN(n5772) );
  CLKBUF_X2 U5022 ( .A(n6181), .Z(n6224) );
  CLKBUF_X2 U5023 ( .A(n6043), .Z(n6228) );
  NAND2_X1 U5024 ( .A1(n5678), .A2(n8801), .ZN(n8748) );
  INV_X1 U5025 ( .A(n6943), .ZN(n5790) );
  INV_X2 U5026 ( .A(n5209), .ZN(n5379) );
  CLKBUF_X2 U5027 ( .A(n6738), .Z(n6286) );
  XNOR2_X1 U5028 ( .A(n5227), .B(SI_5_), .ZN(n5225) );
  INV_X1 U5029 ( .A(n8748), .ZN(n8753) );
  NAND2_X1 U5030 ( .A1(n5790), .A2(n8759), .ZN(n6942) );
  NAND2_X1 U5031 ( .A1(n6699), .A2(n6507), .ZN(n6511) );
  INV_X1 U5032 ( .A(n5967), .ZN(n6050) );
  INV_X1 U5033 ( .A(n5740), .ZN(n8759) );
  OAI21_X1 U5034 ( .B1(n5772), .B2(P2_D_REG_0__SCAN_IN), .A(n6762), .ZN(n6941)
         );
  OAI21_X1 U5035 ( .B1(n5333), .B2(n5005), .A(n5003), .ZN(n8271) );
  INV_X1 U5036 ( .A(n6507), .ZN(n6702) );
  CLKBUF_X2 U5037 ( .A(n7132), .Z(n8838) );
  OR2_X1 U5038 ( .A1(n5614), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5634) );
  OR2_X1 U5039 ( .A1(n5559), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5577) );
  INV_X2 U5040 ( .A(n8799), .ZN(n8049) );
  INV_X2 U5041 ( .A(n6702), .ZN(n6681) );
  AND2_X1 U5042 ( .A1(n5077), .A2(n5076), .ZN(n6463) );
  NAND2_X1 U5043 ( .A1(n6502), .A2(n6504), .ZN(n7216) );
  NAND2_X1 U5044 ( .A1(n5680), .A2(n4509), .ZN(n6736) );
  INV_X1 U5045 ( .A(n5162), .ZN(n6743) );
  INV_X1 U5046 ( .A(n10095), .ZN(n10143) );
  CLKBUF_X3 U5047 ( .A(n5342), .Z(n5470) );
  XNOR2_X1 U5048 ( .A(n4747), .B(n4746), .ZN(n10113) );
  INV_X1 U5049 ( .A(n6039), .ZN(n5949) );
  AOI21_X2 U5050 ( .B1(n8405), .B2(n8403), .A(n8404), .ZN(n8506) );
  XNOR2_X2 U5051 ( .A(n5440), .B(n5371), .ZN(n6848) );
  CLKBUF_X1 U5052 ( .A(n10113), .Z(n4507) );
  INV_X1 U5053 ( .A(n6525), .ZN(n6704) );
  INV_X1 U5054 ( .A(n8799), .ZN(n4509) );
  NAND3_X1 U5055 ( .A1(n4715), .A2(n4712), .A3(n4711), .ZN(n8799) );
  AOI22_X2 U5056 ( .A1(n9773), .A2(n9657), .B1(n9894), .B2(n9762), .ZN(n9756)
         );
  AND2_X2 U5057 ( .A1(n5837), .A2(n5834), .ZN(n6039) );
  OR2_X1 U5058 ( .A1(n6271), .A2(n9684), .ZN(n4745) );
  AND2_X1 U5059 ( .A1(n4754), .A2(n4752), .ZN(n9644) );
  OAI21_X1 U5060 ( .B1(n9672), .B2(n9819), .A(n9673), .ZN(n9804) );
  OR2_X1 U5061 ( .A1(n8486), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U5062 ( .A1(n6101), .A2(n6100), .ZN(n8431) );
  NAND2_X1 U5063 ( .A1(n5286), .A2(n5285), .ZN(n10403) );
  NAND2_X1 U5064 ( .A1(n4514), .A2(n4513), .ZN(n5337) );
  NAND2_X1 U5065 ( .A1(n9511), .A2(n7334), .ZN(n7263) );
  NAND2_X1 U5066 ( .A1(n6393), .A2(n6391), .ZN(n7271) );
  NAND2_X1 U5067 ( .A1(n9512), .A2(n10150), .ZN(n6391) );
  INV_X1 U5068 ( .A(n7273), .ZN(n9511) );
  NAND2_X1 U5069 ( .A1(n9513), .A2(n10143), .ZN(n6390) );
  XNOR2_X2 U5070 ( .A(n5981), .B(n5982), .ZN(n6306) );
  AND3_X1 U5071 ( .A1(n4788), .A2(n4787), .A3(n4786), .ZN(n8647) );
  INV_X1 U5072 ( .A(n5188), .ZN(n4657) );
  INV_X4 U5073 ( .A(n6503), .ZN(n4510) );
  INV_X1 U5074 ( .A(n6736), .ZN(n5342) );
  NAND2_X1 U5075 ( .A1(n6736), .A2(n6743), .ZN(n5205) );
  AND2_X1 U5076 ( .A1(n6736), .A2(n6286), .ZN(n5206) );
  INV_X1 U5077 ( .A(n6505), .ZN(n6502) );
  CLKBUF_X3 U5078 ( .A(n6738), .Z(n6744) );
  OR2_X1 U5079 ( .A1(n9359), .A2(n6712), .ZN(n6732) );
  AND2_X1 U5080 ( .A1(n9469), .A2(n6698), .ZN(n9359) );
  NAND2_X1 U5081 ( .A1(n4905), .A2(n4904), .ZN(n9469) );
  AND2_X1 U5082 ( .A1(n9701), .A2(n9700), .ZN(n9867) );
  AOI21_X1 U5083 ( .B1(n4614), .B2(n6297), .A(n6464), .ZN(n5076) );
  NOR2_X1 U5084 ( .A1(n9719), .A2(n9718), .ZN(n9717) );
  NAND2_X1 U5085 ( .A1(n4515), .A2(n9677), .ZN(n9744) );
  NAND2_X1 U5086 ( .A1(n9757), .A2(n4516), .ZN(n4515) );
  NAND2_X1 U5087 ( .A1(n5054), .A2(n5053), .ZN(n8869) );
  NAND2_X1 U5088 ( .A1(n9776), .A2(n9775), .ZN(n9757) );
  XNOR2_X1 U5089 ( .A(n5660), .B(n5659), .ZN(n8360) );
  NOR2_X1 U5090 ( .A1(n4899), .A2(n4896), .ZN(n4895) );
  NAND2_X1 U5091 ( .A1(n9791), .A2(n9676), .ZN(n9776) );
  OAI21_X1 U5092 ( .B1(n5647), .B2(n4630), .A(n5646), .ZN(n5660) );
  NAND2_X1 U5093 ( .A1(n9804), .A2(n9675), .ZN(n4831) );
  AND2_X1 U5094 ( .A1(n5858), .A2(n5857), .ZN(n9739) );
  AND2_X1 U5095 ( .A1(n9760), .A2(n9758), .ZN(n4516) );
  NAND2_X1 U5096 ( .A1(n6350), .A2(n6426), .ZN(n9672) );
  OR2_X1 U5097 ( .A1(n6594), .A2(n6593), .ZN(n6604) );
  OR2_X1 U5098 ( .A1(n6586), .A2(n8523), .ZN(n6597) );
  OAI21_X1 U5099 ( .B1(n8330), .B2(n8329), .A(n6417), .ZN(n8488) );
  NAND2_X1 U5100 ( .A1(n5576), .A2(n5575), .ZN(n5597) );
  AOI21_X1 U5101 ( .B1(n8284), .B2(n6349), .A(n6348), .ZN(n8330) );
  OAI211_X1 U5102 ( .C1(n6347), .C2(n4830), .A(n4520), .B(n8311), .ZN(n8284)
         );
  NAND2_X1 U5103 ( .A1(n8073), .A2(n4529), .ZN(n4520) );
  AND2_X1 U5104 ( .A1(n6412), .A2(n8285), .ZN(n8311) );
  INV_X1 U5105 ( .A(n8291), .ZN(n8119) );
  AND2_X1 U5106 ( .A1(n5515), .A2(n4600), .ZN(n4960) );
  NAND2_X1 U5107 ( .A1(n5878), .A2(n5877), .ZN(n9398) );
  NAND2_X1 U5108 ( .A1(n6317), .A2(n8304), .ZN(n8291) );
  OR2_X1 U5109 ( .A1(n8001), .A2(n8070), .ZN(n8073) );
  AND2_X1 U5110 ( .A1(n6346), .A2(n8304), .ZN(n4529) );
  INV_X1 U5111 ( .A(n7505), .ZN(n6548) );
  NAND2_X1 U5112 ( .A1(n6140), .A2(n6139), .ZN(n9911) );
  NAND2_X1 U5113 ( .A1(n8442), .A2(n9504), .ZN(n8304) );
  NAND2_X1 U5114 ( .A1(n6112), .A2(n6111), .ZN(n8442) );
  NAND2_X1 U5115 ( .A1(n7226), .A2(n7225), .ZN(n7224) );
  XNOR2_X1 U5116 ( .A(n4512), .B(n5353), .ZN(n6836) );
  NAND2_X1 U5117 ( .A1(n5337), .A2(n5336), .ZN(n4512) );
  NAND2_X1 U5118 ( .A1(n6073), .A2(n6072), .ZN(n9430) );
  INV_X1 U5119 ( .A(n5335), .ZN(n4514) );
  INV_X1 U5120 ( .A(n10179), .ZN(n7499) );
  NAND2_X1 U5121 ( .A1(n5986), .A2(n6304), .ZN(n7206) );
  AND2_X1 U5122 ( .A1(n4784), .A2(n4782), .ZN(n10179) );
  NAND2_X1 U5123 ( .A1(n5255), .A2(n5254), .ZN(n4948) );
  NAND2_X1 U5124 ( .A1(n4521), .A2(n5239), .ZN(n5255) );
  INV_X1 U5125 ( .A(n6066), .ZN(n9508) );
  NAND2_X2 U5126 ( .A1(n6947), .A2(n6946), .ZN(n7132) );
  AND4_X1 U5127 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n7273)
         );
  OAI211_X1 U5128 ( .C1(n5961), .C2(n6746), .A(n5948), .B(n5947), .ZN(n7219)
         );
  AND4_X1 U5129 ( .A1(n5148), .A2(n5147), .A3(n5146), .A4(n5145), .ZN(n6844)
         );
  OR2_X1 U5130 ( .A1(n6942), .A2(n6941), .ZN(n6947) );
  OAI211_X1 U5131 ( .C1(n5205), .C2(n6748), .A(n5165), .B(n5164), .ZN(n7067)
         );
  INV_X2 U5132 ( .A(n7233), .ZN(P1_U3973) );
  NAND4_X1 U5133 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n6991)
         );
  AND2_X1 U5134 ( .A1(n5196), .A2(n5195), .ZN(n4790) );
  OAI211_X1 U5135 ( .C1(n5205), .C2(n6745), .A(n5143), .B(n5142), .ZN(n7157)
         );
  OAI211_X1 U5136 ( .C1(n5205), .C2(n6746), .A(n5182), .B(n5181), .ZN(n10369)
         );
  NAND2_X2 U5137 ( .A1(n10028), .A2(n6452), .ZN(n5980) );
  XNOR2_X1 U5138 ( .A(n5673), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6943) );
  INV_X1 U5139 ( .A(n5334), .ZN(n4513) );
  NOR2_X1 U5140 ( .A1(n5275), .A2(n4947), .ZN(n4946) );
  AND2_X2 U5141 ( .A1(n5130), .A2(n9353), .ZN(n5636) );
  OR3_X2 U5142 ( .A1(n8303), .A2(n8178), .A3(n8216), .ZN(n6775) );
  INV_X1 U5143 ( .A(n5130), .ZN(n8501) );
  NAND2_X1 U5144 ( .A1(n4524), .A2(n5176), .ZN(n4937) );
  NAND2_X1 U5145 ( .A1(n5041), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U5146 ( .A(n5747), .B(n5746), .ZN(n6759) );
  XNOR2_X1 U5147 ( .A(n5124), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U5148 ( .A1(n5833), .A2(n5832), .ZN(n9950) );
  NAND2_X1 U5149 ( .A1(n6150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4747) );
  NAND2_X1 U5150 ( .A1(n5824), .A2(n5823), .ZN(n10028) );
  NAND2_X1 U5151 ( .A1(n5225), .A2(n5228), .ZN(n4522) );
  NAND2_X1 U5152 ( .A1(n5755), .A2(n5754), .ZN(n8181) );
  NAND2_X1 U5153 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5747) );
  AND2_X1 U5154 ( .A1(n5751), .A2(n5750), .ZN(n8243) );
  NAND2_X1 U5155 ( .A1(n4525), .A2(n5161), .ZN(n5174) );
  NAND2_X1 U5156 ( .A1(n5832), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U5157 ( .A1(n5831), .A2(n5830), .ZN(n5833) );
  NAND2_X1 U5158 ( .A1(n5034), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5135) );
  XNOR2_X1 U5159 ( .A(n6380), .B(n6379), .ZN(n7352) );
  AND2_X1 U5160 ( .A1(n6454), .A2(n5089), .ZN(n5829) );
  OR2_X1 U5161 ( .A1(n5122), .A2(n4560), .ZN(n4711) );
  NAND2_X1 U5162 ( .A1(n5916), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5879) );
  INV_X1 U5163 ( .A(n5038), .ZN(n5037) );
  NAND2_X1 U5164 ( .A1(n5162), .A2(n5137), .ZN(n5978) );
  AND2_X1 U5165 ( .A1(n5809), .A2(n6379), .ZN(n5074) );
  AND4_X1 U5166 ( .A1(n4989), .A2(n5118), .A3(n4991), .A4(n5303), .ZN(n4988)
         );
  AND2_X1 U5167 ( .A1(n5466), .A2(n5423), .ZN(n4991) );
  AND3_X1 U5168 ( .A1(n5422), .A2(n4708), .A3(n5675), .ZN(n4989) );
  NAND2_X1 U5169 ( .A1(n5827), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5830) );
  INV_X1 U5170 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5466) );
  AND2_X1 U5171 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4519) );
  INV_X1 U5172 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9634) );
  INV_X4 U5173 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5174 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6298) );
  NOR2_X1 U5175 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5112) );
  NOR2_X1 U5176 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5113) );
  INV_X1 U5177 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5423) );
  INV_X1 U5178 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5422) );
  OAI21_X2 U5179 ( .B1(n5320), .B2(n5319), .A(n5318), .ZN(n5335) );
  OAI21_X1 U5180 ( .B1(n5162), .B2(n4519), .A(n4517), .ZN(n5158) );
  NAND2_X1 U5181 ( .A1(n5162), .A2(n4518), .ZN(n4517) );
  INV_X1 U5182 ( .A(n5137), .ZN(n4518) );
  NAND2_X2 U5183 ( .A1(n4951), .A2(n4949), .ZN(n5162) );
  NAND3_X1 U5184 ( .A1(n4523), .A2(n5236), .A3(n4522), .ZN(n4521) );
  NAND2_X1 U5185 ( .A1(n4563), .A2(n5204), .ZN(n4523) );
  NAND2_X1 U5186 ( .A1(n5201), .A2(n5200), .ZN(n5204) );
  NAND2_X1 U5187 ( .A1(n5174), .A2(n5173), .ZN(n4524) );
  NAND2_X1 U5188 ( .A1(n5157), .A2(SI_1_), .ZN(n4525) );
  NAND2_X1 U5189 ( .A1(n10113), .A2(n7352), .ZN(n6989) );
  NAND2_X4 U5190 ( .A1(n6775), .A2(n6502), .ZN(n6503) );
  AOI21_X2 U5191 ( .B1(n7547), .B2(n7546), .A(n7545), .ZN(n7566) );
  NAND2_X2 U5192 ( .A1(n7308), .A2(n7307), .ZN(n7547) );
  XNOR2_X2 U5193 ( .A(n9293), .B(n8843), .ZN(n9121) );
  OAI211_X2 U5194 ( .C1(n8859), .C2(n5046), .A(n5045), .B(n5047), .ZN(n8941)
         );
  XNOR2_X2 U5195 ( .A(n8829), .B(n8828), .ZN(n8859) );
  INV_X1 U5196 ( .A(n7132), .ZN(n4526) );
  INV_X1 U5197 ( .A(n8838), .ZN(n4527) );
  NAND2_X1 U5198 ( .A1(n5259), .A2(n5258), .ZN(n5274) );
  NOR2_X1 U5199 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5803) );
  NOR2_X1 U5200 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5804) );
  AND2_X1 U5201 ( .A1(n4992), .A2(n5120), .ZN(n4985) );
  INV_X1 U5202 ( .A(n9950), .ZN(n5834) );
  OAI21_X1 U5203 ( .B1(n5501), .B2(n5502), .A(n5503), .ZN(n5514) );
  INV_X1 U5204 ( .A(n10348), .ZN(n10326) );
  NAND2_X2 U5205 ( .A1(n8607), .A2(n5735), .ZN(n10350) );
  AND2_X1 U5206 ( .A1(n7369), .A2(n9858), .ZN(n5088) );
  AOI21_X1 U5207 ( .B1(n4739), .B2(n6032), .A(n4575), .ZN(n4738) );
  NAND2_X1 U5208 ( .A1(n8694), .A2(n5000), .ZN(n4999) );
  NAND2_X1 U5209 ( .A1(n8687), .A2(n4565), .ZN(n4998) );
  AOI211_X1 U5210 ( .C1(n6122), .C2(n8116), .A(n4830), .B(n6121), .ZN(n4749)
         );
  NOR2_X1 U5211 ( .A1(n5443), .A2(SI_16_), .ZN(n5442) );
  INV_X1 U5212 ( .A(n5437), .ZN(n5443) );
  NAND2_X1 U5213 ( .A1(n9054), .A2(n4726), .ZN(n9059) );
  NAND2_X1 U5214 ( .A1(n9055), .A2(n9067), .ZN(n4726) );
  INV_X1 U5215 ( .A(n5722), .ZN(n4803) );
  OR2_X1 U5216 ( .A1(n6599), .A2(n6598), .ZN(n6601) );
  AND2_X1 U5217 ( .A1(n8518), .A2(n6597), .ZN(n6598) );
  OR2_X1 U5218 ( .A1(n5783), .A2(n5671), .ZN(n8791) );
  NAND2_X1 U5219 ( .A1(n5731), .A2(n8843), .ZN(n4808) );
  NAND2_X1 U5220 ( .A1(n4809), .A2(n4806), .ZN(n4805) );
  INV_X1 U5221 ( .A(n4810), .ZN(n4806) );
  OR2_X1 U5222 ( .A1(n5730), .A2(n5732), .ZN(n4804) );
  OR2_X1 U5223 ( .A1(n9293), .A2(n8843), .ZN(n8738) );
  NOR2_X1 U5224 ( .A1(n9299), .A2(n9143), .ZN(n8734) );
  NOR2_X1 U5225 ( .A1(n4822), .A2(n5726), .ZN(n4820) );
  NAND2_X1 U5226 ( .A1(n8923), .A2(n9188), .ZN(n4826) );
  OR2_X1 U5227 ( .A1(n9324), .A2(n9188), .ZN(n8718) );
  OR2_X1 U5228 ( .A1(n9191), .A2(n8825), .ZN(n8716) );
  NAND2_X1 U5229 ( .A1(n4817), .A2(n4532), .ZN(n4816) );
  INV_X1 U5230 ( .A(n8471), .ZN(n4817) );
  OR2_X1 U5231 ( .A1(n8231), .A2(n5719), .ZN(n5721) );
  NOR3_X1 U5232 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5121) );
  INV_X1 U5233 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5357) );
  NOR2_X1 U5234 ( .A1(n5179), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4986) );
  INV_X1 U5235 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U5236 ( .A1(n8415), .A2(n6575), .ZN(n8421) );
  OR3_X1 U5237 ( .A1(n6443), .A2(n6372), .A3(n6326), .ZN(n6375) );
  NAND2_X1 U5238 ( .A1(n6276), .A2(n6275), .ZN(n6285) );
  OR2_X1 U5239 ( .A1(n6274), .A2(n6273), .ZN(n6275) );
  OR2_X1 U5240 ( .A1(n6272), .A2(n7697), .ZN(n6276) );
  NAND2_X1 U5241 ( .A1(n4613), .A2(n5587), .ZN(n5605) );
  NAND2_X1 U5242 ( .A1(n4622), .A2(n4621), .ZN(n5515) );
  AOI21_X1 U5243 ( .B1(n5502), .B2(n5503), .A(SI_20_), .ZN(n4621) );
  NAND2_X1 U5244 ( .A1(n5501), .A2(n5503), .ZN(n4622) );
  OAI21_X1 U5245 ( .B1(n5462), .B2(n5461), .A(n5460), .ZN(n5481) );
  INV_X1 U5246 ( .A(n5316), .ZN(n5319) );
  NAND2_X1 U5247 ( .A1(n5274), .A2(n5261), .ZN(n5275) );
  NAND2_X1 U5248 ( .A1(n8915), .A2(n8827), .ZN(n8829) );
  NAND2_X1 U5249 ( .A1(n5059), .A2(n8814), .ZN(n5058) );
  INV_X1 U5250 ( .A(n5056), .ZN(n5055) );
  OAI21_X1 U5251 ( .B1(n4542), .B2(n4528), .A(n8925), .ZN(n5056) );
  NOR2_X1 U5252 ( .A1(n4545), .A2(n8828), .ZN(n5042) );
  OAI22_X1 U5253 ( .A1(n8883), .A2(n5050), .B1(n9153), .B2(n8833), .ZN(n5048)
         );
  INV_X1 U5254 ( .A(n5636), .ZN(n5287) );
  CLKBUF_X1 U5255 ( .A(n5188), .Z(n5683) );
  NAND2_X1 U5256 ( .A1(n5130), .A2(n5132), .ZN(n5218) );
  OR2_X1 U5257 ( .A1(n7017), .A2(n7016), .ZN(n4710) );
  AND2_X1 U5258 ( .A1(n8508), .A2(n8541), .ZN(n8685) );
  XNOR2_X1 U5259 ( .A(n9114), .B(n9123), .ZN(n9104) );
  OR2_X1 U5260 ( .A1(n4553), .A2(n7491), .ZN(n4902) );
  NAND2_X1 U5261 ( .A1(n4598), .A2(n6647), .ZN(n4881) );
  INV_X1 U5262 ( .A(n7352), .ZN(n9857) );
  AND4_X1 U5263 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n7213)
         );
  AOI21_X1 U5264 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n10027), .A(n10023), .ZN(
        n9520) );
  NAND2_X1 U5265 ( .A1(n4765), .A2(n4763), .ZN(n9699) );
  AOI21_X1 U5266 ( .B1(n9718), .B2(n4764), .A(n4572), .ZN(n4763) );
  INV_X1 U5267 ( .A(n4766), .ZN(n4764) );
  OAI21_X1 U5268 ( .B1(n9743), .B2(n4848), .A(n4847), .ZN(n9719) );
  NAND2_X1 U5269 ( .A1(n6429), .A2(n6360), .ZN(n4848) );
  NAND2_X1 U5270 ( .A1(n9729), .A2(n6429), .ZN(n4847) );
  INV_X1 U5271 ( .A(n4833), .ZN(n4832) );
  OAI21_X1 U5272 ( .B1(n9674), .B2(n4834), .A(n9792), .ZN(n4833) );
  OR2_X1 U5273 ( .A1(n9916), .A2(n9501), .ZN(n8485) );
  AND2_X1 U5274 ( .A1(n8018), .A2(n4547), .ZN(n4775) );
  INV_X1 U5275 ( .A(n5091), .ZN(n4837) );
  NAND2_X1 U5276 ( .A1(n5895), .A2(n5812), .ZN(n4838) );
  OAI21_X1 U5277 ( .B1(n5514), .B2(n5513), .A(n5512), .ZN(n5516) );
  XNOR2_X1 U5278 ( .A(n5399), .B(n5398), .ZN(n6968) );
  AND2_X1 U5279 ( .A1(n4713), .A2(n4714), .ZN(n4712) );
  NAND3_X1 U5280 ( .A1(n5739), .A2(n5738), .A3(n5737), .ZN(n8806) );
  OR2_X1 U5281 ( .A1(n8813), .A2(n10353), .ZN(n5739) );
  NAND2_X1 U5282 ( .A1(n9285), .A2(n10440), .ZN(n9236) );
  OR2_X1 U5283 ( .A1(n8643), .A2(n8642), .ZN(n4678) );
  AOI21_X1 U5284 ( .B1(n6038), .B2(n5088), .A(n4731), .ZN(n4730) );
  NAND2_X1 U5285 ( .A1(n4735), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U5286 ( .A1(n6037), .A2(n5088), .ZN(n4732) );
  INV_X1 U5287 ( .A(n4738), .ZN(n4737) );
  OAI21_X1 U5288 ( .B1(n4672), .B2(n4669), .A(n4533), .ZN(n5020) );
  NOR2_X1 U5289 ( .A1(n9177), .A2(n5019), .ZN(n5018) );
  AND2_X1 U5290 ( .A1(n8717), .A2(n8753), .ZN(n5019) );
  NOR2_X1 U5291 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  AOI21_X1 U5292 ( .B1(n4661), .B2(n8748), .A(n9147), .ZN(n4660) );
  NAND2_X1 U5293 ( .A1(n4662), .A2(n8762), .ZN(n4661) );
  OAI21_X1 U5294 ( .B1(n8727), .B2(n8726), .A(n4663), .ZN(n4662) );
  NAND2_X1 U5295 ( .A1(n8728), .A2(n8753), .ZN(n4666) );
  INV_X1 U5296 ( .A(n8727), .ZN(n8725) );
  AOI21_X1 U5297 ( .B1(n4630), .B2(n5646), .A(n4629), .ZN(n4628) );
  INV_X1 U5298 ( .A(n5659), .ZN(n4629) );
  INV_X1 U5299 ( .A(n5646), .ZN(n4626) );
  INV_X1 U5300 ( .A(n6575), .ZN(n4898) );
  INV_X1 U5301 ( .A(n6600), .ZN(n4899) );
  OR2_X1 U5302 ( .A1(n7392), .A2(n9857), .ZN(n6505) );
  NAND2_X1 U5303 ( .A1(n4866), .A2(n9739), .ZN(n4865) );
  INV_X1 U5304 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4950) );
  INV_X1 U5305 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4953) );
  OR2_X1 U5306 ( .A1(n10417), .A2(n8168), .ZN(n8667) );
  OR2_X1 U5307 ( .A1(n6897), .A2(n10286), .ZN(n4926) );
  NAND2_X1 U5308 ( .A1(n4917), .A2(n7032), .ZN(n4918) );
  INV_X1 U5309 ( .A(n7023), .ZN(n4917) );
  NAND3_X1 U5310 ( .A1(n10296), .A2(n4918), .A3(P2_REG1_REG_5__SCAN_IN), .ZN(
        n10298) );
  OR2_X1 U5311 ( .A1(n7036), .A2(n7257), .ZN(n4707) );
  INV_X1 U5312 ( .A(n9000), .ZN(n4929) );
  AND2_X1 U5313 ( .A1(n5522), .A2(n7923), .ZN(n5524) );
  OR2_X1 U5314 ( .A1(n9334), .A2(n9219), .ZN(n8714) );
  NAND2_X1 U5315 ( .A1(n10375), .A2(n8647), .ZN(n7237) );
  OAI22_X1 U5316 ( .A1(n5184), .A2(n5218), .B1(n5188), .B2(n7020), .ZN(n4789)
         );
  NAND2_X1 U5317 ( .A1(n5692), .A2(n7157), .ZN(n8615) );
  OR2_X1 U5318 ( .A1(n9317), .A2(n8919), .ZN(n8764) );
  NAND2_X1 U5319 ( .A1(n4997), .A2(n8710), .ZN(n4995) );
  NOR2_X1 U5320 ( .A1(n8717), .A2(n8711), .ZN(n4996) );
  AND2_X1 U5321 ( .A1(n8924), .A2(n9218), .ZN(n8690) );
  OR2_X1 U5322 ( .A1(n9339), .A2(n8934), .ZN(n8707) );
  INV_X1 U5323 ( .A(n8671), .ZN(n5005) );
  NOR2_X1 U5324 ( .A1(n8780), .A2(n5007), .ZN(n5006) );
  INV_X1 U5325 ( .A(n8665), .ZN(n5007) );
  AND2_X1 U5326 ( .A1(n5486), .A2(n5040), .ZN(n5039) );
  OR2_X1 U5327 ( .A1(n5179), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5198) );
  OR2_X1 U5328 ( .A1(n6606), .A2(n6605), .ZN(n6608) );
  INV_X1 U5329 ( .A(n7491), .ZN(n4901) );
  INV_X1 U5330 ( .A(n4891), .ZN(n4890) );
  OAI21_X1 U5331 ( .B1(n9390), .B2(n4892), .A(n9404), .ZN(n4891) );
  NAND2_X1 U5332 ( .A1(n4956), .A2(n6328), .ZN(n6443) );
  AND2_X1 U5333 ( .A1(n4957), .A2(n9636), .ZN(n6372) );
  OR2_X1 U5334 ( .A1(n9870), .A2(n9721), .ZN(n6329) );
  OR2_X1 U5335 ( .A1(n9874), .A2(n9732), .ZN(n6352) );
  OR2_X1 U5336 ( .A1(n9879), .A2(n9748), .ZN(n6351) );
  AND2_X1 U5337 ( .A1(n9652), .A2(n4546), .ZN(n4780) );
  NOR2_X1 U5338 ( .A1(n9850), .A2(n9645), .ZN(n4860) );
  OAI21_X1 U5339 ( .B1(n8488), .B2(n4849), .A(n4573), .ZN(n9832) );
  NAND2_X1 U5340 ( .A1(n4850), .A2(n6423), .ZN(n4849) );
  NAND2_X1 U5341 ( .A1(n4551), .A2(n6423), .ZN(n4852) );
  OR2_X1 U5342 ( .A1(n4757), .A2(n4549), .ZN(n4755) );
  OR2_X1 U5343 ( .A1(n9990), .A2(n9430), .ZN(n8016) );
  NAND2_X1 U5344 ( .A1(n9509), .A2(n10179), .ZN(n6065) );
  NOR2_X1 U5345 ( .A1(n4871), .A2(n10083), .ZN(n4870) );
  INV_X1 U5346 ( .A(n7332), .ZN(n4869) );
  NAND2_X1 U5347 ( .A1(n9778), .A2(n9770), .ZN(n9764) );
  NAND2_X1 U5348 ( .A1(n4612), .A2(n5606), .ZN(n5622) );
  NAND2_X1 U5349 ( .A1(n5569), .A2(n5568), .ZN(n5586) );
  NAND2_X1 U5350 ( .A1(n4634), .A2(n4632), .ZN(n5569) );
  AOI21_X1 U5351 ( .B1(n4539), .B2(n5552), .A(n4633), .ZN(n4632) );
  OAI21_X1 U5352 ( .B1(n5481), .B2(n5480), .A(n5479), .ZN(n5501) );
  NAND2_X1 U5353 ( .A1(n4967), .A2(n4969), .ZN(n4964) );
  INV_X1 U5354 ( .A(n4620), .ZN(n5441) );
  AND2_X1 U5355 ( .A1(n5413), .A2(n5414), .ZN(n5439) );
  AND2_X1 U5356 ( .A1(n5393), .A2(n5394), .ZN(n5413) );
  XNOR2_X1 U5357 ( .A(n5354), .B(n5338), .ZN(n5353) );
  NAND2_X1 U5358 ( .A1(n5336), .A2(n5323), .ZN(n5334) );
  OAI21_X1 U5359 ( .B1(n4948), .B2(n4945), .A(n4943), .ZN(n5301) );
  INV_X1 U5360 ( .A(n4944), .ZN(n4943) );
  OAI21_X1 U5361 ( .B1(n4946), .B2(n4945), .A(n5100), .ZN(n4944) );
  XNOR2_X1 U5362 ( .A(n5256), .B(SI_7_), .ZN(n5253) );
  XNOR2_X1 U5363 ( .A(n5238), .B(SI_6_), .ZN(n5235) );
  INV_X1 U5364 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4741) );
  OAI21_X1 U5365 ( .B1(n5162), .B2(n5139), .A(n5138), .ZN(n5160) );
  NAND2_X1 U5366 ( .A1(n5162), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5138) );
  NOR2_X1 U5367 ( .A1(n5069), .A2(n5068), .ZN(n5067) );
  INV_X1 U5368 ( .A(n7565), .ZN(n5068) );
  AND2_X1 U5369 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  NOR2_X1 U5370 ( .A1(n7540), .A2(n7550), .ZN(n7544) );
  AND2_X1 U5371 ( .A1(n8165), .A2(n8965), .ZN(n5069) );
  AND2_X1 U5372 ( .A1(n8798), .A2(n8797), .ZN(n4683) );
  AND2_X1 U5373 ( .A1(n5032), .A2(n5136), .ZN(n5031) );
  NAND2_X1 U5374 ( .A1(n5636), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5147) );
  OR2_X1 U5375 ( .A1(n10289), .A2(n10290), .ZN(n4719) );
  NOR2_X1 U5376 ( .A1(n7461), .A2(n7460), .ZN(n7462) );
  NOR2_X1 U5377 ( .A1(n7466), .A2(n5269), .ZN(n7460) );
  NAND2_X1 U5378 ( .A1(n4723), .A2(n4725), .ZN(n4722) );
  INV_X1 U5379 ( .A(n7481), .ZN(n4725) );
  XNOR2_X1 U5380 ( .A(n8138), .B(n8147), .ZN(n8045) );
  NAND2_X1 U5381 ( .A1(n8045), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U5382 ( .A1(n8198), .A2(n8199), .ZN(n8369) );
  NOR2_X1 U5383 ( .A1(n9084), .A2(n9060), .ZN(n9061) );
  NOR2_X1 U5384 ( .A1(n4568), .A2(n5061), .ZN(n5060) );
  INV_X1 U5385 ( .A(n5062), .ZN(n5061) );
  AOI21_X1 U5386 ( .B1(n5729), .B2(n5728), .A(n5727), .ZN(n9140) );
  NAND2_X1 U5387 ( .A1(n9311), .A2(n9167), .ZN(n5728) );
  INV_X1 U5388 ( .A(n5597), .ZN(n5596) );
  INV_X1 U5389 ( .A(n8714), .ZN(n4997) );
  NOR2_X1 U5390 ( .A1(n9200), .A2(n9199), .ZN(n9202) );
  OR2_X1 U5391 ( .A1(n5473), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5493) );
  OR2_X1 U5392 ( .A1(n5430), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5455) );
  NOR2_X1 U5393 ( .A1(n8336), .A2(n8229), .ZN(n5014) );
  OR2_X1 U5394 ( .A1(n5327), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5346) );
  AND2_X1 U5395 ( .A1(n5314), .A2(n8639), .ZN(n5008) );
  OR2_X1 U5396 ( .A1(n5308), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5327) );
  OR2_X1 U5397 ( .A1(n10403), .A2(n7567), .ZN(n8639) );
  AND2_X1 U5398 ( .A1(n5691), .A2(n5690), .ZN(n5707) );
  INV_X1 U5399 ( .A(n4978), .ZN(n4977) );
  OAI21_X1 U5400 ( .B1(n4981), .B2(n8653), .A(n8657), .ZN(n4978) );
  OR2_X1 U5401 ( .A1(n5106), .A2(n5689), .ZN(n7430) );
  AND2_X1 U5402 ( .A1(n7320), .A2(n5688), .ZN(n5689) );
  OR2_X1 U5403 ( .A1(n10400), .A2(n8967), .ZN(n5688) );
  OR2_X1 U5404 ( .A1(n5267), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5291) );
  OR2_X1 U5405 ( .A1(n5219), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U5406 ( .A1(n5186), .A2(n5185), .ZN(n5212) );
  INV_X1 U5407 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5186) );
  INV_X1 U5408 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U5409 ( .A1(n5211), .A2(n5210), .ZN(n5219) );
  INV_X1 U5410 ( .A(n5212), .ZN(n5211) );
  NAND2_X1 U5411 ( .A1(n8620), .A2(n8619), .ZN(n10344) );
  NAND2_X1 U5412 ( .A1(n5665), .A2(n5664), .ZN(n5783) );
  NAND2_X1 U5413 ( .A1(n5643), .A2(n8738), .ZN(n9103) );
  INV_X1 U5414 ( .A(n5024), .ZN(n5023) );
  NOR2_X1 U5415 ( .A1(n8734), .A2(n5025), .ZN(n5024) );
  INV_X1 U5416 ( .A(n8731), .ZN(n5025) );
  OR2_X1 U5417 ( .A1(n9305), .A2(n8949), .ZN(n8731) );
  NAND2_X1 U5418 ( .A1(n9146), .A2(n8732), .ZN(n5026) );
  AND2_X1 U5419 ( .A1(n4826), .A2(n4827), .ZN(n4821) );
  NAND2_X1 U5420 ( .A1(n4576), .A2(n4826), .ZN(n4822) );
  NAND2_X1 U5421 ( .A1(n9189), .A2(n4827), .ZN(n4824) );
  AND2_X1 U5422 ( .A1(n8764), .A2(n9158), .ZN(n9165) );
  NAND2_X1 U5423 ( .A1(n4828), .A2(n8825), .ZN(n4827) );
  AND2_X1 U5424 ( .A1(n4816), .A2(n4555), .ZN(n9217) );
  NAND2_X1 U5425 ( .A1(n4816), .A2(n4815), .ZN(n9215) );
  INV_X1 U5426 ( .A(n4802), .ZN(n4801) );
  OR2_X1 U5427 ( .A1(n8889), .A2(n8815), .ZN(n8468) );
  NAND2_X1 U5428 ( .A1(n5721), .A2(n5720), .ZN(n8337) );
  NAND2_X1 U5429 ( .A1(n8685), .A2(n8691), .ZN(n5013) );
  NAND2_X1 U5430 ( .A1(n5429), .A2(n5428), .ZN(n9274) );
  NAND2_X1 U5431 ( .A1(n4793), .A2(n4794), .ZN(n8231) );
  AND2_X1 U5432 ( .A1(n4795), .A2(n5718), .ZN(n4794) );
  INV_X1 U5433 ( .A(n10346), .ZN(n10328) );
  NAND2_X1 U5434 ( .A1(n5361), .A2(n5360), .ZN(n5714) );
  AND4_X1 U5435 ( .A1(n5351), .A2(n5350), .A3(n5349), .A4(n5348), .ZN(n8668)
         );
  NAND2_X1 U5436 ( .A1(n5716), .A2(n5715), .ZN(n8182) );
  OR2_X1 U5437 ( .A1(n8748), .A2(n6938), .ZN(n10346) );
  NAND2_X1 U5438 ( .A1(n5333), .A2(n5006), .ZN(n8089) );
  XNOR2_X1 U5439 ( .A(n5128), .B(n5127), .ZN(n5132) );
  INV_X1 U5440 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U5441 ( .A1(n5122), .A2(n5121), .ZN(n5748) );
  AND2_X1 U5442 ( .A1(n5121), .A2(n5033), .ZN(n5032) );
  INV_X1 U5443 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5033) );
  NOR2_X1 U5444 ( .A1(n5116), .A2(n5179), .ZN(n5302) );
  XNOR2_X1 U5445 ( .A(n5163), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6903) );
  NAND2_X1 U5446 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6906), .ZN(n5163) );
  NAND2_X1 U5447 ( .A1(n9448), .A2(n6658), .ZN(n6659) );
  AND2_X1 U5448 ( .A1(n4601), .A2(n4881), .ZN(n4877) );
  INV_X1 U5449 ( .A(n6647), .ZN(n4880) );
  AND2_X1 U5450 ( .A1(n4881), .A2(n6636), .ZN(n4879) );
  INV_X1 U5451 ( .A(n9501), .ZN(n9395) );
  NAND2_X1 U5452 ( .A1(n9389), .A2(n9391), .ZN(n4893) );
  AND2_X1 U5453 ( .A1(n9424), .A2(n9426), .ZN(n6565) );
  NOR2_X1 U5454 ( .A1(n6640), .A2(n6641), .ZN(n4883) );
  NAND2_X1 U5455 ( .A1(n9455), .A2(n9458), .ZN(n4886) );
  NAND2_X1 U5456 ( .A1(n6637), .A2(n6636), .ZN(n9456) );
  INV_X1 U5457 ( .A(n9502), .ZN(n9489) );
  AND4_X1 U5458 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(n8123)
         );
  OR2_X1 U5459 ( .A1(n9520), .A2(n9519), .ZN(n4653) );
  NOR2_X1 U5460 ( .A1(n8261), .A2(n8260), .ZN(n9552) );
  NOR2_X1 U5461 ( .A1(n9552), .A2(n4649), .ZN(n9575) );
  AND2_X1 U5462 ( .A1(n9553), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4649) );
  AND2_X1 U5463 ( .A1(n6329), .A2(n9683), .ZN(n9702) );
  NOR2_X1 U5464 ( .A1(n9717), .A2(n9681), .ZN(n9703) );
  INV_X1 U5465 ( .A(n9663), .ZN(n4771) );
  NAND2_X1 U5466 ( .A1(n4767), .A2(n4768), .ZN(n4766) );
  NAND2_X1 U5467 ( .A1(n4769), .A2(n9665), .ZN(n4768) );
  INV_X1 U5468 ( .A(n9664), .ZN(n4767) );
  NAND2_X1 U5469 ( .A1(n6352), .A2(n9680), .ZN(n9718) );
  AND2_X1 U5470 ( .A1(n9889), .A2(n9658), .ZN(n9659) );
  NAND2_X1 U5471 ( .A1(n4835), .A2(n9674), .ZN(n9802) );
  INV_X1 U5472 ( .A(n9804), .ZN(n4835) );
  AOI21_X1 U5473 ( .B1(n9966), .B2(n9837), .A(n9647), .ZN(n9841) );
  NOR2_X1 U5474 ( .A1(n8552), .A2(n9645), .ZN(n9846) );
  NOR2_X1 U5475 ( .A1(n8488), .A2(n8547), .ZN(n4854) );
  OR2_X1 U5476 ( .A1(n4761), .A2(n4559), .ZN(n4757) );
  OR2_X1 U5477 ( .A1(n4759), .A2(n4559), .ZN(n4756) );
  INV_X1 U5478 ( .A(n4760), .ZN(n4759) );
  OAI21_X1 U5479 ( .B1(n4761), .B2(n8485), .A(n8547), .ZN(n4760) );
  AOI21_X1 U5480 ( .B1(n8292), .B2(n8291), .A(n8290), .ZN(n8312) );
  NAND2_X1 U5481 ( .A1(n4776), .A2(n4547), .ZN(n4774) );
  NAND2_X1 U5482 ( .A1(n4550), .A2(n8070), .ZN(n4776) );
  AOI21_X1 U5483 ( .B1(n8013), .B2(n8012), .A(n5096), .ZN(n8035) );
  NOR2_X1 U5484 ( .A1(n8011), .A2(n10069), .ZN(n5096) );
  AND2_X1 U5485 ( .A1(n10068), .A2(n10071), .ZN(n8013) );
  OR2_X1 U5486 ( .A1(n10073), .A2(n10067), .ZN(n10074) );
  NAND2_X1 U5487 ( .A1(n7215), .A2(n7214), .ZN(n7272) );
  NAND2_X1 U5488 ( .A1(n6992), .A2(n5983), .ZN(n10090) );
  NAND2_X1 U5489 ( .A1(n6390), .A2(n6304), .ZN(n10098) );
  NAND2_X1 U5490 ( .A1(n6306), .A2(n6993), .ZN(n6992) );
  INV_X1 U5491 ( .A(n9770), .ZN(n9889) );
  INV_X1 U5492 ( .A(n9645), .ZN(n9966) );
  XNOR2_X1 U5493 ( .A(n4963), .B(n6289), .ZN(n9345) );
  OAI21_X1 U5494 ( .B1(n6285), .B2(n6284), .A(n6283), .ZN(n4963) );
  XNOR2_X1 U5495 ( .A(n6285), .B(n6284), .ZN(n9351) );
  NOR2_X1 U5496 ( .A1(n5091), .A2(n5090), .ZN(n5089) );
  NAND2_X1 U5497 ( .A1(n5816), .A2(n6456), .ZN(n5090) );
  XNOR2_X1 U5498 ( .A(n5622), .B(n5621), .ZN(n8242) );
  NAND2_X1 U5499 ( .A1(n4959), .A2(n5533), .ZN(n5550) );
  NAND2_X1 U5500 ( .A1(n4960), .A2(n5516), .ZN(n4959) );
  NOR2_X2 U5501 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(n5810), .ZN(n5811) );
  XNOR2_X1 U5502 ( .A(n5374), .B(n4623), .ZN(n6965) );
  INV_X1 U5503 ( .A(n5391), .ZN(n4623) );
  INV_X1 U5504 ( .A(n4942), .ZN(n5299) );
  AOI21_X1 U5505 ( .B1(n4948), .B2(n4946), .A(n4945), .ZN(n4942) );
  XNOR2_X1 U5506 ( .A(n5276), .B(n5275), .ZN(n6771) );
  NAND2_X1 U5507 ( .A1(n4948), .A2(n5257), .ZN(n5276) );
  AOI21_X1 U5508 ( .B1(n5055), .B2(n4528), .A(n4599), .ZN(n5053) );
  INV_X1 U5509 ( .A(n8966), .ZN(n7567) );
  INV_X1 U5510 ( .A(n10327), .ZN(n7075) );
  INV_X1 U5511 ( .A(n9153), .ZN(n8949) );
  INV_X1 U5512 ( .A(n5048), .ZN(n5047) );
  OR2_X1 U5513 ( .A1(n4545), .A2(n9179), .ZN(n5046) );
  NAND2_X1 U5514 ( .A1(n5043), .A2(n5042), .ZN(n5045) );
  NAND2_X1 U5515 ( .A1(n4684), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U5516 ( .A1(n4686), .A2(n4685), .ZN(n4684) );
  NOR2_X1 U5517 ( .A1(n8796), .A2(n4683), .ZN(n4682) );
  NOR2_X1 U5518 ( .A1(n8758), .A2(n8759), .ZN(n4685) );
  XNOR2_X1 U5519 ( .A(n6885), .B(n6871), .ZN(n6886) );
  NOR2_X1 U5520 ( .A1(n10314), .A2(n7014), .ZN(n7017) );
  XNOR2_X1 U5521 ( .A(n7462), .B(n7468), .ZN(n7516) );
  OR2_X1 U5522 ( .A1(n8042), .A2(n10438), .ZN(n4923) );
  OAI21_X1 U5523 ( .B1(n9061), .B2(n4729), .A(n4728), .ZN(n4727) );
  NAND2_X1 U5524 ( .A1(n10272), .A2(n9083), .ZN(n4729) );
  AOI21_X1 U5525 ( .B1(n10248), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9065), .ZN(
        n4728) );
  NOR2_X1 U5526 ( .A1(n4696), .A2(n4690), .ZN(n4689) );
  NOR2_X1 U5527 ( .A1(n9051), .A2(n9050), .ZN(n9053) );
  NOR2_X1 U5528 ( .A1(n10283), .A2(n4910), .ZN(n4909) );
  INV_X1 U5529 ( .A(n4911), .ZN(n4910) );
  OAI21_X1 U5530 ( .B1(n9085), .B2(n9077), .A(n4912), .ZN(n4911) );
  INV_X1 U5531 ( .A(n9278), .ZN(n9100) );
  NAND2_X1 U5532 ( .A1(n5649), .A2(n5648), .ZN(n9114) );
  NOR2_X1 U5533 ( .A1(n8806), .A2(n5742), .ZN(n5802) );
  NAND2_X1 U5534 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  NAND2_X1 U5535 ( .A1(n9134), .A2(n10326), .ZN(n9108) );
  XOR2_X1 U5536 ( .A(n9104), .B(n9103), .Z(n9287) );
  INV_X1 U5537 ( .A(n9774), .ZN(n9894) );
  NAND2_X1 U5538 ( .A1(n8572), .A2(n6524), .ZN(n7175) );
  NAND2_X1 U5539 ( .A1(n6193), .A2(n6192), .ZN(n9906) );
  NAND2_X1 U5540 ( .A1(n6250), .A2(n6249), .ZN(n9884) );
  INV_X1 U5541 ( .A(n9790), .ZN(n9900) );
  INV_X1 U5542 ( .A(n9739), .ZN(n9879) );
  NAND2_X1 U5543 ( .A1(n5883), .A2(n5882), .ZN(n9916) );
  OR3_X1 U5544 ( .A1(n6377), .A2(n6376), .A3(n6504), .ZN(n4939) );
  INV_X1 U5545 ( .A(n6804), .ZN(n10014) );
  AND2_X1 U5546 ( .A1(n5958), .A2(n5957), .ZN(n10027) );
  XNOR2_X1 U5547 ( .A(n9625), .B(n9843), .ZN(n4642) );
  NOR2_X1 U5548 ( .A1(n4548), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5549 ( .A1(n9629), .A2(n6504), .ZN(n4641) );
  OAI21_X1 U5550 ( .B1(n4638), .B2(n10022), .A(n4636), .ZN(n4635) );
  INV_X1 U5551 ( .A(n4637), .ZN(n4636) );
  INV_X1 U5552 ( .A(n4642), .ZN(n4638) );
  OAI21_X1 U5553 ( .B1(n9630), .B2(n9631), .A(n4507), .ZN(n4637) );
  OAI21_X1 U5554 ( .B1(n9636), .B2(n10219), .A(n9855), .ZN(n6475) );
  NAND2_X1 U5555 ( .A1(n9871), .A2(n4844), .ZN(n9926) );
  NOR2_X1 U5556 ( .A1(n9868), .A2(n4845), .ZN(n4844) );
  OR2_X1 U5557 ( .A1(n9869), .A2(n4846), .ZN(n4845) );
  INV_X1 U5558 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U5559 ( .A1(n8610), .A2(n8753), .ZN(n4976) );
  NAND2_X1 U5560 ( .A1(n8611), .A2(n8748), .ZN(n4975) );
  NAND2_X1 U5561 ( .A1(n4972), .A2(n4785), .ZN(n8628) );
  OAI21_X1 U5562 ( .B1(n8624), .B2(n4974), .A(n4973), .ZN(n4972) );
  NAND2_X1 U5563 ( .A1(n4976), .A2(n4975), .ZN(n4974) );
  INV_X1 U5564 ( .A(n8623), .ZN(n4973) );
  NAND2_X1 U5565 ( .A1(n4677), .A2(n4676), .ZN(n4675) );
  NOR2_X1 U5566 ( .A1(n4567), .A2(n8753), .ZN(n4676) );
  NAND2_X1 U5567 ( .A1(n4678), .A2(n4558), .ZN(n4677) );
  AND2_X1 U5568 ( .A1(n7369), .A2(n6307), .ZN(n4739) );
  INV_X1 U5569 ( .A(n8676), .ZN(n5027) );
  NOR2_X1 U5570 ( .A1(n8676), .A2(n5029), .ZN(n5028) );
  AOI21_X1 U5571 ( .B1(n4738), .B2(n4736), .A(n7382), .ZN(n4735) );
  INV_X1 U5572 ( .A(n4739), .ZN(n4736) );
  NAND2_X1 U5573 ( .A1(n4750), .A2(n5988), .ZN(n6002) );
  NAND2_X1 U5574 ( .A1(n5985), .A2(n5984), .ZN(n4750) );
  NOR2_X1 U5575 ( .A1(n5002), .A2(n5001), .ZN(n5000) );
  NAND2_X1 U5576 ( .A1(n8695), .A2(n8753), .ZN(n5001) );
  AOI21_X1 U5577 ( .B1(n4734), .B2(n5087), .A(n6082), .ZN(n6126) );
  INV_X1 U5578 ( .A(n6068), .ZN(n5087) );
  AOI21_X1 U5579 ( .B1(n8703), .B2(n8785), .A(n8702), .ZN(n8704) );
  INV_X1 U5580 ( .A(n8713), .ZN(n4673) );
  NAND2_X1 U5581 ( .A1(n6125), .A2(n9398), .ZN(n4748) );
  NOR2_X1 U5582 ( .A1(n4665), .A2(n4664), .ZN(n4663) );
  INV_X1 U5583 ( .A(n8764), .ZN(n4664) );
  INV_X1 U5584 ( .A(n8763), .ZN(n4665) );
  NAND2_X1 U5585 ( .A1(n5017), .A2(n5016), .ZN(n8727) );
  INV_X1 U5586 ( .A(n8722), .ZN(n5016) );
  NAND2_X1 U5587 ( .A1(n5020), .A2(n5018), .ZN(n5017) );
  NAND2_X1 U5588 ( .A1(n4659), .A2(n4658), .ZN(n8737) );
  AND2_X1 U5589 ( .A1(n9130), .A2(n8733), .ZN(n4658) );
  NAND2_X1 U5590 ( .A1(n4666), .A2(n4660), .ZN(n4659) );
  NAND2_X1 U5591 ( .A1(n10262), .A2(n6907), .ZN(n6909) );
  OR2_X1 U5592 ( .A1(n6568), .A2(n6567), .ZN(n6569) );
  INV_X1 U5593 ( .A(n9405), .ZN(n4892) );
  NOR2_X1 U5594 ( .A1(n4892), .A2(n4889), .ZN(n4888) );
  INV_X1 U5595 ( .A(n9391), .ZN(n4889) );
  NAND2_X1 U5596 ( .A1(n6471), .A2(n5984), .ZN(n5081) );
  INV_X1 U5597 ( .A(n6271), .ZN(n4616) );
  NOR2_X1 U5598 ( .A1(n6114), .A2(n6113), .ZN(n5906) );
  OAI21_X1 U5599 ( .B1(n5647), .B2(n4627), .A(n4625), .ZN(n6274) );
  AOI21_X1 U5600 ( .B1(n4628), .B2(n4626), .A(n4606), .ZN(n4625) );
  INV_X1 U5601 ( .A(n4628), .ZN(n4627) );
  INV_X1 U5602 ( .A(n5566), .ZN(n4633) );
  NOR2_X1 U5603 ( .A1(n4569), .A2(n4968), .ZN(n4967) );
  NOR2_X1 U5604 ( .A1(n4970), .A2(n4969), .ZN(n4968) );
  INV_X1 U5605 ( .A(n5355), .ZN(n4969) );
  INV_X1 U5606 ( .A(n5412), .ZN(n5415) );
  OR2_X1 U5607 ( .A1(n5392), .A2(n5391), .ZN(n5394) );
  NOR2_X1 U5608 ( .A1(n5356), .A2(n4971), .ZN(n4970) );
  INV_X1 U5609 ( .A(n5336), .ZN(n4971) );
  INV_X1 U5610 ( .A(n5353), .ZN(n5356) );
  INV_X1 U5611 ( .A(n8890), .ZN(n5059) );
  INV_X1 U5612 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4708) );
  OR2_X1 U5613 ( .A1(n6906), .A2(n4668), .ZN(n6894) );
  XNOR2_X1 U5614 ( .A(n6909), .B(n6908), .ZN(n10277) );
  AOI21_X1 U5615 ( .B1(n10298), .B2(n10296), .A(n10297), .ZN(n10295) );
  INV_X1 U5616 ( .A(n4724), .ZN(n4723) );
  AOI21_X1 U5617 ( .B1(n7474), .B2(n7521), .A(n7475), .ZN(n4724) );
  NAND2_X1 U5618 ( .A1(n8043), .A2(n4604), .ZN(n8138) );
  INV_X1 U5619 ( .A(n9059), .ZN(n9056) );
  AND2_X1 U5620 ( .A1(n5357), .A2(n5375), .ZN(n5062) );
  OR2_X1 U5621 ( .A1(n5704), .A2(n7430), .ZN(n5691) );
  NAND2_X1 U5622 ( .A1(n8633), .A2(n4982), .ZN(n4981) );
  NAND2_X1 U5623 ( .A1(n8653), .A2(n4983), .ZN(n4982) );
  INV_X1 U5624 ( .A(n8652), .ZN(n4983) );
  INV_X1 U5625 ( .A(n4981), .ZN(n4980) );
  OR2_X1 U5626 ( .A1(n8653), .A2(n5106), .ZN(n7428) );
  OAI21_X1 U5627 ( .B1(n7255), .B2(n7250), .A(n7249), .ZN(n7429) );
  AND2_X1 U5628 ( .A1(n7144), .A2(n5698), .ZN(n5697) );
  AND2_X1 U5629 ( .A1(n8767), .A2(n7143), .ZN(n7144) );
  NAND2_X1 U5630 ( .A1(n7075), .A2(n7067), .ZN(n8620) );
  NAND2_X1 U5631 ( .A1(n5024), .A2(n5022), .ZN(n5021) );
  INV_X1 U5632 ( .A(n8732), .ZN(n5022) );
  AND2_X1 U5633 ( .A1(n8731), .A2(n8732), .ZN(n8729) );
  OR2_X1 U5634 ( .A1(n9311), .A2(n9142), .ZN(n8763) );
  AND2_X1 U5635 ( .A1(n8699), .A2(n8468), .ZN(n8785) );
  OAI21_X1 U5636 ( .B1(n8336), .B2(n4803), .A(n8696), .ZN(n4802) );
  NOR2_X1 U5637 ( .A1(n4803), .A2(n4799), .ZN(n4798) );
  INV_X1 U5638 ( .A(n5720), .ZN(n4799) );
  NOR2_X1 U5639 ( .A1(n8777), .A2(n4796), .ZN(n4792) );
  INV_X1 U5640 ( .A(n5717), .ZN(n4796) );
  NAND2_X1 U5641 ( .A1(n5717), .A2(n5029), .ZN(n4795) );
  OAI21_X1 U5642 ( .B1(n5039), .B2(n9346), .A(n5675), .ZN(n5038) );
  OR2_X1 U5643 ( .A1(n5240), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5283) );
  INV_X1 U5644 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U5645 ( .A1(n6600), .A2(n4898), .ZN(n4897) );
  OR2_X1 U5646 ( .A1(n9636), .A2(n4957), .ZN(n4956) );
  NAND2_X1 U5647 ( .A1(n4745), .A2(n4742), .ZN(n5075) );
  NOR2_X1 U5648 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  INV_X1 U5649 ( .A(n6270), .ZN(n4744) );
  OR2_X1 U5650 ( .A1(n6471), .A2(n9858), .ZN(n5078) );
  NAND2_X1 U5651 ( .A1(n5079), .A2(n4615), .ZN(n4614) );
  INV_X1 U5652 ( .A(n5080), .ZN(n5079) );
  NAND2_X1 U5653 ( .A1(n4616), .A2(n4530), .ZN(n4615) );
  OAI21_X1 U5654 ( .B1(n6270), .B2(n6471), .A(n5081), .ZN(n5080) );
  NOR2_X1 U5655 ( .A1(n9870), .A2(n4865), .ZN(n4864) );
  NAND2_X1 U5656 ( .A1(n5825), .A2(n6191), .ZN(n4619) );
  NAND2_X1 U5657 ( .A1(n4619), .A2(n4617), .ZN(n6330) );
  NOR2_X1 U5658 ( .A1(n7234), .A2(n4618), .ZN(n4617) );
  INV_X1 U5659 ( .A(n5826), .ZN(n4618) );
  INV_X1 U5660 ( .A(n9662), .ZN(n4769) );
  OR2_X1 U5661 ( .A1(n9884), .A2(n9763), .ZN(n6335) );
  OR2_X1 U5662 ( .A1(n9889), .A2(n9747), .ZN(n9677) );
  INV_X1 U5663 ( .A(n6226), .ZN(n6216) );
  NAND2_X1 U5664 ( .A1(n9955), .A2(n4860), .ZN(n4859) );
  OR2_X1 U5665 ( .A1(n8553), .A2(n9911), .ZN(n8552) );
  OR2_X1 U5666 ( .A1(n5908), .A2(n5888), .ZN(n5890) );
  NOR2_X1 U5667 ( .A1(n8442), .A2(n8528), .ZN(n4856) );
  NAND2_X1 U5668 ( .A1(n9508), .A2(n10187), .ZN(n8006) );
  NOR2_X1 U5669 ( .A1(n6007), .A2(n6006), .ZN(n6005) );
  INV_X1 U5670 ( .A(n4865), .ZN(n4863) );
  NOR2_X1 U5671 ( .A1(n9764), .A2(n9884), .ZN(n9749) );
  AND2_X1 U5672 ( .A1(n9787), .A2(n9894), .ZN(n9778) );
  NAND2_X1 U5673 ( .A1(n8127), .A2(n10213), .ZN(n8314) );
  NOR2_X1 U5674 ( .A1(n10074), .A2(n9430), .ZN(n8029) );
  XNOR2_X1 U5675 ( .A(n6274), .B(n6273), .ZN(n6272) );
  INV_X1 U5676 ( .A(n5645), .ZN(n4630) );
  INV_X1 U5677 ( .A(n5644), .ZN(n5647) );
  NAND2_X1 U5678 ( .A1(n5093), .A2(n5092), .ZN(n5091) );
  INV_X1 U5679 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5092) );
  INV_X1 U5680 ( .A(n5814), .ZN(n5093) );
  NAND2_X1 U5681 ( .A1(n5624), .A2(n5623), .ZN(n5644) );
  NAND2_X1 U5682 ( .A1(n5622), .A2(n5621), .ZN(n5624) );
  NAND2_X1 U5683 ( .A1(n5895), .A2(n4840), .ZN(n4839) );
  AND2_X1 U5684 ( .A1(n5812), .A2(n6456), .ZN(n4840) );
  AND3_X1 U5685 ( .A1(n6298), .A2(n6446), .A3(n5873), .ZN(n5812) );
  INV_X1 U5686 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U5687 ( .A1(n5867), .A2(n7748), .ZN(n5916) );
  XNOR2_X1 U5688 ( .A(n5390), .B(n4624), .ZN(n5391) );
  INV_X1 U5689 ( .A(SI_14_), .ZN(n4624) );
  INV_X1 U5690 ( .A(n5371), .ZN(n5393) );
  XNOR2_X1 U5691 ( .A(n5372), .B(SI_13_), .ZN(n5371) );
  XNOR2_X1 U5692 ( .A(n5317), .B(n7727), .ZN(n5316) );
  INV_X1 U5693 ( .A(n5257), .ZN(n4947) );
  INV_X1 U5694 ( .A(n5274), .ZN(n4945) );
  INV_X1 U5695 ( .A(n5805), .ZN(n4740) );
  NAND2_X1 U5696 ( .A1(n5804), .A2(n5803), .ZN(n5994) );
  OAI21_X1 U5697 ( .B1(n6738), .B2(n5178), .A(n5177), .ZN(n5190) );
  NAND2_X1 U5698 ( .A1(n6738), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5177) );
  INV_X1 U5699 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4952) );
  NAND2_X1 U5700 ( .A1(n8537), .A2(n8534), .ZN(n8892) );
  XNOR2_X1 U5701 ( .A(n7157), .B(n7132), .ZN(n6950) );
  INV_X1 U5702 ( .A(n8902), .ZN(n5049) );
  AND2_X1 U5703 ( .A1(n6939), .A2(n6937), .ZN(n8944) );
  NAND2_X1 U5704 ( .A1(n8760), .A2(n8761), .ZN(n4686) );
  OR2_X1 U5705 ( .A1(n5032), .A2(n4560), .ZN(n4713) );
  NAND2_X1 U5706 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n9346), .ZN(n4714) );
  AND2_X1 U5707 ( .A1(n5117), .A2(n5119), .ZN(n4992) );
  INV_X1 U5708 ( .A(n5179), .ZN(n4987) );
  AND3_X1 U5709 ( .A1(n5459), .A2(n5458), .A3(n5457), .ZN(n8815) );
  NAND2_X1 U5710 ( .A1(n5636), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4655) );
  OR2_X1 U5711 ( .A1(n6858), .A2(n5131), .ZN(n6895) );
  NAND2_X1 U5712 ( .A1(n4700), .A2(n4699), .ZN(n10264) );
  OR2_X1 U5713 ( .A1(n6903), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4700) );
  NAND2_X1 U5714 ( .A1(n6903), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U5715 ( .A1(n4701), .A2(n6862), .ZN(n10263) );
  NAND2_X1 U5716 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  NAND2_X1 U5717 ( .A1(n4926), .A2(n6900), .ZN(n4925) );
  AND2_X1 U5718 ( .A1(n4719), .A2(n4718), .ZN(n7007) );
  NOR2_X1 U5719 ( .A1(n6890), .A2(n6891), .ZN(n4718) );
  NAND2_X1 U5720 ( .A1(n4918), .A2(n10296), .ZN(n4919) );
  XNOR2_X1 U5721 ( .A(n7196), .B(n4706), .ZN(n7198) );
  OAI21_X1 U5722 ( .B1(n7198), .B2(n7406), .A(n4705), .ZN(n7200) );
  NAND2_X1 U5723 ( .A1(n7196), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U5724 ( .A1(n7200), .A2(n7199), .ZN(n7465) );
  OR2_X1 U5725 ( .A1(n7473), .A2(n7474), .ZN(n7520) );
  NAND2_X1 U5726 ( .A1(n7520), .A2(n7521), .ZN(n7519) );
  NAND2_X1 U5727 ( .A1(n7470), .A2(n7471), .ZN(n8043) );
  NOR2_X1 U5728 ( .A1(n8048), .A2(n8047), .ZN(n8051) );
  AOI21_X1 U5729 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8197), .A(n8194), .ZN(
        n8363) );
  NAND2_X1 U5730 ( .A1(n8370), .A2(n8371), .ZN(n8983) );
  XNOR2_X1 U5731 ( .A(n4704), .B(n9002), .ZN(n8987) );
  INV_X1 U5732 ( .A(n9012), .ZN(n4704) );
  OAI21_X1 U5733 ( .B1(n8987), .B2(n4703), .A(n4702), .ZN(n9035) );
  NAND2_X1 U5734 ( .A1(n9016), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U5735 ( .A1(n9015), .A2(n9016), .ZN(n4702) );
  NOR2_X1 U5736 ( .A1(n8987), .A2(n8986), .ZN(n9014) );
  NOR2_X1 U5737 ( .A1(n9037), .A2(n9038), .ZN(n9068) );
  NAND2_X1 U5738 ( .A1(n9032), .A2(n9033), .ZN(n9054) );
  NAND2_X1 U5739 ( .A1(n4544), .A2(n4697), .ZN(n4696) );
  INV_X1 U5740 ( .A(n9094), .ZN(n4697) );
  INV_X1 U5741 ( .A(n4693), .ZN(n4691) );
  AOI21_X1 U5742 ( .B1(n9070), .B2(n4608), .A(n4694), .ZN(n4693) );
  NOR2_X1 U5743 ( .A1(n9087), .A2(n9080), .ZN(n4694) );
  INV_X1 U5744 ( .A(n9087), .ZN(n4695) );
  NAND2_X1 U5745 ( .A1(n4927), .A2(n4928), .ZN(n4930) );
  AOI21_X1 U5746 ( .B1(n8997), .B2(n4929), .A(n9024), .ZN(n4928) );
  NAND2_X1 U5747 ( .A1(n9085), .A2(n4913), .ZN(n4912) );
  NAND2_X1 U5748 ( .A1(n9052), .A2(n9076), .ZN(n4913) );
  NAND2_X1 U5749 ( .A1(n5658), .A2(n5657), .ZN(n8600) );
  NAND2_X1 U5750 ( .A1(n4807), .A2(n4564), .ZN(n5734) );
  OR2_X1 U5751 ( .A1(n5650), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U5752 ( .A1(n5633), .A2(n5632), .ZN(n5650) );
  INV_X1 U5753 ( .A(n5634), .ZN(n5633) );
  INV_X1 U5754 ( .A(n5577), .ZN(n5576) );
  NAND2_X1 U5755 ( .A1(n5524), .A2(n5523), .ZN(n5542) );
  INV_X1 U5756 ( .A(n9168), .ZN(n9188) );
  AOI21_X1 U5757 ( .B1(n4815), .B2(n4814), .A(n4597), .ZN(n4813) );
  INV_X1 U5758 ( .A(n4532), .ZN(n4814) );
  AND2_X1 U5759 ( .A1(n8714), .A2(n8710), .ZN(n9199) );
  NAND2_X1 U5760 ( .A1(n5492), .A2(n5491), .ZN(n5521) );
  NAND2_X1 U5761 ( .A1(n5454), .A2(n5453), .ZN(n5473) );
  INV_X1 U5762 ( .A(n5455), .ZN(n5454) );
  NAND2_X1 U5763 ( .A1(n5405), .A2(n5404), .ZN(n5430) );
  INV_X1 U5764 ( .A(n5406), .ZN(n5405) );
  OR2_X1 U5765 ( .A1(n5380), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U5766 ( .A1(n5363), .A2(n5362), .ZN(n5380) );
  INV_X1 U5767 ( .A(n5364), .ZN(n5363) );
  NAND2_X1 U5768 ( .A1(n5345), .A2(n8154), .ZN(n5364) );
  INV_X1 U5769 ( .A(n5346), .ZN(n5345) );
  NAND2_X1 U5770 ( .A1(n5290), .A2(n5289), .ZN(n5308) );
  INV_X1 U5771 ( .A(n5291), .ZN(n5290) );
  OR2_X1 U5772 ( .A1(n7393), .A2(n7341), .ZN(n7318) );
  NAND2_X1 U5773 ( .A1(n5234), .A2(n8652), .ZN(n7395) );
  NAND2_X1 U5774 ( .A1(n7395), .A2(n8653), .ZN(n7394) );
  NAND2_X1 U5775 ( .A1(n5246), .A2(n5245), .ZN(n5267) );
  INV_X1 U5776 ( .A(n5247), .ZN(n5246) );
  INV_X1 U5777 ( .A(n8967), .ZN(n7536) );
  OR2_X1 U5778 ( .A1(n5209), .A2(n7087), .ZN(n4786) );
  NAND2_X1 U5779 ( .A1(n5636), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4787) );
  CLKBUF_X1 U5780 ( .A(n6943), .Z(n5678) );
  INV_X1 U5781 ( .A(n8612), .ZN(n5150) );
  AND2_X1 U5782 ( .A1(n9097), .A2(n9096), .ZN(n9279) );
  NAND2_X1 U5783 ( .A1(n9107), .A2(n10328), .ZN(n9109) );
  NAND2_X1 U5784 ( .A1(n4811), .A2(n9143), .ZN(n4810) );
  NAND2_X1 U5785 ( .A1(n4818), .A2(n4531), .ZN(n9152) );
  OR2_X1 U5786 ( .A1(n8717), .A2(n4995), .ZN(n4994) );
  NAND2_X1 U5787 ( .A1(n5010), .A2(n5009), .ZN(n8469) );
  NOR2_X1 U5788 ( .A1(n5012), .A2(n8689), .ZN(n5009) );
  OR2_X1 U5789 ( .A1(n8229), .A2(n8685), .ZN(n8781) );
  INV_X1 U5790 ( .A(n5004), .ZN(n5003) );
  OAI21_X1 U5791 ( .B1(n5006), .B2(n5005), .A(n5370), .ZN(n5004) );
  INV_X1 U5792 ( .A(n8961), .ZN(n8512) );
  AND4_X1 U5793 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n8168)
         );
  AND2_X2 U5794 ( .A1(n4791), .A2(n4790), .ZN(n10375) );
  OR2_X1 U5795 ( .A1(n6750), .A2(n5205), .ZN(n4791) );
  AND2_X1 U5796 ( .A1(n5792), .A2(n5791), .ZN(n6958) );
  INV_X1 U5797 ( .A(n7157), .ZN(n10360) );
  NAND2_X1 U5798 ( .A1(n5745), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5799 ( .A1(n5036), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5676) );
  AND2_X1 U5800 ( .A1(n5358), .A2(n5357), .ZN(n5376) );
  XNOR2_X1 U5801 ( .A(n5231), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7036) );
  INV_X1 U5802 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U5803 ( .A1(n7502), .A2(n6540), .ZN(n6547) );
  NAND2_X1 U5804 ( .A1(n8421), .A2(n6600), .ZN(n6609) );
  AND2_X1 U5805 ( .A1(n6691), .A2(n6690), .ZN(n6713) );
  NOR2_X1 U5806 ( .A1(n5890), .A2(n9561), .ZN(n5921) );
  XNOR2_X1 U5807 ( .A(n6527), .B(n6702), .ZN(n6528) );
  OR2_X1 U5808 ( .A1(n6052), .A2(n6051), .ZN(n6075) );
  INV_X1 U5809 ( .A(n5981), .ZN(n8577) );
  AND2_X1 U5810 ( .A1(n6544), .A2(n6543), .ZN(n7502) );
  NOR2_X1 U5811 ( .A1(n4906), .A2(n4570), .ZN(n4904) );
  AND2_X1 U5812 ( .A1(n4905), .A2(n6678), .ZN(n9468) );
  NAND2_X1 U5813 ( .A1(n6327), .A2(n6375), .ZN(n4941) );
  INV_X1 U5814 ( .A(n4956), .ZN(n6464) );
  INV_X1 U5815 ( .A(n6372), .ZN(n6465) );
  AND4_X1 U5816 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n8428)
         );
  AND4_X1 U5817 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n9992)
         );
  NOR2_X1 U5818 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  NOR2_X1 U5819 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5954) );
  NAND2_X1 U5820 ( .A1(n4653), .A2(n4652), .ZN(n10044) );
  NAND2_X1 U5821 ( .A1(n6801), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U5822 ( .A1(n10044), .A2(n10045), .ZN(n10042) );
  AND2_X1 U5823 ( .A1(n9528), .A2(n6795), .ZN(n6798) );
  AOI21_X1 U5824 ( .B1(n6822), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6821), .ZN(
        n6824) );
  NOR2_X1 U5825 ( .A1(n7042), .A2(n4646), .ZN(n9542) );
  AND2_X1 U5826 ( .A1(n7043), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4646) );
  NOR2_X1 U5827 ( .A1(n9542), .A2(n9541), .ZN(n9540) );
  NOR2_X1 U5828 ( .A1(n9540), .A2(n4643), .ZN(n7045) );
  NOR2_X1 U5829 ( .A1(n4645), .A2(n4644), .ZN(n4643) );
  INV_X1 U5830 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U5831 ( .A1(n7045), .A2(n7046), .ZN(n7289) );
  NOR2_X1 U5832 ( .A1(n7358), .A2(n4648), .ZN(n7362) );
  AND2_X1 U5833 ( .A1(n7359), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4648) );
  NOR2_X1 U5834 ( .A1(n7362), .A2(n7361), .ZN(n7442) );
  NOR2_X1 U5835 ( .A1(n7442), .A2(n4647), .ZN(n7447) );
  AND2_X1 U5836 ( .A1(n7443), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U5837 ( .A1(n7447), .A2(n7446), .ZN(n8103) );
  NOR2_X1 U5838 ( .A1(n8257), .A2(n4650), .ZN(n8261) );
  AND2_X1 U5839 ( .A1(n8258), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5840 ( .A1(n9577), .A2(n9576), .ZN(n9580) );
  NAND2_X1 U5841 ( .A1(n9590), .A2(n4611), .ZN(n9612) );
  AND2_X1 U5842 ( .A1(n9612), .A2(n9611), .ZN(n9616) );
  NAND2_X1 U5843 ( .A1(n9616), .A2(n9615), .ZN(n9624) );
  AND2_X1 U5844 ( .A1(n9749), .A2(n4861), .ZN(n9691) );
  NOR2_X1 U5845 ( .A1(n9861), .A2(n4862), .ZN(n4861) );
  INV_X1 U5846 ( .A(n4864), .ZN(n4862) );
  NAND2_X1 U5847 ( .A1(n4619), .A2(n5826), .ZN(n9861) );
  AND4_X1 U5848 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n9732)
         );
  AND4_X1 U5849 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n9748)
         );
  NOR2_X1 U5850 ( .A1(n9744), .A2(n9745), .ZN(n9743) );
  AND2_X1 U5851 ( .A1(n9677), .A2(n6357), .ZN(n9760) );
  AND2_X1 U5852 ( .A1(n6300), .A2(n9758), .ZN(n9775) );
  NOR2_X1 U5853 ( .A1(n9809), .A2(n9900), .ZN(n9787) );
  NAND2_X1 U5854 ( .A1(n4779), .A2(n4778), .ZN(n9786) );
  AOI21_X1 U5855 ( .B1(n4780), .B2(n4592), .A(n4534), .ZN(n4778) );
  AND4_X1 U5856 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(n9808)
         );
  NOR2_X1 U5857 ( .A1(n8552), .A2(n4858), .ZN(n9844) );
  INV_X1 U5858 ( .A(n4860), .ZN(n4858) );
  NAND2_X1 U5859 ( .A1(n4851), .A2(n6423), .ZN(n8561) );
  OR2_X1 U5860 ( .A1(n4854), .A2(n4551), .ZN(n4851) );
  INV_X1 U5861 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U5862 ( .B1(n4756), .B2(n4549), .A(n4535), .ZN(n4753) );
  AND2_X1 U5863 ( .A1(n9831), .A2(n6303), .ZN(n8559) );
  INV_X1 U5864 ( .A(n4854), .ZN(n8490) );
  AND2_X1 U5865 ( .A1(n8127), .A2(n4855), .ZN(n8494) );
  AND2_X1 U5866 ( .A1(n4537), .A2(n8487), .ZN(n4855) );
  NAND2_X1 U5867 ( .A1(n8127), .A2(n4856), .ZN(n8315) );
  AND4_X1 U5868 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n9504)
         );
  NAND2_X1 U5869 ( .A1(n8117), .A2(n6347), .ZN(n8306) );
  OR2_X1 U5870 ( .A1(n8431), .A2(n9505), .ZN(n8124) );
  OR2_X1 U5871 ( .A1(n6102), .A2(n8426), .ZN(n6114) );
  AND2_X1 U5872 ( .A1(n8029), .A2(n10199), .ZN(n8082) );
  AND2_X1 U5873 ( .A1(n8082), .A2(n10204), .ZN(n8127) );
  NAND2_X1 U5874 ( .A1(n8073), .A2(n6346), .ZN(n8117) );
  NAND2_X1 U5875 ( .A1(n8007), .A2(n8006), .ZN(n10071) );
  INV_X1 U5876 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6040) );
  NOR2_X1 U5877 ( .A1(n4868), .A2(n7499), .ZN(n4867) );
  INV_X1 U5878 ( .A(n4870), .ZN(n4868) );
  AND4_X1 U5879 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n6066)
         );
  NAND2_X1 U5880 ( .A1(n6342), .A2(n6398), .ZN(n10079) );
  NAND2_X1 U5881 ( .A1(n4869), .A2(n4870), .ZN(n10085) );
  INV_X1 U5882 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6006) );
  NOR2_X1 U5883 ( .A1(n7332), .A2(n4871), .ZN(n10086) );
  NOR2_X1 U5884 ( .A1(n7332), .A2(n10157), .ZN(n7331) );
  OR2_X1 U5885 ( .A1(n10100), .A2(n7219), .ZN(n7332) );
  NOR2_X1 U5886 ( .A1(n5982), .A2(n6976), .ZN(n10101) );
  INV_X1 U5887 ( .A(n6976), .ZN(n10111) );
  INV_X1 U5888 ( .A(n6991), .ZN(n4829) );
  AND2_X1 U5889 ( .A1(n9861), .A2(n10158), .ZN(n9862) );
  AND2_X1 U5890 ( .A1(n9870), .A2(n10158), .ZN(n4846) );
  INV_X1 U5891 ( .A(n9398), .ZN(n9972) );
  INV_X1 U5892 ( .A(n4783), .ZN(n4782) );
  NAND2_X1 U5893 ( .A1(n6767), .A2(n6191), .ZN(n4784) );
  OAI21_X1 U5894 ( .B1(n6050), .B2(n6768), .A(n6049), .ZN(n4783) );
  XNOR2_X1 U5895 ( .A(n6272), .B(SI_29_), .ZN(n5825) );
  NOR2_X1 U5896 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n5814), .ZN(n4873) );
  XNOR2_X1 U5897 ( .A(n5644), .B(n5645), .ZN(n8321) );
  INV_X1 U5898 ( .A(n5533), .ZN(n4958) );
  INV_X1 U5899 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U5900 ( .A1(n5516), .A2(n5515), .ZN(n5534) );
  NAND2_X1 U5901 ( .A1(n5871), .A2(n5102), .ZN(n6150) );
  INV_X1 U5902 ( .A(n6138), .ZN(n5871) );
  XNOR2_X1 U5903 ( .A(n5420), .B(n5419), .ZN(n6972) );
  INV_X1 U5904 ( .A(n5225), .ZN(n4955) );
  INV_X1 U5905 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U5906 ( .A1(n5057), .A2(n5058), .ZN(n8927) );
  NAND2_X1 U5907 ( .A1(n8537), .A2(n4542), .ZN(n5057) );
  NAND2_X1 U5908 ( .A1(n5043), .A2(n5044), .ZN(n5051) );
  AOI22_X1 U5909 ( .A1(n8875), .A2(n8876), .B1(n8825), .B2(n8824), .ZN(n8917)
         );
  OAI21_X1 U5910 ( .B1(n5069), .B2(n5070), .A(n5065), .ZN(n5064) );
  AOI21_X1 U5911 ( .B1(n5071), .B2(n5070), .A(n5069), .ZN(n8224) );
  AND4_X1 U5912 ( .A1(n5172), .A2(n5171), .A3(n5170), .A4(n5169), .ZN(n10347)
         );
  OR2_X1 U5913 ( .A1(n8537), .A2(n4528), .ZN(n5052) );
  INV_X1 U5914 ( .A(n8968), .ZN(n7341) );
  OR2_X1 U5915 ( .A1(n6931), .A2(n6930), .ZN(n8945) );
  NAND2_X1 U5916 ( .A1(n5603), .A2(n5602), .ZN(n9153) );
  NAND4_X1 U5917 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n8970)
         );
  INV_X1 U5918 ( .A(n10347), .ZN(n8971) );
  NAND4_X1 U5919 ( .A1(n5156), .A2(n5155), .A3(n5154), .A4(n5153), .ZN(n10327)
         );
  OAI21_X1 U5920 ( .B1(n10270), .B2(n10271), .A(n4720), .ZN(n10289) );
  OR2_X1 U5921 ( .A1(n6888), .A2(n6903), .ZN(n4720) );
  INV_X1 U5922 ( .A(n4719), .ZN(n10288) );
  NOR2_X1 U5923 ( .A1(n7007), .A2(n4716), .ZN(n7111) );
  NOR2_X1 U5924 ( .A1(n4717), .A2(n7029), .ZN(n4716) );
  INV_X1 U5925 ( .A(n7009), .ZN(n4717) );
  NOR2_X1 U5926 ( .A1(n10316), .A2(n10315), .ZN(n10314) );
  INV_X1 U5927 ( .A(n4710), .ZN(n7182) );
  NAND2_X1 U5928 ( .A1(n7183), .A2(n7197), .ZN(n4709) );
  NOR2_X1 U5929 ( .A1(n7516), .A2(n10434), .ZN(n7515) );
  NAND2_X1 U5930 ( .A1(n4933), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U5931 ( .A1(n7463), .A2(n4933), .ZN(n4931) );
  INV_X1 U5932 ( .A(n7464), .ZN(n4933) );
  INV_X1 U5933 ( .A(n8135), .ZN(n4922) );
  OAI21_X1 U5934 ( .B1(n8042), .B2(n4921), .A(n4920), .ZN(n8194) );
  NAND2_X1 U5935 ( .A1(n4924), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U5936 ( .A1(n8135), .A2(n4924), .ZN(n4920) );
  INV_X1 U5937 ( .A(n8137), .ZN(n4924) );
  XNOR2_X1 U5938 ( .A(n8369), .B(n8364), .ZN(n8200) );
  NAND2_X1 U5939 ( .A1(n8200), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8370) );
  XNOR2_X1 U5940 ( .A(n8363), .B(n8364), .ZN(n8195) );
  NOR2_X1 U5941 ( .A1(n8195), .A2(n8196), .ZN(n8365) );
  OAI21_X1 U5942 ( .B1(n8195), .B2(n4935), .A(n4934), .ZN(n8974) );
  NAND2_X1 U5943 ( .A1(n4936), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U5944 ( .A1(n8366), .A2(n4936), .ZN(n4934) );
  INV_X1 U5945 ( .A(n8368), .ZN(n4936) );
  NOR2_X1 U5946 ( .A1(n8998), .A2(n8997), .ZN(n9001) );
  NOR2_X1 U5947 ( .A1(n9001), .A2(n9000), .ZN(n9025) );
  XNOR2_X1 U5948 ( .A(n4930), .B(n9028), .ZN(n9026) );
  NAND2_X1 U5949 ( .A1(n9086), .A2(n4916), .ZN(n4915) );
  INV_X1 U5950 ( .A(n9052), .ZN(n4916) );
  XNOR2_X1 U5951 ( .A(n8600), .B(n5733), .ZN(n8813) );
  OAI21_X1 U5952 ( .B1(n9197), .B2(n4997), .A(n8710), .ZN(n9190) );
  OR2_X1 U5953 ( .A1(n8230), .A2(n8685), .ZN(n5015) );
  NAND2_X1 U5954 ( .A1(n8089), .A2(n8671), .ZN(n8187) );
  NAND2_X1 U5955 ( .A1(n5326), .A2(n5325), .ZN(n10417) );
  NAND2_X1 U5956 ( .A1(n7433), .A2(n8639), .ZN(n7555) );
  NAND2_X1 U5957 ( .A1(n6069), .A2(n5421), .ZN(n5286) );
  NAND2_X1 U5958 ( .A1(n5265), .A2(n5264), .ZN(n10400) );
  OR2_X1 U5959 ( .A1(n6933), .A2(n6932), .ZN(n10343) );
  INV_X1 U5960 ( .A(n10334), .ZN(n9226) );
  NAND2_X1 U5961 ( .A1(n8596), .A2(n8595), .ZN(n9231) );
  NAND2_X1 U5962 ( .A1(n8598), .A2(n8597), .ZN(n9278) );
  NAND2_X1 U5963 ( .A1(n5026), .A2(n5024), .ZN(n9119) );
  NAND2_X1 U5964 ( .A1(n5026), .A2(n8731), .ZN(n9131) );
  NAND2_X1 U5965 ( .A1(n5594), .A2(n5593), .ZN(n9305) );
  NAND2_X1 U5966 ( .A1(n4819), .A2(n4822), .ZN(n9166) );
  NAND2_X1 U5967 ( .A1(n9185), .A2(n4821), .ZN(n4819) );
  NAND2_X1 U5968 ( .A1(n5541), .A2(n5540), .ZN(n9324) );
  NAND2_X1 U5969 ( .A1(n4823), .A2(n4827), .ZN(n9178) );
  OR2_X1 U5970 ( .A1(n9185), .A2(n9189), .ZN(n4823) );
  OR2_X1 U5971 ( .A1(n9266), .A2(n9265), .ZN(n9332) );
  NAND2_X1 U5972 ( .A1(n5506), .A2(n5505), .ZN(n9334) );
  NAND2_X1 U5973 ( .A1(n5490), .A2(n5489), .ZN(n9339) );
  AND2_X1 U5974 ( .A1(n9222), .A2(n9221), .ZN(n9337) );
  NAND2_X1 U5975 ( .A1(n5472), .A2(n5471), .ZN(n8924) );
  NAND2_X1 U5976 ( .A1(n5452), .A2(n5451), .ZN(n8889) );
  NAND2_X1 U5977 ( .A1(n4800), .A2(n5722), .ZN(n8446) );
  NAND2_X1 U5978 ( .A1(n8337), .A2(n8336), .ZN(n4800) );
  AND2_X1 U5979 ( .A1(n5010), .A2(n5011), .ZN(n8445) );
  NAND2_X1 U5980 ( .A1(n5403), .A2(n5402), .ZN(n8508) );
  NAND2_X1 U5981 ( .A1(n5378), .A2(n5377), .ZN(n8402) );
  NAND2_X1 U5982 ( .A1(n8182), .A2(n8677), .ZN(n8267) );
  NAND2_X1 U5983 ( .A1(n5344), .A2(n5343), .ZN(n8669) );
  AND2_X1 U5984 ( .A1(n5125), .A2(n5136), .ZN(n5126) );
  INV_X1 U5985 ( .A(n5132), .ZN(n9353) );
  NAND2_X1 U5986 ( .A1(n5122), .A2(n5032), .ZN(n5751) );
  INV_X1 U5987 ( .A(n6903), .ZN(n10256) );
  NAND2_X1 U5988 ( .A1(n6906), .A2(n5141), .ZN(n6884) );
  MUX2_X1 U5989 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5140), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5141) );
  NOR2_X1 U5990 ( .A1(n7492), .A2(n7491), .ZN(n7490) );
  AND2_X1 U5991 ( .A1(n4903), .A2(n4553), .ZN(n7492) );
  NAND2_X1 U5992 ( .A1(n6548), .A2(n6547), .ZN(n4903) );
  NAND2_X1 U5993 ( .A1(n4886), .A2(n9456), .ZN(n9365) );
  INV_X1 U5994 ( .A(n6560), .ZN(n6558) );
  AND2_X1 U5995 ( .A1(n4881), .A2(n9458), .ZN(n4878) );
  NAND2_X1 U5996 ( .A1(n9403), .A2(n9405), .ZN(n9402) );
  INV_X1 U5997 ( .A(n4883), .ZN(n4882) );
  INV_X1 U5998 ( .A(n6522), .ZN(n4874) );
  AND2_X1 U5999 ( .A1(n6721), .A2(n6709), .ZN(n10000) );
  NAND2_X1 U6000 ( .A1(n6157), .A2(n6156), .ZN(n9645) );
  INV_X1 U6001 ( .A(n10000), .ZN(n9494) );
  NAND4_X1 U6002 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n9648)
         );
  AND4_X1 U6003 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n9990)
         );
  NAND2_X1 U6004 ( .A1(n6227), .A2(n10082), .ZN(n6023) );
  INV_X1 U6005 ( .A(n4653), .ZN(n9518) );
  XNOR2_X1 U6006 ( .A(n9575), .B(n9574), .ZN(n9554) );
  AND2_X1 U6007 ( .A1(n6778), .A2(n6788), .ZN(n10049) );
  NAND2_X1 U6008 ( .A1(n6290), .A2(n5980), .ZN(n9636) );
  NAND2_X1 U6009 ( .A1(n4962), .A2(n4961), .ZN(n6290) );
  NAND2_X1 U6010 ( .A1(n6743), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U6011 ( .A1(n9345), .A2(n6744), .ZN(n4962) );
  OAI21_X1 U6012 ( .B1(n9705), .B2(n10129), .A(n9704), .ZN(n9868) );
  AND2_X1 U6013 ( .A1(n5852), .A2(n5851), .ZN(n9723) );
  NAND2_X1 U6014 ( .A1(n4762), .A2(n4766), .ZN(n9716) );
  NAND2_X1 U6015 ( .A1(n9742), .A2(n4770), .ZN(n4762) );
  AOI21_X1 U6016 ( .B1(n9742), .B2(n9663), .A(n9662), .ZN(n9728) );
  AND2_X1 U6017 ( .A1(n6237), .A2(n6236), .ZN(n9770) );
  NAND2_X1 U6018 ( .A1(n6223), .A2(n6222), .ZN(n9774) );
  NAND2_X1 U6019 ( .A1(n9802), .A2(n9675), .ZN(n9793) );
  AND2_X1 U6020 ( .A1(n6214), .A2(n6213), .ZN(n9790) );
  AND2_X1 U6021 ( .A1(n4781), .A2(n4546), .ZN(n9801) );
  OR2_X1 U6022 ( .A1(n9818), .A2(n4592), .ZN(n4781) );
  OR2_X1 U6023 ( .A1(n4854), .A2(n4853), .ZN(n8550) );
  NAND2_X1 U6024 ( .A1(n4751), .A2(n4756), .ZN(n8558) );
  OR2_X1 U6025 ( .A1(n8486), .A2(n4757), .ZN(n4751) );
  NAND2_X1 U6026 ( .A1(n4758), .A2(n5098), .ZN(n8548) );
  NAND2_X1 U6027 ( .A1(n4774), .A2(n4773), .ZN(n8126) );
  AND2_X1 U6028 ( .A1(n4777), .A2(n4550), .ZN(n8071) );
  NAND2_X1 U6029 ( .A1(n8035), .A2(n8018), .ZN(n4777) );
  OAI211_X1 U6030 ( .C1(n5961), .C2(n6748), .A(n5960), .B(n5959), .ZN(n10095)
         );
  INV_X1 U6031 ( .A(n9815), .ZN(n10094) );
  NAND2_X1 U6032 ( .A1(n7002), .A2(n10108), .ZN(n10118) );
  NAND2_X1 U6033 ( .A1(n5816), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5817) );
  XNOR2_X1 U6034 ( .A(n5567), .B(n5566), .ZN(n8065) );
  OAI211_X1 U6035 ( .C1(n4960), .C2(n4539), .A(n5552), .B(n4631), .ZN(n5567)
         );
  OR2_X1 U6036 ( .A1(n5516), .A2(n4539), .ZN(n4631) );
  NAND2_X1 U6037 ( .A1(n5867), .A2(n5811), .ZN(n6378) );
  INV_X1 U6038 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7772) );
  XNOR2_X1 U6039 ( .A(n5201), .B(n5200), .ZN(n6750) );
  XNOR2_X1 U6040 ( .A(n5966), .B(n4651), .ZN(n6804) );
  INV_X1 U6041 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4651) );
  XNOR2_X1 U6042 ( .A(n4681), .B(n9093), .ZN(n8805) );
  INV_X1 U6043 ( .A(n4923), .ZN(n8134) );
  AOI21_X1 U6044 ( .B1(n9064), .B2(n9063), .A(n4727), .ZN(n9074) );
  NAND2_X1 U6045 ( .A1(n4909), .A2(n4915), .ZN(n4908) );
  NAND2_X1 U6046 ( .A1(n9236), .A2(n9235), .ZN(n9238) );
  INV_X1 U6047 ( .A(n5800), .ZN(n5801) );
  OAI22_X1 U6048 ( .A1(n8808), .A2(n9331), .B1(n10421), .B2(n5799), .ZN(n5800)
         );
  NAND2_X1 U6049 ( .A1(n4639), .A2(n4635), .ZN(n9633) );
  OAI21_X1 U6050 ( .B1(n4642), .B2(n10022), .A(n4640), .ZN(n4639) );
  NAND2_X1 U6051 ( .A1(n4843), .A2(n4607), .ZN(P1_U3550) );
  NAND2_X1 U6052 ( .A1(n9926), .A2(n10247), .ZN(n4843) );
  INV_X1 U6053 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U6054 ( .A1(n9854), .A2(n10226), .ZN(n6498) );
  NAND2_X1 U6055 ( .A1(n4667), .A2(n10255), .ZN(n6906) );
  AND2_X1 U6056 ( .A1(n5980), .A2(n6744), .ZN(n6097) );
  NAND2_X1 U6057 ( .A1(n5058), .A2(n8819), .ZN(n4528) );
  OAI21_X1 U6058 ( .B1(n8336), .B2(n5013), .A(n8695), .ZN(n5012) );
  AOI21_X1 U6059 ( .B1(n8901), .B2(n8902), .A(n8831), .ZN(n8882) );
  NAND2_X1 U6060 ( .A1(n6282), .A2(n6281), .ZN(n6471) );
  INV_X1 U6061 ( .A(n6471), .ZN(n4743) );
  NAND2_X1 U6062 ( .A1(n5641), .A2(n5640), .ZN(n9134) );
  INV_X1 U6063 ( .A(n9134), .ZN(n8843) );
  NAND2_X1 U6064 ( .A1(n5620), .A2(n5619), .ZN(n9124) );
  INV_X1 U6065 ( .A(n9124), .ZN(n9143) );
  AND2_X1 U6066 ( .A1(n9670), .A2(n4743), .ZN(n4530) );
  NOR2_X1 U6067 ( .A1(n4820), .A2(n4590), .ZN(n4531) );
  NAND2_X1 U6068 ( .A1(n8924), .A2(n8957), .ZN(n4532) );
  NOR2_X1 U6069 ( .A1(n8715), .A2(n4670), .ZN(n4533) );
  NOR2_X1 U6070 ( .A1(n9651), .A2(n9653), .ZN(n4534) );
  OR2_X1 U6071 ( .A1(n9911), .A2(n9499), .ZN(n4535) );
  AND4_X1 U6072 ( .A1(n5941), .A2(n5940), .A3(n6417), .A4(n5939), .ZN(n4536)
         );
  AND2_X1 U6073 ( .A1(n4856), .A2(n8324), .ZN(n4537) );
  NAND2_X1 U6074 ( .A1(n10304), .A2(n4707), .ZN(n7196) );
  AND2_X1 U6075 ( .A1(n4805), .A2(n4808), .ZN(n4538) );
  OR2_X1 U6076 ( .A1(n5551), .A2(n4958), .ZN(n4539) );
  OR2_X1 U6077 ( .A1(n8552), .A2(n4859), .ZN(n4540) );
  AND2_X1 U6078 ( .A1(n5015), .A2(n8691), .ZN(n4541) );
  INV_X1 U6079 ( .A(n5982), .ZN(n10137) );
  NAND3_X1 U6080 ( .A1(n5971), .A2(n5970), .A3(n5969), .ZN(n5982) );
  INV_X1 U6081 ( .A(n6144), .ZN(n6196) );
  INV_X2 U6082 ( .A(n6196), .ZN(n6227) );
  INV_X1 U6083 ( .A(n4785), .ZN(n8767) );
  OAI21_X1 U6084 ( .B1(n10375), .B2(n8647), .A(n7237), .ZN(n4785) );
  INV_X1 U6085 ( .A(n9824), .ZN(n9955) );
  NAND2_X1 U6086 ( .A1(n6178), .A2(n6177), .ZN(n9824) );
  AND2_X1 U6087 ( .A1(n8534), .A2(n5059), .ZN(n4542) );
  OR4_X1 U6088 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6994), .ZN(n4543) );
  OR2_X1 U6089 ( .A1(n9090), .A2(n10317), .ZN(n4544) );
  OR2_X1 U6090 ( .A1(n8883), .A2(n5049), .ZN(n4545) );
  INV_X1 U6091 ( .A(n8784), .ZN(n5002) );
  OAI21_X1 U6092 ( .B1(n8859), .B2(n9179), .A(n5051), .ZN(n8901) );
  OR2_X1 U6093 ( .A1(n9824), .A2(n9835), .ZN(n4546) );
  NAND2_X2 U6094 ( .A1(n5132), .A2(n8501), .ZN(n5188) );
  OR2_X1 U6095 ( .A1(n8069), .A2(n9506), .ZN(n4547) );
  INV_X1 U6096 ( .A(n6420), .ZN(n4853) );
  AND2_X1 U6097 ( .A1(n10053), .A2(n9630), .ZN(n4548) );
  AND2_X1 U6098 ( .A1(n9911), .A2(n9499), .ZN(n4549) );
  INV_X1 U6099 ( .A(n8304), .ZN(n4830) );
  XNOR2_X1 U6100 ( .A(n5158), .B(n5160), .ZN(n5157) );
  INV_X1 U6101 ( .A(n8547), .ZN(n4850) );
  OR2_X1 U6102 ( .A1(n8017), .A2(n8036), .ZN(n4550) );
  OR2_X1 U6103 ( .A1(n8549), .A2(n4853), .ZN(n4551) );
  NAND3_X1 U6104 ( .A1(n10255), .A2(n4667), .A3(n5115), .ZN(n5179) );
  INV_X1 U6105 ( .A(n8549), .ZN(n5083) );
  NAND2_X1 U6106 ( .A1(n5919), .A2(n5918), .ZN(n9920) );
  OR2_X1 U6107 ( .A1(n9863), .A2(n9862), .ZN(n4552) );
  XNOR2_X1 U6108 ( .A(n5299), .B(n5100), .ZN(n6069) );
  NOR2_X1 U6109 ( .A1(n4836), .A2(n4839), .ZN(n5819) );
  INV_X1 U6110 ( .A(n10083), .ZN(n10174) );
  OAI211_X1 U6111 ( .C1(n5961), .C2(n6755), .A(n6031), .B(n6030), .ZN(n10083)
         );
  NOR2_X1 U6112 ( .A1(n4841), .A2(n4838), .ZN(n6454) );
  AND2_X1 U6113 ( .A1(n6546), .A2(n6545), .ZN(n4553) );
  NAND2_X1 U6114 ( .A1(n6167), .A2(n6166), .ZN(n9850) );
  NAND4_X1 U6115 ( .A1(n4988), .A2(n4990), .A3(n4987), .A4(n4992), .ZN(n4554)
         );
  OR2_X1 U6116 ( .A1(n8924), .A2(n8957), .ZN(n4555) );
  AND2_X2 U6117 ( .A1(n5980), .A2(n6743), .ZN(n5967) );
  AND2_X1 U6118 ( .A1(n4710), .A2(n4709), .ZN(n4556) );
  OR2_X1 U6119 ( .A1(n9114), .A2(n9123), .ZN(n4557) );
  NAND2_X1 U6120 ( .A1(n4893), .A2(n9390), .ZN(n9403) );
  AND2_X1 U6121 ( .A1(n8776), .A2(n8641), .ZN(n4558) );
  AND2_X1 U6122 ( .A1(n9398), .A2(n9500), .ZN(n4559) );
  OR2_X1 U6123 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n9346), .ZN(n4560) );
  OR2_X1 U6124 ( .A1(n8508), .A2(n8541), .ZN(n8691) );
  OR2_X1 U6125 ( .A1(n5714), .A2(n8962), .ZN(n8677) );
  INV_X1 U6126 ( .A(n8677), .ZN(n5029) );
  OR2_X1 U6127 ( .A1(n5994), .A2(n4740), .ZN(n6026) );
  OR2_X1 U6128 ( .A1(n4841), .A2(n4839), .ZN(n4561) );
  NOR2_X1 U6129 ( .A1(n9014), .A2(n9015), .ZN(n4562) );
  AND2_X1 U6130 ( .A1(n5228), .A2(n5203), .ZN(n4563) );
  OR2_X1 U6131 ( .A1(n9290), .A2(n8746), .ZN(n4564) );
  AND2_X1 U6132 ( .A1(n8692), .A2(n8748), .ZN(n4565) );
  NOR2_X1 U6133 ( .A1(n9730), .A2(n9729), .ZN(n4566) );
  NOR2_X1 U6134 ( .A1(n9664), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U6135 ( .A1(n8677), .A2(n8674), .ZN(n8777) );
  AND2_X1 U6136 ( .A1(n8644), .A2(n8667), .ZN(n4567) );
  NAND2_X1 U6137 ( .A1(n5843), .A2(n5842), .ZN(n9870) );
  OR2_X1 U6138 ( .A1(n6906), .A2(n7105), .ZN(n6862) );
  OR2_X1 U6139 ( .A1(n5468), .A2(n5467), .ZN(n4568) );
  NAND2_X1 U6140 ( .A1(n5439), .A2(n5438), .ZN(n4569) );
  OR2_X1 U6141 ( .A1(n6553), .A2(n6552), .ZN(n6556) );
  INV_X1 U6142 ( .A(n5726), .ZN(n4825) );
  NOR2_X1 U6143 ( .A1(n9317), .A2(n9179), .ZN(n5726) );
  NAND2_X1 U6144 ( .A1(n5849), .A2(n5848), .ZN(n9874) );
  INV_X1 U6145 ( .A(n9874), .ZN(n4866) );
  NAND2_X1 U6146 ( .A1(n9470), .A2(n9467), .ZN(n4570) );
  NAND3_X1 U6147 ( .A1(n5074), .A2(n5895), .A3(n5811), .ZN(n4571) );
  INV_X1 U6148 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4746) );
  AND2_X1 U6149 ( .A1(n4866), .A2(n9732), .ZN(n4572) );
  AND2_X1 U6150 ( .A1(n4852), .A2(n8559), .ZN(n4573) );
  NAND2_X1 U6151 ( .A1(n5558), .A2(n5557), .ZN(n9317) );
  OR3_X1 U6152 ( .A1(n4749), .A2(n6124), .A3(n6123), .ZN(n4574) );
  OR2_X1 U6153 ( .A1(n8165), .A2(n8965), .ZN(n5070) );
  AND2_X1 U6154 ( .A1(n6366), .A2(n6330), .ZN(n9670) );
  NAND2_X1 U6155 ( .A1(n5984), .A2(n7370), .ZN(n4575) );
  NAND2_X1 U6156 ( .A1(n4824), .A2(n9177), .ZN(n4576) );
  INV_X1 U6157 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U6158 ( .A1(n4884), .A2(n4882), .ZN(n9435) );
  AND2_X1 U6159 ( .A1(n6547), .A2(n4901), .ZN(n4577) );
  AND2_X1 U6160 ( .A1(n9718), .A2(n4770), .ZN(n4578) );
  INV_X1 U6161 ( .A(n9675), .ZN(n4834) );
  NOR2_X1 U6162 ( .A1(n9380), .A2(n6677), .ZN(n4579) );
  AND2_X1 U6163 ( .A1(n5032), .A2(n5126), .ZN(n4580) );
  AND2_X1 U6164 ( .A1(n5032), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4581) );
  AND2_X1 U6165 ( .A1(n10255), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4582) );
  AND2_X1 U6166 ( .A1(n8116), .A2(n6311), .ZN(n8125) );
  NAND2_X1 U6167 ( .A1(n5396), .A2(n5395), .ZN(n4583) );
  AND2_X1 U6168 ( .A1(n5105), .A2(n5078), .ZN(n4584) );
  INV_X1 U6169 ( .A(n5732), .ZN(n4809) );
  NOR2_X1 U6170 ( .A1(n5731), .A2(n8843), .ZN(n5732) );
  AND2_X1 U6171 ( .A1(n5642), .A2(n5021), .ZN(n4585) );
  AND2_X1 U6172 ( .A1(n4994), .A2(n8716), .ZN(n4586) );
  AND2_X1 U6173 ( .A1(n4825), .A2(n4821), .ZN(n4587) );
  INV_X1 U6174 ( .A(n9916), .ZN(n8487) );
  AND2_X1 U6175 ( .A1(n4538), .A2(n4557), .ZN(n4588) );
  AND2_X1 U6176 ( .A1(n6608), .A2(n4897), .ZN(n4589) );
  AND2_X1 U6177 ( .A1(n9317), .A2(n9179), .ZN(n4590) );
  AND2_X1 U6178 ( .A1(n4902), .A2(n6556), .ZN(n4591) );
  AND2_X1 U6179 ( .A1(n9216), .A2(n4555), .ZN(n4815) );
  INV_X1 U6180 ( .A(n6678), .ZN(n4906) );
  OR2_X1 U6181 ( .A1(n6677), .A2(n9381), .ZN(n6678) );
  INV_X1 U6182 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5303) );
  INV_X1 U6183 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5675) );
  AND2_X1 U6184 ( .A1(n9824), .A2(n9835), .ZN(n4592) );
  INV_X1 U6185 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n4668) );
  AND2_X1 U6186 ( .A1(n7318), .A2(n8656), .ZN(n8653) );
  INV_X1 U6187 ( .A(n8653), .ZN(n4984) );
  AND2_X1 U6188 ( .A1(n5262), .A2(n5242), .ZN(n7197) );
  INV_X1 U6189 ( .A(n7197), .ZN(n4706) );
  INV_X1 U6190 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5040) );
  NOR3_X1 U6191 ( .A1(n8552), .A2(n9906), .A3(n4859), .ZN(n4857) );
  INV_X1 U6192 ( .A(n9366), .ZN(n4885) );
  NAND2_X1 U6193 ( .A1(n5358), .A2(n5062), .ZN(n5464) );
  NOR2_X1 U6194 ( .A1(n8365), .A2(n8366), .ZN(n4593) );
  NAND2_X1 U6195 ( .A1(n5613), .A2(n5612), .ZN(n9299) );
  AND2_X1 U6196 ( .A1(n5052), .A2(n5055), .ZN(n4594) );
  AND2_X1 U6197 ( .A1(n4923), .A2(n4922), .ZN(n4595) );
  NAND2_X1 U6198 ( .A1(n5015), .A2(n5014), .ZN(n4596) );
  AND2_X1 U6199 ( .A1(n9339), .A2(n9203), .ZN(n4597) );
  NAND2_X1 U6200 ( .A1(n5631), .A2(n5630), .ZN(n9293) );
  NOR2_X1 U6201 ( .A1(n5339), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5358) );
  OR2_X1 U6202 ( .A1(n6648), .A2(n4883), .ZN(n4598) );
  AND2_X1 U6203 ( .A1(n8820), .A2(n9218), .ZN(n4599) );
  INV_X1 U6204 ( .A(n8831), .ZN(n5050) );
  AND2_X1 U6205 ( .A1(n8830), .A2(n9142), .ZN(n8831) );
  NAND2_X1 U6206 ( .A1(n6001), .A2(n6000), .ZN(n10157) );
  INV_X1 U6207 ( .A(n10157), .ZN(n7334) );
  OR2_X1 U6208 ( .A1(n5532), .A2(SI_21_), .ZN(n4600) );
  NAND2_X1 U6209 ( .A1(n5574), .A2(n5573), .ZN(n9311) );
  OR2_X1 U6210 ( .A1(n9366), .A2(n4880), .ZN(n4601) );
  NAND2_X1 U6211 ( .A1(n5520), .A2(n5519), .ZN(n9191) );
  INV_X1 U6212 ( .A(n9191), .ZN(n4828) );
  AND2_X1 U6213 ( .A1(n8127), .A2(n4537), .ZN(n4602) );
  XNOR2_X1 U6214 ( .A(n5071), .B(n8965), .ZN(n8166) );
  AND2_X1 U6215 ( .A1(n5333), .A2(n8665), .ZN(n4603) );
  NAND2_X1 U6216 ( .A1(n5298), .A2(n5297), .ZN(n7433) );
  OR2_X1 U6217 ( .A1(n8044), .A2(n7477), .ZN(n4604) );
  NOR2_X1 U6218 ( .A1(n7515), .A2(n7463), .ZN(n4605) );
  AND2_X1 U6219 ( .A1(n5662), .A2(n7892), .ZN(n4606) );
  INV_X1 U6220 ( .A(n6474), .ZN(n4957) );
  INV_X1 U6221 ( .A(n5012), .ZN(n5011) );
  XNOR2_X1 U6222 ( .A(n5135), .B(n5134), .ZN(n5680) );
  INV_X1 U6223 ( .A(n6034), .ZN(n7494) );
  OR2_X1 U6224 ( .A1(n10247), .A2(n4842), .ZN(n4607) );
  AND2_X1 U6225 ( .A1(n9087), .A2(n9080), .ZN(n4608) );
  NAND2_X1 U6226 ( .A1(n9085), .A2(n9076), .ZN(n4914) );
  INV_X1 U6227 ( .A(n9070), .ZN(n4698) );
  AND2_X1 U6228 ( .A1(n4909), .A2(n4914), .ZN(n4609) );
  AND2_X1 U6229 ( .A1(n4698), .A2(n4695), .ZN(n4610) );
  INV_X1 U6230 ( .A(n9544), .ZN(n4645) );
  AND2_X1 U6231 ( .A1(n9611), .A2(n9587), .ZN(n4611) );
  INV_X2 U6232 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U6233 ( .A1(n5605), .A2(n5604), .ZN(n4612) );
  NAND2_X1 U6234 ( .A1(n5586), .A2(n5585), .ZN(n4613) );
  NAND3_X1 U6235 ( .A1(n5444), .A2(n4965), .A3(n4964), .ZN(n5462) );
  AOI21_X1 U6236 ( .B1(n5416), .B2(n5097), .A(n5417), .ZN(n4620) );
  NAND2_X1 U6237 ( .A1(n5394), .A2(n4583), .ZN(n5416) );
  NAND3_X1 U6238 ( .A1(n4960), .A2(n5516), .A3(n5552), .ZN(n4634) );
  MUX2_X1 U6239 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6790), .S(n6804), .Z(n10012)
         );
  INV_X1 U6240 ( .A(n6948), .ZN(n5692) );
  NAND4_X2 U6241 ( .A1(n5133), .A2(n4656), .A3(n4655), .A4(n4654), .ZN(n6948)
         );
  OR2_X1 U6242 ( .A1(n5209), .A2(n6867), .ZN(n4654) );
  NAND2_X1 U6243 ( .A1(n4657), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4656) );
  NAND2_X1 U6244 ( .A1(n4582), .A2(n6906), .ZN(n6863) );
  AND2_X1 U6245 ( .A1(n8705), .A2(n8753), .ZN(n4669) );
  NOR2_X1 U6246 ( .A1(n8712), .A2(n4671), .ZN(n4670) );
  INV_X1 U6247 ( .A(n8716), .ZN(n4671) );
  NAND3_X1 U6248 ( .A1(n4674), .A2(n8716), .A3(n4673), .ZN(n4672) );
  NAND2_X1 U6249 ( .A1(n8704), .A2(n8748), .ZN(n4674) );
  NAND2_X1 U6250 ( .A1(n5122), .A2(n4580), .ZN(n9348) );
  INV_X2 U6251 ( .A(n5744), .ZN(n5122) );
  NAND3_X1 U6252 ( .A1(n4679), .A2(n5352), .A3(n4675), .ZN(n8673) );
  NAND4_X1 U6253 ( .A1(n4680), .A2(n8753), .A3(n8666), .A4(n8667), .ZN(n4679)
         );
  NAND4_X1 U6254 ( .A1(n8663), .A2(n8776), .A3(n8661), .A4(n8662), .ZN(n4680)
         );
  NAND3_X1 U6255 ( .A1(n9071), .A2(n4608), .A3(n10308), .ZN(n4688) );
  INV_X1 U6256 ( .A(n4687), .ZN(n9095) );
  OAI211_X1 U6257 ( .C1(n9071), .C2(n4692), .A(n4689), .B(n4688), .ZN(n4687)
         );
  AND2_X1 U6258 ( .A1(n10308), .A2(n4691), .ZN(n4690) );
  NAND2_X1 U6259 ( .A1(n10308), .A2(n4610), .ZN(n4692) );
  NOR2_X1 U6260 ( .A1(n9071), .A2(n9070), .ZN(n9081) );
  NAND2_X1 U6261 ( .A1(n6905), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U6262 ( .A1(n5122), .A2(n4581), .ZN(n4715) );
  NAND2_X1 U6263 ( .A1(n4721), .A2(n4722), .ZN(n8048) );
  NAND3_X1 U6264 ( .A1(n7473), .A2(n7521), .A3(n4725), .ZN(n4721) );
  NAND2_X1 U6265 ( .A1(n4733), .A2(n4730), .ZN(n4734) );
  OR2_X1 U6266 ( .A1(n6033), .A2(n4737), .ZN(n4733) );
  AND4_X2 U6267 ( .A1(n5805), .A2(n5803), .A3(n5804), .A4(n4741), .ZN(n5895)
         );
  INV_X2 U6268 ( .A(n10113), .ZN(n6504) );
  NAND4_X1 U6269 ( .A1(n6137), .A2(n4536), .A3(n4574), .A4(n4748), .ZN(n5086)
         );
  AND2_X2 U6270 ( .A1(n6504), .A2(n7985), .ZN(n5984) );
  NAND2_X1 U6271 ( .A1(n8486), .A2(n8485), .ZN(n4758) );
  INV_X1 U6272 ( .A(n5098), .ZN(n4761) );
  NAND2_X1 U6273 ( .A1(n9742), .A2(n4578), .ZN(n4765) );
  NAND2_X1 U6274 ( .A1(n4772), .A2(n8124), .ZN(n8292) );
  NAND3_X1 U6275 ( .A1(n4773), .A2(n8074), .A3(n4774), .ZN(n4772) );
  NAND2_X1 U6276 ( .A1(n8035), .A2(n4775), .ZN(n4773) );
  NAND2_X1 U6277 ( .A1(n9818), .A2(n4780), .ZN(n4779) );
  INV_X1 U6278 ( .A(n10375), .ZN(n8646) );
  INV_X1 U6279 ( .A(n4789), .ZN(n4788) );
  NAND2_X1 U6280 ( .A1(n5716), .A2(n4792), .ZN(n4793) );
  NAND2_X1 U6281 ( .A1(n4797), .A2(n4801), .ZN(n5724) );
  NAND2_X1 U6282 ( .A1(n5721), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U6283 ( .A1(n4804), .A2(n4538), .ZN(n9106) );
  NAND2_X1 U6284 ( .A1(n4804), .A2(n4588), .ZN(n4807) );
  NAND2_X1 U6285 ( .A1(n5730), .A2(n4810), .ZN(n9122) );
  INV_X1 U6286 ( .A(n9299), .ZN(n4811) );
  NAND2_X1 U6287 ( .A1(n8471), .A2(n4815), .ZN(n4812) );
  NAND2_X1 U6288 ( .A1(n4812), .A2(n4813), .ZN(n9200) );
  NAND2_X1 U6289 ( .A1(n9185), .A2(n4587), .ZN(n4818) );
  NOR2_X2 U6290 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5868) );
  OAI211_X1 U6291 ( .C1(n9053), .C2(n4908), .A(n4907), .B(n9095), .ZN(P2_U3201) );
  AOI21_X1 U6292 ( .B1(n8147), .B2(n8146), .A(n8145), .ZN(n8204) );
  AND2_X1 U6293 ( .A1(n6976), .A2(n4829), .ZN(n6993) );
  NAND2_X1 U6294 ( .A1(n4831), .A2(n4832), .ZN(n9791) );
  NAND3_X1 U6295 ( .A1(n5074), .A2(n4837), .A3(n5811), .ZN(n4836) );
  NAND2_X1 U6296 ( .A1(n5074), .A2(n5811), .ZN(n4841) );
  NOR2_X1 U6297 ( .A1(n9743), .A2(n9678), .ZN(n9730) );
  INV_X1 U6298 ( .A(n4857), .ZN(n9809) );
  AND2_X1 U6299 ( .A1(n9749), .A2(n4863), .ZN(n9722) );
  NAND2_X1 U6300 ( .A1(n9749), .A2(n4864), .ZN(n9706) );
  NAND2_X1 U6301 ( .A1(n9749), .A2(n9739), .ZN(n9733) );
  NAND2_X1 U6302 ( .A1(n4869), .A2(n4867), .ZN(n10073) );
  NAND2_X1 U6303 ( .A1(n10166), .A2(n7334), .ZN(n4871) );
  NAND2_X1 U6304 ( .A1(n6454), .A2(n4873), .ZN(n4872) );
  NAND2_X1 U6305 ( .A1(n4872), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5822) );
  INV_X2 U6306 ( .A(n5980), .ZN(n6165) );
  NAND3_X1 U6307 ( .A1(n10028), .A2(n6452), .A3(n10014), .ZN(n5971) );
  XNOR2_X1 U6308 ( .A(n6523), .B(n4874), .ZN(n8574) );
  AOI21_X2 U6309 ( .B1(n7176), .B2(n7175), .A(n6531), .ZN(n7226) );
  NAND2_X1 U6310 ( .A1(n8573), .A2(n8574), .ZN(n8572) );
  AOI21_X2 U6311 ( .B1(n6879), .B2(n6876), .A(n6878), .ZN(n8573) );
  NAND2_X1 U6312 ( .A1(n4876), .A2(n4875), .ZN(n9373) );
  AOI21_X2 U6313 ( .B1(n6637), .B2(n4879), .A(n4877), .ZN(n4875) );
  NAND2_X1 U6314 ( .A1(n9455), .A2(n4878), .ZN(n4876) );
  NAND3_X1 U6315 ( .A1(n4886), .A2(n9456), .A3(n4885), .ZN(n4884) );
  NAND2_X1 U6316 ( .A1(n4887), .A2(n4890), .ZN(n6634) );
  NAND2_X1 U6317 ( .A1(n9389), .A2(n4888), .ZN(n4887) );
  NAND2_X1 U6318 ( .A1(n9425), .A2(n6569), .ZN(n8415) );
  NAND2_X1 U6319 ( .A1(n4894), .A2(n4589), .ZN(n6610) );
  NAND2_X1 U6320 ( .A1(n9425), .A2(n4895), .ZN(n4894) );
  INV_X1 U6321 ( .A(n6569), .ZN(n4896) );
  NAND2_X1 U6322 ( .A1(n6548), .A2(n4577), .ZN(n4900) );
  NAND2_X1 U6323 ( .A1(n4900), .A2(n4591), .ZN(n6560) );
  NAND2_X1 U6324 ( .A1(n6660), .A2(n6659), .ZN(n8585) );
  NAND3_X1 U6325 ( .A1(n6660), .A2(n6659), .A3(n4579), .ZN(n4905) );
  AND2_X2 U6326 ( .A1(n5895), .A2(n5809), .ZN(n5867) );
  NAND2_X1 U6327 ( .A1(n9053), .A2(n4609), .ZN(n4907) );
  NOR2_X1 U6328 ( .A1(n9053), .A2(n9052), .ZN(n9078) );
  NAND2_X1 U6329 ( .A1(n4919), .A2(n10429), .ZN(n7113) );
  XNOR2_X1 U6330 ( .A(n8133), .B(n8147), .ZN(n8042) );
  NAND3_X1 U6331 ( .A1(n4926), .A2(P2_REG1_REG_3__SCAN_IN), .A3(n6900), .ZN(
        n10281) );
  NAND2_X1 U6332 ( .A1(n4925), .A2(n5167), .ZN(n10280) );
  NAND2_X1 U6333 ( .A1(n8998), .A2(n4929), .ZN(n4927) );
  INV_X1 U6334 ( .A(n4930), .ZN(n9049) );
  OAI21_X1 U6335 ( .B1(n7516), .B2(n4932), .A(n4931), .ZN(n8040) );
  NAND2_X1 U6336 ( .A1(n4937), .A2(n5189), .ZN(n5192) );
  XNOR2_X1 U6337 ( .A(n4937), .B(n5189), .ZN(n6746) );
  NAND2_X1 U6338 ( .A1(n4938), .A2(n9857), .ZN(n5073) );
  NAND2_X1 U6339 ( .A1(n4940), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U6340 ( .A1(n4941), .A2(n6504), .ZN(n4940) );
  NAND3_X1 U6341 ( .A1(n4950), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4949) );
  NAND3_X1 U6342 ( .A1(n9634), .A2(n4953), .A3(n4952), .ZN(n4951) );
  NAND2_X1 U6343 ( .A1(n5204), .A2(n5203), .ZN(n5226) );
  NAND2_X1 U6344 ( .A1(n4954), .A2(n5228), .ZN(n5237) );
  NAND2_X1 U6345 ( .A1(n5226), .A2(n4955), .ZN(n4954) );
  NAND2_X1 U6346 ( .A1(n5337), .A2(n4967), .ZN(n4965) );
  NAND2_X1 U6347 ( .A1(n5337), .A2(n4970), .ZN(n4966) );
  NAND2_X2 U6348 ( .A1(n4966), .A2(n5355), .ZN(n5440) );
  INV_X1 U6349 ( .A(n8628), .ZN(n8650) );
  NAND2_X1 U6350 ( .A1(n4979), .A2(n4977), .ZN(n7434) );
  NAND2_X1 U6351 ( .A1(n5234), .A2(n4980), .ZN(n4979) );
  NAND4_X1 U6352 ( .A1(n4988), .A2(n4990), .A3(n4987), .A4(n4985), .ZN(n5744)
         );
  NAND2_X1 U6353 ( .A1(n4990), .A2(n4986), .ZN(n5339) );
  INV_X1 U6354 ( .A(n5116), .ZN(n4990) );
  NAND2_X1 U6355 ( .A1(n9197), .A2(n4996), .ZN(n4993) );
  NAND2_X1 U6356 ( .A1(n4993), .A2(n4586), .ZN(n9176) );
  NAND3_X1 U6357 ( .A1(n4999), .A2(n4998), .A3(n8698), .ZN(n8703) );
  NAND2_X1 U6358 ( .A1(n7433), .A2(n5008), .ZN(n5315) );
  NAND2_X1 U6359 ( .A1(n8230), .A2(n5014), .ZN(n5010) );
  OAI21_X1 U6360 ( .B1(n9146), .B2(n5023), .A(n4585), .ZN(n5643) );
  OAI22_X1 U6361 ( .A1(n8678), .A2(n5028), .B1(n5027), .B2(n8675), .ZN(n5030)
         );
  NAND2_X1 U6362 ( .A1(n5030), .A2(n8679), .ZN(n8684) );
  NAND2_X1 U6363 ( .A1(n5122), .A2(n5031), .ZN(n5034) );
  OR2_X1 U6364 ( .A1(n5487), .A2(n9346), .ZN(n5035) );
  NAND2_X1 U6365 ( .A1(n5487), .A2(n5039), .ZN(n5036) );
  NAND2_X1 U6366 ( .A1(n5035), .A2(n5037), .ZN(n5041) );
  NAND2_X1 U6367 ( .A1(n5487), .A2(n5486), .ZN(n5672) );
  INV_X1 U6368 ( .A(n8829), .ZN(n5043) );
  INV_X1 U6369 ( .A(n8828), .ZN(n5044) );
  NAND2_X1 U6370 ( .A1(n8537), .A2(n5055), .ZN(n5054) );
  NAND2_X1 U6371 ( .A1(n5358), .A2(n5060), .ZN(n5485) );
  NAND2_X1 U6372 ( .A1(n7566), .A2(n7565), .ZN(n5071) );
  AND2_X2 U6373 ( .A1(n5066), .A2(n5063), .ZN(n8223) );
  INV_X1 U6374 ( .A(n5064), .ZN(n5063) );
  INV_X1 U6375 ( .A(n8225), .ZN(n5065) );
  NAND2_X1 U6376 ( .A1(n7566), .A2(n5067), .ZN(n5066) );
  NAND2_X1 U6377 ( .A1(n5073), .A2(n5072), .ZN(n6470) );
  INV_X1 U6378 ( .A(n6451), .ZN(n5072) );
  NAND2_X1 U6379 ( .A1(n5075), .A2(n4584), .ZN(n5077) );
  NAND2_X1 U6380 ( .A1(n5082), .A2(n6176), .ZN(n6204) );
  NAND2_X1 U6381 ( .A1(n6205), .A2(n6164), .ZN(n5082) );
  NAND2_X1 U6382 ( .A1(n5084), .A2(n5083), .ZN(n6205) );
  NAND2_X1 U6383 ( .A1(n5086), .A2(n5085), .ZN(n5084) );
  NAND2_X1 U6384 ( .A1(n6136), .A2(n6135), .ZN(n5085) );
  OAI21_X2 U6385 ( .B1(n6535), .B2(n6534), .A(n7224), .ZN(n7505) );
  NAND2_X1 U6386 ( .A1(n9639), .A2(n6476), .ZN(n9854) );
  NAND2_X1 U6387 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5140) );
  NAND2_X1 U6388 ( .A1(n5821), .A2(n5820), .ZN(n6452) );
  NAND2_X1 U6389 ( .A1(n5818), .A2(n5817), .ZN(n5821) );
  NAND2_X1 U6390 ( .A1(n8494), .A2(n9972), .ZN(n8553) );
  INV_X1 U6392 ( .A(n5218), .ZN(n5129) );
  AOI21_X2 U6393 ( .B1(n7326), .B2(n7278), .A(n7277), .ZN(n7377) );
  NAND2_X2 U6394 ( .A1(n8510), .A2(n8509), .ZN(n8537) );
  NOR2_X1 U6395 ( .A1(n8813), .A2(n5741), .ZN(n5742) );
  OAI21_X2 U6396 ( .B1(n8869), .B2(n8865), .A(n8866), .ZN(n8908) );
  MUX2_X1 U6397 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9953), .S(n5980), .Z(n6976) );
  NAND4_X1 U6398 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n5981)
         );
  NAND2_X1 U6399 ( .A1(n6043), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U6400 ( .A1(n5829), .A2(n5827), .ZN(n5832) );
  NAND2_X1 U6401 ( .A1(n6391), .A2(n7206), .ZN(n5985) );
  OAI22_X2 U6402 ( .A1(n8941), .A2(n8835), .B1(n9143), .B2(n8834), .ZN(n8853)
         );
  NAND2_X1 U6403 ( .A1(n6976), .A2(n6511), .ZN(n6513) );
  INV_X1 U6404 ( .A(n6306), .ZN(n7210) );
  AOI21_X2 U6405 ( .B1(n9786), .B2(n9656), .A(n9655), .ZN(n9773) );
  OAI22_X2 U6406 ( .A1(n8908), .A2(n8909), .B1(n8823), .B2(n8956), .ZN(n8875)
         );
  AOI21_X2 U6407 ( .B1(n8964), .B2(n8225), .A(n8223), .ZN(n8344) );
  OR3_X1 U6408 ( .A1(n6462), .A2(n6461), .A3(n6473), .ZN(n5094) );
  OR2_X1 U6409 ( .A1(n9961), .A2(n9649), .ZN(n5095) );
  OR2_X1 U6410 ( .A1(n5415), .A2(n7762), .ZN(n5097) );
  OR2_X1 U6411 ( .A1(n8487), .A2(n9395), .ZN(n5098) );
  NAND2_X1 U6412 ( .A1(n8009), .A2(n8008), .ZN(n5099) );
  INV_X1 U6413 ( .A(n9504), .ZN(n8289) );
  AND2_X1 U6414 ( .A1(n5300), .A2(n5279), .ZN(n5100) );
  INV_X1 U6415 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5178) );
  INV_X1 U6416 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5139) );
  OR2_X1 U6417 ( .A1(n10226), .A2(n6497), .ZN(n5101) );
  NAND2_X1 U6418 ( .A1(n8791), .A2(n8603), .ZN(n8742) );
  NOR2_X1 U6419 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5102) );
  INV_X1 U6420 ( .A(n9167), .ZN(n9142) );
  AND2_X1 U6421 ( .A1(n5443), .A2(SI_16_), .ZN(n5103) );
  NOR2_X1 U6422 ( .A1(n5442), .A2(n5441), .ZN(n5104) );
  NOR2_X1 U6423 ( .A1(n9636), .A2(n9686), .ZN(n5105) );
  AND2_X1 U6424 ( .A1(n10400), .A2(n8967), .ZN(n5106) );
  INV_X1 U6425 ( .A(n9906), .ZN(n9651) );
  OR2_X1 U6426 ( .A1(n9675), .A2(n5984), .ZN(n5107) );
  AND3_X1 U6427 ( .A1(n6714), .A2(n6713), .A3(n10000), .ZN(n5108) );
  OR2_X1 U6428 ( .A1(n10440), .A2(n5784), .ZN(n5109) );
  NOR4_X1 U6429 ( .A1(n9819), .A2(n9805), .A3(n9840), .A4(n6322), .ZN(n5110)
         );
  INV_X1 U6430 ( .A(n6426), .ZN(n6175) );
  INV_X1 U6431 ( .A(n8442), .ZN(n10213) );
  INV_X1 U6432 ( .A(n8780), .ZN(n5352) );
  NAND2_X1 U6433 ( .A1(n5987), .A2(n9858), .ZN(n5988) );
  NAND2_X1 U6434 ( .A1(n6303), .A2(n5984), .ZN(n6174) );
  AND2_X1 U6435 ( .A1(n6428), .A2(n9858), .ZN(n6207) );
  INV_X1 U6436 ( .A(n6364), .ZN(n6436) );
  INV_X1 U6437 ( .A(n7237), .ZN(n5699) );
  NOR2_X1 U6438 ( .A1(n7428), .A2(n5704), .ZN(n5705) );
  INV_X1 U6439 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5111) );
  INV_X1 U6440 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5813) );
  NOR2_X1 U6441 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5805) );
  OR2_X1 U6442 ( .A1(n8826), .A2(n9188), .ZN(n8827) );
  AND2_X1 U6443 ( .A1(n8762), .A2(n9158), .ZN(n8723) );
  OR2_X1 U6444 ( .A1(n8416), .A2(n8417), .ZN(n6575) );
  INV_X1 U6445 ( .A(n9805), .ZN(n9674) );
  NAND2_X1 U6446 ( .A1(n7972), .A2(n5813), .ZN(n5814) );
  INV_X1 U6447 ( .A(n5235), .ZN(n5236) );
  INV_X1 U6448 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5245) );
  NOR2_X1 U6449 ( .A1(n9311), .A2(n9167), .ZN(n5727) );
  INV_X1 U6450 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5210) );
  INV_X1 U6451 ( .A(n8742), .ZN(n5733) );
  OR2_X1 U6452 ( .A1(n7393), .A2(n8968), .ZN(n7320) );
  AND2_X1 U6453 ( .A1(n6666), .A2(n6665), .ZN(n6668) );
  OAI21_X1 U6454 ( .B1(n5961), .B2(n6750), .A(n5998), .ZN(n5999) );
  INV_X1 U6455 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5816) );
  INV_X1 U6456 ( .A(n5253), .ZN(n5254) );
  AND2_X1 U6457 ( .A1(n8535), .A2(n8536), .ZN(n8534) );
  OAI22_X1 U6458 ( .A1(n8600), .A2(n8599), .B1(n9284), .B2(n9278), .ZN(n8606)
         );
  AOI21_X1 U6459 ( .B1(n4706), .B2(n7190), .A(n7189), .ZN(n7192) );
  AND2_X1 U6460 ( .A1(n9036), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9024) );
  INV_X1 U6461 ( .A(n5493), .ZN(n5492) );
  INV_X1 U6462 ( .A(n8773), .ZN(n5297) );
  OAI22_X1 U6463 ( .A1(n9140), .A2(n8729), .B1(n9153), .B2(n9305), .ZN(n9133)
         );
  NAND2_X1 U6464 ( .A1(n5744), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6465 ( .A1(n6542), .A2(n6541), .ZN(n6546) );
  INV_X1 U6466 ( .A(n6528), .ZN(n6530) );
  NOR2_X1 U6467 ( .A1(n6075), .A2(n7047), .ZN(n6074) );
  OR2_X1 U6468 ( .A1(n9739), .A2(n6503), .ZN(n6680) );
  OR2_X1 U6469 ( .A1(n6168), .A2(n9368), .ZN(n6179) );
  OAI22_X1 U6470 ( .A1(n9721), .A2(n9991), .B1(n9687), .B2(n9686), .ZN(n9688)
         );
  INV_X1 U6471 ( .A(n9670), .ZN(n9684) );
  AND2_X1 U6472 ( .A1(n9900), .A2(n9654), .ZN(n9655) );
  INV_X1 U6473 ( .A(n5999), .ZN(n6000) );
  NAND2_X1 U6474 ( .A1(n6390), .A2(n10090), .ZN(n5986) );
  NOR2_X1 U6475 ( .A1(n8442), .A2(n8289), .ZN(n8290) );
  NOR2_X1 U6476 ( .A1(n5104), .A2(n5103), .ZN(n5444) );
  NAND2_X1 U6477 ( .A1(n5321), .A2(n7904), .ZN(n5336) );
  INV_X1 U6478 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7935) );
  XNOR2_X1 U6479 ( .A(n7132), .B(n8646), .ZN(n7125) );
  AOI21_X1 U6480 ( .B1(n7166), .B2(n7165), .A(n7164), .ZN(n7167) );
  NAND2_X1 U6481 ( .A1(n5596), .A2(n5595), .ZN(n5614) );
  AND2_X1 U6482 ( .A1(n8716), .A2(n5725), .ZN(n9189) );
  INV_X1 U6483 ( .A(n8164), .ZN(n8776) );
  AND2_X1 U6484 ( .A1(n8748), .A2(n5778), .ZN(n7096) );
  INV_X1 U6485 ( .A(n5783), .ZN(n8808) );
  NAND2_X1 U6486 ( .A1(n8321), .A2(n5421), .ZN(n5631) );
  INV_X1 U6487 ( .A(n8729), .ZN(n9147) );
  AND2_X1 U6488 ( .A1(n6609), .A2(n6608), .ZN(n8389) );
  OR2_X1 U6489 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  OR2_X1 U6490 ( .A1(n6041), .A2(n6040), .ZN(n6052) );
  NOR2_X1 U6491 ( .A1(n6142), .A2(n6141), .ZN(n6158) );
  INV_X1 U6492 ( .A(n9648), .ZN(n9649) );
  NOR2_X1 U6493 ( .A1(n6179), .A2(n9440), .ZN(n6194) );
  NOR2_X1 U6494 ( .A1(n6798), .A2(n6797), .ZN(n6821) );
  INV_X1 U6495 ( .A(n9646), .ZN(n9837) );
  INV_X1 U6496 ( .A(n7271), .ZN(n7205) );
  INV_X1 U6497 ( .A(n9850), .ZN(n9961) );
  AND2_X1 U6498 ( .A1(n6413), .A2(n6415), .ZN(n8293) );
  INV_X1 U6499 ( .A(n9834), .ZN(n9989) );
  INV_X1 U6500 ( .A(n9179), .ZN(n8919) );
  INV_X1 U6501 ( .A(n8601), .ZN(n9097) );
  OAI21_X1 U6502 ( .B1(n8808), .B2(n9263), .A(n5109), .ZN(n5785) );
  INV_X1 U6503 ( .A(n9263), .ZN(n9270) );
  INV_X1 U6504 ( .A(n9331), .ZN(n9338) );
  AND2_X1 U6505 ( .A1(n7141), .A2(n7984), .ZN(n10404) );
  NAND2_X1 U6506 ( .A1(n6711), .A2(n6710), .ZN(n6712) );
  AND4_X1 U6507 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n9721)
         );
  AND4_X1 U6508 ( .A1(n6244), .A2(n6243), .A3(n6242), .A4(n6241), .ZN(n9747)
         );
  AND4_X1 U6509 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n9486)
         );
  AND4_X1 U6510 ( .A1(n5912), .A2(n5911), .A3(n5910), .A4(n5909), .ZN(n8288)
         );
  AND2_X1 U6511 ( .A1(n6986), .A2(n7352), .ZN(n10099) );
  NOR2_X1 U6512 ( .A1(n9864), .A2(n4552), .ZN(n9865) );
  NAND2_X1 U6513 ( .A1(n9859), .A2(n10134), .ZN(n10222) );
  AND2_X1 U6514 ( .A1(n6479), .A2(n6478), .ZN(n9937) );
  INV_X1 U6515 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6456) );
  AND2_X1 U6516 ( .A1(n6086), .A2(n6098), .ZN(n7359) );
  XNOR2_X1 U6517 ( .A(n5202), .B(n5193), .ZN(n5200) );
  INV_X1 U6518 ( .A(n8944), .ZN(n8933) );
  AND2_X1 U6519 ( .A1(n6961), .A2(n6960), .ZN(n8953) );
  NAND2_X1 U6520 ( .A1(n5656), .A2(n5655), .ZN(n9123) );
  OR2_X1 U6521 ( .A1(P2_U3150), .A2(n6860), .ZN(n10321) );
  INV_X1 U6522 ( .A(n5785), .ZN(n5786) );
  INV_X1 U6523 ( .A(n10440), .ZN(n10437) );
  INV_X1 U6524 ( .A(n9231), .ZN(n9284) );
  AND2_X1 U6525 ( .A1(n5798), .A2(n5797), .ZN(n10423) );
  INV_X1 U6526 ( .A(n7466), .ZN(n7459) );
  INV_X1 U6527 ( .A(n6908), .ZN(n10286) );
  NOR2_X1 U6528 ( .A1(n5108), .A2(n6729), .ZN(n6730) );
  AND4_X1 U6529 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n7234)
         );
  INV_X1 U6530 ( .A(n9808), .ZN(n9654) );
  INV_X1 U6531 ( .A(n10247), .ZN(n10244) );
  INV_X1 U6532 ( .A(n10226), .ZN(n10224) );
  INV_X1 U6533 ( .A(n10127), .ZN(n10122) );
  INV_X1 U6534 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U6535 ( .A1(n6498), .A2(n5101), .ZN(P1_U3521) );
  NOR2_X1 U6536 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5114) );
  NAND4_X1 U6537 ( .A1(n5114), .A2(n5113), .A3(n5112), .A4(n5111), .ZN(n5116)
         );
  NOR2_X1 U6538 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5119) );
  NOR2_X1 U6539 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5118) );
  NOR2_X1 U6540 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5117) );
  INV_X1 U6541 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6542 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5123) );
  NAND2_X1 U6543 ( .A1(n5135), .A2(n5123), .ZN(n5124) );
  NOR2_X1 U6544 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5125) );
  NAND2_X1 U6545 ( .A1(n9348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6546 ( .A1(n5129), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5133) );
  INV_X1 U6547 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5131) );
  INV_X1 U6548 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6867) );
  INV_X1 U6549 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5134) );
  INV_X1 U6550 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5136) );
  AND2_X1 U6551 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5137) );
  XNOR2_X1 U6552 ( .A(n5157), .B(SI_1_), .ZN(n6745) );
  INV_X1 U6553 ( .A(n6884), .ZN(n6871) );
  NAND2_X1 U6554 ( .A1(n5342), .A2(n6871), .ZN(n5143) );
  NAND2_X1 U6555 ( .A1(n5206), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6556 ( .A1(n10360), .A2(n6948), .ZN(n8608) );
  NAND2_X1 U6557 ( .A1(n8615), .A2(n8608), .ZN(n8766) );
  INV_X1 U6558 ( .A(n8766), .ZN(n5151) );
  NAND2_X1 U6559 ( .A1(n5379), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5148) );
  OR2_X1 U6560 ( .A1(n5188), .A2(n4668), .ZN(n5146) );
  INV_X1 U6561 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6562 ( .A1(n5218), .A2(n5144), .ZN(n5145) );
  NAND2_X1 U6563 ( .A1(n6743), .A2(SI_0_), .ZN(n5149) );
  XNOR2_X1 U6564 ( .A(n5149), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9356) );
  MUX2_X1 U6565 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9356), .S(n6736), .Z(n8582) );
  NAND2_X1 U6566 ( .A1(n6844), .A2(n8582), .ZN(n8612) );
  NAND2_X1 U6567 ( .A1(n5151), .A2(n5150), .ZN(n7152) );
  NAND2_X1 U6568 ( .A1(n7152), .A2(n8615), .ZN(n10340) );
  NAND2_X1 U6569 ( .A1(n5636), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6570 ( .A1(n4657), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5155) );
  INV_X1 U6571 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10342) );
  OR2_X1 U6572 ( .A1(n5209), .A2(n10342), .ZN(n5154) );
  INV_X1 U6573 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5152) );
  OR2_X1 U6574 ( .A1(n5218), .A2(n5152), .ZN(n5153) );
  INV_X1 U6575 ( .A(n5158), .ZN(n5159) );
  NAND2_X1 U6576 ( .A1(n5160), .A2(n5159), .ZN(n5161) );
  MUX2_X1 U6577 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5162), .Z(n5175) );
  INV_X1 U6578 ( .A(SI_2_), .ZN(n7704) );
  XNOR2_X1 U6579 ( .A(n5175), .B(n7704), .ZN(n5173) );
  XNOR2_X1 U6580 ( .A(n5174), .B(n5173), .ZN(n6748) );
  NAND2_X1 U6581 ( .A1(n5206), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6582 ( .A1(n5470), .A2(n6903), .ZN(n5164) );
  INV_X1 U6583 ( .A(n7067), .ZN(n10365) );
  NAND2_X1 U6584 ( .A1(n10365), .A2(n10327), .ZN(n8619) );
  INV_X1 U6585 ( .A(n10344), .ZN(n8617) );
  NAND2_X1 U6586 ( .A1(n10340), .A2(n8617), .ZN(n5166) );
  NAND2_X1 U6587 ( .A1(n5166), .A2(n8620), .ZN(n10331) );
  NAND2_X1 U6588 ( .A1(n5636), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5172) );
  OR2_X1 U6589 ( .A1(n5209), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5171) );
  INV_X1 U6590 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5167) );
  OR2_X1 U6591 ( .A1(n5188), .A2(n5167), .ZN(n5170) );
  INV_X1 U6592 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5168) );
  OR2_X1 U6593 ( .A1(n5218), .A2(n5168), .ZN(n5169) );
  NAND2_X1 U6594 ( .A1(n5175), .A2(SI_2_), .ZN(n5176) );
  INV_X2 U6595 ( .A(n6743), .ZN(n6738) );
  INV_X1 U6596 ( .A(SI_3_), .ZN(n7754) );
  XNOR2_X1 U6597 ( .A(n5190), .B(n7754), .ZN(n5189) );
  NAND2_X1 U6598 ( .A1(n5206), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6599 ( .A1(n5179), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5180) );
  XNOR2_X1 U6600 ( .A(n5180), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U6601 ( .A1(n5342), .A2(n6908), .ZN(n5181) );
  INV_X1 U6602 ( .A(n10369), .ZN(n10333) );
  XNOR2_X1 U6603 ( .A(n10347), .B(n10333), .ZN(n10332) );
  NAND2_X1 U6604 ( .A1(n10331), .A2(n10332), .ZN(n5183) );
  NAND2_X1 U6605 ( .A1(n10347), .A2(n10369), .ZN(n8649) );
  NAND2_X1 U6606 ( .A1(n5183), .A2(n8649), .ZN(n7140) );
  INV_X1 U6607 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6608 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5187) );
  AND2_X1 U6609 ( .A1(n5212), .A2(n5187), .ZN(n7087) );
  INV_X1 U6610 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7020) );
  NAND2_X1 U6611 ( .A1(n5190), .A2(SI_3_), .ZN(n5191) );
  NAND2_X1 U6612 ( .A1(n5192), .A2(n5191), .ZN(n5201) );
  MUX2_X1 U6613 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6738), .Z(n5202) );
  INV_X1 U6614 ( .A(SI_4_), .ZN(n5193) );
  NAND2_X1 U6615 ( .A1(n5206), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6616 ( .A1(n5198), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6617 ( .A(n5194), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U6618 ( .A1(n5342), .A2(n7029), .ZN(n5195) );
  NAND2_X1 U6619 ( .A1(n7140), .A2(n4785), .ZN(n5197) );
  NAND2_X1 U6620 ( .A1(n8647), .A2(n8646), .ZN(n8626) );
  NAND2_X1 U6621 ( .A1(n5197), .A2(n8626), .ZN(n7235) );
  NOR2_X1 U6622 ( .A1(n5198), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5230) );
  OR2_X1 U6623 ( .A1(n5230), .A2(n9346), .ZN(n5199) );
  XNOR2_X1 U6624 ( .A(n5199), .B(n5229), .ZN(n7118) );
  NAND2_X1 U6625 ( .A1(n5202), .A2(SI_4_), .ZN(n5203) );
  MUX2_X1 U6626 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6744), .Z(n5227) );
  XNOR2_X1 U6627 ( .A(n5226), .B(n5225), .ZN(n6013) );
  INV_X2 U6628 ( .A(n5205), .ZN(n5421) );
  NAND2_X1 U6629 ( .A1(n6013), .A2(n5421), .ZN(n5208) );
  NAND2_X1 U6630 ( .A1(n5539), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5207) );
  OAI211_X1 U6631 ( .C1(n6736), .C2(n7118), .A(n5208), .B(n5207), .ZN(n7246)
         );
  INV_X1 U6632 ( .A(n7246), .ZN(n10379) );
  NAND2_X1 U6633 ( .A1(n7420), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6634 ( .A1(n5636), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6635 ( .A1(n5212), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5213) );
  AND2_X1 U6636 ( .A1(n5219), .A2(n5213), .ZN(n7243) );
  OR2_X1 U6637 ( .A1(n5209), .A2(n7243), .ZN(n5215) );
  OR2_X1 U6638 ( .A1(n5188), .A2(n10429), .ZN(n5214) );
  NAND2_X1 U6639 ( .A1(n10379), .A2(n8970), .ZN(n8645) );
  NAND2_X1 U6640 ( .A1(n7235), .A2(n8645), .ZN(n7253) );
  NAND2_X1 U6641 ( .A1(n7420), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6642 ( .A1(n5636), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6643 ( .A1(n5219), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5220) );
  AND2_X1 U6644 ( .A1(n5247), .A2(n5220), .ZN(n7169) );
  OR2_X1 U6645 ( .A1(n5209), .A2(n7169), .ZN(n5222) );
  INV_X1 U6646 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7024) );
  OR2_X1 U6647 ( .A1(n5683), .A2(n7024), .ZN(n5221) );
  NAND4_X1 U6648 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n8969)
         );
  INV_X1 U6649 ( .A(n8969), .ZN(n7398) );
  NAND2_X1 U6650 ( .A1(n5227), .A2(SI_5_), .ZN(n5228) );
  MUX2_X1 U6651 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6744), .Z(n5238) );
  XNOR2_X1 U6652 ( .A(n5237), .B(n5235), .ZN(n6025) );
  NAND2_X1 U6653 ( .A1(n6025), .A2(n5421), .ZN(n5233) );
  NAND2_X1 U6654 ( .A1(n5230), .A2(n5229), .ZN(n5240) );
  NAND2_X1 U6655 ( .A1(n5240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5231) );
  AOI22_X1 U6656 ( .A1(n5539), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5470), .B2(
        n7036), .ZN(n5232) );
  NAND2_X1 U6657 ( .A1(n5233), .A2(n5232), .ZN(n7259) );
  NAND2_X1 U6658 ( .A1(n7398), .A2(n7259), .ZN(n8629) );
  INV_X1 U6659 ( .A(n8970), .ZN(n7162) );
  NAND2_X1 U6660 ( .A1(n7162), .A2(n7246), .ZN(n7252) );
  AND2_X1 U6661 ( .A1(n8629), .A2(n7252), .ZN(n8651) );
  NAND2_X1 U6662 ( .A1(n7253), .A2(n8651), .ZN(n5234) );
  INV_X1 U6663 ( .A(n7259), .ZN(n10386) );
  NAND2_X1 U6664 ( .A1(n10386), .A2(n8969), .ZN(n8652) );
  NAND2_X1 U6665 ( .A1(n5238), .A2(SI_6_), .ZN(n5239) );
  MUX2_X1 U6666 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6744), .Z(n5256) );
  XNOR2_X1 U6667 ( .A(n5255), .B(n5253), .ZN(n6767) );
  NAND2_X1 U6668 ( .A1(n6767), .A2(n5421), .ZN(n5244) );
  NAND2_X1 U6669 ( .A1(n5283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  INV_X1 U6670 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6671 ( .A1(n5241), .A2(n5281), .ZN(n5262) );
  OR2_X1 U6672 ( .A1(n5241), .A2(n5281), .ZN(n5242) );
  AOI22_X1 U6673 ( .A1(n5539), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5470), .B2(
        n7197), .ZN(n5243) );
  NAND2_X1 U6674 ( .A1(n5244), .A2(n5243), .ZN(n7393) );
  NAND2_X1 U6675 ( .A1(n7420), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6676 ( .A1(n5636), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6677 ( .A1(n5247), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5248) );
  AND2_X1 U6678 ( .A1(n5267), .A2(n5248), .ZN(n7402) );
  OR2_X1 U6679 ( .A1(n5209), .A2(n7402), .ZN(n5250) );
  INV_X1 U6680 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7015) );
  OR2_X1 U6681 ( .A1(n5188), .A2(n7015), .ZN(n5249) );
  NAND4_X1 U6682 ( .A1(n5252), .A2(n5251), .A3(n5250), .A4(n5249), .ZN(n8968)
         );
  NAND2_X1 U6683 ( .A1(n7393), .A2(n7341), .ZN(n8656) );
  NAND2_X1 U6684 ( .A1(n5256), .A2(SI_7_), .ZN(n5257) );
  INV_X1 U6685 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6772) );
  MUX2_X1 U6686 ( .A(n6772), .B(n7772), .S(n6744), .Z(n5259) );
  INV_X1 U6687 ( .A(SI_8_), .ZN(n5258) );
  INV_X1 U6688 ( .A(n5259), .ZN(n5260) );
  NAND2_X1 U6689 ( .A1(n5260), .A2(SI_8_), .ZN(n5261) );
  NAND2_X1 U6690 ( .A1(n6771), .A2(n5421), .ZN(n5265) );
  NAND2_X1 U6691 ( .A1(n5262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5263) );
  XNOR2_X1 U6692 ( .A(n5263), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7466) );
  AOI22_X1 U6693 ( .A1(n5539), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5470), .B2(
        n7466), .ZN(n5264) );
  NAND2_X1 U6694 ( .A1(n7420), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5273) );
  INV_X1 U6695 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6696 ( .A1(n5287), .A2(n5266), .ZN(n5272) );
  NAND2_X1 U6697 ( .A1(n5267), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5268) );
  AND2_X1 U6698 ( .A1(n5291), .A2(n5268), .ZN(n7344) );
  OR2_X1 U6699 ( .A1(n5209), .A2(n7344), .ZN(n5271) );
  INV_X1 U6700 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5269) );
  OR2_X1 U6701 ( .A1(n5188), .A2(n5269), .ZN(n5270) );
  NAND4_X1 U6702 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n8967)
         );
  OR2_X1 U6703 ( .A1(n10400), .A2(n7536), .ZN(n8636) );
  AND2_X1 U6704 ( .A1(n8636), .A2(n7318), .ZN(n8633) );
  NAND2_X1 U6705 ( .A1(n10400), .A2(n7536), .ZN(n8657) );
  INV_X1 U6706 ( .A(n7434), .ZN(n5298) );
  INV_X1 U6707 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6779) );
  MUX2_X1 U6708 ( .A(n6779), .B(n7881), .S(n6744), .Z(n5277) );
  INV_X1 U6709 ( .A(SI_9_), .ZN(n7922) );
  NAND2_X1 U6710 ( .A1(n5277), .A2(n7922), .ZN(n5300) );
  INV_X1 U6711 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6712 ( .A1(n5278), .A2(SI_9_), .ZN(n5279) );
  INV_X1 U6713 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6714 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  OAI21_X1 U6715 ( .B1(n5283), .B2(n5282), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5284) );
  XNOR2_X1 U6716 ( .A(n5284), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7468) );
  AOI22_X1 U6717 ( .A1(n5539), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5470), .B2(
        n7468), .ZN(n5285) );
  NAND2_X1 U6718 ( .A1(n7420), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6719 ( .A1(n4657), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5295) );
  INV_X1 U6720 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5288) );
  OR2_X1 U6721 ( .A1(n5287), .A2(n5288), .ZN(n5294) );
  INV_X1 U6722 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6723 ( .A1(n5291), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5292) );
  AND2_X1 U6724 ( .A1(n5308), .A2(n5292), .ZN(n7531) );
  OR2_X1 U6725 ( .A1(n5209), .A2(n7531), .ZN(n5293) );
  NAND4_X1 U6726 ( .A1(n5296), .A2(n5295), .A3(n5294), .A4(n5293), .ZN(n8966)
         );
  NAND2_X1 U6727 ( .A1(n10403), .A2(n7567), .ZN(n8662) );
  NAND2_X1 U6728 ( .A1(n8639), .A2(n8662), .ZN(n8773) );
  NAND2_X1 U6729 ( .A1(n5301), .A2(n5300), .ZN(n5320) );
  MUX2_X1 U6730 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6744), .Z(n5317) );
  INV_X1 U6731 ( .A(SI_10_), .ZN(n7727) );
  XNOR2_X1 U6732 ( .A(n5320), .B(n5316), .ZN(n6781) );
  NAND2_X1 U6733 ( .A1(n6781), .A2(n5421), .ZN(n5307) );
  OR2_X1 U6734 ( .A1(n5302), .A2(n9346), .ZN(n5304) );
  MUX2_X1 U6735 ( .A(n5304), .B(P2_IR_REG_31__SCAN_IN), .S(n5303), .Z(n5305)
         );
  AND2_X1 U6736 ( .A1(n5339), .A2(n5305), .ZN(n8044) );
  AOI22_X1 U6737 ( .A1(n5539), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5470), .B2(
        n8044), .ZN(n5306) );
  NAND2_X1 U6738 ( .A1(n5307), .A2(n5306), .ZN(n10412) );
  NAND2_X1 U6739 ( .A1(n7420), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5313) );
  INV_X1 U6740 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7477) );
  OR2_X1 U6741 ( .A1(n5287), .A2(n7477), .ZN(n5312) );
  NAND2_X1 U6742 ( .A1(n5308), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5309) );
  AND2_X1 U6743 ( .A1(n5327), .A2(n5309), .ZN(n7571) );
  OR2_X1 U6744 ( .A1(n5209), .A2(n7571), .ZN(n5311) );
  INV_X1 U6745 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7476) );
  OR2_X1 U6746 ( .A1(n5683), .A2(n7476), .ZN(n5310) );
  NAND4_X1 U6747 ( .A1(n5313), .A2(n5312), .A3(n5311), .A4(n5310), .ZN(n8965)
         );
  INV_X1 U6748 ( .A(n8965), .ZN(n8217) );
  NOR2_X1 U6749 ( .A1(n10412), .A2(n8217), .ZN(n8664) );
  INV_X1 U6750 ( .A(n8664), .ZN(n5314) );
  NAND2_X1 U6751 ( .A1(n10412), .A2(n8217), .ZN(n8661) );
  NAND2_X1 U6752 ( .A1(n5315), .A2(n8661), .ZN(n7988) );
  NAND2_X1 U6753 ( .A1(n5317), .A2(SI_10_), .ZN(n5318) );
  INV_X1 U6754 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6818) );
  INV_X1 U6755 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6820) );
  MUX2_X1 U6756 ( .A(n6818), .B(n6820), .S(n6744), .Z(n5321) );
  INV_X1 U6757 ( .A(SI_11_), .ZN(n7904) );
  INV_X1 U6758 ( .A(n5321), .ZN(n5322) );
  NAND2_X1 U6759 ( .A1(n5322), .A2(SI_11_), .ZN(n5323) );
  XNOR2_X1 U6760 ( .A(n5335), .B(n5334), .ZN(n6817) );
  NAND2_X1 U6761 ( .A1(n6817), .A2(n5421), .ZN(n5326) );
  NAND2_X1 U6762 ( .A1(n5339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5324) );
  XNOR2_X1 U6763 ( .A(n5324), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8147) );
  AOI22_X1 U6764 ( .A1(n5539), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5470), .B2(
        n8147), .ZN(n5325) );
  NAND2_X1 U6765 ( .A1(n7420), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5332) );
  INV_X1 U6766 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7996) );
  OR2_X1 U6767 ( .A1(n5287), .A2(n7996), .ZN(n5331) );
  NAND2_X1 U6768 ( .A1(n5327), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5328) );
  AND2_X1 U6769 ( .A1(n5346), .A2(n5328), .ZN(n8222) );
  OR2_X1 U6770 ( .A1(n5209), .A2(n8222), .ZN(n5330) );
  OR2_X1 U6771 ( .A1(n5683), .A2(n10438), .ZN(n5329) );
  NAND2_X1 U6772 ( .A1(n10417), .A2(n8168), .ZN(n8665) );
  NAND2_X1 U6773 ( .A1(n8667), .A2(n8665), .ZN(n8164) );
  NAND2_X1 U6774 ( .A1(n7988), .A2(n8776), .ZN(n5333) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6744), .Z(n5354) );
  INV_X1 U6776 ( .A(SI_12_), .ZN(n5338) );
  NAND2_X1 U6777 ( .A1(n6836), .A2(n5421), .ZN(n5344) );
  INV_X1 U6778 ( .A(n5358), .ZN(n5340) );
  NAND2_X1 U6779 ( .A1(n5340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5341) );
  XNOR2_X1 U6780 ( .A(n5341), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8157) );
  AOI22_X1 U6781 ( .A1(n5539), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5342), .B2(
        n8157), .ZN(n5343) );
  NAND2_X1 U6782 ( .A1(n7420), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5351) );
  INV_X1 U6783 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8149) );
  OR2_X1 U6784 ( .A1(n5287), .A2(n8149), .ZN(n5350) );
  INV_X1 U6785 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U6786 ( .A1(n5346), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5347) );
  AND2_X1 U6787 ( .A1(n5364), .A2(n5347), .ZN(n8172) );
  OR2_X1 U6788 ( .A1(n5209), .A2(n8172), .ZN(n5349) );
  INV_X1 U6789 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8148) );
  OR2_X1 U6790 ( .A1(n5683), .A2(n8148), .ZN(n5348) );
  XNOR2_X1 U6791 ( .A(n8669), .B(n8668), .ZN(n8780) );
  OR2_X1 U6792 ( .A1(n8669), .A2(n8668), .ZN(n8671) );
  NAND2_X1 U6793 ( .A1(n5354), .A2(SI_12_), .ZN(n5355) );
  MUX2_X1 U6794 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6744), .Z(n5372) );
  NAND2_X1 U6795 ( .A1(n6848), .A2(n5421), .ZN(n5361) );
  OR2_X1 U6796 ( .A1(n5376), .A2(n9346), .ZN(n5359) );
  XNOR2_X1 U6797 ( .A(n5359), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8364) );
  AOI22_X1 U6798 ( .A1(n5539), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5470), .B2(
        n8364), .ZN(n5360) );
  NAND2_X1 U6799 ( .A1(n7420), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5369) );
  INV_X1 U6800 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8190) );
  OR2_X1 U6801 ( .A1(n5287), .A2(n8190), .ZN(n5368) );
  INV_X1 U6802 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6803 ( .A1(n5364), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5365) );
  AND2_X1 U6804 ( .A1(n5380), .A2(n5365), .ZN(n8350) );
  OR2_X1 U6805 ( .A1(n5209), .A2(n8350), .ZN(n5367) );
  INV_X1 U6806 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8196) );
  OR2_X1 U6807 ( .A1(n5188), .A2(n8196), .ZN(n5366) );
  NAND4_X1 U6808 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n8962)
         );
  INV_X1 U6809 ( .A(n8962), .ZN(n8409) );
  NAND2_X1 U6810 ( .A1(n5714), .A2(n8409), .ZN(n5370) );
  NAND2_X1 U6811 ( .A1(n5440), .A2(n5393), .ZN(n5373) );
  NAND2_X1 U6812 ( .A1(n5372), .A2(SI_13_), .ZN(n5396) );
  NAND2_X1 U6813 ( .A1(n5373), .A2(n5396), .ZN(n5374) );
  MUX2_X1 U6814 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6286), .Z(n5390) );
  NAND2_X1 U6815 ( .A1(n6965), .A2(n5421), .ZN(n5378) );
  INV_X1 U6816 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6817 ( .A1(n5464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U6818 ( .A(n5425), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8373) );
  AOI22_X1 U6819 ( .A1(n5539), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5470), .B2(
        n8373), .ZN(n5377) );
  NAND2_X1 U6820 ( .A1(n7420), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6821 ( .A1(n5380), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6822 ( .A1(n5406), .A2(n5381), .ZN(n8411) );
  NAND2_X1 U6823 ( .A1(n5379), .A2(n8411), .ZN(n5385) );
  INV_X1 U6824 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5382) );
  OR2_X1 U6825 ( .A1(n5287), .A2(n5382), .ZN(n5384) );
  INV_X1 U6826 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8269) );
  OR2_X1 U6827 ( .A1(n5188), .A2(n8269), .ZN(n5383) );
  NAND4_X1 U6828 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n8961)
         );
  NOR2_X1 U6829 ( .A1(n8402), .A2(n8512), .ZN(n8680) );
  INV_X1 U6830 ( .A(n8680), .ZN(n5387) );
  OR2_X1 U6831 ( .A1(n5714), .A2(n8409), .ZN(n8270) );
  AND2_X1 U6832 ( .A1(n5387), .A2(n8270), .ZN(n5388) );
  NAND2_X1 U6833 ( .A1(n8271), .A2(n5388), .ZN(n5389) );
  NAND2_X1 U6834 ( .A1(n8402), .A2(n8512), .ZN(n8266) );
  NAND2_X1 U6835 ( .A1(n5389), .A2(n8266), .ZN(n8230) );
  NAND2_X1 U6836 ( .A1(n5390), .A2(SI_14_), .ZN(n5395) );
  INV_X1 U6837 ( .A(n5395), .ZN(n5392) );
  NAND2_X1 U6838 ( .A1(n5440), .A2(n5413), .ZN(n5397) );
  NAND2_X1 U6839 ( .A1(n5397), .A2(n5416), .ZN(n5399) );
  MUX2_X1 U6840 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6286), .Z(n5412) );
  XNOR2_X1 U6841 ( .A(n5412), .B(SI_15_), .ZN(n5398) );
  NAND2_X1 U6842 ( .A1(n6968), .A2(n5421), .ZN(n5403) );
  NAND2_X1 U6843 ( .A1(n5425), .A2(n5423), .ZN(n5400) );
  NAND2_X1 U6844 ( .A1(n5400), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U6845 ( .A(n5401), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9013) );
  AOI22_X1 U6846 ( .A1(n5539), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5470), .B2(
        n9013), .ZN(n5402) );
  NAND2_X1 U6847 ( .A1(n7420), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5411) );
  INV_X1 U6848 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6849 ( .A1(n5406), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6850 ( .A1(n5430), .A2(n5407), .ZN(n8514) );
  NAND2_X1 U6851 ( .A1(n5379), .A2(n8514), .ZN(n5410) );
  INV_X1 U6852 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8986) );
  OR2_X1 U6853 ( .A1(n5287), .A2(n8986), .ZN(n5409) );
  INV_X1 U6854 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8976) );
  OR2_X1 U6855 ( .A1(n5188), .A2(n8976), .ZN(n5408) );
  NAND4_X1 U6856 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n8960)
         );
  INV_X1 U6857 ( .A(n8960), .ZN(n8541) );
  INV_X1 U6858 ( .A(SI_15_), .ZN(n7762) );
  NAND2_X1 U6859 ( .A1(n5415), .A2(n7762), .ZN(n5414) );
  NAND2_X1 U6860 ( .A1(n5440), .A2(n5439), .ZN(n5418) );
  INV_X1 U6861 ( .A(n5414), .ZN(n5417) );
  AND2_X1 U6862 ( .A1(n5418), .A2(n5441), .ZN(n5420) );
  INV_X1 U6863 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6973) );
  INV_X1 U6864 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6975) );
  MUX2_X1 U6865 ( .A(n6973), .B(n6975), .S(n6286), .Z(n5437) );
  XNOR2_X1 U6866 ( .A(n5437), .B(SI_16_), .ZN(n5419) );
  NAND2_X1 U6867 ( .A1(n6972), .A2(n5421), .ZN(n5429) );
  NAND2_X1 U6868 ( .A1(n5423), .A2(n5422), .ZN(n5468) );
  NAND2_X1 U6869 ( .A1(n5468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6870 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  OR2_X1 U6871 ( .A1(n5426), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6872 ( .A1(n5426), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5427) );
  AND2_X1 U6873 ( .A1(n5449), .A2(n5427), .ZN(n9021) );
  AOI22_X1 U6874 ( .A1(n5539), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5470), .B2(
        n9021), .ZN(n5428) );
  NAND2_X1 U6875 ( .A1(n5430), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6876 ( .A1(n5455), .A2(n5431), .ZN(n8543) );
  NAND2_X1 U6877 ( .A1(n8543), .A2(n5379), .ZN(n5436) );
  NAND2_X1 U6878 ( .A1(n7420), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5435) );
  INV_X1 U6879 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5432) );
  OR2_X1 U6880 ( .A1(n5287), .A2(n5432), .ZN(n5434) );
  INV_X1 U6881 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8999) );
  OR2_X1 U6882 ( .A1(n5683), .A2(n8999), .ZN(n5433) );
  NAND4_X1 U6883 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), .ZN(n8959)
         );
  INV_X1 U6884 ( .A(n8959), .ZN(n8895) );
  OR2_X1 U6885 ( .A1(n9274), .A2(n8895), .ZN(n8692) );
  NAND2_X1 U6886 ( .A1(n9274), .A2(n8895), .ZN(n8695) );
  NAND2_X1 U6887 ( .A1(n8692), .A2(n8695), .ZN(n8336) );
  INV_X1 U6888 ( .A(n5442), .ZN(n5438) );
  INV_X1 U6889 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7108) );
  INV_X1 U6890 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5445) );
  MUX2_X1 U6891 ( .A(n7108), .B(n5445), .S(n6286), .Z(n5446) );
  INV_X1 U6892 ( .A(SI_17_), .ZN(n7866) );
  NAND2_X1 U6893 ( .A1(n5446), .A2(n7866), .ZN(n5460) );
  INV_X1 U6894 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6895 ( .A1(n5447), .A2(SI_17_), .ZN(n5448) );
  NAND2_X1 U6896 ( .A1(n5460), .A2(n5448), .ZN(n5461) );
  XNOR2_X1 U6897 ( .A(n5462), .B(n5461), .ZN(n7063) );
  NAND2_X1 U6898 ( .A1(n7063), .A2(n5421), .ZN(n5452) );
  NAND2_X1 U6899 ( .A1(n5449), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5450) );
  XNOR2_X1 U6900 ( .A(n5450), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9067) );
  AOI22_X1 U6901 ( .A1(n5539), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5470), .B2(
        n9067), .ZN(n5451) );
  INV_X1 U6902 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6903 ( .A1(n5455), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6904 ( .A1(n5473), .A2(n5456), .ZN(n8897) );
  NAND2_X1 U6905 ( .A1(n8897), .A2(n5379), .ZN(n5459) );
  AOI22_X1 U6906 ( .A1(n7420), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n5636), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5458) );
  INV_X1 U6907 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9027) );
  OR2_X1 U6908 ( .A1(n5188), .A2(n9027), .ZN(n5457) );
  NAND2_X1 U6909 ( .A1(n8889), .A2(n8815), .ZN(n8688) );
  MUX2_X1 U6910 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6286), .Z(n5478) );
  INV_X1 U6911 ( .A(SI_18_), .ZN(n5463) );
  XNOR2_X1 U6912 ( .A(n5478), .B(n5463), .ZN(n5477) );
  XNOR2_X1 U6913 ( .A(n5481), .B(n5477), .ZN(n7123) );
  NAND2_X1 U6914 ( .A1(n7123), .A2(n5421), .ZN(n5472) );
  INV_X1 U6915 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6916 ( .A1(n5466), .A2(n5465), .ZN(n5467) );
  NAND2_X1 U6917 ( .A1(n5485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5469) );
  XNOR2_X1 U6918 ( .A(n5469), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9063) );
  AOI22_X1 U6919 ( .A1(n5539), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5470), .B2(
        n9063), .ZN(n5471) );
  INV_X1 U6920 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U6921 ( .A1(n5473), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6922 ( .A1(n5493), .A2(n5474), .ZN(n8936) );
  NAND2_X1 U6923 ( .A1(n8936), .A2(n5379), .ZN(n5476) );
  AOI22_X1 U6924 ( .A1(n7420), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n5636), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n5475) );
  OAI211_X1 U6925 ( .C1(n5683), .C2(n8477), .A(n5476), .B(n5475), .ZN(n8957)
         );
  INV_X1 U6926 ( .A(n8957), .ZN(n9218) );
  OR2_X1 U6927 ( .A1(n8924), .A2(n9218), .ZN(n8699) );
  AOI21_X1 U6928 ( .B1(n8469), .B2(n8785), .A(n8690), .ZN(n9214) );
  INV_X1 U6929 ( .A(n5477), .ZN(n5480) );
  NAND2_X1 U6930 ( .A1(n5478), .A2(SI_18_), .ZN(n5479) );
  INV_X1 U6931 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7285) );
  INV_X1 U6932 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8848) );
  MUX2_X1 U6933 ( .A(n7285), .B(n8848), .S(n6286), .Z(n5482) );
  NAND2_X1 U6934 ( .A1(n5482), .A2(n7902), .ZN(n5503) );
  INV_X1 U6935 ( .A(n5482), .ZN(n5483) );
  NAND2_X1 U6936 ( .A1(n5483), .A2(SI_19_), .ZN(n5484) );
  NAND2_X1 U6937 ( .A1(n5503), .A2(n5484), .ZN(n5502) );
  XNOR2_X1 U6938 ( .A(n5501), .B(n5502), .ZN(n7284) );
  NAND2_X1 U6939 ( .A1(n7284), .A2(n5421), .ZN(n5490) );
  INV_X1 U6940 ( .A(n5485), .ZN(n5487) );
  INV_X1 U6941 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6942 ( .A1(n5672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5488) );
  XNOR2_X1 U6943 ( .A(n5488), .B(n5040), .ZN(n9093) );
  INV_X1 U6944 ( .A(n9093), .ZN(n9079) );
  AOI22_X1 U6945 ( .A1(n5539), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9079), .B2(
        n5470), .ZN(n5489) );
  INV_X1 U6946 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6947 ( .A1(n5493), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6948 ( .A1(n5521), .A2(n5494), .ZN(n9224) );
  NAND2_X1 U6949 ( .A1(n9224), .A2(n5379), .ZN(n5499) );
  INV_X1 U6950 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U6951 ( .A1(n7420), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6952 ( .A1(n4657), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5495) );
  OAI211_X1 U6953 ( .C1(n5287), .C2(n9223), .A(n5496), .B(n5495), .ZN(n5497)
         );
  INV_X1 U6954 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U6955 ( .A1(n5499), .A2(n5498), .ZN(n9203) );
  INV_X1 U6956 ( .A(n9203), .ZN(n8934) );
  NAND2_X1 U6957 ( .A1(n9339), .A2(n8934), .ZN(n8706) );
  NAND2_X1 U6958 ( .A1(n9214), .A2(n8706), .ZN(n5500) );
  NAND2_X1 U6959 ( .A1(n5500), .A2(n8707), .ZN(n9197) );
  MUX2_X1 U6960 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6286), .Z(n5511) );
  INV_X1 U6961 ( .A(SI_20_), .ZN(n5513) );
  XNOR2_X1 U6962 ( .A(n5511), .B(n5513), .ZN(n5504) );
  XNOR2_X1 U6963 ( .A(n5514), .B(n5504), .ZN(n7338) );
  NAND2_X1 U6964 ( .A1(n7338), .A2(n5421), .ZN(n5506) );
  NAND2_X1 U6965 ( .A1(n5539), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5505) );
  XNOR2_X1 U6966 ( .A(n5521), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n9207) );
  INV_X1 U6967 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U6968 ( .A1(n7420), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U6969 ( .A1(n5636), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5507) );
  OAI211_X1 U6970 ( .C1(n5509), .C2(n5683), .A(n5508), .B(n5507), .ZN(n5510)
         );
  AOI21_X1 U6971 ( .B1(n9207), .B2(n5379), .A(n5510), .ZN(n9219) );
  NAND2_X1 U6972 ( .A1(n9334), .A2(n9219), .ZN(n8710) );
  INV_X1 U6973 ( .A(n5511), .ZN(n5512) );
  MUX2_X1 U6974 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6286), .Z(n5532) );
  INV_X1 U6975 ( .A(SI_21_), .ZN(n5517) );
  XNOR2_X1 U6976 ( .A(n5532), .B(n5517), .ZN(n5518) );
  XNOR2_X1 U6977 ( .A(n5534), .B(n5518), .ZN(n7390) );
  NAND2_X1 U6978 ( .A1(n7390), .A2(n5421), .ZN(n5520) );
  NAND2_X1 U6979 ( .A1(n5539), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5519) );
  INV_X1 U6980 ( .A(n5521), .ZN(n5522) );
  INV_X1 U6981 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7923) );
  INV_X1 U6982 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5523) );
  INV_X1 U6983 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U6984 ( .A1(n5525), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6985 ( .A1(n5542), .A2(n5526), .ZN(n9192) );
  NAND2_X1 U6986 ( .A1(n9192), .A2(n5379), .ZN(n5531) );
  INV_X1 U6987 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U6988 ( .A1(n7420), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U6989 ( .A1(n5636), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5527) );
  OAI211_X1 U6990 ( .C1(n9261), .C2(n5188), .A(n5528), .B(n5527), .ZN(n5529)
         );
  INV_X1 U6991 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U6992 ( .A1(n5531), .A2(n5530), .ZN(n9204) );
  INV_X1 U6993 ( .A(n9204), .ZN(n8825) );
  NAND2_X1 U6994 ( .A1(n9191), .A2(n8825), .ZN(n5725) );
  INV_X1 U6995 ( .A(n5725), .ZN(n8717) );
  NAND2_X1 U6996 ( .A1(n5532), .A2(SI_21_), .ZN(n5533) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7983) );
  INV_X1 U6998 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7987) );
  MUX2_X1 U6999 ( .A(n7983), .B(n7987), .S(n6286), .Z(n5536) );
  INV_X1 U7000 ( .A(SI_22_), .ZN(n5535) );
  NAND2_X1 U7001 ( .A1(n5536), .A2(n5535), .ZN(n5552) );
  INV_X1 U7002 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7003 ( .A1(n5537), .A2(SI_22_), .ZN(n5538) );
  NAND2_X1 U7004 ( .A1(n5552), .A2(n5538), .ZN(n5551) );
  XNOR2_X1 U7005 ( .A(n5550), .B(n5551), .ZN(n7982) );
  NAND2_X1 U7006 ( .A1(n7982), .A2(n5421), .ZN(n5541) );
  NAND2_X1 U7007 ( .A1(n5539), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5540) );
  OR2_X2 U7008 ( .A1(n5542), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7009 ( .A1(n5542), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7010 ( .A1(n5559), .A2(n5543), .ZN(n9182) );
  NAND2_X1 U7011 ( .A1(n9182), .A2(n5379), .ZN(n5548) );
  INV_X1 U7012 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U7013 ( .A1(n7420), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7014 ( .A1(n5636), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U7015 ( .C1(n9256), .C2(n5683), .A(n5545), .B(n5544), .ZN(n5546)
         );
  INV_X1 U7016 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7017 ( .A1(n5548), .A2(n5547), .ZN(n9168) );
  NAND2_X1 U7018 ( .A1(n9324), .A2(n9188), .ZN(n8719) );
  INV_X1 U7019 ( .A(n8718), .ZN(n5549) );
  AOI21_X1 U7020 ( .B1(n9176), .B2(n8719), .A(n5549), .ZN(n9164) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5553) );
  INV_X1 U7022 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8068) );
  MUX2_X1 U7023 ( .A(n5553), .B(n8068), .S(n6286), .Z(n5554) );
  NAND2_X1 U7024 ( .A1(n5554), .A2(n7868), .ZN(n5568) );
  INV_X1 U7025 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7026 ( .A1(n5555), .A2(SI_23_), .ZN(n5556) );
  AND2_X1 U7027 ( .A1(n5568), .A2(n5556), .ZN(n5566) );
  NAND2_X1 U7028 ( .A1(n8065), .A2(n5421), .ZN(n5558) );
  NAND2_X1 U7029 ( .A1(n5539), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7030 ( .A1(n5559), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7031 ( .A1(n5577), .A2(n5560), .ZN(n9171) );
  NAND2_X1 U7032 ( .A1(n9171), .A2(n5379), .ZN(n5565) );
  INV_X1 U7033 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U7034 ( .A1(n5636), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7035 ( .A1(n7420), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5561) );
  OAI211_X1 U7036 ( .C1(n5683), .C2(n9252), .A(n5562), .B(n5561), .ZN(n5563)
         );
  INV_X1 U7037 ( .A(n5563), .ZN(n5564) );
  NAND2_X1 U7038 ( .A1(n5565), .A2(n5564), .ZN(n9179) );
  NAND2_X1 U7039 ( .A1(n9164), .A2(n8764), .ZN(n9159) );
  INV_X1 U7040 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8179) );
  INV_X1 U7041 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8177) );
  MUX2_X1 U7042 ( .A(n8179), .B(n8177), .S(n6286), .Z(n5570) );
  NAND2_X1 U7043 ( .A1(n5570), .A2(n7889), .ZN(n5587) );
  INV_X1 U7044 ( .A(n5570), .ZN(n5571) );
  NAND2_X1 U7045 ( .A1(n5571), .A2(SI_24_), .ZN(n5572) );
  AND2_X1 U7046 ( .A1(n5587), .A2(n5572), .ZN(n5585) );
  XNOR2_X1 U7047 ( .A(n5586), .B(n5585), .ZN(n8176) );
  NAND2_X1 U7048 ( .A1(n8176), .A2(n5421), .ZN(n5574) );
  NAND2_X1 U7049 ( .A1(n5539), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5573) );
  INV_X1 U7050 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7051 ( .A1(n5577), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7052 ( .A1(n5597), .A2(n5578), .ZN(n9157) );
  NAND2_X1 U7053 ( .A1(n9157), .A2(n5379), .ZN(n5583) );
  INV_X1 U7054 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U7055 ( .A1(n7420), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7056 ( .A1(n5636), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5579) );
  OAI211_X1 U7057 ( .C1(n9249), .C2(n5188), .A(n5580), .B(n5579), .ZN(n5581)
         );
  INV_X1 U7058 ( .A(n5581), .ZN(n5582) );
  NAND2_X1 U7059 ( .A1(n5583), .A2(n5582), .ZN(n9167) );
  NAND2_X1 U7060 ( .A1(n9311), .A2(n9142), .ZN(n8762) );
  NAND2_X1 U7061 ( .A1(n9317), .A2(n8919), .ZN(n9158) );
  NAND2_X1 U7062 ( .A1(n9159), .A2(n8723), .ZN(n5584) );
  NAND2_X1 U7063 ( .A1(n5584), .A2(n8763), .ZN(n9146) );
  INV_X1 U7064 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5588) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8214) );
  MUX2_X1 U7066 ( .A(n5588), .B(n8214), .S(n6286), .Z(n5590) );
  INV_X1 U7067 ( .A(SI_25_), .ZN(n5589) );
  NAND2_X1 U7068 ( .A1(n5590), .A2(n5589), .ZN(n5606) );
  INV_X1 U7069 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U7070 ( .A1(n5591), .A2(SI_25_), .ZN(n5592) );
  AND2_X1 U7071 ( .A1(n5606), .A2(n5592), .ZN(n5604) );
  XNOR2_X1 U7072 ( .A(n5605), .B(n5604), .ZN(n8191) );
  NAND2_X1 U7073 ( .A1(n8191), .A2(n5421), .ZN(n5594) );
  NAND2_X1 U7074 ( .A1(n5539), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5593) );
  INV_X1 U7075 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7076 ( .A1(n5597), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7077 ( .A1(n5614), .A2(n5598), .ZN(n9145) );
  NAND2_X1 U7078 ( .A1(n9145), .A2(n5379), .ZN(n5603) );
  INV_X1 U7079 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U7080 ( .A1(n5636), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7081 ( .A1(n7420), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5599) );
  OAI211_X1 U7082 ( .C1(n9246), .C2(n5683), .A(n5600), .B(n5599), .ZN(n5601)
         );
  INV_X1 U7083 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7084 ( .A1(n9305), .A2(n8949), .ZN(n8732) );
  INV_X1 U7085 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5607) );
  INV_X1 U7086 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8301) );
  MUX2_X1 U7087 ( .A(n5607), .B(n8301), .S(n6738), .Z(n5609) );
  INV_X1 U7088 ( .A(SI_26_), .ZN(n5608) );
  NAND2_X1 U7089 ( .A1(n5609), .A2(n5608), .ZN(n5623) );
  INV_X1 U7090 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U7091 ( .A1(n5610), .A2(SI_26_), .ZN(n5611) );
  AND2_X1 U7092 ( .A1(n5623), .A2(n5611), .ZN(n5621) );
  NAND2_X1 U7093 ( .A1(n8242), .A2(n5421), .ZN(n5613) );
  NAND2_X1 U7094 ( .A1(n5539), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7095 ( .A1(n5614), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7096 ( .A1(n5634), .A2(n5615), .ZN(n9137) );
  NAND2_X1 U7097 ( .A1(n9137), .A2(n5379), .ZN(n5620) );
  INV_X1 U7098 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U7099 ( .A1(n5129), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7100 ( .A1(n5636), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5616) );
  OAI211_X1 U7101 ( .C1(n9242), .C2(n5188), .A(n5617), .B(n5616), .ZN(n5618)
         );
  INV_X1 U7102 ( .A(n5618), .ZN(n5619) );
  INV_X1 U7103 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5625) );
  INV_X1 U7104 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8359) );
  MUX2_X1 U7105 ( .A(n5625), .B(n8359), .S(n6286), .Z(n5627) );
  INV_X1 U7106 ( .A(SI_27_), .ZN(n5626) );
  NAND2_X1 U7107 ( .A1(n5627), .A2(n5626), .ZN(n5646) );
  INV_X1 U7108 ( .A(n5627), .ZN(n5628) );
  NAND2_X1 U7109 ( .A1(n5628), .A2(SI_27_), .ZN(n5629) );
  AND2_X1 U7110 ( .A1(n5646), .A2(n5629), .ZN(n5645) );
  NAND2_X1 U7111 ( .A1(n5539), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5630) );
  INV_X1 U7112 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7113 ( .A1(n5634), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7114 ( .A1(n5650), .A2(n5635), .ZN(n9127) );
  NAND2_X1 U7115 ( .A1(n9127), .A2(n5379), .ZN(n5641) );
  INV_X1 U7116 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U7117 ( .A1(n5636), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7118 ( .A1(n7420), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5637) );
  OAI211_X1 U7119 ( .C1(n9239), .C2(n5683), .A(n5638), .B(n5637), .ZN(n5639)
         );
  INV_X1 U7120 ( .A(n5639), .ZN(n5640) );
  INV_X1 U7121 ( .A(n9121), .ZN(n8789) );
  NAND2_X1 U7122 ( .A1(n9299), .A2(n9143), .ZN(n9118) );
  AND2_X1 U7123 ( .A1(n8789), .A2(n9118), .ZN(n5642) );
  MUX2_X1 U7124 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6286), .Z(n5661) );
  INV_X1 U7125 ( .A(SI_28_), .ZN(n7892) );
  XNOR2_X1 U7126 ( .A(n5661), .B(n7892), .ZN(n5659) );
  NAND2_X1 U7127 ( .A1(n8360), .A2(n5421), .ZN(n5649) );
  NAND2_X1 U7128 ( .A1(n5539), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7129 ( .A1(n5650), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7130 ( .A1(n8807), .A2(n5651), .ZN(n9113) );
  NAND2_X1 U7131 ( .A1(n9113), .A2(n5379), .ZN(n5656) );
  INV_X1 U7132 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U7133 ( .A1(n5636), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7134 ( .A1(n7420), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5652) );
  OAI211_X1 U7135 ( .C1(n9234), .C2(n5188), .A(n5653), .B(n5652), .ZN(n5654)
         );
  INV_X1 U7136 ( .A(n5654), .ZN(n5655) );
  NAND2_X1 U7137 ( .A1(n9103), .A2(n9104), .ZN(n5658) );
  INV_X1 U7138 ( .A(n9123), .ZN(n8746) );
  OR2_X1 U7139 ( .A1(n9114), .A2(n8746), .ZN(n5657) );
  INV_X1 U7140 ( .A(n5661), .ZN(n5662) );
  INV_X1 U7141 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5663) );
  INV_X1 U7142 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9951) );
  MUX2_X1 U7143 ( .A(n5663), .B(n9951), .S(n6286), .Z(n6273) );
  NAND2_X1 U7144 ( .A1(n5825), .A2(n5421), .ZN(n5665) );
  NAND2_X1 U7145 ( .A1(n5539), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5664) );
  INV_X1 U7146 ( .A(n8807), .ZN(n5666) );
  NAND2_X1 U7147 ( .A1(n5666), .A2(n5379), .ZN(n7426) );
  INV_X1 U7148 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7149 ( .A1(n5636), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7150 ( .A1(n5129), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5667) );
  OAI211_X1 U7151 ( .C1(n5188), .C2(n5784), .A(n5668), .B(n5667), .ZN(n5669)
         );
  INV_X1 U7152 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U7153 ( .A1(n7426), .A2(n5670), .ZN(n9107) );
  INV_X1 U7154 ( .A(n9107), .ZN(n5671) );
  NAND2_X1 U7155 ( .A1(n5783), .A2(n5671), .ZN(n8603) );
  NAND2_X1 U7156 ( .A1(n4554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5674) );
  XNOR2_X1 U7157 ( .A(n5674), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8801) );
  INV_X1 U7158 ( .A(n8801), .ZN(n7984) );
  NAND2_X1 U7159 ( .A1(n5790), .A2(n7984), .ZN(n10390) );
  XNOR2_X1 U7160 ( .A(n5676), .B(n5675), .ZN(n5740) );
  AOI21_X1 U7161 ( .B1(n8759), .B2(n7984), .A(n9079), .ZN(n5677) );
  AND2_X1 U7162 ( .A1(n10390), .A2(n5677), .ZN(n5679) );
  NAND2_X1 U7163 ( .A1(n5740), .A2(n9093), .ZN(n6944) );
  OR2_X1 U7164 ( .A1(n8748), .A2(n6944), .ZN(n6935) );
  NAND2_X1 U7165 ( .A1(n5679), .A2(n6935), .ZN(n10353) );
  INV_X1 U7166 ( .A(n5680), .ZN(n6872) );
  XNOR2_X1 U7167 ( .A(n6872), .B(n8799), .ZN(n6937) );
  OR2_X1 U7168 ( .A1(n8748), .A2(n6937), .ZN(n10348) );
  INV_X1 U7169 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7170 ( .A1(n7420), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7171 ( .A1(n5636), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5681) );
  OAI211_X1 U7172 ( .C1(n5684), .C2(n5683), .A(n5682), .B(n5681), .ZN(n5685)
         );
  INV_X1 U7173 ( .A(n5685), .ZN(n5686) );
  NAND2_X1 U7174 ( .A1(n7426), .A2(n5686), .ZN(n8955) );
  INV_X1 U7175 ( .A(n6937), .ZN(n6938) );
  AND2_X1 U7176 ( .A1(n6736), .A2(P2_B_REG_SCAN_IN), .ZN(n5687) );
  NOR2_X1 U7177 ( .A1(n10346), .A2(n5687), .ZN(n9096) );
  AOI22_X1 U7178 ( .A1(n10326), .A2(n9123), .B1(n8955), .B2(n9096), .ZN(n5738)
         );
  INV_X1 U7179 ( .A(n9334), .ZN(n9209) );
  AND2_X1 U7180 ( .A1(n10403), .A2(n8966), .ZN(n5704) );
  OR2_X1 U7181 ( .A1(n10403), .A2(n8966), .ZN(n5690) );
  INV_X1 U7182 ( .A(n6844), .ZN(n8973) );
  NAND2_X1 U7183 ( .A1(n8973), .A2(n8582), .ZN(n7154) );
  NAND2_X1 U7184 ( .A1(n8766), .A2(n7154), .ZN(n5694) );
  NAND2_X1 U7185 ( .A1(n5692), .A2(n10360), .ZN(n5693) );
  NAND2_X1 U7186 ( .A1(n5694), .A2(n5693), .ZN(n10345) );
  NAND2_X1 U7187 ( .A1(n10345), .A2(n10344), .ZN(n10324) );
  NAND2_X1 U7188 ( .A1(n7075), .A2(n10365), .ZN(n10323) );
  NAND2_X1 U7189 ( .A1(n10347), .A2(n10333), .ZN(n5695) );
  AND2_X1 U7190 ( .A1(n10323), .A2(n5695), .ZN(n5696) );
  NAND2_X1 U7191 ( .A1(n10324), .A2(n5696), .ZN(n7145) );
  NAND2_X1 U7192 ( .A1(n8971), .A2(n10369), .ZN(n7143) );
  NAND2_X1 U7193 ( .A1(n8970), .A2(n7246), .ZN(n5698) );
  NAND2_X1 U7194 ( .A1(n7145), .A2(n5697), .ZN(n5703) );
  INV_X1 U7195 ( .A(n5698), .ZN(n5701) );
  AOI21_X1 U7196 ( .B1(n7162), .B2(n10379), .A(n5699), .ZN(n5700) );
  OR2_X1 U7197 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  NAND2_X1 U7198 ( .A1(n5703), .A2(n5702), .ZN(n7255) );
  NOR2_X1 U7199 ( .A1(n7259), .A2(n8969), .ZN(n7250) );
  NAND2_X1 U7200 ( .A1(n7259), .A2(n8969), .ZN(n7249) );
  INV_X1 U7201 ( .A(n7429), .ZN(n7397) );
  NAND2_X1 U7202 ( .A1(n7397), .A2(n5705), .ZN(n5706) );
  NAND2_X1 U7203 ( .A1(n5707), .A2(n5706), .ZN(n7557) );
  NAND2_X1 U7204 ( .A1(n10412), .A2(n8965), .ZN(n5708) );
  NAND2_X1 U7205 ( .A1(n7557), .A2(n5708), .ZN(n7990) );
  OR2_X1 U7206 ( .A1(n10412), .A2(n8965), .ZN(n7989) );
  AND2_X1 U7207 ( .A1(n8164), .A2(n7989), .ZN(n5709) );
  NAND2_X1 U7208 ( .A1(n7990), .A2(n5709), .ZN(n7993) );
  INV_X1 U7209 ( .A(n8168), .ZN(n8964) );
  NAND2_X1 U7210 ( .A1(n10417), .A2(n8964), .ZN(n5710) );
  NAND2_X1 U7211 ( .A1(n7993), .A2(n5710), .ZN(n8090) );
  INV_X1 U7212 ( .A(n8668), .ZN(n8963) );
  OR2_X1 U7213 ( .A1(n8669), .A2(n8963), .ZN(n5711) );
  NAND2_X1 U7214 ( .A1(n8090), .A2(n5711), .ZN(n5713) );
  NAND2_X1 U7215 ( .A1(n8669), .A2(n8963), .ZN(n5712) );
  NAND2_X1 U7216 ( .A1(n5713), .A2(n5712), .ZN(n8184) );
  INV_X1 U7217 ( .A(n8184), .ZN(n5716) );
  NAND2_X1 U7218 ( .A1(n5714), .A2(n8962), .ZN(n8674) );
  INV_X1 U7219 ( .A(n8777), .ZN(n5715) );
  NAND2_X1 U7220 ( .A1(n8402), .A2(n8961), .ZN(n5717) );
  OR2_X1 U7221 ( .A1(n8402), .A2(n8961), .ZN(n5718) );
  NOR2_X1 U7222 ( .A1(n8508), .A2(n8960), .ZN(n5719) );
  NAND2_X1 U7223 ( .A1(n8508), .A2(n8960), .ZN(n5720) );
  NAND2_X1 U7224 ( .A1(n9274), .A2(n8959), .ZN(n5722) );
  NAND2_X1 U7225 ( .A1(n8468), .A2(n8688), .ZN(n8696) );
  INV_X1 U7226 ( .A(n8815), .ZN(n8958) );
  NAND2_X1 U7227 ( .A1(n8889), .A2(n8958), .ZN(n5723) );
  NAND2_X1 U7228 ( .A1(n5724), .A2(n5723), .ZN(n8471) );
  NAND2_X1 U7229 ( .A1(n8707), .A2(n8706), .ZN(n9216) );
  AOI21_X2 U7230 ( .B1(n9209), .B2(n9219), .A(n9202), .ZN(n9185) );
  NAND2_X1 U7231 ( .A1(n8718), .A2(n8719), .ZN(n9177) );
  INV_X1 U7232 ( .A(n9324), .ZN(n8923) );
  INV_X1 U7233 ( .A(n9152), .ZN(n5729) );
  INV_X1 U7234 ( .A(n9311), .ZN(n9151) );
  OAI21_X1 U7235 ( .B1(n9143), .B2(n4811), .A(n9133), .ZN(n5730) );
  INV_X1 U7236 ( .A(n9293), .ZN(n5731) );
  INV_X1 U7237 ( .A(n9114), .ZN(n9290) );
  XNOR2_X1 U7238 ( .A(n5734), .B(n5733), .ZN(n5736) );
  NAND2_X1 U7239 ( .A1(n5678), .A2(n8759), .ZN(n8607) );
  AND2_X1 U7240 ( .A1(n9079), .A2(n8801), .ZN(n5791) );
  INV_X1 U7241 ( .A(n5791), .ZN(n5735) );
  NAND2_X1 U7242 ( .A1(n5736), .A2(n10350), .ZN(n5737) );
  AND2_X1 U7243 ( .A1(n5740), .A2(n9079), .ZN(n7141) );
  INV_X1 U7244 ( .A(n10404), .ZN(n5741) );
  INV_X1 U7245 ( .A(n6944), .ZN(n5743) );
  OR2_X1 U7246 ( .A1(n8748), .A2(n5743), .ZN(n6922) );
  INV_X1 U7247 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7248 ( .A1(n5757), .A2(n5758), .ZN(n5745) );
  INV_X1 U7249 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7250 ( .A1(n5753), .A2(n5752), .ZN(n5755) );
  INV_X1 U7251 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5746) );
  INV_X1 U7252 ( .A(n6759), .ZN(n8192) );
  NAND2_X1 U7253 ( .A1(n5748), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5749) );
  MUX2_X1 U7254 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5749), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5750) );
  INV_X1 U7255 ( .A(n8243), .ZN(n5773) );
  OR2_X1 U7256 ( .A1(n5753), .A2(n5752), .ZN(n5754) );
  NOR2_X1 U7257 ( .A1(n5773), .A2(n8181), .ZN(n5756) );
  NAND2_X1 U7258 ( .A1(n8192), .A2(n5756), .ZN(n6921) );
  XNOR2_X1 U7259 ( .A(n5757), .B(n5758), .ZN(n6920) );
  AND2_X1 U7260 ( .A1(n6920), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6764) );
  NAND2_X1 U7261 ( .A1(n6921), .A2(n6764), .ZN(n6932) );
  INV_X1 U7262 ( .A(n6932), .ZN(n6757) );
  XNOR2_X1 U7263 ( .A(n8181), .B(P2_B_REG_SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7264 ( .A1(n6759), .A2(n5759), .ZN(n5760) );
  NOR2_X1 U7265 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5764) );
  NOR4_X1 U7266 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5763) );
  NOR4_X1 U7267 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5762) );
  NOR4_X1 U7268 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5761) );
  NAND4_X1 U7269 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n5770)
         );
  NOR4_X1 U7270 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5768) );
  NOR4_X1 U7271 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5767) );
  NOR4_X1 U7272 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5766) );
  NOR4_X1 U7273 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5765) );
  NAND4_X1 U7274 ( .A1(n5768), .A2(n5767), .A3(n5766), .A4(n5765), .ZN(n5769)
         );
  NOR2_X1 U7275 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  OR2_X1 U7276 ( .A1(n5772), .A2(n5771), .ZN(n5796) );
  AND2_X1 U7277 ( .A1(n6757), .A2(n5796), .ZN(n5776) );
  NAND2_X1 U7278 ( .A1(n5773), .A2(n8181), .ZN(n6762) );
  OR2_X1 U7279 ( .A1(n5772), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7280 ( .A1(n6759), .A2(n5773), .ZN(n5774) );
  NAND2_X1 U7281 ( .A1(n5775), .A2(n5774), .ZN(n7093) );
  OR2_X1 U7282 ( .A1(n6941), .A2(n7093), .ZN(n5787) );
  AND3_X1 U7283 ( .A1(n6922), .A2(n5776), .A3(n5787), .ZN(n7095) );
  NAND2_X1 U7284 ( .A1(n10404), .A2(n5790), .ZN(n6933) );
  INV_X1 U7285 ( .A(n6941), .ZN(n7097) );
  NAND2_X1 U7286 ( .A1(n6933), .A2(n7097), .ZN(n5779) );
  NAND2_X1 U7287 ( .A1(n9093), .A2(n8801), .ZN(n5777) );
  OR2_X1 U7288 ( .A1(n5777), .A2(n5740), .ZN(n5778) );
  NAND2_X1 U7289 ( .A1(n5779), .A2(n7096), .ZN(n5782) );
  INV_X1 U7290 ( .A(n7096), .ZN(n5780) );
  NAND2_X1 U7291 ( .A1(n5780), .A2(n7093), .ZN(n5781) );
  AND3_X2 U7292 ( .A1(n7095), .A2(n5782), .A3(n5781), .ZN(n10440) );
  INV_X1 U7293 ( .A(n10390), .ZN(n10416) );
  NAND2_X1 U7294 ( .A1(n10440), .A2(n10416), .ZN(n9263) );
  OAI21_X1 U7295 ( .B1(n5802), .B2(n10437), .A(n5786), .ZN(P2_U3488) );
  INV_X1 U7296 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7297 ( .A1(n5788), .A2(n5796), .ZN(n6924) );
  INV_X1 U7298 ( .A(n6924), .ZN(n5789) );
  NAND2_X1 U7299 ( .A1(n5789), .A2(n6757), .ZN(n6957) );
  INV_X1 U7300 ( .A(n6935), .ZN(n7099) );
  INV_X1 U7301 ( .A(n6942), .ZN(n5792) );
  NOR2_X1 U7302 ( .A1(n7099), .A2(n6958), .ZN(n5793) );
  OR2_X1 U7303 ( .A1(n6957), .A2(n5793), .ZN(n5798) );
  AND2_X1 U7304 ( .A1(n8748), .A2(n10390), .ZN(n5795) );
  INV_X1 U7305 ( .A(n6958), .ZN(n5794) );
  NAND2_X1 U7306 ( .A1(n5795), .A2(n5794), .ZN(n6956) );
  OR2_X1 U7307 ( .A1(n10390), .A2(n7141), .ZN(n10341) );
  NAND2_X1 U7308 ( .A1(n6956), .A2(n10341), .ZN(n6925) );
  NAND3_X1 U7309 ( .A1(n6941), .A2(n7093), .A3(n5796), .ZN(n6928) );
  OR2_X1 U7310 ( .A1(n6928), .A2(n6932), .ZN(n6936) );
  INV_X1 U7311 ( .A(n6936), .ZN(n6959) );
  NAND2_X1 U7312 ( .A1(n6925), .A2(n6959), .ZN(n5797) );
  INV_X2 U7313 ( .A(n10423), .ZN(n10421) );
  NAND2_X1 U7314 ( .A1(n10421), .A2(n10416), .ZN(n9331) );
  INV_X1 U7315 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5799) );
  OAI21_X1 U7316 ( .B1(n5802), .B2(n10423), .A(n5801), .ZN(P2_U3456) );
  NOR2_X1 U7317 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5897) );
  NOR2_X1 U7318 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5808) );
  NOR2_X1 U7319 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5807) );
  INV_X1 U7320 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5806) );
  AND4_X1 U7321 ( .A1(n5897), .A2(n5808), .A3(n5807), .A4(n5806), .ZN(n5809)
         );
  INV_X1 U7322 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7776) );
  INV_X1 U7323 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6152) );
  NAND4_X1 U7324 ( .A1(n5868), .A2(n4746), .A3(n7776), .A4(n6152), .ZN(n5810)
         );
  OAI21_X1 U7325 ( .B1(n5819), .B2(n5815), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n5818) );
  INV_X1 U7326 ( .A(n5829), .ZN(n5820) );
  MUX2_X1 U7327 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5822), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5824) );
  INV_X1 U7328 ( .A(n5819), .ZN(n5823) );
  NAND2_X1 U7329 ( .A1(n5967), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5826) );
  INV_X1 U7330 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5827) );
  XNOR2_X2 U7331 ( .A(n5828), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9944) );
  OAI21_X1 U7332 ( .B1(n5829), .B2(n5815), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5831) );
  AND2_X2 U7333 ( .A1(n9944), .A2(n9950), .ZN(n6181) );
  NAND2_X1 U7334 ( .A1(n6224), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5841) );
  INV_X1 U7335 ( .A(n9944), .ZN(n5837) );
  INV_X2 U7336 ( .A(n5949), .ZN(n6215) );
  NAND2_X1 U7337 ( .A1(n6215), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5840) );
  AND2_X2 U7338 ( .A1(n9944), .A2(n5834), .ZN(n6144) );
  NAND2_X1 U7339 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6007) );
  NAND2_X1 U7340 ( .A1(n6005), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6041) );
  INV_X1 U7341 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6051) );
  INV_X1 U7342 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U7343 ( .A1(n6074), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6102) );
  INV_X1 U7344 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8426) );
  INV_X1 U7345 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7346 ( .A1(n5906), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5908) );
  INV_X1 U7347 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5888) );
  INV_X1 U7348 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U7349 ( .A1(n5921), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6142) );
  INV_X1 U7350 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7351 ( .A1(n6158), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6168) );
  INV_X1 U7352 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9368) );
  INV_X1 U7353 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U7354 ( .A1(n6194), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6217) );
  INV_X1 U7355 ( .A(n6217), .ZN(n5835) );
  NAND2_X1 U7356 ( .A1(n5835), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7357 ( .A1(n6216), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6239) );
  INV_X1 U7358 ( .A(n6239), .ZN(n6225) );
  NAND2_X1 U7359 ( .A1(n6225), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6252) );
  INV_X1 U7360 ( .A(n6252), .ZN(n6238) );
  NAND2_X1 U7361 ( .A1(n6238), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5859) );
  INV_X1 U7362 ( .A(n5859), .ZN(n6251) );
  NAND2_X1 U7363 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6251), .ZN(n5861) );
  INV_X1 U7364 ( .A(n5861), .ZN(n5836) );
  NAND2_X1 U7365 ( .A1(n5836), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5852) );
  INV_X1 U7366 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6720) );
  NOR2_X1 U7367 ( .A1(n5852), .A2(n6720), .ZN(n9692) );
  NAND2_X1 U7368 ( .A1(n6144), .A2(n9692), .ZN(n5839) );
  AND2_X2 U7369 ( .A1(n5837), .A2(n9950), .ZN(n6043) );
  NAND2_X1 U7370 ( .A1(n6228), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7371 ( .A1(n9861), .A2(n7234), .ZN(n6366) );
  NAND2_X1 U7372 ( .A1(n8360), .A2(n6191), .ZN(n5843) );
  NAND2_X1 U7373 ( .A1(n5967), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7374 ( .A1(n6224), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7375 ( .A1(n6228), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U7376 ( .A(n5852), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U7377 ( .A1(n6227), .A2(n9709), .ZN(n5845) );
  NAND2_X1 U7378 ( .A1(n6215), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7379 ( .A1(n9870), .A2(n9721), .ZN(n9683) );
  NAND2_X1 U7380 ( .A1(n8321), .A2(n6191), .ZN(n5849) );
  NAND2_X1 U7381 ( .A1(n5967), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7382 ( .A1(n6224), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7383 ( .A1(n6228), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5855) );
  INV_X1 U7384 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7385 ( .A1(n5861), .A2(n5850), .ZN(n5851) );
  NAND2_X1 U7386 ( .A1(n6144), .A2(n9723), .ZN(n5854) );
  NAND2_X1 U7387 ( .A1(n6215), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7388 ( .A1(n9874), .A2(n9732), .ZN(n9680) );
  AND2_X1 U7389 ( .A1(n9683), .A2(n9680), .ZN(n6364) );
  NAND2_X1 U7390 ( .A1(n8242), .A2(n6191), .ZN(n5858) );
  NAND2_X1 U7391 ( .A1(n6062), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7392 ( .A1(n6224), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7393 ( .A1(n6215), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5865) );
  INV_X1 U7394 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7395 ( .A1(n5860), .A2(n5859), .ZN(n5862) );
  AND2_X1 U7396 ( .A1(n5862), .A2(n5861), .ZN(n9736) );
  NAND2_X1 U7397 ( .A1(n6227), .A2(n9736), .ZN(n5864) );
  NAND2_X1 U7398 ( .A1(n6228), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5863) );
  INV_X1 U7399 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7748) );
  INV_X1 U7400 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U7401 ( .A1(n5869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7402 ( .A1(n5879), .A2(n5870), .ZN(n6138) );
  NAND2_X1 U7403 ( .A1(n4571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7404 ( .A1(n6299), .A2(n6298), .ZN(n5872) );
  NAND2_X1 U7405 ( .A1(n5872), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7406 ( .A1(n5874), .A2(n5873), .ZN(n6445) );
  OR2_X1 U7407 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  NAND2_X1 U7408 ( .A1(n6445), .A2(n5875), .ZN(n7985) );
  OAI21_X1 U7409 ( .B1(n6351), .B2(n9858), .A(n6352), .ZN(n6261) );
  INV_X1 U7410 ( .A(n6329), .ZN(n9682) );
  NAND2_X1 U7411 ( .A1(n6972), .A2(n6191), .ZN(n5878) );
  INV_X1 U7412 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U7413 ( .A1(n5879), .A2(n7753), .ZN(n5881) );
  NAND2_X1 U7414 ( .A1(n5881), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U7415 ( .A(n5876), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9589) );
  AOI22_X1 U7416 ( .A1(n6062), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6165), .B2(
        n9589), .ZN(n5877) );
  NAND2_X1 U7417 ( .A1(n6968), .A2(n6191), .ZN(n5883) );
  OR2_X1 U7418 ( .A1(n5879), .A2(n7753), .ZN(n5880) );
  AND2_X1 U7419 ( .A1(n5881), .A2(n5880), .ZN(n9568) );
  AOI22_X1 U7420 ( .A1(n6062), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6165), .B2(
        n9568), .ZN(n5882) );
  NAND2_X1 U7421 ( .A1(n6181), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7422 ( .A1(n6228), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7423 ( .A1(n6215), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5885) );
  AOI21_X1 U7424 ( .B1(n5890), .B2(n9561), .A(n5921), .ZN(n9484) );
  NAND2_X1 U7425 ( .A1(n6144), .A2(n9484), .ZN(n5884) );
  NAND4_X1 U7426 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n9501)
         );
  NAND2_X1 U7427 ( .A1(n9916), .A2(n9395), .ZN(n6416) );
  NAND2_X1 U7428 ( .A1(n6215), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7429 ( .A1(n6224), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7430 ( .A1(n5908), .A2(n5888), .ZN(n5889) );
  AND2_X1 U7431 ( .A1(n5890), .A2(n5889), .ZN(n8394) );
  NAND2_X1 U7432 ( .A1(n6227), .A2(n8394), .ZN(n5892) );
  NAND2_X1 U7433 ( .A1(n6228), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5891) );
  NAND4_X1 U7434 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n9502)
         );
  NAND2_X1 U7435 ( .A1(n6848), .A2(n6191), .ZN(n5905) );
  INV_X1 U7436 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5896) );
  AND2_X1 U7437 ( .A1(n5895), .A2(n5896), .ZN(n6058) );
  AND2_X1 U7438 ( .A1(n6058), .A2(n5897), .ZN(n6083) );
  INV_X1 U7439 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7440 ( .A1(n6083), .A2(n5898), .ZN(n6098) );
  INV_X1 U7441 ( .A(n6098), .ZN(n5900) );
  INV_X1 U7442 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5899) );
  AOI21_X1 U7443 ( .B1(n5900), .B2(n5899), .A(n5815), .ZN(n6108) );
  INV_X1 U7444 ( .A(n6108), .ZN(n5902) );
  INV_X1 U7445 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7446 ( .A1(n5902), .A2(n5901), .ZN(n6109) );
  NAND2_X1 U7447 ( .A1(n6109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5903) );
  XNOR2_X1 U7448 ( .A(n5903), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8258) );
  AOI22_X1 U7449 ( .A1(n6062), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6165), .B2(
        n8258), .ZN(n5904) );
  NAND2_X2 U7450 ( .A1(n5905), .A2(n5904), .ZN(n8528) );
  NAND2_X1 U7451 ( .A1(n6215), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7452 ( .A1(n6224), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5911) );
  INV_X1 U7453 ( .A(n5906), .ZN(n6116) );
  INV_X1 U7454 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U7455 ( .A1(n6116), .A2(n8524), .ZN(n5907) );
  AND2_X1 U7456 ( .A1(n5908), .A2(n5907), .ZN(n8313) );
  NAND2_X1 U7457 ( .A1(n6144), .A2(n8313), .ZN(n5910) );
  NAND2_X1 U7458 ( .A1(n6228), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5909) );
  AND2_X1 U7459 ( .A1(n8288), .A2(n5984), .ZN(n5926) );
  NAND2_X1 U7460 ( .A1(n8528), .A2(n5926), .ZN(n5913) );
  OAI21_X1 U7461 ( .B1(n9858), .B2(n9502), .A(n5913), .ZN(n5920) );
  NAND2_X1 U7462 ( .A1(n6965), .A2(n6191), .ZN(n5919) );
  NOR2_X1 U7463 ( .A1(n5867), .A2(n5815), .ZN(n5914) );
  MUX2_X1 U7464 ( .A(n5815), .B(n5914), .S(P1_IR_REG_14__SCAN_IN), .Z(n5915)
         );
  INV_X1 U7465 ( .A(n5915), .ZN(n5917) );
  AND2_X1 U7466 ( .A1(n5917), .A2(n5916), .ZN(n9553) );
  AOI22_X1 U7467 ( .A1(n6062), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6165), .B2(
        n9553), .ZN(n5918) );
  NAND2_X1 U7468 ( .A1(n5920), .A2(n9920), .ZN(n5928) );
  NAND2_X1 U7469 ( .A1(n6224), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7470 ( .A1(n6215), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7471 ( .A1(n6228), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5923) );
  OAI21_X1 U7472 ( .B1(n5921), .B2(P1_REG3_REG_16__SCAN_IN), .A(n6142), .ZN(
        n9394) );
  INV_X1 U7473 ( .A(n9394), .ZN(n8495) );
  NAND2_X1 U7474 ( .A1(n6227), .A2(n8495), .ZN(n5922) );
  AND2_X1 U7475 ( .A1(n9486), .A2(n5984), .ZN(n5938) );
  INV_X1 U7476 ( .A(n5938), .ZN(n5931) );
  NAND3_X1 U7477 ( .A1(n8528), .A2(n9489), .A3(n5926), .ZN(n5927) );
  NAND4_X1 U7478 ( .A1(n6416), .A2(n5928), .A3(n5931), .A4(n5927), .ZN(n6125)
         );
  OR3_X1 U7479 ( .A1(n9398), .A2(n9486), .A3(n5984), .ZN(n5941) );
  INV_X1 U7480 ( .A(n9920), .ZN(n8324) );
  OR2_X1 U7481 ( .A1(n8288), .A2(n5984), .ZN(n5933) );
  OAI22_X1 U7482 ( .A1(n8528), .A2(n5933), .B1(n9489), .B2(n5984), .ZN(n5929)
         );
  NAND2_X1 U7483 ( .A1(n8324), .A2(n5929), .ZN(n5937) );
  NAND3_X1 U7484 ( .A1(n8528), .A2(n8288), .A3(n5938), .ZN(n5930) );
  OAI21_X1 U7485 ( .B1(n5931), .B2(n9502), .A(n5930), .ZN(n5932) );
  NAND2_X1 U7486 ( .A1(n5932), .A2(n9920), .ZN(n5936) );
  NAND4_X1 U7487 ( .A1(n8528), .A2(n9489), .A3(n8288), .A4(n5938), .ZN(n5935)
         );
  OR3_X1 U7488 ( .A1(n8528), .A2(n9489), .A3(n5933), .ZN(n5934) );
  AND4_X1 U7489 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(n5940)
         );
  OR2_X1 U7490 ( .A1(n9916), .A2(n9395), .ZN(n6417) );
  NAND3_X1 U7491 ( .A1(n9916), .A2(n9395), .A3(n5938), .ZN(n5939) );
  INV_X1 U7492 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U7493 ( .A1(n6144), .A2(n9514), .ZN(n5945) );
  NAND2_X1 U7494 ( .A1(n6215), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7495 ( .A1(n6043), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7496 ( .A1(n6181), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5942) );
  AND4_X2 U7497 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n8576)
         );
  INV_X2 U7498 ( .A(n8576), .ZN(n9512) );
  NAND2_X1 U7499 ( .A1(n5967), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7500 ( .A1(n7935), .A2(n5954), .ZN(n5957) );
  NAND2_X1 U7501 ( .A1(n5957), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U7502 ( .A(n5946), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U7503 ( .A1(n6165), .A2(n6801), .ZN(n5947) );
  INV_X1 U7504 ( .A(n7219), .ZN(n10150) );
  INV_X1 U7505 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6803) );
  OR2_X1 U7506 ( .A1(n5949), .A2(n6803), .ZN(n5953) );
  NAND2_X1 U7507 ( .A1(n6144), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U7508 ( .A1(n6043), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7509 ( .A1(n6181), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5950) );
  INV_X1 U7510 ( .A(n7213), .ZN(n9513) );
  INV_X1 U7511 ( .A(n6097), .ZN(n5961) );
  NAND2_X1 U7512 ( .A1(n5967), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5960) );
  INV_X1 U7513 ( .A(n5954), .ZN(n5955) );
  NAND2_X1 U7514 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5955), .ZN(n5956) );
  MUX2_X1 U7515 ( .A(n5956), .B(P1_IR_REG_31__SCAN_IN), .S(n7935), .Z(n5958)
         );
  NAND2_X1 U7516 ( .A1(n6165), .A2(n10027), .ZN(n5959) );
  NAND2_X1 U7517 ( .A1(n6144), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7518 ( .A1(n6043), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7519 ( .A1(n6039), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7520 ( .A1(n6181), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7521 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5966) );
  NAND2_X1 U7522 ( .A1(n5967), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5970) );
  INV_X1 U7523 ( .A(n6745), .ZN(n5968) );
  NAND2_X1 U7524 ( .A1(n6097), .A2(n5968), .ZN(n5969) );
  NAND2_X1 U7525 ( .A1(n6181), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7526 ( .A1(n6144), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7527 ( .A1(n6039), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7528 ( .A1(n6744), .A2(SI_0_), .ZN(n5977) );
  INV_X1 U7529 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7530 ( .A1(n5977), .A2(n5976), .ZN(n5979) );
  AND2_X1 U7531 ( .A1(n5979), .A2(n5978), .ZN(n9953) );
  NAND2_X1 U7532 ( .A1(n8577), .A2(n5982), .ZN(n5983) );
  NAND2_X1 U7533 ( .A1(n7213), .A2(n10095), .ZN(n6304) );
  NAND2_X1 U7534 ( .A1(n8576), .A2(n7219), .ZN(n6393) );
  AND2_X1 U7535 ( .A1(n6393), .A2(n6304), .ZN(n6389) );
  NAND2_X1 U7536 ( .A1(n5986), .A2(n6389), .ZN(n5987) );
  NAND2_X1 U7537 ( .A1(n6039), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7538 ( .A1(n6181), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5992) );
  INV_X1 U7539 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U7540 ( .A1(n9514), .A2(n10041), .ZN(n5989) );
  AND2_X1 U7541 ( .A1(n5989), .A2(n6007), .ZN(n7227) );
  NAND2_X1 U7542 ( .A1(n6144), .A2(n7227), .ZN(n5991) );
  NAND2_X1 U7543 ( .A1(n6043), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5990) );
  INV_X4 U7544 ( .A(n6050), .ZN(n6062) );
  NAND2_X1 U7545 ( .A1(n6062), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7546 ( .A1(n5994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7547 ( .A1(n5996), .A2(n5995), .ZN(n6014) );
  OR2_X1 U7548 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  AND2_X1 U7549 ( .A1(n6014), .A2(n5997), .ZN(n10050) );
  NAND2_X1 U7550 ( .A1(n6165), .A2(n10050), .ZN(n5998) );
  NAND2_X1 U7551 ( .A1(n6002), .A2(n7263), .ZN(n6035) );
  NAND2_X1 U7552 ( .A1(n7273), .A2(n10157), .ZN(n7264) );
  INV_X1 U7553 ( .A(n7264), .ZN(n6004) );
  INV_X1 U7554 ( .A(n6393), .ZN(n6003) );
  NOR3_X1 U7555 ( .A1(n6035), .A2(n6004), .A3(n6003), .ZN(n6033) );
  NAND2_X1 U7556 ( .A1(n6215), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7557 ( .A1(n6224), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6011) );
  INV_X1 U7558 ( .A(n6005), .ZN(n6019) );
  NAND2_X1 U7559 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  AND2_X1 U7560 ( .A1(n6019), .A2(n6008), .ZN(n7411) );
  NAND2_X1 U7561 ( .A1(n6144), .A2(n7411), .ZN(n6010) );
  NAND2_X1 U7562 ( .A1(n6228), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6009) );
  AND4_X2 U7563 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n7509)
         );
  INV_X1 U7564 ( .A(n7509), .ZN(n9510) );
  INV_X1 U7565 ( .A(n6013), .ZN(n6753) );
  NAND2_X1 U7566 ( .A1(n6062), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7567 ( .A1(n6014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6015) );
  XNOR2_X1 U7568 ( .A(n6015), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U7569 ( .A1(n6165), .A2(n9535), .ZN(n6016) );
  OAI211_X1 U7570 ( .C1(n5961), .C2(n6753), .A(n6017), .B(n6016), .ZN(n7413)
         );
  NAND2_X1 U7571 ( .A1(n9510), .A2(n10166), .ZN(n6340) );
  AND2_X1 U7572 ( .A1(n6340), .A2(n7263), .ZN(n6396) );
  INV_X1 U7573 ( .A(n6396), .ZN(n6032) );
  NAND2_X1 U7574 ( .A1(n6228), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6024) );
  INV_X1 U7575 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7576 ( .A1(n6019), .A2(n6018), .ZN(n6020) );
  AND2_X1 U7577 ( .A1(n6041), .A2(n6020), .ZN(n10082) );
  NAND2_X1 U7578 ( .A1(n6181), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7579 ( .A1(n6215), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6021) );
  NAND4_X1 U7580 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n6034)
         );
  INV_X1 U7581 ( .A(n6025), .ZN(n6755) );
  NAND2_X1 U7582 ( .A1(n6062), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7583 ( .A1(n6026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6027) );
  MUX2_X1 U7584 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6027), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6028) );
  INV_X1 U7585 ( .A(n6028), .ZN(n6029) );
  NOR2_X1 U7586 ( .A1(n6029), .A2(n5895), .ZN(n6822) );
  NAND2_X1 U7587 ( .A1(n6165), .A2(n6822), .ZN(n6030) );
  NAND2_X1 U7588 ( .A1(n7494), .A2(n10083), .ZN(n7369) );
  NAND2_X1 U7589 ( .A1(n7509), .A2(n7413), .ZN(n6307) );
  NAND2_X1 U7590 ( .A1(n6034), .A2(n10174), .ZN(n7370) );
  INV_X1 U7591 ( .A(n6035), .ZN(n6036) );
  NAND2_X1 U7592 ( .A1(n7264), .A2(n6307), .ZN(n6341) );
  AOI21_X1 U7593 ( .B1(n6036), .B2(n6391), .A(n6341), .ZN(n6038) );
  NAND2_X1 U7594 ( .A1(n7370), .A2(n6340), .ZN(n6037) );
  NAND2_X1 U7595 ( .A1(n6215), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7596 ( .A1(n6181), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7597 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  AND2_X1 U7598 ( .A1(n6052), .A2(n6042), .ZN(n7493) );
  NAND2_X1 U7599 ( .A1(n6144), .A2(n7493), .ZN(n6045) );
  NAND2_X1 U7600 ( .A1(n6043), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6044) );
  INV_X1 U7601 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6768) );
  OR2_X1 U7602 ( .A1(n5895), .A2(n5815), .ZN(n6048) );
  XNOR2_X1 U7603 ( .A(n6048), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U7604 ( .A1(n6165), .A2(n7043), .ZN(n6049) );
  NAND2_X1 U7605 ( .A1(n9992), .A2(n7499), .ZN(n8025) );
  INV_X1 U7606 ( .A(n9992), .ZN(n9509) );
  NAND2_X1 U7607 ( .A1(n8025), .A2(n6065), .ZN(n7382) );
  INV_X1 U7608 ( .A(n7382), .ZN(n8005) );
  NAND2_X1 U7609 ( .A1(n6224), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7610 ( .A1(n6215), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7611 ( .A1(n6228), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7612 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  NAND2_X1 U7613 ( .A1(n6075), .A2(n6053), .ZN(n10004) );
  INV_X1 U7614 ( .A(n10004), .ZN(n10066) );
  NAND2_X1 U7615 ( .A1(n6227), .A2(n10066), .ZN(n6054) );
  NAND2_X1 U7616 ( .A1(n6771), .A2(n6191), .ZN(n6064) );
  NOR2_X1 U7617 ( .A1(n6058), .A2(n5815), .ZN(n6059) );
  NAND2_X1 U7618 ( .A1(n6059), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6061) );
  INV_X1 U7619 ( .A(n6059), .ZN(n6060) );
  INV_X1 U7620 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U7621 ( .A1(n6060), .A2(n7931), .ZN(n6070) );
  AND2_X1 U7622 ( .A1(n6061), .A2(n6070), .ZN(n9544) );
  AOI22_X1 U7623 ( .A1(n6062), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6165), .B2(
        n9544), .ZN(n6063) );
  NAND2_X1 U7624 ( .A1(n6064), .A2(n6063), .ZN(n10067) );
  INV_X1 U7625 ( .A(n10067), .ZN(n10187) );
  AND2_X1 U7626 ( .A1(n8006), .A2(n6065), .ZN(n6309) );
  INV_X1 U7627 ( .A(n6309), .ZN(n6067) );
  NAND2_X1 U7628 ( .A1(n6066), .A2(n10067), .ZN(n8007) );
  NAND2_X1 U7629 ( .A1(n8025), .A2(n8007), .ZN(n6312) );
  MUX2_X1 U7630 ( .A(n6067), .B(n6312), .S(n9858), .Z(n6068) );
  INV_X1 U7631 ( .A(n8006), .ZN(n8026) );
  NAND2_X1 U7632 ( .A1(n6069), .A2(n6191), .ZN(n6073) );
  NAND2_X1 U7633 ( .A1(n6070), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7634 ( .A(n6071), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7295) );
  AOI22_X1 U7635 ( .A1(n6062), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6165), .B2(
        n7295), .ZN(n6072) );
  NAND2_X1 U7636 ( .A1(n6224), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7637 ( .A1(n6228), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6079) );
  INV_X1 U7638 ( .A(n6074), .ZN(n6090) );
  NAND2_X1 U7639 ( .A1(n6075), .A2(n7047), .ZN(n6076) );
  AND2_X1 U7640 ( .A1(n6090), .A2(n6076), .ZN(n9429) );
  NAND2_X1 U7641 ( .A1(n6227), .A2(n9429), .ZN(n6078) );
  NAND2_X1 U7642 ( .A1(n6215), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7643 ( .A1(n9430), .A2(n9990), .ZN(n8015) );
  NAND2_X1 U7644 ( .A1(n8015), .A2(n8007), .ZN(n6081) );
  MUX2_X1 U7645 ( .A(n8026), .B(n6081), .S(n5984), .Z(n6082) );
  NAND2_X1 U7646 ( .A1(n6781), .A2(n6191), .ZN(n6088) );
  NOR2_X1 U7647 ( .A1(n6083), .A2(n5815), .ZN(n6084) );
  MUX2_X1 U7648 ( .A(n5815), .B(n6084), .S(P1_IR_REG_10__SCAN_IN), .Z(n6085)
         );
  INV_X1 U7649 ( .A(n6085), .ZN(n6086) );
  AOI22_X1 U7650 ( .A1(n6062), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6165), .B2(
        n7359), .ZN(n6087) );
  NAND2_X1 U7651 ( .A1(n6088), .A2(n6087), .ZN(n8069) );
  NAND2_X1 U7652 ( .A1(n6224), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7653 ( .A1(n6228), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6094) );
  INV_X1 U7654 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7655 ( .A1(n6090), .A2(n6089), .ZN(n6091) );
  AND2_X1 U7656 ( .A1(n6102), .A2(n6091), .ZN(n8461) );
  NAND2_X1 U7657 ( .A1(n6227), .A2(n8461), .ZN(n6093) );
  NAND2_X1 U7658 ( .A1(n6215), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7659 ( .A1(n8069), .A2(n8428), .ZN(n6401) );
  NAND2_X1 U7660 ( .A1(n6401), .A2(n8016), .ZN(n6096) );
  NAND2_X1 U7661 ( .A1(n8069), .A2(n8428), .ZN(n8072) );
  OAI21_X1 U7662 ( .B1(n6126), .B2(n6096), .A(n8072), .ZN(n6122) );
  NAND2_X1 U7663 ( .A1(n6817), .A2(n6191), .ZN(n6101) );
  NAND2_X1 U7664 ( .A1(n6098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7665 ( .A(n6099), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7443) );
  AOI22_X1 U7666 ( .A1(n6062), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6165), .B2(
        n7443), .ZN(n6100) );
  NAND2_X1 U7667 ( .A1(n6215), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7668 ( .A1(n6224), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7669 ( .A1(n6102), .A2(n8426), .ZN(n6103) );
  AND2_X1 U7670 ( .A1(n6114), .A2(n6103), .ZN(n8425) );
  NAND2_X1 U7671 ( .A1(n6144), .A2(n8425), .ZN(n6105) );
  NAND2_X1 U7672 ( .A1(n6228), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7673 ( .A1(n8431), .A2(n8123), .ZN(n8116) );
  NAND2_X1 U7674 ( .A1(n6836), .A2(n6191), .ZN(n6112) );
  NAND2_X1 U7675 ( .A1(n6108), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6110) );
  AND2_X1 U7676 ( .A1(n6110), .A2(n6109), .ZN(n8107) );
  AOI22_X1 U7677 ( .A1(n6062), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6165), .B2(
        n8107), .ZN(n6111) );
  NAND2_X1 U7678 ( .A1(n6215), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7679 ( .A1(n6224), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7680 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  AND2_X1 U7681 ( .A1(n6116), .A2(n6115), .ZN(n8436) );
  NAND2_X1 U7682 ( .A1(n6227), .A2(n8436), .ZN(n6118) );
  NAND2_X1 U7683 ( .A1(n6228), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7684 ( .A1(n8431), .A2(n8123), .ZN(n6311) );
  INV_X1 U7685 ( .A(n6311), .ZN(n6121) );
  OR2_X1 U7686 ( .A1(n9398), .A2(n9486), .ZN(n6422) );
  INV_X1 U7687 ( .A(n6422), .ZN(n6124) );
  OR2_X1 U7688 ( .A1(n9920), .A2(n9489), .ZN(n6413) );
  OR2_X1 U7689 ( .A1(n8528), .A2(n8288), .ZN(n6412) );
  OR2_X1 U7690 ( .A1(n8442), .A2(n9504), .ZN(n6317) );
  NAND4_X1 U7691 ( .A1(n6413), .A2(n5984), .A3(n6412), .A4(n6317), .ZN(n6123)
         );
  INV_X1 U7692 ( .A(n6126), .ZN(n6128) );
  INV_X1 U7693 ( .A(n8016), .ZN(n6127) );
  OAI21_X1 U7694 ( .B1(n6128), .B2(n6127), .A(n8015), .ZN(n6129) );
  NAND2_X1 U7695 ( .A1(n6311), .A2(n8072), .ZN(n6404) );
  AOI21_X1 U7696 ( .B1(n6129), .B2(n6401), .A(n6404), .ZN(n6132) );
  NAND2_X1 U7697 ( .A1(n6317), .A2(n8116), .ZN(n6407) );
  NAND2_X1 U7698 ( .A1(n8528), .A2(n8288), .ZN(n8285) );
  INV_X1 U7699 ( .A(n8285), .ZN(n6130) );
  NOR3_X1 U7700 ( .A1(n6130), .A2(n4830), .A3(n5984), .ZN(n6131) );
  NAND2_X1 U7701 ( .A1(n9920), .A2(n9489), .ZN(n6415) );
  OAI211_X1 U7702 ( .C1(n6132), .C2(n6407), .A(n6131), .B(n6415), .ZN(n6137)
         );
  INV_X1 U7703 ( .A(n6416), .ZN(n6133) );
  NAND2_X1 U7704 ( .A1(n6422), .A2(n6133), .ZN(n6134) );
  NAND2_X1 U7705 ( .A1(n9398), .A2(n9486), .ZN(n6420) );
  OAI211_X1 U7706 ( .C1(n9916), .C2(n9858), .A(n6134), .B(n6420), .ZN(n6136)
         );
  OAI21_X1 U7707 ( .B1(n4853), .B2(n9395), .A(n5984), .ZN(n6135) );
  NAND2_X1 U7708 ( .A1(n7063), .A2(n6191), .ZN(n6140) );
  XNOR2_X1 U7709 ( .A(n6138), .B(n7776), .ZN(n9605) );
  AOI22_X1 U7710 ( .A1(n6062), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6165), .B2(
        n9605), .ZN(n6139) );
  NAND2_X1 U7711 ( .A1(n6215), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7712 ( .A1(n6224), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6147) );
  AND2_X1 U7713 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  NOR2_X1 U7714 ( .A1(n6158), .A2(n6143), .ZN(n9409) );
  NAND2_X1 U7715 ( .A1(n6144), .A2(n9409), .ZN(n6146) );
  NAND2_X1 U7716 ( .A1(n6228), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6145) );
  NAND4_X1 U7717 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n9499)
         );
  INV_X1 U7718 ( .A(n9499), .ZN(n9462) );
  OR2_X1 U7719 ( .A1(n9911), .A2(n9462), .ZN(n6423) );
  NAND2_X1 U7720 ( .A1(n9911), .A2(n9462), .ZN(n6206) );
  NAND2_X1 U7721 ( .A1(n6423), .A2(n6206), .ZN(n8549) );
  NAND2_X1 U7722 ( .A1(n7123), .A2(n6191), .ZN(n6157) );
  OR2_X1 U7723 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6149) );
  AND2_X1 U7724 ( .A1(n6150), .A2(n6149), .ZN(n6155) );
  OR2_X1 U7725 ( .A1(n6138), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7726 ( .A1(n6151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6153) );
  OR2_X1 U7727 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  AND2_X1 U7728 ( .A1(n6155), .A2(n6154), .ZN(n9622) );
  AOI22_X1 U7729 ( .A1(n6062), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6165), .B2(
        n9622), .ZN(n6156) );
  NAND2_X1 U7730 ( .A1(n6215), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7731 ( .A1(n6181), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6162) );
  OR2_X1 U7732 ( .A1(n6158), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6159) );
  AND2_X1 U7733 ( .A1(n6168), .A2(n6159), .ZN(n9459) );
  NAND2_X1 U7734 ( .A1(n6227), .A2(n9459), .ZN(n6161) );
  NAND2_X1 U7735 ( .A1(n6228), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6160) );
  NAND4_X1 U7736 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n9646)
         );
  OR2_X1 U7737 ( .A1(n9645), .A2(n9837), .ZN(n9831) );
  AND2_X1 U7738 ( .A1(n9831), .A2(n6423), .ZN(n6164) );
  NAND2_X1 U7739 ( .A1(n7284), .A2(n6191), .ZN(n6167) );
  AOI22_X1 U7740 ( .A1(n6062), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6165), .B2(
        n6504), .ZN(n6166) );
  NAND2_X1 U7741 ( .A1(n6215), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7742 ( .A1(n6224), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7743 ( .A1(n6168), .A2(n9368), .ZN(n6169) );
  AND2_X1 U7744 ( .A1(n6179), .A2(n6169), .ZN(n9367) );
  NAND2_X1 U7745 ( .A1(n6227), .A2(n9367), .ZN(n6171) );
  NAND2_X1 U7746 ( .A1(n6228), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7747 ( .A1(n9850), .A2(n9649), .ZN(n6426) );
  NAND2_X1 U7748 ( .A1(n9645), .A2(n9837), .ZN(n6303) );
  NAND2_X1 U7749 ( .A1(n7338), .A2(n6191), .ZN(n6178) );
  NAND2_X1 U7750 ( .A1(n6062), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6177) );
  AND2_X1 U7751 ( .A1(n6179), .A2(n9440), .ZN(n6180) );
  OR2_X1 U7752 ( .A1(n6180), .A2(n6194), .ZN(n9822) );
  INV_X1 U7753 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7754 ( .A1(n6181), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7755 ( .A1(n6228), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6182) );
  OAI211_X1 U7756 ( .C1(n6184), .C2(n5949), .A(n6183), .B(n6182), .ZN(n6185)
         );
  INV_X1 U7757 ( .A(n6185), .ZN(n6186) );
  OAI21_X1 U7758 ( .B1(n9822), .B2(n6196), .A(n6186), .ZN(n9835) );
  INV_X1 U7759 ( .A(n9835), .ZN(n9807) );
  OR2_X1 U7760 ( .A1(n9824), .A2(n9807), .ZN(n9673) );
  INV_X1 U7761 ( .A(n9673), .ZN(n6190) );
  OR2_X1 U7762 ( .A1(n9850), .A2(n9649), .ZN(n6302) );
  INV_X1 U7763 ( .A(n6302), .ZN(n6189) );
  NAND2_X1 U7764 ( .A1(n9824), .A2(n9807), .ZN(n6301) );
  AOI21_X1 U7765 ( .B1(n6301), .B2(n9961), .A(n5984), .ZN(n6188) );
  INV_X1 U7766 ( .A(n6301), .ZN(n6187) );
  OAI33_X1 U7767 ( .A1(n6190), .A2(n6189), .A3(n6188), .B1(n6187), .B2(n9649), 
        .B3(n5984), .ZN(n6203) );
  NAND2_X1 U7768 ( .A1(n7390), .A2(n6191), .ZN(n6193) );
  NAND2_X1 U7769 ( .A1(n6062), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7770 ( .A1(n6194), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7771 ( .A1(n6195), .A2(n6217), .ZN(n9811) );
  OR2_X1 U7772 ( .A1(n9811), .A2(n6196), .ZN(n6202) );
  INV_X1 U7773 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7774 ( .A1(n6228), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7775 ( .A1(n6224), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6197) );
  OAI211_X1 U7776 ( .C1(n5949), .C2(n6199), .A(n6198), .B(n6197), .ZN(n6200)
         );
  INV_X1 U7777 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7778 ( .A1(n6202), .A2(n6201), .ZN(n9795) );
  INV_X1 U7779 ( .A(n9795), .ZN(n9653) );
  NAND2_X1 U7780 ( .A1(n9906), .A2(n9653), .ZN(n9675) );
  NAND2_X1 U7781 ( .A1(n9675), .A2(n6301), .ZN(n6353) );
  AOI22_X1 U7782 ( .A1(n6204), .A2(n6203), .B1(n5984), .B2(n6353), .ZN(n6211)
         );
  INV_X1 U7783 ( .A(n6205), .ZN(n6208) );
  NAND2_X1 U7784 ( .A1(n6303), .A2(n6206), .ZN(n6384) );
  AND2_X1 U7785 ( .A1(n6302), .A2(n9831), .ZN(n6428) );
  OAI21_X1 U7786 ( .B1(n6208), .B2(n6384), .A(n6207), .ZN(n6209) );
  OR2_X1 U7787 ( .A1(n9906), .A2(n9653), .ZN(n6354) );
  NAND2_X1 U7788 ( .A1(n6209), .A2(n6354), .ZN(n6210) );
  AND2_X1 U7789 ( .A1(n9673), .A2(n6354), .ZN(n6336) );
  OAI22_X1 U7790 ( .A1(n6211), .A2(n6210), .B1(n6336), .B2(n5984), .ZN(n6212)
         );
  NAND2_X1 U7791 ( .A1(n6212), .A2(n5107), .ZN(n6235) );
  NAND2_X1 U7792 ( .A1(n7982), .A2(n6191), .ZN(n6214) );
  NAND2_X1 U7793 ( .A1(n6062), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7794 ( .A1(n6224), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7795 ( .A1(n6215), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6220) );
  INV_X1 U7796 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9449) );
  AOI21_X1 U7797 ( .B1(n9449), .B2(n6217), .A(n6216), .ZN(n9788) );
  NAND2_X1 U7798 ( .A1(n6227), .A2(n9788), .ZN(n6219) );
  NAND2_X1 U7799 ( .A1(n6228), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6218) );
  XNOR2_X1 U7800 ( .A(n9900), .B(n9654), .ZN(n9792) );
  NAND2_X1 U7801 ( .A1(n8065), .A2(n6191), .ZN(n6223) );
  NAND2_X1 U7802 ( .A1(n6062), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7803 ( .A1(n6215), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7804 ( .A1(n6224), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6231) );
  INV_X1 U7805 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8590) );
  AOI21_X1 U7806 ( .B1(n8590), .B2(n6226), .A(n6225), .ZN(n9780) );
  NAND2_X1 U7807 ( .A1(n6227), .A2(n9780), .ZN(n6230) );
  NAND2_X1 U7808 ( .A1(n6228), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6229) );
  NAND4_X1 U7809 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n9796)
         );
  INV_X1 U7810 ( .A(n9796), .ZN(n9762) );
  OR2_X1 U7811 ( .A1(n9774), .A2(n9762), .ZN(n6300) );
  NAND2_X1 U7812 ( .A1(n9790), .A2(n9654), .ZN(n6233) );
  NAND2_X1 U7813 ( .A1(n6300), .A2(n6233), .ZN(n6331) );
  NAND2_X1 U7814 ( .A1(n9774), .A2(n9762), .ZN(n9758) );
  NAND2_X1 U7815 ( .A1(n9900), .A2(n9808), .ZN(n9676) );
  NAND2_X1 U7816 ( .A1(n9758), .A2(n9676), .ZN(n6355) );
  MUX2_X1 U7817 ( .A(n6331), .B(n6355), .S(n9858), .Z(n6234) );
  AOI21_X1 U7818 ( .B1(n6235), .B2(n9792), .A(n6234), .ZN(n6248) );
  NAND2_X1 U7819 ( .A1(n8176), .A2(n6191), .ZN(n6237) );
  NAND2_X1 U7820 ( .A1(n6062), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7821 ( .A1(n6215), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7822 ( .A1(n6224), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6243) );
  INV_X1 U7823 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6240) );
  AOI21_X1 U7824 ( .B1(n6240), .B2(n6239), .A(n6238), .ZN(n9767) );
  NAND2_X1 U7825 ( .A1(n6227), .A2(n9767), .ZN(n6242) );
  NAND2_X1 U7826 ( .A1(n6228), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7827 ( .A1(n9889), .A2(n9747), .ZN(n6357) );
  MUX2_X1 U7828 ( .A(n9758), .B(n6300), .S(n9858), .Z(n6245) );
  NAND2_X1 U7829 ( .A1(n9760), .A2(n6245), .ZN(n6247) );
  MUX2_X1 U7830 ( .A(n9677), .B(n6357), .S(n9858), .Z(n6246) );
  OAI21_X1 U7831 ( .B1(n6248), .B2(n6247), .A(n6246), .ZN(n6265) );
  NAND2_X1 U7832 ( .A1(n8191), .A2(n6191), .ZN(n6250) );
  NAND2_X1 U7833 ( .A1(n5967), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7834 ( .A1(n6215), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7835 ( .A1(n6224), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6256) );
  INV_X1 U7836 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6253) );
  AOI21_X1 U7837 ( .B1(n6253), .B2(n6252), .A(n6251), .ZN(n9750) );
  NAND2_X1 U7838 ( .A1(n6227), .A2(n9750), .ZN(n6255) );
  NAND2_X1 U7839 ( .A1(n6228), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6254) );
  NAND4_X1 U7840 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6254), .ZN(n9661)
         );
  INV_X1 U7841 ( .A(n9661), .ZN(n9763) );
  NAND2_X1 U7842 ( .A1(n9879), .A2(n9748), .ZN(n6429) );
  NAND2_X1 U7843 ( .A1(n9884), .A2(n9763), .ZN(n6360) );
  NAND2_X1 U7844 ( .A1(n6429), .A2(n6360), .ZN(n6262) );
  AOI21_X1 U7845 ( .B1(n6265), .B2(n6335), .A(n6262), .ZN(n6259) );
  INV_X1 U7846 ( .A(n6351), .ZN(n6258) );
  NOR3_X1 U7847 ( .A1(n6259), .A2(n6258), .A3(n5984), .ZN(n6260) );
  AOI211_X1 U7848 ( .C1(n6364), .C2(n6261), .A(n9682), .B(n6260), .ZN(n6269)
         );
  INV_X1 U7849 ( .A(n6335), .ZN(n6264) );
  INV_X1 U7850 ( .A(n6262), .ZN(n6263) );
  OAI211_X1 U7851 ( .C1(n6265), .C2(n6264), .A(n5984), .B(n6263), .ZN(n6266)
         );
  MUX2_X1 U7852 ( .A(n6266), .B(n5984), .S(n6436), .Z(n6268) );
  OAI21_X1 U7853 ( .B1(n6436), .B2(n6352), .A(n6329), .ZN(n6267) );
  AOI22_X1 U7854 ( .A1(n6269), .A2(n6268), .B1(n9858), .B2(n6267), .ZN(n6271)
         );
  MUX2_X1 U7855 ( .A(n6366), .B(n6330), .S(n9858), .Z(n6270) );
  INV_X1 U7856 ( .A(SI_29_), .ZN(n7697) );
  INV_X1 U7857 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6277) );
  INV_X1 U7858 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7869) );
  MUX2_X1 U7859 ( .A(n6277), .B(n7869), .S(n6738), .Z(n6278) );
  NAND2_X1 U7860 ( .A1(n6278), .A2(n7920), .ZN(n6283) );
  INV_X1 U7861 ( .A(n6278), .ZN(n6279) );
  NAND2_X1 U7862 ( .A1(n6279), .A2(SI_30_), .ZN(n6280) );
  NAND2_X1 U7863 ( .A1(n6283), .A2(n6280), .ZN(n6284) );
  NAND2_X1 U7864 ( .A1(n9351), .A2(n6191), .ZN(n6282) );
  NAND2_X1 U7865 ( .A1(n5967), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6281) );
  MUX2_X1 U7866 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6286), .Z(n6288) );
  INV_X1 U7867 ( .A(SI_31_), .ZN(n6287) );
  XNOR2_X1 U7868 ( .A(n6288), .B(n6287), .ZN(n6289) );
  NAND2_X1 U7869 ( .A1(n6215), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7870 ( .A1(n6224), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7871 ( .A1(n6228), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6291) );
  AND3_X1 U7872 ( .A1(n6293), .A2(n6292), .A3(n6291), .ZN(n9686) );
  INV_X1 U7873 ( .A(n9686), .ZN(n9496) );
  NAND2_X1 U7874 ( .A1(n6215), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7875 ( .A1(n6224), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7876 ( .A1(n6228), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6294) );
  AND3_X1 U7877 ( .A1(n6296), .A2(n6295), .A3(n6294), .ZN(n6474) );
  OAI21_X1 U7878 ( .B1(n9636), .B2(n9496), .A(n4957), .ZN(n6297) );
  XNOR2_X1 U7879 ( .A(n6299), .B(n6298), .ZN(n7392) );
  INV_X1 U7880 ( .A(n7392), .ZN(n6466) );
  OAI21_X1 U7881 ( .B1(n6463), .B2(n7985), .A(n6466), .ZN(n6327) );
  OR2_X1 U7882 ( .A1(n6471), .A2(n9686), .ZN(n6328) );
  NAND2_X1 U7883 ( .A1(n6471), .A2(n9686), .ZN(n6367) );
  NAND2_X1 U7884 ( .A1(n6351), .A2(n6429), .ZN(n9729) );
  NAND2_X1 U7885 ( .A1(n9673), .A2(n6301), .ZN(n9819) );
  XNOR2_X1 U7886 ( .A(n9906), .B(n9653), .ZN(n9805) );
  NAND2_X1 U7887 ( .A1(n6302), .A2(n6426), .ZN(n9840) );
  NAND2_X1 U7888 ( .A1(n6422), .A2(n6420), .ZN(n8547) );
  NAND2_X1 U7889 ( .A1(n6417), .A2(n6416), .ZN(n8329) );
  NOR2_X1 U7890 ( .A1(n7271), .A2(n10098), .ZN(n6305) );
  NAND2_X1 U7891 ( .A1(n7264), .A2(n7263), .ZN(n7276) );
  INV_X1 U7892 ( .A(n7276), .ZN(n7329) );
  AND2_X1 U7893 ( .A1(n6991), .A2(n10111), .ZN(n6385) );
  NOR2_X1 U7894 ( .A1(n6993), .A2(n6385), .ZN(n10128) );
  NAND4_X1 U7895 ( .A1(n6305), .A2(n7329), .A3(n10128), .A4(n7392), .ZN(n6308)
         );
  NAND2_X1 U7896 ( .A1(n6307), .A2(n6340), .ZN(n7376) );
  OR3_X1 U7897 ( .A1(n6308), .A2(n7210), .A3(n7376), .ZN(n6310) );
  NAND3_X1 U7898 ( .A1(n6309), .A2(n8016), .A3(n7370), .ZN(n6343) );
  NOR2_X1 U7899 ( .A1(n6310), .A2(n6343), .ZN(n6316) );
  NAND2_X1 U7900 ( .A1(n6401), .A2(n8072), .ZN(n8070) );
  INV_X1 U7901 ( .A(n8070), .ZN(n6315) );
  NAND3_X1 U7902 ( .A1(n6312), .A2(n8016), .A3(n8006), .ZN(n6313) );
  AND2_X1 U7903 ( .A1(n6313), .A2(n8015), .ZN(n6344) );
  NAND2_X1 U7904 ( .A1(n6344), .A2(n7369), .ZN(n6402) );
  INV_X1 U7905 ( .A(n6402), .ZN(n6314) );
  NAND4_X1 U7906 ( .A1(n6316), .A2(n8125), .A3(n6315), .A4(n6314), .ZN(n6318)
         );
  NOR2_X1 U7907 ( .A1(n6318), .A2(n8291), .ZN(n6319) );
  NAND3_X1 U7908 ( .A1(n8293), .A2(n8311), .A3(n6319), .ZN(n6320) );
  NOR2_X1 U7909 ( .A1(n8329), .A2(n6320), .ZN(n6321) );
  NAND4_X1 U7910 ( .A1(n8559), .A2(n5083), .A3(n4850), .A4(n6321), .ZN(n6322)
         );
  NAND4_X1 U7911 ( .A1(n9760), .A2(n9775), .A3(n5110), .A4(n9792), .ZN(n6323)
         );
  NAND2_X1 U7912 ( .A1(n6335), .A2(n6360), .ZN(n9745) );
  OR3_X1 U7913 ( .A1(n9729), .A2(n6323), .A3(n9745), .ZN(n6324) );
  NOR2_X1 U7914 ( .A1(n9718), .A2(n6324), .ZN(n6325) );
  NAND4_X1 U7915 ( .A1(n9670), .A2(n9702), .A3(n6367), .A4(n6325), .ZN(n6326)
         );
  INV_X1 U7916 ( .A(n6328), .ZN(n6370) );
  AND2_X1 U7917 ( .A1(n6330), .A2(n6329), .ZN(n6381) );
  NAND2_X1 U7918 ( .A1(n6331), .A2(n9758), .ZN(n6332) );
  NAND2_X1 U7919 ( .A1(n9677), .A2(n6332), .ZN(n6333) );
  NAND2_X1 U7920 ( .A1(n6333), .A2(n6357), .ZN(n6334) );
  AND2_X1 U7921 ( .A1(n6335), .A2(n6334), .ZN(n6362) );
  INV_X1 U7922 ( .A(n6362), .ZN(n6338) );
  INV_X1 U7923 ( .A(n6336), .ZN(n6337) );
  NOR2_X1 U7924 ( .A1(n6338), .A2(n6337), .ZN(n6383) );
  NAND2_X1 U7925 ( .A1(n7206), .A2(n7205), .ZN(n6339) );
  NAND2_X1 U7926 ( .A1(n6339), .A2(n6393), .ZN(n7262) );
  NAND2_X1 U7927 ( .A1(n7262), .A2(n6396), .ZN(n6342) );
  NAND2_X1 U7928 ( .A1(n6341), .A2(n6340), .ZN(n6398) );
  NAND2_X1 U7929 ( .A1(n6344), .A2(n6343), .ZN(n6400) );
  OAI21_X1 U7930 ( .B1(n10079), .B2(n6402), .A(n6400), .ZN(n8001) );
  INV_X1 U7931 ( .A(n8125), .ZN(n8074) );
  INV_X1 U7932 ( .A(n8072), .ZN(n6345) );
  NOR2_X1 U7933 ( .A1(n8074), .A2(n6345), .ZN(n6346) );
  AND2_X1 U7934 ( .A1(n8119), .A2(n8116), .ZN(n6347) );
  AND2_X1 U7935 ( .A1(n8285), .A2(n6415), .ZN(n6349) );
  INV_X1 U7936 ( .A(n6413), .ZN(n6348) );
  NAND2_X1 U7937 ( .A1(n9832), .A2(n6428), .ZN(n6350) );
  INV_X1 U7938 ( .A(n6429), .ZN(n9679) );
  AOI21_X1 U7939 ( .B1(n6383), .B2(n9672), .A(n9679), .ZN(n6365) );
  NAND2_X1 U7940 ( .A1(n6352), .A2(n6351), .ZN(n6382) );
  INV_X1 U7941 ( .A(n6353), .ZN(n6359) );
  INV_X1 U7942 ( .A(n6354), .ZN(n6358) );
  INV_X1 U7943 ( .A(n6355), .ZN(n6356) );
  OAI211_X1 U7944 ( .C1(n6359), .C2(n6358), .A(n6357), .B(n6356), .ZN(n6361)
         );
  INV_X1 U7945 ( .A(n6360), .ZN(n9678) );
  AOI21_X1 U7946 ( .B1(n6362), .B2(n6361), .A(n9678), .ZN(n6363) );
  OR2_X1 U7947 ( .A1(n6382), .A2(n6363), .ZN(n6434) );
  OAI211_X1 U7948 ( .C1(n6365), .C2(n6382), .A(n6364), .B(n6434), .ZN(n6368)
         );
  NAND2_X1 U7949 ( .A1(n6367), .A2(n6366), .ZN(n6440) );
  AOI21_X1 U7950 ( .B1(n6381), .B2(n6368), .A(n6440), .ZN(n6369) );
  AOI21_X1 U7951 ( .B1(n6370), .B2(n4957), .A(n6369), .ZN(n6371) );
  AOI21_X1 U7952 ( .B1(n6474), .B2(n6471), .A(n6371), .ZN(n6374) );
  INV_X1 U7953 ( .A(n7985), .ZN(n6499) );
  AND2_X1 U7954 ( .A1(n6499), .A2(n6466), .ZN(n6985) );
  INV_X1 U7955 ( .A(n6985), .ZN(n6373) );
  AOI211_X1 U7956 ( .C1(n6374), .C2(n6465), .A(n6464), .B(n6373), .ZN(n6377)
         );
  INV_X1 U7957 ( .A(n6375), .ZN(n6376) );
  NAND2_X1 U7958 ( .A1(n6378), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6380) );
  INV_X1 U7959 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6379) );
  INV_X1 U7960 ( .A(n6381), .ZN(n6439) );
  INV_X1 U7961 ( .A(n6382), .ZN(n6433) );
  INV_X1 U7962 ( .A(n6383), .ZN(n6431) );
  INV_X1 U7963 ( .A(n6384), .ZN(n6425) );
  INV_X1 U7964 ( .A(n6385), .ZN(n6387) );
  NAND2_X1 U7965 ( .A1(n5981), .A2(n10137), .ZN(n6386) );
  NAND3_X1 U7966 ( .A1(n6387), .A2(n6466), .A3(n6386), .ZN(n6388) );
  NAND2_X1 U7967 ( .A1(n6389), .A2(n6388), .ZN(n6397) );
  INV_X1 U7968 ( .A(n6390), .ZN(n6394) );
  INV_X1 U7969 ( .A(n6391), .ZN(n6392) );
  AOI21_X1 U7970 ( .B1(n6394), .B2(n6393), .A(n6392), .ZN(n6395) );
  OAI211_X1 U7971 ( .C1(n10090), .C2(n6397), .A(n6396), .B(n6395), .ZN(n6399)
         );
  NAND2_X1 U7972 ( .A1(n6399), .A2(n6398), .ZN(n6403) );
  OAI211_X1 U7973 ( .C1(n6403), .C2(n6402), .A(n6401), .B(n6400), .ZN(n6406)
         );
  INV_X1 U7974 ( .A(n6404), .ZN(n6405) );
  NAND2_X1 U7975 ( .A1(n6406), .A2(n6405), .ZN(n6409) );
  INV_X1 U7976 ( .A(n6407), .ZN(n6408) );
  NAND2_X1 U7977 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  NAND3_X1 U7978 ( .A1(n6410), .A2(n8285), .A3(n8304), .ZN(n6411) );
  NAND3_X1 U7979 ( .A1(n6413), .A2(n6412), .A3(n6411), .ZN(n6414) );
  NAND3_X1 U7980 ( .A1(n6416), .A2(n6415), .A3(n6414), .ZN(n6418) );
  NAND2_X1 U7981 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  NAND2_X1 U7982 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  NAND3_X1 U7983 ( .A1(n6423), .A2(n6422), .A3(n6421), .ZN(n6424) );
  NAND2_X1 U7984 ( .A1(n6425), .A2(n6424), .ZN(n6427) );
  AOI21_X1 U7985 ( .B1(n6428), .B2(n6427), .A(n6175), .ZN(n6430) );
  OAI21_X1 U7986 ( .B1(n6431), .B2(n6430), .A(n6429), .ZN(n6432) );
  NAND2_X1 U7987 ( .A1(n6433), .A2(n6432), .ZN(n6435) );
  NAND2_X1 U7988 ( .A1(n6435), .A2(n6434), .ZN(n6437) );
  NOR2_X1 U7989 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  NOR2_X1 U7990 ( .A1(n6439), .A2(n6438), .ZN(n6441) );
  NOR2_X1 U7991 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  OR2_X1 U7992 ( .A1(n6443), .A2(n6442), .ZN(n6444) );
  NAND2_X1 U7993 ( .A1(n6444), .A2(n6465), .ZN(n6450) );
  NAND3_X1 U7994 ( .A1(n6450), .A2(n6504), .A3(n7352), .ZN(n6449) );
  NAND2_X1 U7995 ( .A1(n6445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6447) );
  XNOR2_X1 U7996 ( .A(n6447), .B(n6446), .ZN(n6776) );
  OR2_X1 U7997 ( .A1(n6776), .A2(P1_U3086), .ZN(n8066) );
  INV_X1 U7998 ( .A(n8066), .ZN(n6448) );
  OAI211_X1 U7999 ( .C1(n6450), .C2(n6989), .A(n6449), .B(n6448), .ZN(n6451)
         );
  INV_X1 U8000 ( .A(n6452), .ZN(n10031) );
  NAND2_X1 U8001 ( .A1(n10031), .A2(n6985), .ZN(n9991) );
  NAND2_X1 U8002 ( .A1(n4561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6458) );
  INV_X1 U8003 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U8004 ( .A1(n6458), .A2(n7972), .ZN(n6460) );
  NAND2_X1 U8005 ( .A1(n6460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6453) );
  XNOR2_X1 U8006 ( .A(n6453), .B(n5813), .ZN(n8303) );
  INV_X1 U8007 ( .A(n6454), .ZN(n6455) );
  NAND2_X1 U8008 ( .A1(n6455), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6457) );
  XNOR2_X1 U8009 ( .A(n6457), .B(n6456), .ZN(n8178) );
  OR2_X1 U8010 ( .A1(n6458), .A2(n7972), .ZN(n6459) );
  NAND2_X1 U8011 ( .A1(n6460), .A2(n6459), .ZN(n8216) );
  AND2_X1 U8012 ( .A1(n6776), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6733) );
  NAND2_X1 U8013 ( .A1(n6775), .A2(n6733), .ZN(n9939) );
  NOR4_X1 U8014 ( .A1(n9991), .A2(n9939), .A3(n10028), .A4(n6989), .ZN(n6462)
         );
  OR2_X1 U8015 ( .A1(n8066), .A2(n6499), .ZN(n6467) );
  INV_X1 U8016 ( .A(n6467), .ZN(n6461) );
  INV_X1 U8017 ( .A(P1_B_REG_SCAN_IN), .ZN(n6473) );
  AOI21_X1 U8018 ( .B1(n6504), .B2(n6464), .A(n6463), .ZN(n6469) );
  NOR2_X1 U8019 ( .A1(n6465), .A2(n4507), .ZN(n6468) );
  NAND2_X1 U8020 ( .A1(n6466), .A2(n9857), .ZN(n6994) );
  NAND3_X1 U8021 ( .A1(n6470), .A2(n5094), .A3(n4543), .ZN(P1_U3242) );
  NAND2_X1 U8022 ( .A1(n10101), .A2(n10143), .ZN(n10100) );
  INV_X1 U8023 ( .A(n8069), .ZN(n10199) );
  INV_X1 U8024 ( .A(n8431), .ZN(n10204) );
  INV_X1 U8025 ( .A(n9870), .ZN(n6725) );
  NAND2_X1 U8026 ( .A1(n4743), .A2(n9691), .ZN(n9640) );
  XNOR2_X1 U8027 ( .A(n9636), .B(n9640), .ZN(n6472) );
  AND2_X1 U8028 ( .A1(n7985), .A2(n7392), .ZN(n6986) );
  NAND2_X1 U8029 ( .A1(n6472), .A2(n10099), .ZN(n9639) );
  AND2_X1 U8030 ( .A1(n6989), .A2(n6986), .ZN(n10158) );
  INV_X1 U8031 ( .A(n10158), .ZN(n10219) );
  AND2_X1 U8032 ( .A1(n6452), .A2(n6985), .ZN(n9834) );
  OAI21_X1 U8033 ( .B1(n10028), .B2(n6473), .A(n9834), .ZN(n9687) );
  OR2_X1 U8034 ( .A1(n6474), .A2(n9687), .ZN(n9855) );
  INV_X1 U8035 ( .A(n6475), .ZN(n6476) );
  NAND2_X1 U8036 ( .A1(n8216), .A2(P1_B_REG_SCAN_IN), .ZN(n6477) );
  MUX2_X1 U8037 ( .A(P1_B_REG_SCAN_IN), .B(n6477), .S(n8178), .Z(n6479) );
  INV_X1 U8038 ( .A(n8303), .ZN(n6478) );
  INV_X1 U8039 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8040 ( .A1(n9937), .A2(n6480), .ZN(n6481) );
  NAND2_X1 U8041 ( .A1(n8303), .A2(n8216), .ZN(n9938) );
  NAND2_X1 U8042 ( .A1(n6481), .A2(n9938), .ZN(n6708) );
  NAND2_X1 U8043 ( .A1(n10099), .A2(n6504), .ZN(n6722) );
  NAND2_X1 U8044 ( .A1(n6985), .A2(n6989), .ZN(n6977) );
  NAND2_X1 U8045 ( .A1(n6722), .A2(n6977), .ZN(n6482) );
  NOR2_X1 U8046 ( .A1(n9939), .A2(n6482), .ZN(n6493) );
  NOR4_X1 U8047 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6491) );
  NOR4_X1 U8048 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6490) );
  INV_X1 U8049 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10124) );
  INV_X1 U8050 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10126) );
  INV_X1 U8051 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10123) );
  INV_X1 U8052 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10125) );
  NAND4_X1 U8053 ( .A1(n10124), .A2(n10126), .A3(n10123), .A4(n10125), .ZN(
        n6488) );
  NOR4_X1 U8054 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6486) );
  NOR4_X1 U8055 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6485) );
  NOR4_X1 U8056 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6484) );
  NOR4_X1 U8057 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6483) );
  NAND4_X1 U8058 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n6487)
         );
  NOR4_X1 U8059 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6488), .A4(n6487), .ZN(n6489) );
  NAND3_X1 U8060 ( .A1(n6491), .A2(n6490), .A3(n6489), .ZN(n6492) );
  NAND2_X1 U8061 ( .A1(n9937), .A2(n6492), .ZN(n6978) );
  AND3_X1 U8062 ( .A1(n6708), .A2(n6493), .A3(n6978), .ZN(n9853) );
  INV_X1 U8063 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8064 ( .A1(n9937), .A2(n6494), .ZN(n6496) );
  NAND2_X1 U8065 ( .A1(n8303), .A2(n8178), .ZN(n6495) );
  AND2_X1 U8066 ( .A1(n6496), .A2(n6495), .ZN(n9940) );
  INV_X1 U8067 ( .A(n9940), .ZN(n6982) );
  AND2_X2 U8068 ( .A1(n9853), .A2(n6982), .ZN(n10226) );
  INV_X1 U8069 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6497) );
  OAI21_X1 U8070 ( .B1(n6989), .B2(n6499), .A(n7216), .ZN(n6500) );
  INV_X1 U8071 ( .A(n6500), .ZN(n6501) );
  NAND2_X4 U8072 ( .A1(n6501), .A2(n6775), .ZN(n6699) );
  OAI22_X1 U8073 ( .A1(n7273), .A2(n6699), .B1(n7334), .B2(n6503), .ZN(n6533)
         );
  INV_X1 U8074 ( .A(n6533), .ZN(n6535) );
  OR2_X1 U8075 ( .A1(n6504), .A2(n7985), .ZN(n6988) );
  AND2_X1 U8076 ( .A1(n6988), .A2(n6505), .ZN(n6506) );
  NAND2_X1 U8077 ( .A1(n6775), .A2(n6506), .ZN(n6507) );
  INV_X2 U8078 ( .A(n6511), .ZN(n6525) );
  OAI22_X1 U8079 ( .A1(n7273), .A2(n6503), .B1(n7334), .B2(n6525), .ZN(n6508)
         );
  XNOR2_X1 U8080 ( .A(n6508), .B(n6681), .ZN(n6532) );
  INV_X1 U8081 ( .A(n6532), .ZN(n6534) );
  OAI22_X1 U8082 ( .A1(n7213), .A2(n6503), .B1(n10143), .B2(n6525), .ZN(n6509)
         );
  XNOR2_X1 U8083 ( .A(n6509), .B(n6681), .ZN(n6523) );
  OAI22_X1 U8084 ( .A1(n7213), .A2(n6699), .B1(n10143), .B2(n6503), .ZN(n6522)
         );
  INV_X1 U8085 ( .A(n6775), .ZN(n6510) );
  AOI222_X1 U8086 ( .A1(n6991), .A2(n6675), .B1(n6976), .B2(n4510), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(n6510), .ZN(n6839) );
  INV_X1 U8087 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10227) );
  OAI21_X1 U8088 ( .B1(n6775), .B2(n10227), .A(n6513), .ZN(n6512) );
  AOI21_X1 U8089 ( .B1(n4510), .B2(n6991), .A(n6512), .ZN(n6840) );
  INV_X1 U8090 ( .A(n6513), .ZN(n6514) );
  OAI22_X1 U8091 ( .A1(n6839), .A2(n6840), .B1(n6514), .B2(n6681), .ZN(n6879)
         );
  OR2_X1 U8092 ( .A1(n10137), .A2(n6525), .ZN(n6516) );
  NAND2_X1 U8093 ( .A1(n5981), .A2(n4510), .ZN(n6515) );
  NAND2_X1 U8094 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  XNOR2_X1 U8095 ( .A(n6517), .B(n6702), .ZN(n6521) );
  NAND2_X1 U8096 ( .A1(n5981), .A2(n6675), .ZN(n6519) );
  OR2_X1 U8097 ( .A1(n10137), .A2(n6503), .ZN(n6518) );
  AND2_X1 U8098 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  NAND2_X1 U8099 ( .A1(n6521), .A2(n6520), .ZN(n6876) );
  NOR2_X1 U8100 ( .A1(n6521), .A2(n6520), .ZN(n6878) );
  AOI22_X1 U8101 ( .A1(n9512), .A2(n4510), .B1(n7219), .B2(n6704), .ZN(n6526)
         );
  INV_X1 U8102 ( .A(n6526), .ZN(n6527) );
  OAI22_X1 U8103 ( .A1(n8576), .A2(n6699), .B1(n10150), .B2(n6503), .ZN(n6529)
         );
  XNOR2_X1 U8104 ( .A(n6528), .B(n6529), .ZN(n7176) );
  NOR2_X1 U8105 ( .A1(n6530), .A2(n6529), .ZN(n6531) );
  XOR2_X1 U8106 ( .A(n6533), .B(n6532), .Z(n7225) );
  OAI22_X1 U8107 ( .A1(n7494), .A2(n6503), .B1(n10174), .B2(n6525), .ZN(n6536)
         );
  XNOR2_X1 U8108 ( .A(n6536), .B(n6681), .ZN(n6544) );
  OR2_X1 U8109 ( .A1(n7494), .A2(n6699), .ZN(n6538) );
  NAND2_X1 U8110 ( .A1(n10083), .A2(n4510), .ZN(n6537) );
  NAND2_X1 U8111 ( .A1(n6538), .A2(n6537), .ZN(n6543) );
  OAI22_X1 U8112 ( .A1(n7509), .A2(n6503), .B1(n10166), .B2(n6525), .ZN(n6539)
         );
  XNOR2_X1 U8113 ( .A(n6539), .B(n6681), .ZN(n7506) );
  OAI22_X1 U8114 ( .A1(n7509), .A2(n6699), .B1(n10166), .B2(n6503), .ZN(n7408)
         );
  AND2_X1 U8115 ( .A1(n7506), .A2(n7408), .ZN(n6540) );
  NOR2_X1 U8116 ( .A1(n7506), .A2(n7408), .ZN(n6542) );
  INV_X1 U8117 ( .A(n7502), .ZN(n6541) );
  NOR2_X1 U8118 ( .A1(n6544), .A2(n6543), .ZN(n7503) );
  INV_X1 U8119 ( .A(n7503), .ZN(n6545) );
  OAI22_X1 U8120 ( .A1(n9992), .A2(n6503), .B1(n10179), .B2(n6525), .ZN(n6549)
         );
  XNOR2_X1 U8121 ( .A(n6549), .B(n6681), .ZN(n6553) );
  INV_X1 U8122 ( .A(n6553), .ZN(n6555) );
  OR2_X1 U8123 ( .A1(n9992), .A2(n6699), .ZN(n6551) );
  NAND2_X1 U8124 ( .A1(n7499), .A2(n4510), .ZN(n6550) );
  NAND2_X1 U8125 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  INV_X1 U8126 ( .A(n6552), .ZN(n6554) );
  OAI21_X1 U8127 ( .B1(n6555), .B2(n6554), .A(n6556), .ZN(n7491) );
  AOI22_X1 U8128 ( .A1(n9508), .A2(n4510), .B1(n10067), .B2(n4508), .ZN(n6557)
         );
  XNOR2_X1 U8129 ( .A(n6557), .B(n6681), .ZN(n6559) );
  XNOR2_X1 U8130 ( .A(n6558), .B(n6559), .ZN(n9987) );
  AOI22_X1 U8131 ( .A1(n9508), .A2(n6675), .B1(n4510), .B2(n10067), .ZN(n9988)
         );
  NAND2_X1 U8132 ( .A1(n9987), .A2(n9988), .ZN(n9986) );
  NAND2_X1 U8133 ( .A1(n6560), .A2(n6559), .ZN(n9424) );
  NAND2_X1 U8134 ( .A1(n9430), .A2(n4508), .ZN(n6561) );
  OAI21_X1 U8135 ( .B1(n9990), .B2(n6503), .A(n6561), .ZN(n6562) );
  XNOR2_X1 U8136 ( .A(n6562), .B(n6702), .ZN(n6568) );
  OR2_X1 U8137 ( .A1(n9990), .A2(n6699), .ZN(n6564) );
  NAND2_X1 U8138 ( .A1(n9430), .A2(n4510), .ZN(n6563) );
  NAND2_X1 U8139 ( .A1(n6564), .A2(n6563), .ZN(n6566) );
  XNOR2_X1 U8140 ( .A(n6568), .B(n6566), .ZN(n9426) );
  INV_X1 U8142 ( .A(n6566), .ZN(n6567) );
  NAND2_X1 U8143 ( .A1(n8069), .A2(n4508), .ZN(n6571) );
  OR2_X1 U8144 ( .A1(n8428), .A2(n6503), .ZN(n6570) );
  NAND2_X1 U8145 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  XNOR2_X1 U8146 ( .A(n6572), .B(n6681), .ZN(n8416) );
  NAND2_X1 U8147 ( .A1(n8069), .A2(n4510), .ZN(n6574) );
  OR2_X1 U8148 ( .A1(n8428), .A2(n6699), .ZN(n6573) );
  NAND2_X1 U8149 ( .A1(n6574), .A2(n6573), .ZN(n8417) );
  NAND2_X1 U8150 ( .A1(n8431), .A2(n4508), .ZN(n6577) );
  OR2_X1 U8151 ( .A1(n8123), .A2(n6503), .ZN(n6576) );
  NAND2_X1 U8152 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  XNOR2_X1 U8153 ( .A(n6578), .B(n6702), .ZN(n6603) );
  NOR2_X1 U8154 ( .A1(n8123), .A2(n6699), .ZN(n6579) );
  AOI21_X1 U8155 ( .B1(n8431), .B2(n4510), .A(n6579), .ZN(n6602) );
  NOR2_X1 U8156 ( .A1(n6603), .A2(n6602), .ZN(n8418) );
  AOI21_X1 U8157 ( .B1(n8416), .B2(n8417), .A(n8418), .ZN(n8422) );
  NAND2_X1 U8158 ( .A1(n8528), .A2(n4508), .ZN(n6581) );
  OR2_X1 U8159 ( .A1(n8288), .A2(n6503), .ZN(n6580) );
  NAND2_X1 U8160 ( .A1(n6581), .A2(n6580), .ZN(n6582) );
  XNOR2_X1 U8161 ( .A(n6582), .B(n6681), .ZN(n6585) );
  INV_X1 U8162 ( .A(n6585), .ZN(n6583) );
  INV_X1 U8163 ( .A(n8288), .ZN(n9503) );
  AOI22_X1 U8164 ( .A1(n8528), .A2(n4510), .B1(n6675), .B2(n9503), .ZN(n6584)
         );
  NAND2_X1 U8165 ( .A1(n6583), .A2(n6584), .ZN(n6592) );
  INV_X1 U8166 ( .A(n6592), .ZN(n6586) );
  XNOR2_X1 U8167 ( .A(n6585), .B(n6584), .ZN(n8523) );
  INV_X1 U8168 ( .A(n6597), .ZN(n6594) );
  NAND2_X1 U8169 ( .A1(n8442), .A2(n4508), .ZN(n6588) );
  OR2_X1 U8170 ( .A1(n9504), .A2(n6503), .ZN(n6587) );
  NAND2_X1 U8171 ( .A1(n6588), .A2(n6587), .ZN(n6589) );
  XNOR2_X1 U8172 ( .A(n6589), .B(n6681), .ZN(n6595) );
  INV_X1 U8173 ( .A(n6595), .ZN(n6591) );
  OAI22_X1 U8174 ( .A1(n10213), .A2(n6503), .B1(n9504), .B2(n6699), .ZN(n6596)
         );
  INV_X1 U8175 ( .A(n6596), .ZN(n6590) );
  NAND2_X1 U8176 ( .A1(n6591), .A2(n6590), .ZN(n8520) );
  AND2_X1 U8177 ( .A1(n8520), .A2(n6592), .ZN(n6593) );
  INV_X1 U8178 ( .A(n6604), .ZN(n6599) );
  XOR2_X1 U8179 ( .A(n6596), .B(n6595), .Z(n8518) );
  AND2_X1 U8180 ( .A1(n8422), .A2(n6601), .ZN(n6600) );
  INV_X1 U8181 ( .A(n6601), .ZN(n6606) );
  NAND2_X1 U8182 ( .A1(n6603), .A2(n6602), .ZN(n8434) );
  AND2_X1 U8183 ( .A1(n8434), .A2(n6604), .ZN(n6605) );
  AOI22_X1 U8184 ( .A1(n9920), .A2(n4508), .B1(n4510), .B2(n9502), .ZN(n6607)
         );
  XNOR2_X1 U8185 ( .A(n6607), .B(n6681), .ZN(n8391) );
  INV_X1 U8186 ( .A(n8391), .ZN(n6612) );
  AOI22_X1 U8187 ( .A1(n9920), .A2(n4510), .B1(n6675), .B2(n9502), .ZN(n8390)
         );
  OAI21_X1 U8188 ( .B1(n6610), .B2(n8391), .A(n8390), .ZN(n6611) );
  OAI21_X1 U8189 ( .B1(n8389), .B2(n6612), .A(n6611), .ZN(n6613) );
  INV_X1 U8190 ( .A(n6613), .ZN(n9479) );
  AOI22_X1 U8191 ( .A1(n9916), .A2(n4508), .B1(n4510), .B2(n9501), .ZN(n6614)
         );
  XNOR2_X1 U8192 ( .A(n6614), .B(n6681), .ZN(n9481) );
  INV_X1 U8193 ( .A(n9481), .ZN(n6616) );
  NAND2_X1 U8194 ( .A1(n9479), .A2(n6616), .ZN(n6615) );
  AOI22_X1 U8195 ( .A1(n9916), .A2(n4510), .B1(n6675), .B2(n9501), .ZN(n9480)
         );
  NAND2_X1 U8196 ( .A1(n6615), .A2(n9480), .ZN(n6618) );
  NAND2_X1 U8197 ( .A1(n9483), .A2(n9481), .ZN(n6617) );
  NAND2_X1 U8198 ( .A1(n6618), .A2(n6617), .ZN(n9389) );
  INV_X1 U8199 ( .A(n9486), .ZN(n9500) );
  AOI22_X1 U8200 ( .A1(n9398), .A2(n4508), .B1(n4510), .B2(n9500), .ZN(n6619)
         );
  XOR2_X1 U8201 ( .A(n6681), .B(n6619), .Z(n6620) );
  OAI22_X1 U8202 ( .A1(n9972), .A2(n6503), .B1(n9486), .B2(n6699), .ZN(n6621)
         );
  NAND2_X1 U8203 ( .A1(n6620), .A2(n6621), .ZN(n9391) );
  INV_X1 U8204 ( .A(n6620), .ZN(n6623) );
  INV_X1 U8205 ( .A(n6621), .ZN(n6622) );
  NAND2_X1 U8206 ( .A1(n6623), .A2(n6622), .ZN(n9390) );
  NAND2_X1 U8207 ( .A1(n9911), .A2(n4508), .ZN(n6625) );
  NAND2_X1 U8208 ( .A1(n9499), .A2(n4510), .ZN(n6624) );
  NAND2_X1 U8209 ( .A1(n6625), .A2(n6624), .ZN(n6626) );
  XNOR2_X1 U8210 ( .A(n6626), .B(n6681), .ZN(n6629) );
  NAND2_X1 U8211 ( .A1(n9911), .A2(n4510), .ZN(n6628) );
  NAND2_X1 U8212 ( .A1(n9499), .A2(n6675), .ZN(n6627) );
  NAND2_X1 U8213 ( .A1(n6628), .A2(n6627), .ZN(n6630) );
  NAND2_X1 U8214 ( .A1(n6629), .A2(n6630), .ZN(n9405) );
  INV_X1 U8215 ( .A(n6629), .ZN(n6632) );
  INV_X1 U8216 ( .A(n6630), .ZN(n6631) );
  NAND2_X1 U8217 ( .A1(n6632), .A2(n6631), .ZN(n9404) );
  AOI22_X1 U8218 ( .A1(n9645), .A2(n4508), .B1(n4510), .B2(n9646), .ZN(n6633)
         );
  XNOR2_X1 U8219 ( .A(n6633), .B(n6681), .ZN(n6635) );
  NAND2_X1 U8220 ( .A1(n6634), .A2(n6635), .ZN(n9455) );
  OAI22_X1 U8221 ( .A1(n9966), .A2(n6503), .B1(n9837), .B2(n6699), .ZN(n9458)
         );
  INV_X1 U8222 ( .A(n6634), .ZN(n6637) );
  INV_X1 U8223 ( .A(n6635), .ZN(n6636) );
  OAI22_X1 U8224 ( .A1(n9961), .A2(n6503), .B1(n9649), .B2(n6699), .ZN(n6641)
         );
  AOI22_X1 U8225 ( .A1(n9850), .A2(n4508), .B1(n4510), .B2(n9648), .ZN(n6638)
         );
  XNOR2_X1 U8226 ( .A(n6638), .B(n6681), .ZN(n6639) );
  XOR2_X1 U8227 ( .A(n6641), .B(n6639), .Z(n9366) );
  INV_X1 U8228 ( .A(n6639), .ZN(n6640) );
  NAND2_X1 U8229 ( .A1(n9824), .A2(n4508), .ZN(n6643) );
  NAND2_X1 U8230 ( .A1(n9835), .A2(n4510), .ZN(n6642) );
  NAND2_X1 U8231 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  XNOR2_X1 U8232 ( .A(n6644), .B(n6681), .ZN(n9437) );
  NAND2_X1 U8233 ( .A1(n9824), .A2(n4510), .ZN(n6646) );
  NAND2_X1 U8234 ( .A1(n9835), .A2(n6675), .ZN(n6645) );
  NAND2_X1 U8235 ( .A1(n6646), .A2(n6645), .ZN(n9436) );
  NOR2_X1 U8236 ( .A1(n9437), .A2(n9436), .ZN(n6648) );
  NAND2_X1 U8237 ( .A1(n9437), .A2(n9436), .ZN(n6647) );
  AND2_X1 U8238 ( .A1(n9795), .A2(n6675), .ZN(n6649) );
  AOI21_X1 U8239 ( .B1(n9906), .B2(n4510), .A(n6649), .ZN(n6652) );
  AOI22_X1 U8240 ( .A1(n9906), .A2(n4508), .B1(n4510), .B2(n9795), .ZN(n6650)
         );
  XNOR2_X1 U8241 ( .A(n6650), .B(n6681), .ZN(n6651) );
  XOR2_X1 U8242 ( .A(n6652), .B(n6651), .Z(n9374) );
  NAND2_X1 U8243 ( .A1(n9373), .A2(n9374), .ZN(n6656) );
  INV_X1 U8244 ( .A(n6651), .ZN(n6654) );
  INV_X1 U8245 ( .A(n6652), .ZN(n6653) );
  NAND2_X1 U8246 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  NAND2_X1 U8247 ( .A1(n6656), .A2(n6655), .ZN(n9448) );
  AOI22_X1 U8248 ( .A1(n9900), .A2(n4508), .B1(n4510), .B2(n9654), .ZN(n6657)
         );
  XOR2_X1 U8249 ( .A(n6681), .B(n6657), .Z(n6658) );
  OAI22_X1 U8250 ( .A1(n9790), .A2(n6503), .B1(n9808), .B2(n6699), .ZN(n9445)
         );
  OAI21_X2 U8251 ( .B1(n9448), .B2(n6658), .A(n9445), .ZN(n6660) );
  INV_X1 U8252 ( .A(n6658), .ZN(n9446) );
  AOI22_X1 U8253 ( .A1(n9774), .A2(n4508), .B1(n4510), .B2(n9796), .ZN(n6661)
         );
  XNOR2_X1 U8254 ( .A(n6661), .B(n6681), .ZN(n6663) );
  AOI22_X1 U8255 ( .A1(n9774), .A2(n4510), .B1(n6675), .B2(n9796), .ZN(n6662)
         );
  NAND2_X1 U8256 ( .A1(n6663), .A2(n6662), .ZN(n9416) );
  OAI21_X1 U8257 ( .B1(n6663), .B2(n6662), .A(n9416), .ZN(n8587) );
  OAI22_X1 U8258 ( .A1(n9770), .A2(n6525), .B1(n9747), .B2(n6503), .ZN(n6664)
         );
  XNOR2_X1 U8259 ( .A(n6664), .B(n6702), .ZN(n6667) );
  OR2_X1 U8260 ( .A1(n9770), .A2(n6503), .ZN(n6666) );
  OR2_X1 U8261 ( .A1(n9747), .A2(n6699), .ZN(n6665) );
  NAND2_X1 U8262 ( .A1(n6667), .A2(n6668), .ZN(n6676) );
  INV_X1 U8263 ( .A(n6667), .ZN(n6670) );
  INV_X1 U8264 ( .A(n6668), .ZN(n6669) );
  NAND2_X1 U8265 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  NAND2_X1 U8266 ( .A1(n6676), .A2(n6671), .ZN(n9415) );
  OR2_X1 U8267 ( .A1(n8587), .A2(n9415), .ZN(n9380) );
  NAND2_X1 U8268 ( .A1(n9884), .A2(n4508), .ZN(n6673) );
  NAND2_X1 U8269 ( .A1(n9661), .A2(n4510), .ZN(n6672) );
  NAND2_X1 U8270 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  XNOR2_X1 U8271 ( .A(n6674), .B(n6681), .ZN(n6683) );
  AOI22_X1 U8272 ( .A1(n9884), .A2(n4510), .B1(n6675), .B2(n9661), .ZN(n6684)
         );
  XNOR2_X1 U8273 ( .A(n6683), .B(n6684), .ZN(n9383) );
  INV_X1 U8274 ( .A(n9383), .ZN(n6677) );
  OR2_X1 U8275 ( .A1(n9415), .A2(n9416), .ZN(n9413) );
  AND2_X1 U8276 ( .A1(n9413), .A2(n6676), .ZN(n9381) );
  OR2_X1 U8277 ( .A1(n9748), .A2(n6699), .ZN(n6679) );
  NAND2_X1 U8278 ( .A1(n6680), .A2(n6679), .ZN(n6694) );
  OAI22_X1 U8279 ( .A1(n9739), .A2(n6525), .B1(n9748), .B2(n6503), .ZN(n6682)
         );
  XNOR2_X1 U8280 ( .A(n6682), .B(n6681), .ZN(n6695) );
  XOR2_X1 U8281 ( .A(n6694), .B(n6695), .Z(n9470) );
  INV_X1 U8282 ( .A(n6683), .ZN(n6685) );
  NAND2_X1 U8283 ( .A1(n6685), .A2(n6684), .ZN(n9467) );
  NAND2_X1 U8284 ( .A1(n9874), .A2(n4508), .ZN(n6687) );
  OR2_X1 U8285 ( .A1(n9732), .A2(n6503), .ZN(n6686) );
  NAND2_X1 U8286 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  XNOR2_X1 U8287 ( .A(n6688), .B(n6702), .ZN(n6691) );
  INV_X1 U8288 ( .A(n6691), .ZN(n6693) );
  NOR2_X1 U8289 ( .A1(n9732), .A2(n6699), .ZN(n6689) );
  AOI21_X1 U8290 ( .B1(n9874), .B2(n4510), .A(n6689), .ZN(n6690) );
  INV_X1 U8291 ( .A(n6690), .ZN(n6692) );
  AOI21_X1 U8292 ( .B1(n6693), .B2(n6692), .A(n6713), .ZN(n9357) );
  INV_X1 U8293 ( .A(n9357), .ZN(n6697) );
  NAND2_X1 U8294 ( .A1(n6695), .A2(n6694), .ZN(n9358) );
  INV_X1 U8295 ( .A(n9358), .ZN(n6696) );
  NOR2_X1 U8296 ( .A1(n6697), .A2(n6696), .ZN(n6698) );
  NAND2_X1 U8297 ( .A1(n9870), .A2(n4510), .ZN(n6701) );
  OR2_X1 U8298 ( .A1(n9721), .A2(n6699), .ZN(n6700) );
  NAND2_X1 U8299 ( .A1(n6701), .A2(n6700), .ZN(n6703) );
  XNOR2_X1 U8300 ( .A(n6703), .B(n6702), .ZN(n6707) );
  NAND2_X1 U8301 ( .A1(n9870), .A2(n4508), .ZN(n6705) );
  OAI21_X1 U8302 ( .B1(n9721), .B2(n6503), .A(n6705), .ZN(n6706) );
  XNOR2_X1 U8303 ( .A(n6707), .B(n6706), .ZN(n6714) );
  INV_X1 U8304 ( .A(n6714), .ZN(n6711) );
  INV_X1 U8305 ( .A(n6708), .ZN(n6981) );
  NAND3_X1 U8306 ( .A1(n6981), .A2(n9940), .A3(n6978), .ZN(n6715) );
  NOR2_X1 U8307 ( .A1(n6715), .A2(n9939), .ZN(n6721) );
  NOR2_X1 U8308 ( .A1(n10158), .A2(n6985), .ZN(n6709) );
  NOR2_X1 U8309 ( .A1(n6713), .A2(n9494), .ZN(n6710) );
  NAND3_X1 U8310 ( .A1(n9359), .A2(n10000), .A3(n6714), .ZN(n6731) );
  NAND2_X1 U8311 ( .A1(n6715), .A2(n6722), .ZN(n6717) );
  AND3_X1 U8312 ( .A1(n6775), .A2(n6776), .A3(n6977), .ZN(n6716) );
  NAND2_X1 U8313 ( .A1(n6717), .A2(n6716), .ZN(n6841) );
  NAND2_X1 U8314 ( .A1(n6841), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10003) );
  INV_X1 U8315 ( .A(n10003), .ZN(n9472) );
  OR2_X1 U8316 ( .A1(n9732), .A2(n9991), .ZN(n6719) );
  OR2_X1 U8317 ( .A1(n7234), .A2(n9989), .ZN(n6718) );
  AND2_X1 U8318 ( .A1(n6719), .A2(n6718), .ZN(n9704) );
  INV_X1 U8319 ( .A(n6989), .ZN(n6984) );
  AND2_X1 U8320 ( .A1(n6721), .A2(n6984), .ZN(n9996) );
  INV_X1 U8321 ( .A(n9996), .ZN(n9439) );
  OAI22_X1 U8322 ( .A1(n9704), .A2(n9439), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6720), .ZN(n6727) );
  NAND2_X1 U8323 ( .A1(n6986), .A2(n9857), .ZN(n10110) );
  INV_X1 U8324 ( .A(n10110), .ZN(n6999) );
  NAND2_X1 U8325 ( .A1(n6721), .A2(n6999), .ZN(n6724) );
  INV_X1 U8326 ( .A(n9939), .ZN(n6979) );
  INV_X1 U8327 ( .A(n6722), .ZN(n6723) );
  NAND2_X1 U8328 ( .A1(n6979), .A2(n6723), .ZN(n10108) );
  NAND2_X1 U8329 ( .A1(n6724), .A2(n10108), .ZN(n9492) );
  INV_X1 U8330 ( .A(n9492), .ZN(n9998) );
  NOR2_X1 U8331 ( .A1(n6725), .A2(n9998), .ZN(n6726) );
  AOI211_X1 U8332 ( .C1(n9472), .C2(n9709), .A(n6727), .B(n6726), .ZN(n6728)
         );
  INV_X1 U8333 ( .A(n6728), .ZN(n6729) );
  NAND3_X1 U8334 ( .A1(n6732), .A2(n6731), .A3(n6730), .ZN(P1_U3220) );
  INV_X1 U8335 ( .A(n6733), .ZN(n6734) );
  OR2_X1 U8336 ( .A1(n6734), .A2(n6775), .ZN(n7233) );
  NAND2_X1 U8337 ( .A1(n8748), .A2(n6921), .ZN(n6735) );
  NAND2_X1 U8338 ( .A1(n6735), .A2(n6920), .ZN(n6855) );
  NAND2_X1 U8339 ( .A1(n6855), .A2(n6736), .ZN(n6737) );
  NAND2_X1 U8340 ( .A1(n6737), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8341 ( .A(n6764), .ZN(n6758) );
  OR2_X2 U8342 ( .A1(n6921), .A2(n6758), .ZN(n8972) );
  INV_X1 U8343 ( .A(n8972), .ZN(P2_U3893) );
  AND2_X1 U8344 ( .A1(n6738), .A2(P1_U3086), .ZN(n8064) );
  INV_X2 U8345 ( .A(n8064), .ZN(n9949) );
  INV_X1 U8346 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6739) );
  NOR2_X1 U8347 ( .A1(n6738), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9945) );
  INV_X1 U8348 ( .A(n9945), .ZN(n9952) );
  OAI222_X1 U8349 ( .A1(P1_U3086), .A2(n6804), .B1(n9949), .B2(n6745), .C1(
        n6739), .C2(n9952), .ZN(P1_U3354) );
  INV_X1 U8350 ( .A(n10027), .ZN(n6805) );
  INV_X1 U8351 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6740) );
  OAI222_X1 U8352 ( .A1(P1_U3086), .A2(n6805), .B1(n9949), .B2(n6748), .C1(
        n6740), .C2(n9952), .ZN(P1_U3353) );
  INV_X1 U8353 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6741) );
  INV_X1 U8354 ( .A(n6801), .ZN(n9515) );
  OAI222_X1 U8355 ( .A1(n9952), .A2(n6741), .B1(n9949), .B2(n6746), .C1(
        P1_U3086), .C2(n9515), .ZN(P1_U3352) );
  AOI22_X1 U8356 ( .A1(n9945), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10050), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6742) );
  OAI21_X1 U8357 ( .B1(n6750), .B2(n9949), .A(n6742), .ZN(P1_U3351) );
  NAND2_X1 U8358 ( .A1(n6743), .A2(P2_U3151), .ZN(n7286) );
  AND2_X1 U8359 ( .A1(n6744), .A2(P2_U3151), .ZN(n9352) );
  INV_X1 U8360 ( .A(n9352), .ZN(n8849) );
  OAI222_X1 U8361 ( .A1(n6884), .A2(P2_U3151), .B1(n7286), .B2(n6745), .C1(
        n5139), .C2(n8849), .ZN(P2_U3294) );
  CLKBUF_X1 U8362 ( .A(n7286), .Z(n9355) );
  OAI222_X1 U8363 ( .A1(n10286), .A2(P2_U3151), .B1(n9355), .B2(n6746), .C1(
        n5178), .C2(n8849), .ZN(P2_U3292) );
  INV_X1 U8364 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6747) );
  OAI222_X1 U8365 ( .A1(n10256), .A2(P2_U3151), .B1(n9355), .B2(n6748), .C1(
        n6747), .C2(n8849), .ZN(P2_U3293) );
  INV_X1 U8366 ( .A(n7029), .ZN(n7008) );
  INV_X1 U8367 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6749) );
  OAI222_X1 U8368 ( .A1(n7008), .A2(P2_U3151), .B1(n9355), .B2(n6750), .C1(
        n6749), .C2(n8849), .ZN(P2_U3291) );
  AOI22_X1 U8369 ( .A1(n9535), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9945), .ZN(n6751) );
  OAI21_X1 U8370 ( .B1(n6753), .B2(n9949), .A(n6751), .ZN(P1_U3350) );
  INV_X1 U8371 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6752) );
  OAI222_X1 U8372 ( .A1(n7118), .A2(P2_U3151), .B1(n7286), .B2(n6753), .C1(
        n6752), .C2(n8849), .ZN(P2_U3290) );
  INV_X1 U8373 ( .A(n7036), .ZN(n10311) );
  INV_X1 U8374 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6754) );
  OAI222_X1 U8375 ( .A1(n10311), .A2(P2_U3151), .B1(n7286), .B2(n6755), .C1(
        n6754), .C2(n8849), .ZN(P2_U3289) );
  INV_X1 U8376 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6756) );
  INV_X1 U8377 ( .A(n6822), .ZN(n6825) );
  OAI222_X1 U8378 ( .A1(n9952), .A2(n6756), .B1(n9949), .B2(n6755), .C1(
        P1_U3086), .C2(n6825), .ZN(P1_U3349) );
  NAND2_X1 U8379 ( .A1(n6757), .A2(n5772), .ZN(n6766) );
  INV_X1 U8380 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U8381 ( .A1(n6758), .A2(n8243), .ZN(n6760) );
  AOI22_X1 U8382 ( .A1(n6766), .A2(n6761), .B1(n6760), .B2(n6759), .ZN(
        P2_U3377) );
  INV_X1 U8383 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6765) );
  INV_X1 U8384 ( .A(n6762), .ZN(n6763) );
  AOI22_X1 U8385 ( .A1(n6766), .A2(n6765), .B1(n6764), .B2(n6763), .ZN(
        P2_U3376) );
  AND2_X1 U8386 ( .A1(n6766), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8387 ( .A1(n6766), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8388 ( .A1(n6766), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8389 ( .A1(n6766), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8390 ( .A1(n6766), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8391 ( .A1(n6766), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8392 ( .A1(n6766), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8393 ( .A1(n6766), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8394 ( .A1(n6766), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8395 ( .A1(n6766), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8396 ( .A1(n6766), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8397 ( .A1(n6766), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8398 ( .A1(n6766), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8399 ( .A1(n6766), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8400 ( .A1(n6766), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8401 ( .A1(n6766), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8402 ( .A1(n6766), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8403 ( .A1(n6766), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8404 ( .A1(n6766), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8405 ( .A1(n6766), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8406 ( .A1(n6766), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8407 ( .A1(n6766), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8408 ( .A1(n6766), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8409 ( .A1(n6766), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8410 ( .A1(n6766), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8411 ( .A1(n6766), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8412 ( .A1(n6766), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8413 ( .A1(n6766), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8414 ( .A1(n6766), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8415 ( .A1(n6766), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  INV_X1 U8416 ( .A(n6767), .ZN(n6770) );
  INV_X1 U8417 ( .A(n7043), .ZN(n7052) );
  OAI222_X1 U8418 ( .A1(n9952), .A2(n6768), .B1(n9949), .B2(n6770), .C1(
        P1_U3086), .C2(n7052), .ZN(P1_U3348) );
  INV_X1 U8419 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6769) );
  OAI222_X1 U8420 ( .A1(n4706), .A2(P2_U3151), .B1(n7286), .B2(n6770), .C1(
        n6769), .C2(n8849), .ZN(P2_U3288) );
  INV_X1 U8421 ( .A(n6771), .ZN(n6773) );
  OAI222_X1 U8422 ( .A1(n9952), .A2(n7772), .B1(n9949), .B2(n6773), .C1(
        P1_U3086), .C2(n4645), .ZN(P1_U3347) );
  OAI222_X1 U8423 ( .A1(n7459), .A2(P2_U3151), .B1(n7286), .B2(n6773), .C1(
        n6772), .C2(n8849), .ZN(P2_U3287) );
  INV_X1 U8424 ( .A(n6776), .ZN(n6774) );
  OAI21_X1 U8425 ( .B1(n6775), .B2(n6774), .A(P1_STATE_REG_SCAN_IN), .ZN(n6787) );
  INV_X1 U8426 ( .A(n6787), .ZN(n6778) );
  NAND2_X1 U8427 ( .A1(n6776), .A2(n6985), .ZN(n6777) );
  NAND2_X1 U8428 ( .A1(n5980), .A2(n6777), .ZN(n6788) );
  NOR2_X1 U8429 ( .A1(n10049), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8430 ( .A(n6069), .ZN(n6780) );
  INV_X1 U8431 ( .A(n7295), .ZN(n7049) );
  OAI222_X1 U8432 ( .A1(n9952), .A2(n7881), .B1(n9949), .B2(n6780), .C1(n7049), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8433 ( .A(n7468), .ZN(n7525) );
  OAI222_X1 U8434 ( .A1(P2_U3151), .A2(n7525), .B1(n7286), .B2(n6780), .C1(
        n6779), .C2(n8849), .ZN(P2_U3286) );
  INV_X1 U8435 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7767) );
  INV_X1 U8436 ( .A(n6781), .ZN(n6784) );
  INV_X1 U8437 ( .A(n7359), .ZN(n6782) );
  OAI222_X1 U8438 ( .A1(n9952), .A2(n7767), .B1(n9949), .B2(n6784), .C1(n6782), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8439 ( .A(n8044), .ZN(n8041) );
  INV_X1 U8440 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6783) );
  OAI222_X1 U8441 ( .A1(P2_U3151), .A2(n8041), .B1(n7286), .B2(n6784), .C1(
        n6783), .C2(n8849), .ZN(P2_U3285) );
  INV_X1 U8442 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8443 ( .A1(n6991), .A2(P1_U3973), .ZN(n6785) );
  OAI21_X1 U8444 ( .B1(P1_U3973), .B2(n6786), .A(n6785), .ZN(P1_U3554) );
  OR2_X1 U8445 ( .A1(n6788), .A2(n6787), .ZN(n10008) );
  INV_X1 U8446 ( .A(n10008), .ZN(n6799) );
  NAND2_X1 U8447 ( .A1(n6799), .A2(n6452), .ZN(n9629) );
  INV_X1 U8448 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6789) );
  MUX2_X1 U8449 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6789), .S(n10050), .Z(n10045) );
  INV_X1 U8450 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6790) );
  INV_X1 U8451 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10015) );
  INV_X1 U8452 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U8453 ( .A1(n10015), .A2(n10120), .ZN(n10030) );
  INV_X1 U8454 ( .A(n10030), .ZN(n10011) );
  AOI21_X1 U8455 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n10014), .A(n10010), .ZN(
        n10024) );
  INV_X1 U8456 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U8457 ( .A1(n10027), .A2(n6791), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n6805), .ZN(n10025) );
  NOR2_X1 U8458 ( .A1(n10024), .A2(n10025), .ZN(n10023) );
  INV_X1 U8459 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6792) );
  AOI22_X1 U8460 ( .A1(n6801), .A2(n6792), .B1(P1_REG2_REG_3__SCAN_IN), .B2(
        n9515), .ZN(n9519) );
  NAND2_X1 U8461 ( .A1(n10050), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U8462 ( .A1(n10042), .A2(n6793), .ZN(n9529) );
  INV_X1 U8463 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6794) );
  XNOR2_X1 U8464 ( .A(n9535), .B(n6794), .ZN(n9530) );
  NAND2_X1 U8465 ( .A1(n9529), .A2(n9530), .ZN(n9528) );
  NAND2_X1 U8466 ( .A1(n9535), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6795) );
  XNOR2_X1 U8467 ( .A(n6822), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U8468 ( .A1(n6452), .A2(n10028), .ZN(n6796) );
  NAND2_X1 U8469 ( .A1(n6799), .A2(n6796), .ZN(n10022) );
  AOI211_X1 U8470 ( .C1(n6798), .C2(n6797), .A(n6821), .B(n10022), .ZN(n6813)
         );
  NAND2_X1 U8471 ( .A1(n6799), .A2(n10028), .ZN(n9631) );
  INV_X1 U8472 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6800) );
  MUX2_X1 U8473 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6800), .S(n10050), .Z(n10054) );
  NAND2_X1 U8474 ( .A1(n6801), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6806) );
  INV_X1 U8475 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6802) );
  MUX2_X1 U8476 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6802), .S(n6801), .Z(n9523)
         );
  MUX2_X1 U8477 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6803), .S(n10027), .Z(n10036) );
  INV_X1 U8478 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10229) );
  MUX2_X1 U8479 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10229), .S(n10014), .Z(
        n10017) );
  NAND3_X1 U8480 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n10017), .ZN(n10016) );
  OAI21_X1 U8481 ( .B1(n6804), .B2(n10229), .A(n10016), .ZN(n10037) );
  NAND2_X1 U8482 ( .A1(n10036), .A2(n10037), .ZN(n10035) );
  OAI21_X1 U8483 ( .B1(n6805), .B2(n6803), .A(n10035), .ZN(n9524) );
  NAND2_X1 U8484 ( .A1(n9523), .A2(n9524), .ZN(n9522) );
  NAND2_X1 U8485 ( .A1(n6806), .A2(n9522), .ZN(n10055) );
  NAND2_X1 U8486 ( .A1(n10054), .A2(n10055), .ZN(n10052) );
  NAND2_X1 U8487 ( .A1(n10050), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6807) );
  NAND2_X1 U8488 ( .A1(n10052), .A2(n6807), .ZN(n9532) );
  INV_X1 U8489 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6808) );
  MUX2_X1 U8490 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6808), .S(n9535), .Z(n9533)
         );
  NAND2_X1 U8491 ( .A1(n9532), .A2(n9533), .ZN(n9531) );
  NAND2_X1 U8492 ( .A1(n9535), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6810) );
  INV_X1 U8493 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10235) );
  MUX2_X1 U8494 ( .A(n10235), .B(P1_REG1_REG_6__SCAN_IN), .S(n6822), .Z(n6809)
         );
  AOI21_X1 U8495 ( .B1(n9531), .B2(n6810), .A(n6809), .ZN(n6828) );
  AND3_X1 U8496 ( .A1(n9531), .A2(n6810), .A3(n6809), .ZN(n6811) );
  NOR3_X1 U8497 ( .A1(n9631), .A2(n6828), .A3(n6811), .ZN(n6812) );
  NOR2_X1 U8498 ( .A1(n6813), .A2(n6812), .ZN(n6816) );
  AND2_X1 U8499 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6814) );
  AOI21_X1 U8500 ( .B1(n10049), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6814), .ZN(
        n6815) );
  OAI211_X1 U8501 ( .C1(n6825), .C2(n9629), .A(n6816), .B(n6815), .ZN(P1_U3249) );
  INV_X1 U8502 ( .A(n8147), .ZN(n8139) );
  INV_X1 U8503 ( .A(n6817), .ZN(n6819) );
  OAI222_X1 U8504 ( .A1(n8139), .A2(P2_U3151), .B1(n7286), .B2(n6819), .C1(
        n6818), .C2(n8849), .ZN(P2_U3284) );
  INV_X1 U8505 ( .A(n7443), .ZN(n7449) );
  OAI222_X1 U8506 ( .A1(n9952), .A2(n6820), .B1(n9949), .B2(n6819), .C1(
        P1_U3086), .C2(n7449), .ZN(P1_U3344) );
  XNOR2_X1 U8507 ( .A(n7043), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6823) );
  NOR2_X1 U8508 ( .A1(n6824), .A2(n6823), .ZN(n7042) );
  AOI211_X1 U8509 ( .C1(n6824), .C2(n6823), .A(n7042), .B(n10022), .ZN(n6832)
         );
  NOR2_X1 U8510 ( .A1(n6825), .A2(n10235), .ZN(n6827) );
  INV_X1 U8511 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7053) );
  MUX2_X1 U8512 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7053), .S(n7043), .Z(n6826)
         );
  OAI21_X1 U8513 ( .B1(n6828), .B2(n6827), .A(n6826), .ZN(n7051) );
  INV_X1 U8514 ( .A(n7051), .ZN(n6830) );
  NOR3_X1 U8515 ( .A1(n6828), .A2(n6827), .A3(n6826), .ZN(n6829) );
  NOR3_X1 U8516 ( .A1(n9631), .A2(n6830), .A3(n6829), .ZN(n6831) );
  NOR2_X1 U8517 ( .A1(n6832), .A2(n6831), .ZN(n6835) );
  NAND2_X1 U8518 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7495) );
  INV_X1 U8519 ( .A(n7495), .ZN(n6833) );
  AOI21_X1 U8520 ( .B1(n10049), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6833), .ZN(
        n6834) );
  OAI211_X1 U8521 ( .C1(n7052), .C2(n9629), .A(n6835), .B(n6834), .ZN(P1_U3250) );
  INV_X1 U8522 ( .A(n8157), .ZN(n8197) );
  INV_X1 U8523 ( .A(n6836), .ZN(n6838) );
  INV_X1 U8524 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6837) );
  OAI222_X1 U8525 ( .A1(P2_U3151), .A2(n8197), .B1(n9355), .B2(n6838), .C1(
        n6837), .C2(n8849), .ZN(P2_U3283) );
  INV_X1 U8526 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7880) );
  INV_X1 U8527 ( .A(n8107), .ZN(n7458) );
  OAI222_X1 U8528 ( .A1(n9952), .A2(n7880), .B1(n9949), .B2(n6838), .C1(n7458), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  XNOR2_X1 U8529 ( .A(n6839), .B(n6840), .ZN(n10029) );
  NOR2_X1 U8530 ( .A1(n8577), .A2(n9989), .ZN(n10131) );
  OR2_X1 U8531 ( .A1(n6841), .A2(P1_U3086), .ZN(n8578) );
  AOI22_X1 U8532 ( .A1(n10131), .A2(n9996), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8578), .ZN(n6843) );
  NAND2_X1 U8533 ( .A1(n9492), .A2(n6976), .ZN(n6842) );
  OAI211_X1 U8534 ( .C1(n10029), .C2(n9494), .A(n6843), .B(n6842), .ZN(
        P1_U3232) );
  INV_X1 U8535 ( .A(n8582), .ZN(n7107) );
  NAND2_X1 U8536 ( .A1(n10353), .A2(n5741), .ZN(n10414) );
  NOR2_X1 U8537 ( .A1(n6844), .A2(n8582), .ZN(n8609) );
  INV_X1 U8538 ( .A(n8609), .ZN(n8614) );
  NAND2_X1 U8539 ( .A1(n8614), .A2(n8612), .ZN(n8765) );
  OAI21_X1 U8540 ( .B1(n10350), .B2(n10414), .A(n8765), .ZN(n6846) );
  NOR2_X1 U8541 ( .A1(n5692), .A2(n10346), .ZN(n7102) );
  INV_X1 U8542 ( .A(n7102), .ZN(n6845) );
  OAI211_X1 U8543 ( .C1(n7107), .C2(n10390), .A(n6846), .B(n6845), .ZN(n6850)
         );
  NAND2_X1 U8544 ( .A1(n6850), .A2(n10440), .ZN(n6847) );
  OAI21_X1 U8545 ( .B1(n10440), .B2(n4668), .A(n6847), .ZN(P2_U3459) );
  INV_X1 U8546 ( .A(n6848), .ZN(n6853) );
  AOI22_X1 U8547 ( .A1(n8258), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9945), .ZN(n6849) );
  OAI21_X1 U8548 ( .B1(n6853), .B2(n9949), .A(n6849), .ZN(P1_U3342) );
  NAND2_X1 U8549 ( .A1(n10421), .A2(n6850), .ZN(n6851) );
  OAI21_X1 U8550 ( .B1(n10421), .B2(n5144), .A(n6851), .ZN(P2_U3390) );
  INV_X1 U8551 ( .A(n8364), .ZN(n8374) );
  INV_X1 U8552 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6852) );
  OAI222_X1 U8553 ( .A1(n8374), .A2(P2_U3151), .B1(n9355), .B2(n6853), .C1(
        n6852), .C2(n8849), .ZN(P2_U3282) );
  NOR2_X1 U8554 ( .A1(n8049), .A2(P2_U3151), .ZN(n8322) );
  NAND2_X1 U8555 ( .A1(n6855), .A2(n8322), .ZN(n6854) );
  MUX2_X1 U8556 ( .A(n8972), .B(n6854), .S(n5680), .Z(n10312) );
  NOR2_X1 U8557 ( .A1(n5680), .A2(P2_U3151), .ZN(n8361) );
  AND2_X1 U8558 ( .A1(n6855), .A2(n8361), .ZN(n10252) );
  INV_X1 U8559 ( .A(n10252), .ZN(n6856) );
  OR2_X1 U8560 ( .A1(n6856), .A2(n8799), .ZN(n10283) );
  INV_X1 U8561 ( .A(n10283), .ZN(n10303) );
  INV_X1 U8562 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10255) );
  AND2_X1 U8563 ( .A1(n10255), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6857) );
  OAI21_X1 U8564 ( .B1(n6884), .B2(n6857), .A(n6894), .ZN(n6858) );
  NAND2_X1 U8565 ( .A1(n6858), .A2(n5131), .ZN(n6859) );
  NAND2_X1 U8566 ( .A1(n6895), .A2(n6859), .ZN(n6870) );
  INV_X1 U8567 ( .A(n6920), .ZN(n8061) );
  NOR2_X1 U8568 ( .A1(n6921), .A2(n8061), .ZN(n6860) );
  INV_X1 U8569 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6861) );
  NOR2_X1 U8570 ( .A1(n10321), .A2(n6861), .ZN(n6869) );
  AND2_X1 U8571 ( .A1(n10252), .A2(n8799), .ZN(n10308) );
  NAND2_X1 U8572 ( .A1(n6884), .A2(n6862), .ZN(n6864) );
  NAND2_X1 U8573 ( .A1(n6864), .A2(n6863), .ZN(n6905) );
  XNOR2_X1 U8574 ( .A(n6905), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U8575 ( .A1(n10308), .A2(n6865), .ZN(n6866) );
  OAI21_X1 U8576 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6867), .A(n6866), .ZN(n6868) );
  AOI211_X1 U8577 ( .C1(n10303), .C2(n6870), .A(n6869), .B(n6868), .ZN(n6875)
         );
  INV_X1 U8578 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7105) );
  MUX2_X1 U8579 ( .A(n7105), .B(n4668), .S(n8049), .Z(n10250) );
  NAND2_X1 U8580 ( .A1(n10250), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10249) );
  MUX2_X1 U8581 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8049), .Z(n6885) );
  XOR2_X1 U8582 ( .A(n10249), .B(n6886), .Z(n6873) );
  OR2_X1 U8583 ( .A1(n8972), .A2(n6872), .ZN(n10317) );
  INV_X1 U8584 ( .A(n10317), .ZN(n10272) );
  NAND2_X1 U8585 ( .A1(n6873), .A2(n10272), .ZN(n6874) );
  OAI211_X1 U8586 ( .C1(n10312), .C2(n6884), .A(n6875), .B(n6874), .ZN(
        P2_U3183) );
  INV_X1 U8587 ( .A(n6876), .ZN(n6877) );
  NOR2_X1 U8588 ( .A1(n6878), .A2(n6877), .ZN(n6880) );
  XNOR2_X1 U8589 ( .A(n6880), .B(n6879), .ZN(n6883) );
  AOI22_X1 U8590 ( .A1(n9492), .A2(n5982), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8578), .ZN(n6882) );
  AND2_X1 U8591 ( .A1(n9996), .A2(n9834), .ZN(n9473) );
  INV_X1 U8592 ( .A(n9991), .ZN(n9794) );
  AND2_X1 U8593 ( .A1(n9996), .A2(n9794), .ZN(n9474) );
  AOI22_X1 U8594 ( .A1(n9473), .A2(n9513), .B1(n9474), .B2(n6991), .ZN(n6881)
         );
  OAI211_X1 U8595 ( .C1(n6883), .C2(n9494), .A(n6882), .B(n6881), .ZN(P1_U3222) );
  AOI22_X1 U8596 ( .A1(n6886), .A2(n10249), .B1(n6885), .B2(n6884), .ZN(n10270) );
  MUX2_X1 U8597 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8049), .Z(n6887) );
  XNOR2_X1 U8598 ( .A(n6887), .B(n10256), .ZN(n10271) );
  INV_X1 U8599 ( .A(n6887), .ZN(n6888) );
  MUX2_X1 U8600 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8049), .Z(n6889) );
  XOR2_X1 U8601 ( .A(n6908), .B(n6889), .Z(n10290) );
  NOR2_X1 U8602 ( .A1(n6889), .A2(n10286), .ZN(n6891) );
  MUX2_X1 U8603 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8049), .Z(n7009) );
  XNOR2_X1 U8604 ( .A(n7009), .B(n7008), .ZN(n6890) );
  INV_X1 U8605 ( .A(n7007), .ZN(n6893) );
  OAI21_X1 U8606 ( .B1(n10288), .B2(n6891), .A(n6890), .ZN(n6892) );
  NAND3_X1 U8607 ( .A1(n6893), .A2(n10272), .A3(n6892), .ZN(n6919) );
  INV_X1 U8608 ( .A(n10321), .ZN(n10248) );
  NAND2_X1 U8609 ( .A1(n6895), .A2(n6894), .ZN(n10258) );
  XNOR2_X1 U8610 ( .A(n6903), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U8611 ( .A1(n10258), .A2(n10259), .ZN(n10257) );
  NAND2_X1 U8612 ( .A1(n10256), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8613 ( .A1(n10257), .A2(n6896), .ZN(n6897) );
  NAND2_X1 U8614 ( .A1(n6897), .A2(n10286), .ZN(n6900) );
  NAND2_X1 U8615 ( .A1(n10281), .A2(n6900), .ZN(n6898) );
  XNOR2_X1 U8616 ( .A(n7029), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8617 ( .A1(n6898), .A2(n6899), .ZN(n7022) );
  INV_X1 U8618 ( .A(n6899), .ZN(n6901) );
  NAND3_X1 U8619 ( .A1(n10281), .A2(n6901), .A3(n6900), .ZN(n6902) );
  AND2_X1 U8620 ( .A1(n7022), .A2(n6902), .ZN(n6916) );
  INV_X1 U8621 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7148) );
  MUX2_X1 U8622 ( .A(n7148), .B(P2_REG2_REG_4__SCAN_IN), .S(n7029), .Z(n6913)
         );
  INV_X1 U8623 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8624 ( .A1(n10256), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U8625 ( .A1(n10277), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8626 ( .A1(n6909), .A2(n10286), .ZN(n6910) );
  NAND2_X1 U8627 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  NAND2_X1 U8628 ( .A1(n6912), .A2(n6913), .ZN(n7031) );
  OAI21_X1 U8629 ( .B1(n6913), .B2(n6912), .A(n7031), .ZN(n6914) );
  NAND2_X1 U8630 ( .A1(n10308), .A2(n6914), .ZN(n6915) );
  NAND2_X1 U8631 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7088) );
  OAI211_X1 U8632 ( .C1(n6916), .C2(n10283), .A(n6915), .B(n7088), .ZN(n6917)
         );
  AOI21_X1 U8633 ( .B1(n10248), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6917), .ZN(
        n6918) );
  OAI211_X1 U8634 ( .C1(n10312), .C2(n7008), .A(n6919), .B(n6918), .ZN(
        P2_U3186) );
  NAND3_X1 U8635 ( .A1(n6922), .A2(n6921), .A3(n6920), .ZN(n6923) );
  AOI21_X1 U8636 ( .B1(n6958), .B2(n6928), .A(n6923), .ZN(n6927) );
  NAND2_X1 U8637 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  AOI21_X1 U8638 ( .B1(n6927), .B2(n6926), .A(P2_U3151), .ZN(n6931) );
  OR2_X1 U8639 ( .A1(n6935), .A2(n6932), .ZN(n8800) );
  INV_X1 U8640 ( .A(n6928), .ZN(n6929) );
  NOR2_X1 U8641 ( .A1(n8800), .A2(n6929), .ZN(n6930) );
  INV_X1 U8642 ( .A(n8945), .ZN(n8221) );
  OR2_X1 U8643 ( .A1(n6957), .A2(n10390), .ZN(n6934) );
  NAND2_X1 U8644 ( .A1(n6934), .A2(n10343), .ZN(n8951) );
  AND2_X1 U8645 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U8646 ( .A1(n6936), .A2(n6935), .ZN(n6939) );
  NAND2_X1 U8647 ( .A1(n6939), .A2(n6938), .ZN(n8948) );
  OAI22_X1 U8648 ( .A1(n8933), .A2(n8647), .B1(n7075), .B2(n8948), .ZN(n6940)
         );
  AOI211_X1 U8649 ( .C1(n10369), .C2(n8951), .A(n10278), .B(n6940), .ZN(n6964)
         );
  NAND2_X1 U8650 ( .A1(n6943), .A2(n5740), .ZN(n6945) );
  AND2_X1 U8651 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  XNOR2_X1 U8652 ( .A(n6950), .B(n6948), .ZN(n7072) );
  NAND2_X1 U8653 ( .A1(n4526), .A2(n7107), .ZN(n6949) );
  NAND2_X1 U8654 ( .A1(n8612), .A2(n6949), .ZN(n7073) );
  NAND2_X1 U8655 ( .A1(n7072), .A2(n7073), .ZN(n6952) );
  NAND2_X1 U8656 ( .A1(n6950), .A2(n5692), .ZN(n6951) );
  NAND2_X1 U8657 ( .A1(n6952), .A2(n6951), .ZN(n7065) );
  XNOR2_X1 U8658 ( .A(n7132), .B(n7067), .ZN(n6953) );
  XNOR2_X1 U8659 ( .A(n6953), .B(n10327), .ZN(n7066) );
  NAND2_X1 U8660 ( .A1(n7065), .A2(n7066), .ZN(n6955) );
  NAND2_X1 U8661 ( .A1(n6953), .A2(n7075), .ZN(n6954) );
  NAND2_X1 U8662 ( .A1(n6955), .A2(n6954), .ZN(n7130) );
  XNOR2_X1 U8663 ( .A(n7132), .B(n10369), .ZN(n7079) );
  XNOR2_X1 U8664 ( .A(n7079), .B(n10347), .ZN(n7126) );
  OR2_X1 U8665 ( .A1(n6957), .A2(n6956), .ZN(n6961) );
  NAND2_X1 U8666 ( .A1(n6959), .A2(n6958), .ZN(n6960) );
  AOI21_X1 U8667 ( .B1(n7130), .B2(n7126), .A(n8953), .ZN(n6962) );
  OR2_X1 U8668 ( .A1(n7130), .A2(n7126), .ZN(n7083) );
  NAND2_X1 U8669 ( .A1(n6962), .A2(n7083), .ZN(n6963) );
  OAI211_X1 U8670 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8221), .A(n6964), .B(
        n6963), .ZN(P2_U3158) );
  INV_X1 U8671 ( .A(n8373), .ZN(n8985) );
  INV_X1 U8672 ( .A(n6965), .ZN(n6967) );
  INV_X1 U8673 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6966) );
  OAI222_X1 U8674 ( .A1(n8985), .A2(P2_U3151), .B1(n9355), .B2(n6967), .C1(
        n6966), .C2(n8849), .ZN(P2_U3281) );
  INV_X1 U8675 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7917) );
  INV_X1 U8676 ( .A(n9553), .ZN(n9558) );
  OAI222_X1 U8677 ( .A1(n9952), .A2(n7917), .B1(n9949), .B2(n6967), .C1(
        P1_U3086), .C2(n9558), .ZN(P1_U3341) );
  INV_X1 U8678 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6969) );
  INV_X1 U8679 ( .A(n6968), .ZN(n6971) );
  INV_X1 U8680 ( .A(n9568), .ZN(n9574) );
  OAI222_X1 U8681 ( .A1(n9952), .A2(n6969), .B1(n9949), .B2(n6971), .C1(
        P1_U3086), .C2(n9574), .ZN(P1_U3340) );
  INV_X1 U8682 ( .A(n9013), .ZN(n9002) );
  INV_X1 U8683 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6970) );
  OAI222_X1 U8684 ( .A1(n9002), .A2(P2_U3151), .B1(n9355), .B2(n6971), .C1(
        n6970), .C2(n8849), .ZN(P2_U3280) );
  INV_X1 U8685 ( .A(n9021), .ZN(n9036) );
  INV_X1 U8686 ( .A(n6972), .ZN(n6974) );
  OAI222_X1 U8687 ( .A1(P2_U3151), .A2(n9036), .B1(n9355), .B2(n6974), .C1(
        n6973), .C2(n8849), .ZN(P2_U3279) );
  INV_X1 U8688 ( .A(n9589), .ZN(n9595) );
  OAI222_X1 U8689 ( .A1(n9952), .A2(n6975), .B1(n9949), .B2(n6974), .C1(n9595), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  NAND2_X1 U8690 ( .A1(n6991), .A2(n6976), .ZN(n7209) );
  XNOR2_X1 U8691 ( .A(n6306), .B(n7209), .ZN(n10135) );
  AND3_X1 U8692 ( .A1(n6979), .A2(n6978), .A3(n6977), .ZN(n6980) );
  NAND3_X1 U8693 ( .A1(n6982), .A2(n6981), .A3(n6980), .ZN(n7002) );
  INV_X1 U8694 ( .A(n7216), .ZN(n6983) );
  NAND2_X1 U8695 ( .A1(n10118), .A2(n6983), .ZN(n8297) );
  NAND2_X1 U8696 ( .A1(n6985), .A2(n6984), .ZN(n6987) );
  INV_X1 U8697 ( .A(n6986), .ZN(n10107) );
  AND2_X1 U8698 ( .A1(n6987), .A2(n10107), .ZN(n10117) );
  NAND2_X1 U8699 ( .A1(n6989), .A2(n6988), .ZN(n6990) );
  NAND2_X1 U8700 ( .A1(n10117), .A2(n6990), .ZN(n9859) );
  AOI22_X1 U8701 ( .A1(n9513), .A2(n9834), .B1(n9794), .B2(n6991), .ZN(n6998)
         );
  OAI21_X1 U8702 ( .B1(n6306), .B2(n6993), .A(n6992), .ZN(n6996) );
  OR2_X1 U8703 ( .A1(n4507), .A2(n7985), .ZN(n6995) );
  AND2_X1 U8704 ( .A1(n6995), .A2(n6994), .ZN(n10129) );
  INV_X1 U8705 ( .A(n10129), .ZN(n10092) );
  NAND2_X1 U8706 ( .A1(n6996), .A2(n10092), .ZN(n6997) );
  OAI211_X1 U8707 ( .C1(n10135), .C2(n9859), .A(n6998), .B(n6997), .ZN(n10138)
         );
  NAND2_X1 U8708 ( .A1(n10138), .A2(n10118), .ZN(n7006) );
  NAND2_X1 U8709 ( .A1(n10118), .A2(n6999), .ZN(n9815) );
  INV_X1 U8710 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7000) );
  OAI22_X1 U8711 ( .A1(n10118), .A2(n6790), .B1(n7000), .B2(n10108), .ZN(n7004) );
  INV_X1 U8712 ( .A(n10101), .ZN(n7001) );
  OAI211_X1 U8713 ( .C1(n10137), .C2(n10111), .A(n7001), .B(n10099), .ZN(
        n10136) );
  OR2_X1 U8714 ( .A1(n7002), .A2(n6504), .ZN(n9847) );
  NOR2_X1 U8715 ( .A1(n10136), .A2(n9847), .ZN(n7003) );
  AOI211_X1 U8716 ( .C1(n10094), .C2(n5982), .A(n7004), .B(n7003), .ZN(n7005)
         );
  OAI211_X1 U8717 ( .C1(n10135), .C2(n8297), .A(n7006), .B(n7005), .ZN(
        P1_U3292) );
  MUX2_X1 U8718 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8049), .Z(n7010) );
  XNOR2_X1 U8719 ( .A(n7010), .B(n7118), .ZN(n7110) );
  INV_X1 U8720 ( .A(n7118), .ZN(n7032) );
  INV_X1 U8721 ( .A(n7010), .ZN(n7011) );
  OAI22_X1 U8722 ( .A1(n7111), .A2(n7110), .B1(n7032), .B2(n7011), .ZN(n10316)
         );
  INV_X1 U8723 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7257) );
  MUX2_X1 U8724 ( .A(n7257), .B(n7024), .S(n8049), .Z(n7012) );
  NAND2_X1 U8725 ( .A1(n7012), .A2(n7036), .ZN(n7013) );
  OAI21_X1 U8726 ( .B1(n7012), .B2(n7036), .A(n7013), .ZN(n10315) );
  INV_X1 U8727 ( .A(n7013), .ZN(n7014) );
  INV_X1 U8728 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7406) );
  MUX2_X1 U8729 ( .A(n7406), .B(n7015), .S(n8049), .Z(n7183) );
  XNOR2_X1 U8730 ( .A(n7183), .B(n7197), .ZN(n7016) );
  AOI21_X1 U8731 ( .B1(n7017), .B2(n7016), .A(n7182), .ZN(n7040) );
  INV_X1 U8732 ( .A(n10312), .ZN(n9045) );
  INV_X1 U8733 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7019) );
  AND2_X1 U8734 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7313) );
  INV_X1 U8735 ( .A(n7313), .ZN(n7018) );
  OAI21_X1 U8736 ( .B1(n10321), .B2(n7019), .A(n7018), .ZN(n7028) );
  OR2_X1 U8737 ( .A1(n7029), .A2(n7020), .ZN(n7021) );
  NAND2_X1 U8738 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  NAND2_X1 U8739 ( .A1(n7023), .A2(n7118), .ZN(n10296) );
  INV_X1 U8740 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10429) );
  MUX2_X1 U8741 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7024), .S(n7036), .Z(n10297)
         );
  AOI21_X1 U8742 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n10311), .A(n10295), .ZN(
        n7188) );
  XNOR2_X1 U8743 ( .A(n7188), .B(n7197), .ZN(n7025) );
  NOR2_X1 U8744 ( .A1(n7025), .A2(n7015), .ZN(n7189) );
  AOI21_X1 U8745 ( .B1(n7015), .B2(n7025), .A(n7189), .ZN(n7026) );
  NOR2_X1 U8746 ( .A1(n7026), .A2(n10283), .ZN(n7027) );
  AOI211_X1 U8747 ( .C1(n9045), .C2(n7197), .A(n7028), .B(n7027), .ZN(n7039)
         );
  OR2_X1 U8748 ( .A1(n7029), .A2(n7148), .ZN(n7030) );
  NAND2_X1 U8749 ( .A1(n7031), .A2(n7030), .ZN(n7033) );
  XNOR2_X1 U8750 ( .A(n7033), .B(n7032), .ZN(n7112) );
  NAND2_X1 U8751 ( .A1(n7112), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7035) );
  NAND2_X1 U8752 ( .A1(n7033), .A2(n7118), .ZN(n7034) );
  NAND2_X1 U8753 ( .A1(n7035), .A2(n7034), .ZN(n10305) );
  MUX2_X1 U8754 ( .A(n7257), .B(P2_REG2_REG_6__SCAN_IN), .S(n7036), .Z(n10306)
         );
  NAND2_X1 U8755 ( .A1(n10305), .A2(n10306), .ZN(n10304) );
  XNOR2_X1 U8756 ( .A(n7198), .B(n7406), .ZN(n7037) );
  NAND2_X1 U8757 ( .A1(n7037), .A2(n10308), .ZN(n7038) );
  OAI211_X1 U8758 ( .C1(n7040), .C2(n10317), .A(n7039), .B(n7038), .ZN(
        P2_U3189) );
  INV_X1 U8759 ( .A(n10022), .ZN(n10043) );
  NOR2_X1 U8760 ( .A1(n7295), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7041) );
  AOI21_X1 U8761 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7295), .A(n7041), .ZN(
        n7046) );
  NAND2_X1 U8762 ( .A1(n9544), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7044) );
  OAI21_X1 U8763 ( .B1(n9544), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7044), .ZN(
        n9541) );
  OAI21_X1 U8764 ( .B1(n7046), .B2(n7045), .A(n7289), .ZN(n7061) );
  NOR2_X1 U8765 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7047), .ZN(n9428) );
  AOI21_X1 U8766 ( .B1(n10049), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9428), .ZN(
        n7048) );
  OAI21_X1 U8767 ( .B1(n9629), .B2(n7049), .A(n7048), .ZN(n7060) );
  NAND2_X1 U8768 ( .A1(n9544), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7054) );
  INV_X1 U8769 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7050) );
  MUX2_X1 U8770 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7050), .S(n9544), .Z(n9546)
         );
  OAI21_X1 U8771 ( .B1(n7053), .B2(n7052), .A(n7051), .ZN(n9547) );
  NAND2_X1 U8772 ( .A1(n9546), .A2(n9547), .ZN(n9545) );
  NAND2_X1 U8773 ( .A1(n7054), .A2(n9545), .ZN(n7057) );
  INV_X1 U8774 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7055) );
  MUX2_X1 U8775 ( .A(n7055), .B(P1_REG1_REG_9__SCAN_IN), .S(n7295), .Z(n7056)
         );
  NOR2_X1 U8776 ( .A1(n7056), .A2(n7057), .ZN(n7296) );
  AOI21_X1 U8777 ( .B1(n7057), .B2(n7056), .A(n7296), .ZN(n7058) );
  NOR2_X1 U8778 ( .A1(n7058), .A2(n9631), .ZN(n7059) );
  AOI211_X1 U8779 ( .C1(n10043), .C2(n7061), .A(n7060), .B(n7059), .ZN(n7062)
         );
  INV_X1 U8780 ( .A(n7062), .ZN(P1_U3252) );
  INV_X1 U8781 ( .A(n7063), .ZN(n7109) );
  AOI22_X1 U8782 ( .A1(n9605), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9945), .ZN(n7064) );
  OAI21_X1 U8783 ( .B1(n7109), .B2(n9949), .A(n7064), .ZN(P1_U3338) );
  XOR2_X1 U8784 ( .A(n7066), .B(n7065), .Z(n7071) );
  NAND2_X1 U8785 ( .A1(n8221), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8581) );
  INV_X1 U8786 ( .A(n8948), .ZN(n8931) );
  AOI22_X1 U8787 ( .A1(n8931), .A2(n6948), .B1(n8951), .B2(n7067), .ZN(n7068)
         );
  OAI21_X1 U8788 ( .B1(n10347), .B2(n8933), .A(n7068), .ZN(n7069) );
  AOI21_X1 U8789 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n8581), .A(n7069), .ZN(
        n7070) );
  OAI21_X1 U8790 ( .B1(n7071), .B2(n8953), .A(n7070), .ZN(P2_U3177) );
  XOR2_X1 U8791 ( .A(n7073), .B(n7072), .Z(n7078) );
  AOI22_X1 U8792 ( .A1(n8931), .A2(n8973), .B1(n8951), .B2(n7157), .ZN(n7074)
         );
  OAI21_X1 U8793 ( .B1(n7075), .B2(n8933), .A(n7074), .ZN(n7076) );
  AOI21_X1 U8794 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8581), .A(n7076), .ZN(
        n7077) );
  OAI21_X1 U8795 ( .B1(n8953), .B2(n7078), .A(n7077), .ZN(P2_U3162) );
  XNOR2_X1 U8796 ( .A(n7125), .B(n8647), .ZN(n7086) );
  INV_X1 U8797 ( .A(n7079), .ZN(n7080) );
  NAND2_X1 U8798 ( .A1(n7080), .A2(n8971), .ZN(n7082) );
  NAND2_X1 U8799 ( .A1(n7083), .A2(n7082), .ZN(n7085) );
  INV_X1 U8800 ( .A(n7086), .ZN(n7081) );
  AND2_X1 U8801 ( .A1(n7082), .A2(n7081), .ZN(n7128) );
  AND2_X1 U8802 ( .A1(n7083), .A2(n7128), .ZN(n7084) );
  AOI21_X1 U8803 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7092) );
  INV_X1 U8804 ( .A(n7087), .ZN(n7149) );
  AOI22_X1 U8805 ( .A1(n8944), .A2(n8970), .B1(n8951), .B2(n8646), .ZN(n7089)
         );
  OAI211_X1 U8806 ( .C1(n10347), .C2(n8948), .A(n7089), .B(n7088), .ZN(n7090)
         );
  AOI21_X1 U8807 ( .B1(n7149), .B2(n8945), .A(n7090), .ZN(n7091) );
  OAI21_X1 U8808 ( .B1(n7092), .B2(n8953), .A(n7091), .ZN(P2_U3170) );
  NAND2_X1 U8809 ( .A1(n7096), .A2(n7093), .ZN(n7094) );
  OAI211_X1 U8810 ( .C1(n7097), .C2(n7096), .A(n7095), .B(n7094), .ZN(n7103)
         );
  INV_X1 U8811 ( .A(n7103), .ZN(n7098) );
  INV_X1 U8812 ( .A(n10341), .ZN(n9144) );
  NAND2_X1 U8813 ( .A1(n7098), .A2(n9144), .ZN(n10334) );
  INV_X1 U8814 ( .A(n10343), .ZN(n9225) );
  INV_X1 U8815 ( .A(n8765), .ZN(n7100) );
  NOR3_X1 U8816 ( .A1(n7100), .A2(n10416), .A3(n7099), .ZN(n7101) );
  AOI211_X1 U8817 ( .C1(n9225), .C2(P2_REG3_REG_0__SCAN_IN), .A(n7102), .B(
        n7101), .ZN(n7104) );
  NAND2_X1 U8818 ( .A1(n7103), .A2(n10343), .ZN(n9211) );
  INV_X2 U8819 ( .A(n10339), .ZN(n10357) );
  MUX2_X1 U8820 ( .A(n7105), .B(n7104), .S(n10357), .Z(n7106) );
  OAI21_X1 U8821 ( .B1(n10334), .B2(n7107), .A(n7106), .ZN(P2_U3233) );
  INV_X1 U8822 ( .A(n9067), .ZN(n9028) );
  OAI222_X1 U8823 ( .A1(n9028), .A2(P2_U3151), .B1(n7286), .B2(n7109), .C1(
        n7108), .C2(n8849), .ZN(P2_U3278) );
  XNOR2_X1 U8824 ( .A(n7111), .B(n7110), .ZN(n7122) );
  XNOR2_X1 U8825 ( .A(n7112), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U8826 ( .A1(n10298), .A2(n7113), .ZN(n7114) );
  NOR2_X1 U8827 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5210), .ZN(n7133) );
  AOI21_X1 U8828 ( .B1(n10303), .B2(n7114), .A(n7133), .ZN(n7117) );
  INV_X1 U8829 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7115) );
  OR2_X1 U8830 ( .A1(n10321), .A2(n7115), .ZN(n7116) );
  OAI211_X1 U8831 ( .C1(n10312), .C2(n7118), .A(n7117), .B(n7116), .ZN(n7119)
         );
  AOI21_X1 U8832 ( .B1(n10308), .B2(n7120), .A(n7119), .ZN(n7121) );
  OAI21_X1 U8833 ( .B1(n7122), .B2(n10317), .A(n7121), .ZN(P2_U3187) );
  INV_X1 U8834 ( .A(n7123), .ZN(n7161) );
  AOI22_X1 U8835 ( .A1(n9622), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9945), .ZN(n7124) );
  OAI21_X1 U8836 ( .B1(n7161), .B2(n9949), .A(n7124), .ZN(P1_U3337) );
  AND2_X1 U8837 ( .A1(n7125), .A2(n8647), .ZN(n7127) );
  OR2_X1 U8838 ( .A1(n7126), .A2(n7127), .ZN(n7129) );
  OAI22_X1 U8839 ( .A1(n7130), .A2(n7129), .B1(n7128), .B2(n7127), .ZN(n7131)
         );
  INV_X1 U8840 ( .A(n7131), .ZN(n7166) );
  XNOR2_X1 U8841 ( .A(n8838), .B(n7246), .ZN(n7163) );
  XNOR2_X1 U8842 ( .A(n7163), .B(n8970), .ZN(n7165) );
  XOR2_X1 U8843 ( .A(n7166), .B(n7165), .Z(n7139) );
  INV_X1 U8844 ( .A(n8647), .ZN(n10329) );
  AOI21_X1 U8845 ( .B1(n8931), .B2(n10329), .A(n7133), .ZN(n7136) );
  INV_X1 U8846 ( .A(n7243), .ZN(n7134) );
  NAND2_X1 U8847 ( .A1(n8945), .A2(n7134), .ZN(n7135) );
  OAI211_X1 U8848 ( .C1(n7398), .C2(n8933), .A(n7136), .B(n7135), .ZN(n7137)
         );
  AOI21_X1 U8849 ( .B1(n7246), .B2(n8951), .A(n7137), .ZN(n7138) );
  OAI21_X1 U8850 ( .B1(n7139), .B2(n8953), .A(n7138), .ZN(P2_U3167) );
  XNOR2_X1 U8851 ( .A(n7140), .B(n8767), .ZN(n10373) );
  AND2_X1 U8852 ( .A1(n7141), .A2(n5678), .ZN(n10356) );
  INV_X1 U8853 ( .A(n10356), .ZN(n7403) );
  NAND2_X1 U8854 ( .A1(n10353), .A2(n7403), .ZN(n7142) );
  NAND2_X1 U8855 ( .A1(n10357), .A2(n7142), .ZN(n9229) );
  AND2_X1 U8856 ( .A1(n7145), .A2(n7143), .ZN(n7146) );
  NAND2_X1 U8857 ( .A1(n7145), .A2(n7144), .ZN(n7238) );
  OAI21_X1 U8858 ( .B1(n8767), .B2(n7146), .A(n7238), .ZN(n7147) );
  AOI222_X1 U8859 ( .A1(n10350), .A2(n7147), .B1(n8971), .B2(n10326), .C1(
        n8970), .C2(n10328), .ZN(n10374) );
  MUX2_X1 U8860 ( .A(n7148), .B(n10374), .S(n10357), .Z(n7151) );
  AOI22_X1 U8861 ( .A1(n9226), .A2(n8646), .B1(n9225), .B2(n7149), .ZN(n7150)
         );
  OAI211_X1 U8862 ( .C1(n10373), .C2(n9229), .A(n7151), .B(n7150), .ZN(
        P2_U3229) );
  INV_X1 U8863 ( .A(n7152), .ZN(n7153) );
  AOI21_X1 U8864 ( .B1(n8612), .B2(n8766), .A(n7153), .ZN(n10361) );
  INV_X1 U8865 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7156) );
  XNOR2_X1 U8866 ( .A(n8766), .B(n7154), .ZN(n7155) );
  AOI222_X1 U8867 ( .A1(n10350), .A2(n7155), .B1(n8973), .B2(n10326), .C1(
        n10327), .C2(n10328), .ZN(n10359) );
  MUX2_X1 U8868 ( .A(n7156), .B(n10359), .S(n10357), .Z(n7159) );
  AOI22_X1 U8869 ( .A1(n9226), .A2(n7157), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9225), .ZN(n7158) );
  OAI211_X1 U8870 ( .C1(n10361), .C2(n9229), .A(n7159), .B(n7158), .ZN(
        P2_U3232) );
  INV_X1 U8871 ( .A(n9063), .ZN(n9083) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7160) );
  OAI222_X1 U8873 ( .A1(P2_U3151), .A2(n9083), .B1(n9355), .B2(n7161), .C1(
        n7160), .C2(n8849), .ZN(P2_U3277) );
  AND2_X1 U8874 ( .A1(n7163), .A2(n7162), .ZN(n7164) );
  XNOR2_X1 U8875 ( .A(n7259), .B(n8838), .ZN(n7303) );
  XNOR2_X1 U8876 ( .A(n7303), .B(n8969), .ZN(n7168) );
  NAND2_X1 U8877 ( .A1(n7167), .A2(n7168), .ZN(n7306) );
  INV_X1 U8878 ( .A(n8953), .ZN(n8928) );
  OAI211_X1 U8879 ( .C1(n7167), .C2(n7168), .A(n7306), .B(n8928), .ZN(n7174)
         );
  INV_X1 U8880 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7944) );
  NOR2_X1 U8881 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7944), .ZN(n10301) );
  AOI21_X1 U8882 ( .B1(n8931), .B2(n8970), .A(n10301), .ZN(n7171) );
  INV_X1 U8883 ( .A(n7169), .ZN(n7258) );
  NAND2_X1 U8884 ( .A1(n8945), .A2(n7258), .ZN(n7170) );
  OAI211_X1 U8885 ( .C1(n7341), .C2(n8933), .A(n7171), .B(n7170), .ZN(n7172)
         );
  AOI21_X1 U8886 ( .B1(n7259), .B2(n8951), .A(n7172), .ZN(n7173) );
  NAND2_X1 U8887 ( .A1(n7174), .A2(n7173), .ZN(P2_U3179) );
  XOR2_X1 U8888 ( .A(n7176), .B(n7175), .Z(n7181) );
  OR2_X1 U8889 ( .A1(n7213), .A2(n9991), .ZN(n7178) );
  OR2_X1 U8890 ( .A1(n7273), .A2(n9989), .ZN(n7177) );
  NAND2_X1 U8891 ( .A1(n7178), .A2(n7177), .ZN(n7207) );
  AOI22_X1 U8892 ( .A1(n7207), .A2(n9996), .B1(n7219), .B2(n9492), .ZN(n7180)
         );
  MUX2_X1 U8893 ( .A(n10003), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7179) );
  OAI211_X1 U8894 ( .C1(n7181), .C2(n9494), .A(n7180), .B(n7179), .ZN(P1_U3218) );
  MUX2_X1 U8895 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8049), .Z(n7184) );
  NOR2_X1 U8896 ( .A1(n7184), .A2(n7459), .ZN(n7474) );
  AOI21_X1 U8897 ( .B1(n7184), .B2(n7459), .A(n7474), .ZN(n7185) );
  INV_X1 U8898 ( .A(n7185), .ZN(n7186) );
  NOR2_X1 U8899 ( .A1(n4556), .A2(n7186), .ZN(n7473) );
  AOI21_X1 U8900 ( .B1(n4556), .B2(n7186), .A(n7473), .ZN(n7204) );
  INV_X1 U8901 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7590) );
  INV_X1 U8902 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7934) );
  NOR2_X1 U8903 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7934), .ZN(n7343) );
  INV_X1 U8904 ( .A(n7343), .ZN(n7187) );
  OAI21_X1 U8905 ( .B1(n10321), .B2(n7590), .A(n7187), .ZN(n7195) );
  INV_X1 U8906 ( .A(n7188), .ZN(n7190) );
  AOI22_X1 U8907 ( .A1(n7466), .A2(P2_REG1_REG_8__SCAN_IN), .B1(n5269), .B2(
        n7459), .ZN(n7191) );
  NOR2_X1 U8908 ( .A1(n7192), .A2(n7191), .ZN(n7461) );
  AOI21_X1 U8909 ( .B1(n7192), .B2(n7191), .A(n7461), .ZN(n7193) );
  NOR2_X1 U8910 ( .A1(n7193), .A2(n10283), .ZN(n7194) );
  AOI211_X1 U8911 ( .C1(n9045), .C2(n7466), .A(n7195), .B(n7194), .ZN(n7203)
         );
  AOI22_X1 U8912 ( .A1(n7466), .A2(n5266), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n7459), .ZN(n7199) );
  OAI21_X1 U8913 ( .B1(n7200), .B2(n7199), .A(n7465), .ZN(n7201) );
  NAND2_X1 U8914 ( .A1(n7201), .A2(n10308), .ZN(n7202) );
  OAI211_X1 U8915 ( .C1(n7204), .C2(n10317), .A(n7203), .B(n7202), .ZN(
        P2_U3190) );
  XNOR2_X1 U8916 ( .A(n7206), .B(n7205), .ZN(n7208) );
  AOI21_X1 U8917 ( .B1(n7208), .B2(n10092), .A(n7207), .ZN(n10154) );
  INV_X2 U8918 ( .A(n10118), .ZN(n10121) );
  NAND2_X1 U8919 ( .A1(n7210), .A2(n7209), .ZN(n7212) );
  NAND2_X1 U8920 ( .A1(n8577), .A2(n10137), .ZN(n7211) );
  NAND2_X1 U8921 ( .A1(n7212), .A2(n7211), .ZN(n10097) );
  NAND2_X1 U8922 ( .A1(n10097), .A2(n10098), .ZN(n7215) );
  NAND2_X1 U8923 ( .A1(n7213), .A2(n10143), .ZN(n7214) );
  XNOR2_X1 U8924 ( .A(n7272), .B(n7271), .ZN(n10152) );
  NAND2_X1 U8925 ( .A1(n9859), .A2(n7216), .ZN(n7217) );
  NAND2_X1 U8926 ( .A1(n10118), .A2(n7217), .ZN(n9829) );
  INV_X1 U8927 ( .A(n9829), .ZN(n10104) );
  INV_X1 U8928 ( .A(n10099), .ZN(n9810) );
  AOI21_X1 U8929 ( .B1(n10100), .B2(n7219), .A(n9810), .ZN(n7218) );
  NAND2_X1 U8930 ( .A1(n7218), .A2(n7332), .ZN(n10149) );
  INV_X1 U8931 ( .A(n10108), .ZN(n10096) );
  AOI22_X1 U8932 ( .A1(n10121), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10096), .B2(
        n9514), .ZN(n7221) );
  NAND2_X1 U8933 ( .A1(n10094), .A2(n7219), .ZN(n7220) );
  OAI211_X1 U8934 ( .C1(n10149), .C2(n9847), .A(n7221), .B(n7220), .ZN(n7222)
         );
  AOI21_X1 U8935 ( .B1(n10152), .B2(n10104), .A(n7222), .ZN(n7223) );
  OAI21_X1 U8936 ( .B1(n10154), .B2(n10121), .A(n7223), .ZN(P1_U3290) );
  OAI211_X1 U8937 ( .C1(n7226), .C2(n7225), .A(n7224), .B(n10000), .ZN(n7231)
         );
  OAI22_X1 U8938 ( .A1(n9998), .A2(n7334), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10041), .ZN(n7229) );
  INV_X1 U8939 ( .A(n9473), .ZN(n9487) );
  INV_X1 U8940 ( .A(n7227), .ZN(n7333) );
  OAI22_X1 U8941 ( .A1(n9487), .A2(n7509), .B1(n10003), .B2(n7333), .ZN(n7228)
         );
  AOI211_X1 U8942 ( .C1(n9474), .C2(n9512), .A(n7229), .B(n7228), .ZN(n7230)
         );
  NAND2_X1 U8943 ( .A1(n7231), .A2(n7230), .ZN(P1_U3230) );
  NAND2_X1 U8944 ( .A1(n7233), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7232) );
  OAI21_X1 U8945 ( .B1(n7234), .B2(n7233), .A(n7232), .ZN(P1_U3583) );
  XNOR2_X1 U8946 ( .A(n8970), .B(n7246), .ZN(n8769) );
  INV_X1 U8947 ( .A(n8769), .ZN(n7236) );
  XNOR2_X1 U8948 ( .A(n7235), .B(n7236), .ZN(n10378) );
  NAND2_X1 U8949 ( .A1(n10357), .A2(n10356), .ZN(n8812) );
  NAND2_X1 U8950 ( .A1(n7238), .A2(n7237), .ZN(n7239) );
  XOR2_X1 U8951 ( .A(n8769), .B(n7239), .Z(n7241) );
  OAI22_X1 U8952 ( .A1(n7398), .A2(n10346), .B1(n8647), .B2(n10348), .ZN(n7240) );
  AOI21_X1 U8953 ( .B1(n7241), .B2(n10350), .A(n7240), .ZN(n7242) );
  OAI21_X1 U8954 ( .B1(n10378), .B2(n10353), .A(n7242), .ZN(n10380) );
  NAND2_X1 U8955 ( .A1(n10380), .A2(n9211), .ZN(n7248) );
  INV_X1 U8956 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7244) );
  OAI22_X1 U8957 ( .A1(n10357), .A2(n7244), .B1(n7243), .B2(n10343), .ZN(n7245) );
  AOI21_X1 U8958 ( .B1(n9226), .B2(n7246), .A(n7245), .ZN(n7247) );
  OAI211_X1 U8959 ( .C1(n10378), .C2(n8812), .A(n7248), .B(n7247), .ZN(
        P2_U3228) );
  INV_X1 U8960 ( .A(n7249), .ZN(n7251) );
  OR2_X1 U8961 ( .A1(n7251), .A2(n7250), .ZN(n8768) );
  NAND2_X1 U8962 ( .A1(n7253), .A2(n7252), .ZN(n7254) );
  XOR2_X1 U8963 ( .A(n8768), .B(n7254), .Z(n10384) );
  XOR2_X1 U8964 ( .A(n8768), .B(n7255), .Z(n7256) );
  AOI222_X1 U8965 ( .A1(n10350), .A2(n7256), .B1(n8968), .B2(n10328), .C1(
        n8970), .C2(n10326), .ZN(n10385) );
  MUX2_X1 U8966 ( .A(n7257), .B(n10385), .S(n10357), .Z(n7261) );
  AOI22_X1 U8967 ( .A1(n9226), .A2(n7259), .B1(n9225), .B2(n7258), .ZN(n7260)
         );
  OAI211_X1 U8968 ( .C1(n10384), .C2(n9229), .A(n7261), .B(n7260), .ZN(
        P2_U3227) );
  NAND2_X1 U8969 ( .A1(n7262), .A2(n7263), .ZN(n7265) );
  NAND2_X1 U8970 ( .A1(n7265), .A2(n7264), .ZN(n7267) );
  INV_X1 U8971 ( .A(n7376), .ZN(n7266) );
  XNOR2_X1 U8972 ( .A(n7267), .B(n7266), .ZN(n7270) );
  OR2_X1 U8973 ( .A1(n7273), .A2(n9991), .ZN(n7269) );
  OR2_X1 U8974 ( .A1(n7494), .A2(n9989), .ZN(n7268) );
  NAND2_X1 U8975 ( .A1(n7269), .A2(n7268), .ZN(n7412) );
  AOI21_X1 U8976 ( .B1(n7270), .B2(n10092), .A(n7412), .ZN(n10170) );
  NAND2_X1 U8977 ( .A1(n7272), .A2(n7271), .ZN(n7326) );
  NAND2_X1 U8978 ( .A1(n8576), .A2(n10150), .ZN(n7327) );
  NAND2_X1 U8979 ( .A1(n7273), .A2(n7334), .ZN(n7274) );
  AND2_X1 U8980 ( .A1(n7327), .A2(n7274), .ZN(n7278) );
  INV_X1 U8981 ( .A(n7274), .ZN(n7275) );
  NOR2_X1 U8982 ( .A1(n7276), .A2(n7275), .ZN(n7277) );
  XNOR2_X1 U8983 ( .A(n7377), .B(n7376), .ZN(n10168) );
  OAI21_X1 U8984 ( .B1(n7331), .B2(n10166), .A(n10099), .ZN(n7279) );
  OR2_X1 U8985 ( .A1(n7279), .A2(n10086), .ZN(n10165) );
  AOI22_X1 U8986 ( .A1(n10121), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7411), .B2(
        n10096), .ZN(n7281) );
  NAND2_X1 U8987 ( .A1(n10094), .A2(n7413), .ZN(n7280) );
  OAI211_X1 U8988 ( .C1(n10165), .C2(n9847), .A(n7281), .B(n7280), .ZN(n7282)
         );
  AOI21_X1 U8989 ( .B1(n10168), .B2(n10104), .A(n7282), .ZN(n7283) );
  OAI21_X1 U8990 ( .B1(n10170), .B2(n10121), .A(n7283), .ZN(P1_U3288) );
  INV_X1 U8991 ( .A(n7284), .ZN(n8847) );
  OAI222_X1 U8992 ( .A1(P2_U3151), .A2(n9093), .B1(n7286), .B2(n8847), .C1(
        n7285), .C2(n8849), .ZN(P2_U3276) );
  INV_X1 U8993 ( .A(n9629), .ZN(n10051) );
  INV_X1 U8994 ( .A(n10049), .ZN(n9635) );
  INV_X1 U8995 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7288) );
  AND2_X1 U8996 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8464) );
  INV_X1 U8997 ( .A(n8464), .ZN(n7287) );
  OAI21_X1 U8998 ( .B1(n9635), .B2(n7288), .A(n7287), .ZN(n7294) );
  OAI21_X1 U8999 ( .B1(n7295), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7289), .ZN(
        n7292) );
  NAND2_X1 U9000 ( .A1(n7359), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7290) );
  OAI21_X1 U9001 ( .B1(n7359), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7290), .ZN(
        n7291) );
  NOR2_X1 U9002 ( .A1(n7291), .A2(n7292), .ZN(n7358) );
  AOI211_X1 U9003 ( .C1(n7292), .C2(n7291), .A(n7358), .B(n10022), .ZN(n7293)
         );
  AOI211_X1 U9004 ( .C1(n10051), .C2(n7359), .A(n7294), .B(n7293), .ZN(n7302)
         );
  NOR2_X1 U9005 ( .A1(n7295), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7297) );
  NOR2_X1 U9006 ( .A1(n7297), .A2(n7296), .ZN(n7300) );
  INV_X1 U9007 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7298) );
  MUX2_X1 U9008 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7298), .S(n7359), .Z(n7299)
         );
  INV_X1 U9009 ( .A(n9631), .ZN(n10053) );
  NAND2_X1 U9010 ( .A1(n7299), .A2(n7300), .ZN(n7353) );
  OAI211_X1 U9011 ( .C1(n7300), .C2(n7299), .A(n10053), .B(n7353), .ZN(n7301)
         );
  NAND2_X1 U9012 ( .A1(n7302), .A2(n7301), .ZN(P1_U3253) );
  XNOR2_X1 U9013 ( .A(n7393), .B(n4527), .ZN(n7340) );
  XNOR2_X1 U9014 ( .A(n7340), .B(n8968), .ZN(n7311) );
  INV_X1 U9015 ( .A(n7303), .ZN(n7304) );
  NAND2_X1 U9016 ( .A1(n7304), .A2(n8969), .ZN(n7305) );
  NAND2_X1 U9017 ( .A1(n7306), .A2(n7305), .ZN(n7310) );
  INV_X1 U9018 ( .A(n7310), .ZN(n7308) );
  INV_X1 U9019 ( .A(n7311), .ZN(n7307) );
  INV_X1 U9020 ( .A(n7547), .ZN(n7309) );
  AOI21_X1 U9021 ( .B1(n7311), .B2(n7310), .A(n7309), .ZN(n7317) );
  NOR2_X1 U9022 ( .A1(n8948), .A2(n7398), .ZN(n7312) );
  AOI211_X1 U9023 ( .C1(n8944), .C2(n8967), .A(n7313), .B(n7312), .ZN(n7314)
         );
  OAI21_X1 U9024 ( .B1(n7402), .B2(n8221), .A(n7314), .ZN(n7315) );
  AOI21_X1 U9025 ( .B1(n7393), .B2(n8951), .A(n7315), .ZN(n7316) );
  OAI21_X1 U9026 ( .B1(n7317), .B2(n8953), .A(n7316), .ZN(P2_U3153) );
  NAND2_X1 U9027 ( .A1(n8636), .A2(n8657), .ZN(n8771) );
  NAND2_X1 U9028 ( .A1(n7394), .A2(n7318), .ZN(n7319) );
  XOR2_X1 U9029 ( .A(n8771), .B(n7319), .Z(n10397) );
  INV_X1 U9030 ( .A(n10350), .ZN(n9187) );
  OR2_X1 U9031 ( .A1(n7429), .A2(n8653), .ZN(n7396) );
  NAND2_X1 U9032 ( .A1(n7396), .A2(n7320), .ZN(n7321) );
  XOR2_X1 U9033 ( .A(n8771), .B(n7321), .Z(n7322) );
  OAI222_X1 U9034 ( .A1(n10346), .A2(n7567), .B1(n10348), .B2(n7341), .C1(
        n9187), .C2(n7322), .ZN(n10398) );
  NAND2_X1 U9035 ( .A1(n10398), .A2(n9211), .ZN(n7325) );
  OAI22_X1 U9036 ( .A1(n10357), .A2(n5266), .B1(n7344), .B2(n10343), .ZN(n7323) );
  AOI21_X1 U9037 ( .B1(n9226), .B2(n10400), .A(n7323), .ZN(n7324) );
  OAI211_X1 U9038 ( .C1(n10397), .C2(n9229), .A(n7325), .B(n7324), .ZN(
        P2_U3225) );
  NAND2_X1 U9039 ( .A1(n7326), .A2(n7327), .ZN(n7328) );
  XNOR2_X1 U9040 ( .A(n7328), .B(n7329), .ZN(n10161) );
  XNOR2_X1 U9041 ( .A(n7262), .B(n7329), .ZN(n7330) );
  AOI222_X1 U9042 ( .A1(n10092), .A2(n7330), .B1(n9510), .B2(n9834), .C1(n9512), .C2(n9794), .ZN(n10160) );
  MUX2_X1 U9043 ( .A(n6789), .B(n10160), .S(n10118), .Z(n7337) );
  AOI211_X1 U9044 ( .C1(n10157), .C2(n7332), .A(n9810), .B(n7331), .ZN(n10156)
         );
  INV_X1 U9045 ( .A(n9847), .ZN(n10103) );
  OAI22_X1 U9046 ( .A1(n9815), .A2(n7334), .B1(n10108), .B2(n7333), .ZN(n7335)
         );
  AOI21_X1 U9047 ( .B1(n10156), .B2(n10103), .A(n7335), .ZN(n7336) );
  OAI211_X1 U9048 ( .C1(n10161), .C2(n9829), .A(n7337), .B(n7336), .ZN(
        P1_U3289) );
  INV_X1 U9049 ( .A(n7338), .ZN(n7351) );
  INV_X1 U9050 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7339) );
  OAI222_X1 U9051 ( .A1(n5740), .A2(P2_U3151), .B1(n9355), .B2(n7351), .C1(
        n7339), .C2(n8849), .ZN(P2_U3275) );
  XNOR2_X1 U9052 ( .A(n10400), .B(n8838), .ZN(n7537) );
  XNOR2_X1 U9053 ( .A(n7537), .B(n8967), .ZN(n7542) );
  INV_X1 U9054 ( .A(n7340), .ZN(n7342) );
  NAND2_X1 U9055 ( .A1(n7342), .A2(n7341), .ZN(n7541) );
  NAND2_X1 U9056 ( .A1(n7547), .A2(n7541), .ZN(n7535) );
  XOR2_X1 U9057 ( .A(n7542), .B(n7535), .Z(n7350) );
  AOI21_X1 U9058 ( .B1(n8931), .B2(n8968), .A(n7343), .ZN(n7347) );
  INV_X1 U9059 ( .A(n7344), .ZN(n7345) );
  NAND2_X1 U9060 ( .A1(n8945), .A2(n7345), .ZN(n7346) );
  OAI211_X1 U9061 ( .C1(n7567), .C2(n8933), .A(n7347), .B(n7346), .ZN(n7348)
         );
  AOI21_X1 U9062 ( .B1(n10400), .B2(n8951), .A(n7348), .ZN(n7349) );
  OAI21_X1 U9063 ( .B1(n7350), .B2(n8953), .A(n7349), .ZN(P2_U3161) );
  INV_X1 U9064 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7932) );
  OAI222_X1 U9065 ( .A1(n9952), .A2(n7932), .B1(P1_U3086), .B2(n7352), .C1(
        n9949), .C2(n7351), .ZN(P1_U3335) );
  NAND2_X1 U9066 ( .A1(n7359), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7354) );
  NAND2_X1 U9067 ( .A1(n7354), .A2(n7353), .ZN(n7357) );
  INV_X1 U9068 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7355) );
  MUX2_X1 U9069 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7355), .S(n7443), .Z(n7356)
         );
  NAND2_X1 U9070 ( .A1(n7356), .A2(n7357), .ZN(n7448) );
  OAI211_X1 U9071 ( .C1(n7357), .C2(n7356), .A(n10053), .B(n7448), .ZN(n7368)
         );
  INV_X1 U9072 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7360) );
  AOI22_X1 U9073 ( .A1(n7443), .A2(n7360), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7449), .ZN(n7361) );
  AOI211_X1 U9074 ( .C1(n7362), .C2(n7361), .A(n7442), .B(n10022), .ZN(n7366)
         );
  NOR2_X1 U9075 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8426), .ZN(n7363) );
  AOI21_X1 U9076 ( .B1(n10049), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7363), .ZN(
        n7364) );
  OAI21_X1 U9077 ( .B1(n9629), .B2(n7449), .A(n7364), .ZN(n7365) );
  NOR2_X1 U9078 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  NAND2_X1 U9079 ( .A1(n7368), .A2(n7367), .ZN(P1_U3254) );
  NAND2_X1 U9080 ( .A1(n7369), .A2(n7370), .ZN(n10084) );
  OR2_X1 U9081 ( .A1(n10079), .A2(n10084), .ZN(n7371) );
  NAND2_X1 U9082 ( .A1(n7371), .A2(n7370), .ZN(n7372) );
  NOR2_X1 U9083 ( .A1(n7372), .A2(n7382), .ZN(n10062) );
  AND2_X1 U9084 ( .A1(n7372), .A2(n7382), .ZN(n7373) );
  OR2_X1 U9085 ( .A1(n10062), .A2(n7373), .ZN(n7375) );
  OAI22_X1 U9086 ( .A1(n6066), .A2(n9989), .B1(n7494), .B2(n9991), .ZN(n7374)
         );
  AOI21_X1 U9087 ( .B1(n7375), .B2(n10092), .A(n7374), .ZN(n7384) );
  NAND2_X1 U9088 ( .A1(n7377), .A2(n7376), .ZN(n7379) );
  NAND2_X1 U9089 ( .A1(n7509), .A2(n10166), .ZN(n7378) );
  NAND2_X1 U9090 ( .A1(n7379), .A2(n7378), .ZN(n8012) );
  NAND2_X1 U9091 ( .A1(n8012), .A2(n10084), .ZN(n7380) );
  NAND2_X1 U9092 ( .A1(n7494), .A2(n10174), .ZN(n8009) );
  NAND2_X1 U9093 ( .A1(n7380), .A2(n8009), .ZN(n7381) );
  XNOR2_X1 U9094 ( .A(n7382), .B(n7381), .ZN(n10181) );
  INV_X1 U9095 ( .A(n9859), .ZN(n8081) );
  NAND2_X1 U9096 ( .A1(n10181), .A2(n8081), .ZN(n7383) );
  AND2_X1 U9097 ( .A1(n7384), .A2(n7383), .ZN(n10183) );
  INV_X1 U9098 ( .A(n8297), .ZN(n8087) );
  AOI21_X1 U9099 ( .B1(n10085), .B2(n7499), .A(n9810), .ZN(n7385) );
  NAND2_X1 U9100 ( .A1(n7385), .A2(n10073), .ZN(n10178) );
  AOI22_X1 U9101 ( .A1(n10121), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7493), .B2(
        n10096), .ZN(n7387) );
  NAND2_X1 U9102 ( .A1(n10094), .A2(n7499), .ZN(n7386) );
  OAI211_X1 U9103 ( .C1(n10178), .C2(n9847), .A(n7387), .B(n7386), .ZN(n7388)
         );
  AOI21_X1 U9104 ( .B1(n10181), .B2(n8087), .A(n7388), .ZN(n7389) );
  OAI21_X1 U9105 ( .B1(n10183), .B2(n10121), .A(n7389), .ZN(P1_U3286) );
  INV_X1 U9106 ( .A(n7390), .ZN(n8851) );
  INV_X1 U9107 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7391) );
  OAI222_X1 U9108 ( .A1(P1_U3086), .A2(n7392), .B1(n9949), .B2(n8851), .C1(
        n7391), .C2(n9952), .ZN(P1_U3334) );
  INV_X1 U9109 ( .A(n7393), .ZN(n10391) );
  OAI21_X1 U9110 ( .B1(n7395), .B2(n8653), .A(n7394), .ZN(n10392) );
  OAI21_X1 U9111 ( .B1(n7397), .B2(n4984), .A(n7396), .ZN(n7400) );
  OAI22_X1 U9112 ( .A1(n7398), .A2(n10348), .B1(n7536), .B2(n10346), .ZN(n7399) );
  AOI21_X1 U9113 ( .B1(n7400), .B2(n10350), .A(n7399), .ZN(n7401) );
  OAI21_X1 U9114 ( .B1(n10353), .B2(n10392), .A(n7401), .ZN(n10394) );
  OAI22_X1 U9115 ( .A1(n10392), .A2(n7403), .B1(n7402), .B2(n10343), .ZN(n7404) );
  NOR2_X1 U9116 ( .A1(n10394), .A2(n7404), .ZN(n7405) );
  MUX2_X1 U9117 ( .A(n7406), .B(n7405), .S(n10357), .Z(n7407) );
  OAI21_X1 U9118 ( .B1(n10391), .B2(n10334), .A(n7407), .ZN(P2_U3226) );
  XOR2_X1 U9119 ( .A(n7506), .B(n7505), .Z(n7410) );
  INV_X1 U9120 ( .A(n7408), .ZN(n7409) );
  NAND2_X1 U9121 ( .A1(n7410), .A2(n7409), .ZN(n7504) );
  OAI21_X1 U9122 ( .B1(n7410), .B2(n7409), .A(n7504), .ZN(n7418) );
  INV_X1 U9123 ( .A(n7411), .ZN(n7416) );
  AOI22_X1 U9124 ( .A1(n7412), .A2(n9996), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n7415) );
  NAND2_X1 U9125 ( .A1(n9492), .A2(n7413), .ZN(n7414) );
  OAI211_X1 U9126 ( .C1(n10003), .C2(n7416), .A(n7415), .B(n7414), .ZN(n7417)
         );
  AOI21_X1 U9127 ( .B1(n7418), .B2(n10000), .A(n7417), .ZN(n7419) );
  INV_X1 U9128 ( .A(n7419), .ZN(P1_U3227) );
  INV_X1 U9129 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7863) );
  INV_X1 U9130 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9131 ( .A1(n5636), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U9132 ( .A1(n7420), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7421) );
  OAI211_X1 U9133 ( .C1(n7423), .C2(n5188), .A(n7422), .B(n7421), .ZN(n7424)
         );
  INV_X1 U9134 ( .A(n7424), .ZN(n7425) );
  AND2_X1 U9135 ( .A1(n7426), .A2(n7425), .ZN(n8601) );
  NAND2_X1 U9136 ( .A1(n9097), .A2(P2_U3893), .ZN(n7427) );
  OAI21_X1 U9137 ( .B1(P2_U3893), .B2(n7863), .A(n7427), .ZN(P2_U3522) );
  OR2_X1 U9138 ( .A1(n7429), .A2(n7428), .ZN(n7431) );
  NAND2_X1 U9139 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  XNOR2_X1 U9140 ( .A(n7432), .B(n8773), .ZN(n7438) );
  NAND2_X1 U9141 ( .A1(n7434), .A2(n8773), .ZN(n7435) );
  NAND2_X1 U9142 ( .A1(n7433), .A2(n7435), .ZN(n10402) );
  AOI22_X1 U9143 ( .A1(n10326), .A2(n8967), .B1(n10328), .B2(n8965), .ZN(n7436) );
  OAI21_X1 U9144 ( .B1(n10402), .B2(n10353), .A(n7436), .ZN(n7437) );
  AOI21_X1 U9145 ( .B1(n7438), .B2(n10350), .A(n7437), .ZN(n10407) );
  OAI22_X1 U9146 ( .A1(n10357), .A2(n5288), .B1(n7531), .B2(n10343), .ZN(n7440) );
  NOR2_X1 U9147 ( .A1(n10402), .A2(n8812), .ZN(n7439) );
  AOI211_X1 U9148 ( .C1(n9226), .C2(n10403), .A(n7440), .B(n7439), .ZN(n7441)
         );
  OAI21_X1 U9149 ( .B1(n10339), .B2(n10407), .A(n7441), .ZN(P2_U3224) );
  INV_X1 U9150 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7444) );
  MUX2_X1 U9151 ( .A(n7444), .B(P1_REG2_REG_12__SCAN_IN), .S(n8107), .Z(n7445)
         );
  INV_X1 U9152 ( .A(n7445), .ZN(n7446) );
  OAI21_X1 U9153 ( .B1(n7447), .B2(n7446), .A(n8103), .ZN(n7454) );
  INV_X1 U9154 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10242) );
  MUX2_X1 U9155 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10242), .S(n8107), .Z(n7452) );
  OAI21_X1 U9156 ( .B1(n7355), .B2(n7449), .A(n7448), .ZN(n7450) );
  INV_X1 U9157 ( .A(n7450), .ZN(n7451) );
  NAND2_X1 U9158 ( .A1(n7452), .A2(n7451), .ZN(n8106) );
  OAI21_X1 U9159 ( .B1(n7452), .B2(n7451), .A(n8106), .ZN(n7453) );
  AOI22_X1 U9160 ( .A1(n10043), .A2(n7454), .B1(n10053), .B2(n7453), .ZN(n7457) );
  NAND2_X1 U9161 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8438) );
  INV_X1 U9162 ( .A(n8438), .ZN(n7455) );
  AOI21_X1 U9163 ( .B1(n10049), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7455), .ZN(
        n7456) );
  OAI211_X1 U9164 ( .C1(n7458), .C2(n9629), .A(n7457), .B(n7456), .ZN(P1_U3255) );
  INV_X1 U9165 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10434) );
  NOR2_X1 U9166 ( .A1(n7468), .A2(n7462), .ZN(n7463) );
  AOI22_X1 U9167 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8044), .B1(n8041), .B2(
        n7476), .ZN(n7464) );
  AOI21_X1 U9168 ( .B1(n4605), .B2(n7464), .A(n8040), .ZN(n7489) );
  AOI22_X1 U9169 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8041), .B1(n8044), .B2(
        n7477), .ZN(n7471) );
  OAI21_X1 U9170 ( .B1(n7466), .B2(n5266), .A(n7465), .ZN(n7467) );
  NAND2_X1 U9171 ( .A1(n7525), .A2(n7467), .ZN(n7469) );
  XNOR2_X1 U9172 ( .A(n7468), .B(n7467), .ZN(n7518) );
  NAND2_X1 U9173 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n7518), .ZN(n7517) );
  NAND2_X1 U9174 ( .A1(n7469), .A2(n7517), .ZN(n7470) );
  OAI21_X1 U9175 ( .B1(n7471), .B2(n7470), .A(n8043), .ZN(n7487) );
  MUX2_X1 U9176 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8049), .Z(n7472) );
  NOR2_X1 U9177 ( .A1(n7472), .A2(n7525), .ZN(n7475) );
  AOI21_X1 U9178 ( .B1(n7472), .B2(n7525), .A(n7475), .ZN(n7521) );
  INV_X1 U9179 ( .A(n7475), .ZN(n7482) );
  MUX2_X1 U9180 ( .A(n7477), .B(n7476), .S(n8049), .Z(n7478) );
  NAND2_X1 U9181 ( .A1(n7478), .A2(n8044), .ZN(n8046) );
  INV_X1 U9182 ( .A(n7478), .ZN(n7479) );
  NAND2_X1 U9183 ( .A1(n7479), .A2(n8041), .ZN(n7480) );
  NAND2_X1 U9184 ( .A1(n8046), .A2(n7480), .ZN(n7481) );
  AND3_X1 U9185 ( .A1(n7519), .A2(n7482), .A3(n7481), .ZN(n7483) );
  OAI21_X1 U9186 ( .B1(n8048), .B2(n7483), .A(n10272), .ZN(n7485) );
  INV_X1 U9187 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7956) );
  NOR2_X1 U9188 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7956), .ZN(n7569) );
  AOI21_X1 U9189 ( .B1(n10248), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7569), .ZN(
        n7484) );
  OAI211_X1 U9190 ( .C1(n10312), .C2(n8041), .A(n7485), .B(n7484), .ZN(n7486)
         );
  AOI21_X1 U9191 ( .B1(n7487), .B2(n10308), .A(n7486), .ZN(n7488) );
  OAI21_X1 U9192 ( .B1(n7489), .B2(n10283), .A(n7488), .ZN(P2_U3192) );
  AOI21_X1 U9193 ( .B1(n7492), .B2(n7491), .A(n7490), .ZN(n7501) );
  INV_X1 U9194 ( .A(n7493), .ZN(n7497) );
  AOI22_X1 U9195 ( .A1(n9473), .A2(n9508), .B1(n9474), .B2(n6034), .ZN(n7496)
         );
  OAI211_X1 U9196 ( .C1(n7497), .C2(n10003), .A(n7496), .B(n7495), .ZN(n7498)
         );
  AOI21_X1 U9197 ( .B1(n7499), .B2(n9492), .A(n7498), .ZN(n7500) );
  OAI21_X1 U9198 ( .B1(n7501), .B2(n9494), .A(n7500), .ZN(P1_U3213) );
  NOR2_X1 U9199 ( .A1(n7503), .A2(n7502), .ZN(n7508) );
  OAI21_X1 U9200 ( .B1(n7506), .B2(n7505), .A(n7504), .ZN(n7507) );
  XOR2_X1 U9201 ( .A(n7508), .B(n7507), .Z(n7514) );
  INV_X1 U9202 ( .A(n10082), .ZN(n7511) );
  OAI22_X1 U9203 ( .A1(n7509), .A2(n9991), .B1(n9992), .B2(n9989), .ZN(n10080)
         );
  AOI22_X1 U9204 ( .A1(n10080), .A2(n9996), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7510) );
  OAI21_X1 U9205 ( .B1(n7511), .B2(n10003), .A(n7510), .ZN(n7512) );
  AOI21_X1 U9206 ( .B1(n10083), .B2(n9492), .A(n7512), .ZN(n7513) );
  OAI21_X1 U9207 ( .B1(n7514), .B2(n9494), .A(n7513), .ZN(P1_U3239) );
  AOI21_X1 U9208 ( .B1(n10434), .B2(n7516), .A(n7515), .ZN(n7529) );
  OAI21_X1 U9209 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7518), .A(n7517), .ZN(
        n7527) );
  OAI21_X1 U9210 ( .B1(n7521), .B2(n7520), .A(n7519), .ZN(n7523) );
  AND2_X1 U9211 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7530) );
  INV_X1 U9212 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7594) );
  NOR2_X1 U9213 ( .A1(n10321), .A2(n7594), .ZN(n7522) );
  AOI211_X1 U9214 ( .C1(n10272), .C2(n7523), .A(n7530), .B(n7522), .ZN(n7524)
         );
  OAI21_X1 U9215 ( .B1(n7525), .B2(n10312), .A(n7524), .ZN(n7526) );
  AOI21_X1 U9216 ( .B1(n7527), .B2(n10308), .A(n7526), .ZN(n7528) );
  OAI21_X1 U9217 ( .B1(n7529), .B2(n10283), .A(n7528), .ZN(P2_U3191) );
  AOI21_X1 U9218 ( .B1(n8931), .B2(n8967), .A(n7530), .ZN(n7534) );
  INV_X1 U9219 ( .A(n7531), .ZN(n7532) );
  NAND2_X1 U9220 ( .A1(n8945), .A2(n7532), .ZN(n7533) );
  OAI211_X1 U9221 ( .C1(n8217), .C2(n8933), .A(n7534), .B(n7533), .ZN(n7552)
         );
  XNOR2_X1 U9222 ( .A(n10403), .B(n4527), .ZN(n7564) );
  XNOR2_X1 U9223 ( .A(n7564), .B(n8966), .ZN(n7550) );
  NAND2_X1 U9224 ( .A1(n7535), .A2(n7542), .ZN(n7538) );
  NAND2_X1 U9225 ( .A1(n7537), .A2(n7536), .ZN(n7539) );
  NAND2_X1 U9226 ( .A1(n7538), .A2(n7539), .ZN(n7549) );
  INV_X1 U9227 ( .A(n7539), .ZN(n7540) );
  AND2_X1 U9228 ( .A1(n7541), .A2(n7544), .ZN(n7546) );
  INV_X1 U9229 ( .A(n7542), .ZN(n7543) );
  INV_X1 U9230 ( .A(n7566), .ZN(n7548) );
  AOI211_X1 U9231 ( .C1(n7550), .C2(n7549), .A(n8953), .B(n7548), .ZN(n7551)
         );
  AOI211_X1 U9232 ( .C1(n10403), .C2(n8951), .A(n7552), .B(n7551), .ZN(n7553)
         );
  INV_X1 U9233 ( .A(n7553), .ZN(P2_U3171) );
  INV_X1 U9234 ( .A(n8661), .ZN(n7554) );
  OR2_X1 U9235 ( .A1(n8664), .A2(n7554), .ZN(n7556) );
  INV_X1 U9236 ( .A(n7556), .ZN(n8775) );
  XNOR2_X1 U9237 ( .A(n7555), .B(n8775), .ZN(n10409) );
  XNOR2_X1 U9238 ( .A(n7557), .B(n7556), .ZN(n7559) );
  OAI22_X1 U9239 ( .A1(n7567), .A2(n10348), .B1(n8168), .B2(n10346), .ZN(n7558) );
  AOI21_X1 U9240 ( .B1(n7559), .B2(n10350), .A(n7558), .ZN(n7560) );
  OAI21_X1 U9241 ( .B1(n10409), .B2(n10353), .A(n7560), .ZN(n10410) );
  NAND2_X1 U9242 ( .A1(n10410), .A2(n9211), .ZN(n7563) );
  OAI22_X1 U9243 ( .A1(n10357), .A2(n7477), .B1(n7571), .B2(n10343), .ZN(n7561) );
  AOI21_X1 U9244 ( .B1(n10412), .B2(n9226), .A(n7561), .ZN(n7562) );
  OAI211_X1 U9245 ( .C1(n10409), .C2(n8812), .A(n7563), .B(n7562), .ZN(
        P2_U3223) );
  NAND2_X1 U9246 ( .A1(n7564), .A2(n8966), .ZN(n7565) );
  XOR2_X1 U9247 ( .A(n8838), .B(n10412), .Z(n8165) );
  XOR2_X1 U9248 ( .A(n8166), .B(n8165), .Z(n7574) );
  NOR2_X1 U9249 ( .A1(n8948), .A2(n7567), .ZN(n7568) );
  AOI211_X1 U9250 ( .C1(n8944), .C2(n8964), .A(n7569), .B(n7568), .ZN(n7570)
         );
  OAI21_X1 U9251 ( .B1(n7571), .B2(n8221), .A(n7570), .ZN(n7572) );
  AOI21_X1 U9252 ( .B1(n10412), .B2(n8951), .A(n7572), .ZN(n7573) );
  OAI21_X1 U9253 ( .B1(n7574), .B2(n8953), .A(n7573), .ZN(P2_U3157) );
  INV_X1 U9254 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10446) );
  NOR2_X1 U9255 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7620) );
  NOR2_X1 U9256 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7617) );
  NOR2_X1 U9257 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7614) );
  NOR2_X1 U9258 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7611) );
  NOR2_X1 U9259 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7608) );
  NOR2_X1 U9260 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7606) );
  NOR2_X1 U9261 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7603) );
  NOR2_X1 U9262 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7600) );
  NOR2_X1 U9263 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7597) );
  NOR2_X1 U9264 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7593) );
  NOR2_X1 U9265 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7589) );
  NOR2_X1 U9266 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7587) );
  NOR2_X1 U9267 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7585) );
  NOR2_X1 U9268 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7583) );
  NAND2_X1 U9269 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7581) );
  INV_X1 U9270 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10294) );
  XNOR2_X1 U9271 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n10294), .ZN(n10477) );
  NAND2_X1 U9272 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7579) );
  AOI21_X1 U9273 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10441) );
  INV_X1 U9274 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U9275 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7575) );
  NOR2_X1 U9276 ( .A1(n7576), .A2(n7575), .ZN(n10442) );
  NOR2_X1 U9277 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10442), .ZN(n7577) );
  NOR2_X1 U9278 ( .A1(n10441), .A2(n7577), .ZN(n10467) );
  INV_X1 U9279 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10276) );
  XNOR2_X1 U9280 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n10276), .ZN(n10466) );
  NAND2_X1 U9281 ( .A1(n10467), .A2(n10466), .ZN(n7578) );
  NAND2_X1 U9282 ( .A1(n7579), .A2(n7578), .ZN(n10476) );
  NAND2_X1 U9283 ( .A1(n10477), .A2(n10476), .ZN(n7580) );
  NAND2_X1 U9284 ( .A1(n7581), .A2(n7580), .ZN(n10479) );
  XNOR2_X1 U9285 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10478) );
  NOR2_X1 U9286 ( .A1(n10479), .A2(n10478), .ZN(n7582) );
  NOR2_X1 U9287 ( .A1(n7583), .A2(n7582), .ZN(n10469) );
  XNOR2_X1 U9288 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10468) );
  NOR2_X1 U9289 ( .A1(n10469), .A2(n10468), .ZN(n7584) );
  NOR2_X1 U9290 ( .A1(n7585), .A2(n7584), .ZN(n10475) );
  INV_X1 U9291 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10322) );
  XOR2_X1 U9292 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10322), .Z(n10474) );
  NOR2_X1 U9293 ( .A1(n10475), .A2(n10474), .ZN(n7586) );
  NOR2_X1 U9294 ( .A1(n7587), .A2(n7586), .ZN(n10471) );
  XNOR2_X1 U9295 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10470) );
  NOR2_X1 U9296 ( .A1(n10471), .A2(n10470), .ZN(n7588) );
  NOR2_X1 U9297 ( .A1(n7589), .A2(n7588), .ZN(n10473) );
  INV_X1 U9298 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7591) );
  AOI22_X1 U9299 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n7591), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n7590), .ZN(n10472) );
  NOR2_X1 U9300 ( .A1(n10473), .A2(n10472), .ZN(n7592) );
  NOR2_X1 U9301 ( .A1(n7593), .A2(n7592), .ZN(n10465) );
  INV_X1 U9302 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7595) );
  AOI22_X1 U9303 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7595), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7594), .ZN(n10464) );
  NOR2_X1 U9304 ( .A1(n10465), .A2(n10464), .ZN(n7596) );
  NOR2_X1 U9305 ( .A1(n7597), .A2(n7596), .ZN(n10463) );
  INV_X1 U9306 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7598) );
  AOI22_X1 U9307 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7288), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7598), .ZN(n10462) );
  NOR2_X1 U9308 ( .A1(n10463), .A2(n10462), .ZN(n7599) );
  NOR2_X1 U9309 ( .A1(n7600), .A2(n7599), .ZN(n10461) );
  INV_X1 U9310 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7601) );
  INV_X1 U9311 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8053) );
  AOI22_X1 U9312 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7601), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n8053), .ZN(n10460) );
  NOR2_X1 U9313 ( .A1(n10461), .A2(n10460), .ZN(n7602) );
  NOR2_X1 U9314 ( .A1(n7603), .A2(n7602), .ZN(n10459) );
  INV_X1 U9315 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7604) );
  INV_X1 U9316 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8155) );
  AOI22_X1 U9317 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7604), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n8155), .ZN(n10458) );
  NOR2_X1 U9318 ( .A1(n10459), .A2(n10458), .ZN(n7605) );
  NOR2_X1 U9319 ( .A1(n7606), .A2(n7605), .ZN(n10457) );
  XNOR2_X1 U9320 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10456) );
  NOR2_X1 U9321 ( .A1(n10457), .A2(n10456), .ZN(n7607) );
  NOR2_X1 U9322 ( .A1(n7608), .A2(n7607), .ZN(n10455) );
  INV_X1 U9323 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7609) );
  INV_X1 U9324 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8381) );
  AOI22_X1 U9325 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7609), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n8381), .ZN(n10454) );
  NOR2_X1 U9326 ( .A1(n10455), .A2(n10454), .ZN(n7610) );
  NOR2_X1 U9327 ( .A1(n7611), .A2(n7610), .ZN(n10453) );
  INV_X1 U9328 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7612) );
  INV_X1 U9329 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8982) );
  AOI22_X1 U9330 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7612), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8982), .ZN(n10452) );
  NOR2_X1 U9331 ( .A1(n10453), .A2(n10452), .ZN(n7613) );
  NOR2_X1 U9332 ( .A1(n7614), .A2(n7613), .ZN(n10451) );
  INV_X1 U9333 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7615) );
  INV_X1 U9334 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9011) );
  AOI22_X1 U9335 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7615), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n9011), .ZN(n10450) );
  NOR2_X1 U9336 ( .A1(n10451), .A2(n10450), .ZN(n7616) );
  NOR2_X1 U9337 ( .A1(n7617), .A2(n7616), .ZN(n10449) );
  INV_X1 U9338 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7618) );
  INV_X1 U9339 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9034) );
  AOI22_X1 U9340 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7618), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n9034), .ZN(n10448) );
  NOR2_X1 U9341 ( .A1(n10449), .A2(n10448), .ZN(n7619) );
  NOR2_X1 U9342 ( .A1(n7620), .A2(n7619), .ZN(n10445) );
  NOR2_X1 U9343 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10445), .ZN(n7621) );
  NAND2_X1 U9344 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10445), .ZN(n10444) );
  OAI21_X1 U9345 ( .B1(n10446), .B2(n7621), .A(n10444), .ZN(n7981) );
  XOR2_X1 U9346 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_f115), .Z(n7977) );
  XOR2_X1 U9347 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f91), .Z(n7628) );
  AOI22_X1 U9348 ( .A1(SI_14_), .A2(keyinput_f18), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_f43), .ZN(n7622) );
  OAI221_X1 U9349 ( .B1(SI_14_), .B2(keyinput_f18), .C1(P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n7622), .ZN(n7627) );
  AOI22_X1 U9350 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_f113), .B1(SI_27_), 
        .B2(keyinput_f5), .ZN(n7623) );
  OAI221_X1 U9351 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_f113), .C1(SI_27_), .C2(keyinput_f5), .A(n7623), .ZN(n7626) );
  AOI22_X1 U9352 ( .A1(SI_6_), .A2(keyinput_f26), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n7624) );
  OAI221_X1 U9353 ( .B1(SI_6_), .B2(keyinput_f26), .C1(P2_REG3_REG_4__SCAN_IN), 
        .C2(keyinput_f52), .A(n7624), .ZN(n7625) );
  NOR4_X1 U9354 ( .A1(n7628), .A2(n7627), .A3(n7626), .A4(n7625), .ZN(n7656)
         );
  AOI22_X1 U9355 ( .A1(SI_20_), .A2(keyinput_f12), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n7629) );
  OAI221_X1 U9356 ( .B1(SI_20_), .B2(keyinput_f12), .C1(SI_21_), .C2(
        keyinput_f11), .A(n7629), .ZN(n7636) );
  AOI22_X1 U9357 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_f111), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .ZN(n7630) );
  OAI221_X1 U9358 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_f111), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_f68), .A(n7630), .ZN(n7635) );
  AOI22_X1 U9359 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_f81), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n7631) );
  OAI221_X1 U9360 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n7631), .ZN(n7634) );
  AOI22_X1 U9361 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n7632) );
  OAI221_X1 U9362 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n7632), .ZN(n7633) );
  NOR4_X1 U9363 ( .A1(n7636), .A2(n7635), .A3(n7634), .A4(n7633), .ZN(n7655)
         );
  AOI22_X1 U9364 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(keyinput_f51), .ZN(n7637) );
  OAI221_X1 U9365 ( .B1(SI_28_), .B2(keyinput_f4), .C1(P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n7637), .ZN(n7644) );
  AOI22_X1 U9366 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f117), .B1(SI_5_), 
        .B2(keyinput_f27), .ZN(n7638) );
  OAI221_X1 U9367 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f117), .C1(SI_5_), 
        .C2(keyinput_f27), .A(n7638), .ZN(n7643) );
  AOI22_X1 U9368 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        SI_22_), .B2(keyinput_f10), .ZN(n7639) );
  OAI221_X1 U9369 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        SI_22_), .C2(keyinput_f10), .A(n7639), .ZN(n7642) );
  AOI22_X1 U9370 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n7640) );
  OAI221_X1 U9371 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n7640), .ZN(n7641) );
  NOR4_X1 U9372 ( .A1(n7644), .A2(n7643), .A3(n7642), .A4(n7641), .ZN(n7654)
         );
  AOI22_X1 U9373 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n7645) );
  OAI221_X1 U9374 ( .B1(SI_25_), .B2(keyinput_f7), .C1(P2_REG3_REG_3__SCAN_IN), 
        .C2(keyinput_f40), .A(n7645), .ZN(n7652) );
  AOI22_X1 U9375 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_f35), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n7646) );
  OAI221_X1 U9376 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n7646), .ZN(n7651) );
  AOI22_X1 U9377 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_f112), .B1(SI_26_), 
        .B2(keyinput_f6), .ZN(n7647) );
  OAI221_X1 U9378 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_f112), .C1(SI_26_), .C2(keyinput_f6), .A(n7647), .ZN(n7650) );
  AOI22_X1 U9379 ( .A1(SI_17_), .A2(keyinput_f15), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n7648) );
  OAI221_X1 U9380 ( .B1(SI_17_), .B2(keyinput_f15), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n7648), .ZN(n7649) );
  NOR4_X1 U9381 ( .A1(n7652), .A2(n7651), .A3(n7650), .A4(n7649), .ZN(n7653)
         );
  NAND4_X1 U9382 ( .A1(n7656), .A2(n7655), .A3(n7654), .A4(n7653), .ZN(n7790)
         );
  AOI22_X1 U9383 ( .A1(SI_8_), .A2(keyinput_f24), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(keyinput_f41), .ZN(n7657) );
  OAI221_X1 U9384 ( .B1(SI_8_), .B2(keyinput_f24), .C1(P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n7657), .ZN(n7664) );
  AOI22_X1 U9385 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f101), .B1(SI_9_), 
        .B2(keyinput_f23), .ZN(n7658) );
  OAI221_X1 U9386 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f101), .C1(SI_9_), 
        .C2(keyinput_f23), .A(n7658), .ZN(n7663) );
  AOI22_X1 U9387 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f123), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_f97), .ZN(n7659) );
  OAI221_X1 U9388 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f123), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_f97), .A(n7659), .ZN(n7662) );
  AOI22_X1 U9389 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f119), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_f98), .ZN(n7660) );
  OAI221_X1 U9390 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f119), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_f98), .A(n7660), .ZN(n7661) );
  NOR4_X1 U9391 ( .A1(n7664), .A2(n7663), .A3(n7662), .A4(n7661), .ZN(n7692)
         );
  AOI22_X1 U9392 ( .A1(SI_13_), .A2(keyinput_f19), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n7665) );
  OAI221_X1 U9393 ( .B1(SI_13_), .B2(keyinput_f19), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n7665), .ZN(n7672) );
  AOI22_X1 U9394 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f103), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_f108), .ZN(n7666) );
  OAI221_X1 U9395 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f103), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_f108), .A(n7666), .ZN(n7671) );
  AOI22_X1 U9396 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_DATAO_REG_7__SCAN_IN), 
        .B2(keyinput_f89), .ZN(n7667) );
  OAI221_X1 U9397 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_f89), .A(n7667), .ZN(n7670) );
  AOI22_X1 U9398 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n7668) );
  OAI221_X1 U9399 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n7668), .ZN(n7669) );
  NOR4_X1 U9400 ( .A1(n7672), .A2(n7671), .A3(n7670), .A4(n7669), .ZN(n7691)
         );
  AOI22_X1 U9401 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f114), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .ZN(n7673) );
  OAI221_X1 U9402 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f114), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_f33), .A(n7673), .ZN(n7680) );
  AOI22_X1 U9403 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_f99), .B1(SI_18_), 
        .B2(keyinput_f14), .ZN(n7674) );
  OAI221_X1 U9404 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_f99), .C1(SI_18_), 
        .C2(keyinput_f14), .A(n7674), .ZN(n7679) );
  AOI22_X1 U9405 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_f126), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n7675) );
  OAI221_X1 U9406 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_f126), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n7675), .ZN(n7678) );
  AOI22_X1 U9407 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P1_IR_REG_10__SCAN_IN), 
        .B2(keyinput_f100), .ZN(n7676) );
  OAI221_X1 U9408 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P1_IR_REG_10__SCAN_IN), 
        .C2(keyinput_f100), .A(n7676), .ZN(n7677) );
  NOR4_X1 U9409 ( .A1(n7680), .A2(n7679), .A3(n7678), .A4(n7677), .ZN(n7690)
         );
  AOI22_X1 U9410 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f118), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n7681) );
  OAI221_X1 U9411 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f118), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n7681), .ZN(n7688) );
  AOI22_X1 U9412 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_f124), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_f122), .ZN(n7682) );
  OAI221_X1 U9413 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_f124), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_f122), .A(n7682), .ZN(n7687) );
  AOI22_X1 U9414 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_f127), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_f92), .ZN(n7683) );
  OAI221_X1 U9415 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_f127), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput_f92), .A(n7683), .ZN(n7686) );
  AOI22_X1 U9416 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_f78), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n7684) );
  OAI221_X1 U9417 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .C1(
        SI_23_), .C2(keyinput_f9), .A(n7684), .ZN(n7685) );
  NOR4_X1 U9418 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n7689)
         );
  NAND4_X1 U9419 ( .A1(n7692), .A2(n7691), .A3(n7690), .A4(n7689), .ZN(n7789)
         );
  AOI22_X1 U9420 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_f106), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n7693) );
  OAI221_X1 U9421 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_f106), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n7693), .ZN(n7702) );
  AOI22_X1 U9422 ( .A1(SI_0_), .A2(keyinput_f32), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(keyinput_f50), .ZN(n7694) );
  OAI221_X1 U9423 ( .B1(SI_0_), .B2(keyinput_f32), .C1(P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n7694), .ZN(n7701) );
  INV_X1 U9424 ( .A(SI_24_), .ZN(n7889) );
  INV_X1 U9425 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8930) );
  AOI22_X1 U9426 ( .A1(n7889), .A2(keyinput_f8), .B1(n8930), .B2(keyinput_f60), 
        .ZN(n7695) );
  OAI221_X1 U9427 ( .B1(n7889), .B2(keyinput_f8), .C1(n8930), .C2(keyinput_f60), .A(n7695), .ZN(n7700) );
  INV_X1 U9428 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7698) );
  AOI22_X1 U9429 ( .A1(n7698), .A2(keyinput_f42), .B1(keyinput_f3), .B2(n7697), 
        .ZN(n7696) );
  OAI221_X1 U9430 ( .B1(n7698), .B2(keyinput_f42), .C1(n7697), .C2(keyinput_f3), .A(n7696), .ZN(n7699) );
  NOR4_X1 U9431 ( .A1(n7702), .A2(n7701), .A3(n7700), .A4(n7699), .ZN(n7737)
         );
  AOI22_X1 U9432 ( .A1(n5210), .A2(keyinput_f49), .B1(keyinput_f72), .B2(n8177), .ZN(n7703) );
  OAI221_X1 U9433 ( .B1(n5210), .B2(keyinput_f49), .C1(n8177), .C2(
        keyinput_f72), .A(n7703), .ZN(n7712) );
  XNOR2_X1 U9434 ( .A(n7704), .B(keyinput_f30), .ZN(n7711) );
  INV_X1 U9435 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7890) );
  XNOR2_X1 U9436 ( .A(keyinput_f38), .B(n7890), .ZN(n7710) );
  XNOR2_X1 U9437 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_f95), .ZN(n7708) );
  XNOR2_X1 U9438 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n7707) );
  XNOR2_X1 U9439 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_f120), .ZN(n7706) );
  XNOR2_X1 U9440 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f110), .ZN(n7705) );
  NAND4_X1 U9441 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n7709)
         );
  NOR4_X1 U9442 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n7736)
         );
  INV_X1 U9443 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8380) );
  INV_X1 U9444 ( .A(SI_19_), .ZN(n7902) );
  AOI22_X1 U9445 ( .A1(n8380), .A2(keyinput_f37), .B1(keyinput_f13), .B2(n7902), .ZN(n7713) );
  OAI221_X1 U9446 ( .B1(n8380), .B2(keyinput_f37), .C1(n7902), .C2(
        keyinput_f13), .A(n7713), .ZN(n7721) );
  AOI22_X1 U9447 ( .A1(n5632), .A2(keyinput_f36), .B1(keyinput_f70), .B2(n8301), .ZN(n7714) );
  OAI221_X1 U9448 ( .B1(n5632), .B2(keyinput_f36), .C1(n8301), .C2(
        keyinput_f70), .A(n7714), .ZN(n7720) );
  XNOR2_X1 U9449 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_f55), .ZN(n7718)
         );
  XNOR2_X1 U9450 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_f102), .ZN(n7717) );
  XNOR2_X1 U9451 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_f77), .ZN(n7716)
         );
  XNOR2_X1 U9452 ( .A(SI_4_), .B(keyinput_f28), .ZN(n7715) );
  NAND4_X1 U9453 ( .A1(n7718), .A2(n7717), .A3(n7716), .A4(n7715), .ZN(n7719)
         );
  NOR3_X1 U9454 ( .A1(n7721), .A2(n7720), .A3(n7719), .ZN(n7735) );
  AOI22_X1 U9455 ( .A1(n9951), .A2(keyinput_f67), .B1(n5595), .B2(keyinput_f47), .ZN(n7722) );
  OAI221_X1 U9456 ( .B1(n9951), .B2(keyinput_f67), .C1(n5595), .C2(
        keyinput_f47), .A(n7722), .ZN(n7733) );
  INV_X1 U9457 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7725) );
  INV_X1 U9458 ( .A(SI_16_), .ZN(n7724) );
  AOI22_X1 U9459 ( .A1(n7725), .A2(keyinput_f93), .B1(n7724), .B2(keyinput_f16), .ZN(n7723) );
  OAI221_X1 U9460 ( .B1(n7725), .B2(keyinput_f93), .C1(n7724), .C2(
        keyinput_f16), .A(n7723), .ZN(n7732) );
  INV_X1 U9461 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7901) );
  AOI22_X1 U9462 ( .A1(n7901), .A2(keyinput_f62), .B1(keyinput_f22), .B2(n7727), .ZN(n7726) );
  OAI221_X1 U9463 ( .B1(n7901), .B2(keyinput_f62), .C1(n7727), .C2(
        keyinput_f22), .A(n7726), .ZN(n7731) );
  XOR2_X1 U9464 ( .A(n5362), .B(keyinput_f56), .Z(n7729) );
  XNOR2_X1 U9465 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f94), .ZN(n7728) );
  NAND2_X1 U9466 ( .A1(n7729), .A2(n7728), .ZN(n7730) );
  NOR4_X1 U9467 ( .A1(n7733), .A2(n7732), .A3(n7731), .A4(n7730), .ZN(n7734)
         );
  NAND4_X1 U9468 ( .A1(n7737), .A2(n7736), .A3(n7735), .A4(n7734), .ZN(n7788)
         );
  AOI22_X1 U9469 ( .A1(n10125), .A2(keyinput_f125), .B1(n7987), .B2(
        keyinput_f74), .ZN(n7738) );
  OAI221_X1 U9470 ( .B1(n10125), .B2(keyinput_f125), .C1(n7987), .C2(
        keyinput_f74), .A(n7738), .ZN(n7746) );
  AOI22_X1 U9471 ( .A1(n8154), .A2(keyinput_f46), .B1(keyinput_f73), .B2(n8068), .ZN(n7739) );
  OAI221_X1 U9472 ( .B1(n8154), .B2(keyinput_f46), .C1(n8068), .C2(
        keyinput_f73), .A(n7739), .ZN(n7745) );
  XNOR2_X1 U9473 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_f69), .ZN(n7743)
         );
  XNOR2_X1 U9474 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f96), .ZN(n7742) );
  XNOR2_X1 U9475 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_f71), .ZN(n7741)
         );
  XNOR2_X1 U9476 ( .A(SI_1_), .B(keyinput_f31), .ZN(n7740) );
  NAND4_X1 U9477 ( .A1(n7743), .A2(n7742), .A3(n7741), .A4(n7740), .ZN(n7744)
         );
  NOR3_X1 U9478 ( .A1(n7746), .A2(n7745), .A3(n7744), .ZN(n7786) );
  AOI22_X1 U9479 ( .A1(n7748), .A2(keyinput_f104), .B1(n7932), .B2(
        keyinput_f76), .ZN(n7747) );
  OAI221_X1 U9480 ( .B1(n7748), .B2(keyinput_f104), .C1(n7932), .C2(
        keyinput_f76), .A(n7747), .ZN(n7758) );
  XNOR2_X1 U9481 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_f116), .ZN(n7752) );
  XNOR2_X1 U9482 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_f85), .ZN(n7751)
         );
  XNOR2_X1 U9483 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f109), .ZN(n7750) );
  XNOR2_X1 U9484 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_f79), .ZN(n7749)
         );
  NAND4_X1 U9485 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n7757)
         );
  XNOR2_X1 U9486 ( .A(n7753), .B(keyinput_f105), .ZN(n7756) );
  XNOR2_X1 U9487 ( .A(n7754), .B(keyinput_f29), .ZN(n7755) );
  NOR4_X1 U9488 ( .A1(n7758), .A2(n7757), .A3(n7756), .A4(n7755), .ZN(n7785)
         );
  INV_X1 U9489 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7760) );
  AOI22_X1 U9490 ( .A1(n7863), .A2(keyinput_f65), .B1(n7760), .B2(keyinput_f54), .ZN(n7759) );
  OAI221_X1 U9491 ( .B1(n7863), .B2(keyinput_f65), .C1(n7760), .C2(
        keyinput_f54), .A(n7759), .ZN(n7770) );
  AOI22_X1 U9492 ( .A1(n7917), .A2(keyinput_f82), .B1(n7762), .B2(keyinput_f17), .ZN(n7761) );
  OAI221_X1 U9493 ( .B1(n7917), .B2(keyinput_f82), .C1(n7762), .C2(
        keyinput_f17), .A(n7761), .ZN(n7765) );
  INV_X1 U9494 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9985) );
  XNOR2_X1 U9495 ( .A(n9985), .B(keyinput_f0), .ZN(n7764) );
  XOR2_X1 U9496 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f121), .Z(n7763) );
  OR3_X1 U9497 ( .A1(n7765), .A2(n7764), .A3(n7763), .ZN(n7769) );
  AOI22_X1 U9498 ( .A1(n10015), .A2(keyinput_f90), .B1(n7767), .B2(
        keyinput_f86), .ZN(n7766) );
  OAI221_X1 U9499 ( .B1(n10015), .B2(keyinput_f90), .C1(n7767), .C2(
        keyinput_f86), .A(n7766), .ZN(n7768) );
  NOR3_X1 U9500 ( .A1(n7770), .A2(n7769), .A3(n7768), .ZN(n7784) );
  AOI22_X1 U9501 ( .A1(n7956), .A2(keyinput_f39), .B1(keyinput_f88), .B2(n7772), .ZN(n7771) );
  OAI221_X1 U9502 ( .B1(n7956), .B2(keyinput_f39), .C1(n7772), .C2(
        keyinput_f88), .A(n7771), .ZN(n7782) );
  INV_X1 U9503 ( .A(SI_7_), .ZN(n7774) );
  AOI22_X1 U9504 ( .A1(n7881), .A2(keyinput_f87), .B1(keyinput_f25), .B2(n7774), .ZN(n7773) );
  OAI221_X1 U9505 ( .B1(n7881), .B2(keyinput_f87), .C1(n7774), .C2(
        keyinput_f25), .A(n7773), .ZN(n7781) );
  AOI22_X1 U9506 ( .A1(n7776), .A2(keyinput_f107), .B1(n7880), .B2(
        keyinput_f84), .ZN(n7775) );
  OAI221_X1 U9507 ( .B1(n7776), .B2(keyinput_f107), .C1(n7880), .C2(
        keyinput_f84), .A(n7775), .ZN(n7780) );
  XNOR2_X1 U9508 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_f59), .ZN(n7778) );
  XNOR2_X1 U9509 ( .A(SI_12_), .B(keyinput_f20), .ZN(n7777) );
  NAND2_X1 U9510 ( .A1(n7778), .A2(n7777), .ZN(n7779) );
  NOR4_X1 U9511 ( .A1(n7782), .A2(n7781), .A3(n7780), .A4(n7779), .ZN(n7783)
         );
  NAND4_X1 U9512 ( .A1(n7786), .A2(n7785), .A3(n7784), .A4(n7783), .ZN(n7787)
         );
  NOR4_X1 U9513 ( .A1(n7790), .A2(n7789), .A3(n7788), .A4(n7787), .ZN(n7976)
         );
  XOR2_X1 U9514 ( .A(keyinput_g121), .B(P1_IR_REG_31__SCAN_IN), .Z(n7797) );
  AOI22_X1 U9515 ( .A1(SI_8_), .A2(keyinput_g24), .B1(SI_16_), .B2(
        keyinput_g16), .ZN(n7791) );
  OAI221_X1 U9516 ( .B1(SI_8_), .B2(keyinput_g24), .C1(SI_16_), .C2(
        keyinput_g16), .A(n7791), .ZN(n7796) );
  AOI22_X1 U9517 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_g127), .B1(SI_7_), 
        .B2(keyinput_g25), .ZN(n7792) );
  OAI221_X1 U9518 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_g127), .C1(SI_7_), 
        .C2(keyinput_g25), .A(n7792), .ZN(n7795) );
  AOI22_X1 U9519 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        SI_20_), .B2(keyinput_g12), .ZN(n7793) );
  OAI221_X1 U9520 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        SI_20_), .C2(keyinput_g12), .A(n7793), .ZN(n7794) );
  NOR4_X1 U9521 ( .A1(n7797), .A2(n7796), .A3(n7795), .A4(n7794), .ZN(n7825)
         );
  AOI22_X1 U9522 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        SI_22_), .B2(keyinput_g10), .ZN(n7798) );
  OAI221_X1 U9523 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        SI_22_), .C2(keyinput_g10), .A(n7798), .ZN(n7805) );
  AOI22_X1 U9524 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g110), .B1(SI_1_), 
        .B2(keyinput_g31), .ZN(n7799) );
  OAI221_X1 U9525 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g110), .C1(SI_1_), 
        .C2(keyinput_g31), .A(n7799), .ZN(n7804) );
  AOI22_X1 U9526 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .ZN(n7800) );
  OAI221_X1 U9527 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_g83), .A(n7800), .ZN(n7803) );
  AOI22_X1 U9528 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_g120), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .ZN(n7801) );
  OAI221_X1 U9529 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_g120), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_g78), .A(n7801), .ZN(n7802) );
  NOR4_X1 U9530 ( .A1(n7805), .A2(n7804), .A3(n7803), .A4(n7802), .ZN(n7824)
         );
  AOI22_X1 U9531 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g104), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .ZN(n7806) );
  OAI221_X1 U9532 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g104), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_g67), .A(n7806), .ZN(n7813) );
  AOI22_X1 U9533 ( .A1(SI_12_), .A2(keyinput_g20), .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n7807) );
  OAI221_X1 U9534 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n7807), .ZN(n7812) );
  AOI22_X1 U9535 ( .A1(SI_26_), .A2(keyinput_g6), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n7808) );
  OAI221_X1 U9536 ( .B1(SI_26_), .B2(keyinput_g6), .C1(P2_REG3_REG_9__SCAN_IN), 
        .C2(keyinput_g53), .A(n7808), .ZN(n7811) );
  AOI22_X1 U9537 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_g118), .B1(SI_29_), 
        .B2(keyinput_g3), .ZN(n7809) );
  OAI221_X1 U9538 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_g118), .C1(SI_29_), .C2(keyinput_g3), .A(n7809), .ZN(n7810) );
  NOR4_X1 U9539 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n7823)
         );
  AOI22_X1 U9540 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_g94), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_g101), .ZN(n7814) );
  OAI221_X1 U9541 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_g94), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_g101), .A(n7814), .ZN(n7821) );
  AOI22_X1 U9542 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g93), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_g89), .ZN(n7815) );
  OAI221_X1 U9543 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g93), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_g89), .A(n7815), .ZN(n7820) );
  AOI22_X1 U9544 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_g114), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_g100), .ZN(n7816) );
  OAI221_X1 U9545 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_g114), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g100), .A(n7816), .ZN(n7819) );
  AOI22_X1 U9546 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .ZN(n7817) );
  OAI221_X1 U9547 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_g35), .A(n7817), .ZN(n7818) );
  NOR4_X1 U9548 ( .A1(n7821), .A2(n7820), .A3(n7819), .A4(n7818), .ZN(n7822)
         );
  NAND4_X1 U9549 ( .A1(n7825), .A2(n7824), .A3(n7823), .A4(n7822), .ZN(n7971)
         );
  AOI22_X1 U9550 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_g80), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .ZN(n7826) );
  OAI221_X1 U9551 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_g52), .A(n7826), .ZN(n7833) );
  AOI22_X1 U9552 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n7827) );
  OAI221_X1 U9553 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n7827), .ZN(n7832) );
  AOI22_X1 U9554 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n7828) );
  OAI221_X1 U9555 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n7828), .ZN(n7831) );
  AOI22_X1 U9556 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n7829) );
  OAI221_X1 U9557 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n7829), .ZN(n7830) );
  NOR4_X1 U9558 ( .A1(n7833), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n7861)
         );
  AOI22_X1 U9559 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_g91), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .ZN(n7834) );
  OAI221_X1 U9560 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_g91), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_g54), .A(n7834), .ZN(n7841) );
  AOI22_X1 U9561 ( .A1(SI_2_), .A2(keyinput_g30), .B1(SI_25_), .B2(keyinput_g7), .ZN(n7835) );
  OAI221_X1 U9562 ( .B1(SI_2_), .B2(keyinput_g30), .C1(SI_25_), .C2(
        keyinput_g7), .A(n7835), .ZN(n7840) );
  AOI22_X1 U9563 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_g107), .B1(SI_18_), 
        .B2(keyinput_g14), .ZN(n7836) );
  OAI221_X1 U9564 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_g107), .C1(SI_18_), .C2(keyinput_g14), .A(n7836), .ZN(n7839) );
  AOI22_X1 U9565 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_g123), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_g122), .ZN(n7837) );
  OAI221_X1 U9566 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_g123), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_g122), .A(n7837), .ZN(n7838) );
  NOR4_X1 U9567 ( .A1(n7841), .A2(n7840), .A3(n7839), .A4(n7838), .ZN(n7860)
         );
  AOI22_X1 U9568 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_g124), .B1(SI_10_), 
        .B2(keyinput_g22), .ZN(n7842) );
  OAI221_X1 U9569 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_g124), .C1(SI_10_), 
        .C2(keyinput_g22), .A(n7842), .ZN(n7849) );
  AOI22_X1 U9570 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g109), .B1(SI_21_), 
        .B2(keyinput_g11), .ZN(n7843) );
  OAI221_X1 U9571 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g109), .C1(SI_21_), .C2(keyinput_g11), .A(n7843), .ZN(n7848) );
  AOI22_X1 U9572 ( .A1(SI_0_), .A2(keyinput_g32), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(keyinput_g42), .ZN(n7844) );
  OAI221_X1 U9573 ( .B1(SI_0_), .B2(keyinput_g32), .C1(P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n7844), .ZN(n7847) );
  AOI22_X1 U9574 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_g126), .B1(SI_27_), 
        .B2(keyinput_g5), .ZN(n7845) );
  OAI221_X1 U9575 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_g126), .C1(SI_27_), 
        .C2(keyinput_g5), .A(n7845), .ZN(n7846) );
  NOR4_X1 U9576 ( .A1(n7849), .A2(n7848), .A3(n7847), .A4(n7846), .ZN(n7859)
         );
  AOI22_X1 U9577 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_g90), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .ZN(n7850) );
  OAI221_X1 U9578 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_g90), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_g70), .A(n7850), .ZN(n7857) );
  AOI22_X1 U9579 ( .A1(SI_15_), .A2(keyinput_g17), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .ZN(n7851) );
  OAI221_X1 U9580 ( .B1(SI_15_), .B2(keyinput_g17), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_g79), .A(n7851), .ZN(n7856) );
  AOI22_X1 U9581 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_g105), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .ZN(n7852) );
  OAI221_X1 U9582 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_g105), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n7852), .ZN(n7855) );
  AOI22_X1 U9583 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_g96), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .ZN(n7853) );
  OAI221_X1 U9584 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_g96), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n7853), .ZN(n7854) );
  NOR4_X1 U9585 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n7858)
         );
  NAND4_X1 U9586 ( .A1(n7861), .A2(n7860), .A3(n7859), .A4(n7858), .ZN(n7970)
         );
  INV_X1 U9587 ( .A(P2_B_REG_SCAN_IN), .ZN(n7864) );
  AOI22_X1 U9588 ( .A1(n7864), .A2(keyinput_g64), .B1(keyinput_g65), .B2(n7863), .ZN(n7862) );
  OAI221_X1 U9589 ( .B1(n7864), .B2(keyinput_g64), .C1(n7863), .C2(
        keyinput_g65), .A(n7862), .ZN(n7876) );
  INV_X1 U9590 ( .A(SI_13_), .ZN(n7867) );
  AOI22_X1 U9591 ( .A1(n7867), .A2(keyinput_g19), .B1(n7866), .B2(keyinput_g15), .ZN(n7865) );
  OAI221_X1 U9592 ( .B1(n7867), .B2(keyinput_g19), .C1(n7866), .C2(
        keyinput_g15), .A(n7865), .ZN(n7875) );
  INV_X1 U9593 ( .A(SI_23_), .ZN(n7868) );
  XOR2_X1 U9594 ( .A(n7868), .B(keyinput_g9), .Z(n7873) );
  XNOR2_X1 U9595 ( .A(n7869), .B(keyinput_g66), .ZN(n7872) );
  XNOR2_X1 U9596 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_g59), .ZN(n7871) );
  XNOR2_X1 U9597 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_g116), .ZN(n7870) );
  NAND4_X1 U9598 ( .A1(n7873), .A2(n7872), .A3(n7871), .A4(n7870), .ZN(n7874)
         );
  NOR3_X1 U9599 ( .A1(n7876), .A2(n7875), .A3(n7874), .ZN(n7915) );
  AOI22_X1 U9600 ( .A1(n9985), .A2(keyinput_g0), .B1(n10125), .B2(
        keyinput_g125), .ZN(n7877) );
  OAI221_X1 U9601 ( .B1(n9985), .B2(keyinput_g0), .C1(n10125), .C2(
        keyinput_g125), .A(n7877), .ZN(n7887) );
  AOI22_X1 U9602 ( .A1(n5595), .A2(keyinput_g47), .B1(P2_U3151), .B2(
        keyinput_g34), .ZN(n7878) );
  OAI221_X1 U9603 ( .B1(n5595), .B2(keyinput_g47), .C1(P2_U3151), .C2(
        keyinput_g34), .A(n7878), .ZN(n7886) );
  AOI22_X1 U9604 ( .A1(n7881), .A2(keyinput_g87), .B1(n7880), .B2(keyinput_g84), .ZN(n7879) );
  OAI221_X1 U9605 ( .B1(n7881), .B2(keyinput_g87), .C1(n7880), .C2(
        keyinput_g84), .A(n7879), .ZN(n7885) );
  XNOR2_X1 U9606 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_g74), .ZN(n7883)
         );
  XNOR2_X1 U9607 ( .A(SI_3_), .B(keyinput_g29), .ZN(n7882) );
  NAND2_X1 U9608 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  NOR4_X1 U9609 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n7914)
         );
  AOI22_X1 U9610 ( .A1(n7890), .A2(keyinput_g38), .B1(keyinput_g8), .B2(n7889), 
        .ZN(n7888) );
  OAI221_X1 U9611 ( .B1(n7890), .B2(keyinput_g38), .C1(n7889), .C2(keyinput_g8), .A(n7888), .ZN(n7899) );
  INV_X1 U9612 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8504) );
  AOI22_X1 U9613 ( .A1(n8504), .A2(keyinput_g68), .B1(n7892), .B2(keyinput_g4), 
        .ZN(n7891) );
  OAI221_X1 U9614 ( .B1(n8504), .B2(keyinput_g68), .C1(n7892), .C2(keyinput_g4), .A(n7891), .ZN(n7898) );
  XNOR2_X1 U9615 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_g63), .ZN(n7896)
         );
  XNOR2_X1 U9616 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g117), .ZN(n7895) );
  XNOR2_X1 U9617 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_g119), .ZN(n7894) );
  XNOR2_X1 U9618 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_g103), .ZN(n7893) );
  NAND4_X1 U9619 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n7897)
         );
  NOR3_X1 U9620 ( .A1(n7899), .A2(n7898), .A3(n7897), .ZN(n7913) );
  AOI22_X1 U9621 ( .A1(n7902), .A2(keyinput_g13), .B1(n7901), .B2(keyinput_g62), .ZN(n7900) );
  OAI221_X1 U9622 ( .B1(n7902), .B2(keyinput_g13), .C1(n7901), .C2(
        keyinput_g62), .A(n7900), .ZN(n7911) );
  AOI22_X1 U9623 ( .A1(n8214), .A2(keyinput_g71), .B1(keyinput_g21), .B2(n7904), .ZN(n7903) );
  OAI221_X1 U9624 ( .B1(n8214), .B2(keyinput_g71), .C1(n7904), .C2(
        keyinput_g21), .A(n7903), .ZN(n7910) );
  XNOR2_X1 U9625 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_g51), .ZN(n7908)
         );
  XNOR2_X1 U9626 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_g113), .ZN(n7907) );
  XNOR2_X1 U9627 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g111), .ZN(n7906) );
  XNOR2_X1 U9628 ( .A(SI_5_), .B(keyinput_g27), .ZN(n7905) );
  NAND4_X1 U9629 ( .A1(n7908), .A2(n7907), .A3(n7906), .A4(n7905), .ZN(n7909)
         );
  NOR3_X1 U9630 ( .A1(n7911), .A2(n7910), .A3(n7909), .ZN(n7912) );
  NAND4_X1 U9631 ( .A1(n7915), .A2(n7914), .A3(n7913), .A4(n7912), .ZN(n7969)
         );
  AOI22_X1 U9632 ( .A1(n5210), .A2(keyinput_g49), .B1(keyinput_g82), .B2(n7917), .ZN(n7916) );
  OAI221_X1 U9633 ( .B1(n5210), .B2(keyinput_g49), .C1(n7917), .C2(
        keyinput_g82), .A(n7916), .ZN(n7929) );
  INV_X1 U9634 ( .A(SI_30_), .ZN(n7920) );
  INV_X1 U9635 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7919) );
  AOI22_X1 U9636 ( .A1(n7920), .A2(keyinput_g2), .B1(n7919), .B2(keyinput_g99), 
        .ZN(n7918) );
  OAI221_X1 U9637 ( .B1(n7920), .B2(keyinput_g2), .C1(n7919), .C2(keyinput_g99), .A(n7918), .ZN(n7928) );
  AOI22_X1 U9638 ( .A1(n7923), .A2(keyinput_g55), .B1(keyinput_g23), .B2(n7922), .ZN(n7921) );
  OAI221_X1 U9639 ( .B1(n7923), .B2(keyinput_g55), .C1(n7922), .C2(
        keyinput_g23), .A(n7921), .ZN(n7927) );
  XNOR2_X1 U9640 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g95), .ZN(n7925) );
  XNOR2_X1 U9641 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_g50), .ZN(n7924)
         );
  NAND2_X1 U9642 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  NOR4_X1 U9643 ( .A1(n7929), .A2(n7928), .A3(n7927), .A4(n7926), .ZN(n7967)
         );
  AOI22_X1 U9644 ( .A1(n7932), .A2(keyinput_g76), .B1(keyinput_g98), .B2(n7931), .ZN(n7930) );
  OAI221_X1 U9645 ( .B1(n7932), .B2(keyinput_g76), .C1(n7931), .C2(
        keyinput_g98), .A(n7930), .ZN(n7942) );
  AOI22_X1 U9646 ( .A1(n7935), .A2(keyinput_g92), .B1(n7934), .B2(keyinput_g43), .ZN(n7933) );
  OAI221_X1 U9647 ( .B1(n7935), .B2(keyinput_g92), .C1(n7934), .C2(
        keyinput_g43), .A(n7933), .ZN(n7941) );
  XNOR2_X1 U9648 ( .A(SI_14_), .B(keyinput_g18), .ZN(n7939) );
  XNOR2_X1 U9649 ( .A(SI_4_), .B(keyinput_g28), .ZN(n7938) );
  XNOR2_X1 U9650 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_g112), .ZN(n7937) );
  XNOR2_X1 U9651 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .ZN(n7936)
         );
  NAND4_X1 U9652 ( .A1(n7939), .A2(n7938), .A3(n7937), .A4(n7936), .ZN(n7940)
         );
  NOR3_X1 U9653 ( .A1(n7942), .A2(n7941), .A3(n7940), .ZN(n7966) );
  INV_X1 U9654 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8052) );
  AOI22_X1 U9655 ( .A1(n8052), .A2(keyinput_g58), .B1(keyinput_g61), .B2(n7944), .ZN(n7943) );
  OAI221_X1 U9656 ( .B1(n8052), .B2(keyinput_g58), .C1(n7944), .C2(
        keyinput_g61), .A(n7943), .ZN(n7952) );
  AOI22_X1 U9657 ( .A1(n8930), .A2(keyinput_g60), .B1(keyinput_g77), .B2(n8848), .ZN(n7945) );
  OAI221_X1 U9658 ( .B1(n8930), .B2(keyinput_g60), .C1(n8848), .C2(
        keyinput_g77), .A(n7945), .ZN(n7951) );
  AOI22_X1 U9659 ( .A1(n8068), .A2(keyinput_g73), .B1(n8359), .B2(keyinput_g69), .ZN(n7946) );
  OAI221_X1 U9660 ( .B1(n8068), .B2(keyinput_g73), .C1(n8359), .C2(
        keyinput_g69), .A(n7946), .ZN(n7950) );
  XNOR2_X1 U9661 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g102), .ZN(n7948) );
  XNOR2_X1 U9662 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_g45), .ZN(n7947)
         );
  NAND2_X1 U9663 ( .A1(n7948), .A2(n7947), .ZN(n7949) );
  NOR4_X1 U9664 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n7965)
         );
  INV_X1 U9665 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7954) );
  AOI22_X1 U9666 ( .A1(n5362), .A2(keyinput_g56), .B1(keyinput_g106), .B2(
        n7954), .ZN(n7953) );
  OAI221_X1 U9667 ( .B1(n5362), .B2(keyinput_g56), .C1(n7954), .C2(
        keyinput_g106), .A(n7953), .ZN(n7963) );
  AOI22_X1 U9668 ( .A1(n8177), .A2(keyinput_g72), .B1(n7956), .B2(keyinput_g39), .ZN(n7955) );
  OAI221_X1 U9669 ( .B1(n8177), .B2(keyinput_g72), .C1(n7956), .C2(
        keyinput_g39), .A(n7955), .ZN(n7962) );
  XNOR2_X1 U9670 ( .A(SI_6_), .B(keyinput_g26), .ZN(n7960) );
  XNOR2_X1 U9671 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_g40), .ZN(n7959) );
  XNOR2_X1 U9672 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g108), .ZN(n7958) );
  XNOR2_X1 U9673 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g97), .ZN(n7957) );
  NAND4_X1 U9674 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n7957), .ZN(n7961)
         );
  NOR3_X1 U9675 ( .A1(n7963), .A2(n7962), .A3(n7961), .ZN(n7964) );
  NAND4_X1 U9676 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n7968)
         );
  NOR4_X1 U9677 ( .A1(n7971), .A2(n7970), .A3(n7969), .A4(n7968), .ZN(n7974)
         );
  XNOR2_X1 U9678 ( .A(n7972), .B(keyinput_g115), .ZN(n7973) );
  NOR2_X1 U9679 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  OAI21_X1 U9680 ( .B1(n7977), .B2(n7976), .A(n7975), .ZN(n7979) );
  XNOR2_X1 U9681 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7978) );
  XNOR2_X1 U9682 ( .A(n7979), .B(n7978), .ZN(n7980) );
  XNOR2_X1 U9683 ( .A(n7981), .B(n7980), .ZN(ADD_1068_U4) );
  INV_X1 U9684 ( .A(n7982), .ZN(n7986) );
  OAI222_X1 U9685 ( .A1(P2_U3151), .A2(n7984), .B1(n9355), .B2(n7986), .C1(
        n7983), .C2(n8849), .ZN(P2_U3273) );
  OAI222_X1 U9686 ( .A1(n9952), .A2(n7987), .B1(n9949), .B2(n7986), .C1(
        P1_U3086), .C2(n7985), .ZN(P1_U3333) );
  XNOR2_X1 U9687 ( .A(n7988), .B(n8776), .ZN(n10415) );
  INV_X1 U9688 ( .A(n10415), .ZN(n8000) );
  NAND2_X1 U9689 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U9690 ( .A1(n7991), .A2(n8776), .ZN(n7992) );
  NAND3_X1 U9691 ( .A1(n7993), .A2(n10350), .A3(n7992), .ZN(n7995) );
  AOI22_X1 U9692 ( .A1(n8963), .A2(n10328), .B1(n10326), .B2(n8965), .ZN(n7994) );
  NAND2_X1 U9693 ( .A1(n7995), .A2(n7994), .ZN(n10420) );
  NAND2_X1 U9694 ( .A1(n10420), .A2(n9211), .ZN(n7999) );
  OAI22_X1 U9695 ( .A1(n10357), .A2(n7996), .B1(n8222), .B2(n10343), .ZN(n7997) );
  AOI21_X1 U9696 ( .B1(n10417), .B2(n9226), .A(n7997), .ZN(n7998) );
  OAI211_X1 U9697 ( .C1(n8000), .C2(n9229), .A(n7999), .B(n7998), .ZN(P2_U3222) );
  XNOR2_X1 U9698 ( .A(n8001), .B(n8070), .ZN(n8004) );
  OR2_X1 U9699 ( .A1(n9990), .A2(n9991), .ZN(n8003) );
  OR2_X1 U9700 ( .A1(n8123), .A2(n9989), .ZN(n8002) );
  NAND2_X1 U9701 ( .A1(n8003), .A2(n8002), .ZN(n8465) );
  AOI21_X1 U9702 ( .B1(n8004), .B2(n10092), .A(n8465), .ZN(n10198) );
  NAND2_X1 U9703 ( .A1(n9992), .A2(n10179), .ZN(n8008) );
  NAND2_X1 U9704 ( .A1(n8005), .A2(n8008), .ZN(n8010) );
  AND2_X1 U9705 ( .A1(n10084), .A2(n8010), .ZN(n10068) );
  INV_X1 U9706 ( .A(n10071), .ZN(n8011) );
  NAND2_X1 U9707 ( .A1(n5099), .A2(n8010), .ZN(n10069) );
  NAND2_X1 U9708 ( .A1(n6066), .A2(n10187), .ZN(n8034) );
  INV_X1 U9709 ( .A(n9430), .ZN(n10193) );
  NAND2_X1 U9710 ( .A1(n10193), .A2(n9990), .ZN(n8014) );
  AND2_X1 U9711 ( .A1(n8034), .A2(n8014), .ZN(n8018) );
  INV_X1 U9712 ( .A(n8014), .ZN(n8017) );
  NAND2_X1 U9713 ( .A1(n8016), .A2(n8015), .ZN(n8036) );
  XNOR2_X1 U9714 ( .A(n8071), .B(n8070), .ZN(n10201) );
  NAND2_X1 U9715 ( .A1(n10201), .A2(n10104), .ZN(n8024) );
  INV_X1 U9716 ( .A(n8082), .ZN(n8019) );
  OAI211_X1 U9717 ( .C1(n10199), .C2(n8029), .A(n8019), .B(n10099), .ZN(n10197) );
  INV_X1 U9718 ( .A(n10197), .ZN(n8022) );
  AOI22_X1 U9719 ( .A1(n10121), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8461), .B2(
        n10096), .ZN(n8020) );
  OAI21_X1 U9720 ( .B1(n10199), .B2(n9815), .A(n8020), .ZN(n8021) );
  AOI21_X1 U9721 ( .B1(n8022), .B2(n10103), .A(n8021), .ZN(n8023) );
  OAI211_X1 U9722 ( .C1(n10121), .C2(n10198), .A(n8024), .B(n8023), .ZN(
        P1_U3283) );
  INV_X1 U9723 ( .A(n8025), .ZN(n10061) );
  NOR3_X1 U9724 ( .A1(n10062), .A2(n10061), .A3(n10071), .ZN(n10060) );
  NOR2_X1 U9725 ( .A1(n10060), .A2(n8026), .ZN(n8027) );
  XOR2_X1 U9726 ( .A(n8036), .B(n8027), .Z(n8028) );
  AOI22_X1 U9727 ( .A1(n8028), .A2(n10092), .B1(n9794), .B2(n9508), .ZN(n10192) );
  INV_X1 U9728 ( .A(n8428), .ZN(n9506) );
  AOI211_X1 U9729 ( .C1(n9430), .C2(n10074), .A(n9810), .B(n8029), .ZN(n8030)
         );
  AOI21_X1 U9730 ( .B1(n9834), .B2(n9506), .A(n8030), .ZN(n10191) );
  INV_X1 U9731 ( .A(n10191), .ZN(n8033) );
  AOI22_X1 U9732 ( .A1(n10121), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9429), .B2(
        n10096), .ZN(n8031) );
  OAI21_X1 U9733 ( .B1(n10193), .B2(n9815), .A(n8031), .ZN(n8032) );
  AOI21_X1 U9734 ( .B1(n8033), .B2(n10103), .A(n8032), .ZN(n8039) );
  NAND2_X1 U9735 ( .A1(n8035), .A2(n8034), .ZN(n8037) );
  XNOR2_X1 U9736 ( .A(n8037), .B(n8036), .ZN(n10195) );
  NAND2_X1 U9737 ( .A1(n10195), .A2(n10104), .ZN(n8038) );
  OAI211_X1 U9738 ( .C1(n10192), .C2(n10121), .A(n8039), .B(n8038), .ZN(
        P1_U3284) );
  INV_X1 U9739 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10438) );
  AOI21_X1 U9740 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n8041), .A(n8040), .ZN(
        n8133) );
  AOI21_X1 U9741 ( .B1(n10438), .B2(n8042), .A(n8134), .ZN(n8060) );
  OAI21_X1 U9742 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n8045), .A(n8140), .ZN(
        n8058) );
  INV_X1 U9743 ( .A(n8046), .ZN(n8047) );
  MUX2_X1 U9744 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8049), .Z(n8144) );
  XNOR2_X1 U9745 ( .A(n8144), .B(n8139), .ZN(n8050) );
  NOR2_X1 U9746 ( .A1(n8051), .A2(n8050), .ZN(n8145) );
  AOI21_X1 U9747 ( .B1(n8051), .B2(n8050), .A(n8145), .ZN(n8056) );
  NOR2_X1 U9748 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8052), .ZN(n8219) );
  NOR2_X1 U9749 ( .A1(n10321), .A2(n8053), .ZN(n8054) );
  AOI211_X1 U9750 ( .C1(n9045), .C2(n8147), .A(n8219), .B(n8054), .ZN(n8055)
         );
  OAI21_X1 U9751 ( .B1(n8056), .B2(n10317), .A(n8055), .ZN(n8057) );
  AOI21_X1 U9752 ( .B1(n8058), .B2(n10308), .A(n8057), .ZN(n8059) );
  OAI21_X1 U9753 ( .B1(n8060), .B2(n10283), .A(n8059), .ZN(P2_U3193) );
  INV_X1 U9754 ( .A(n8065), .ZN(n8063) );
  NAND2_X1 U9755 ( .A1(n8061), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8804) );
  NAND2_X1 U9756 ( .A1(n9352), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8062) );
  OAI211_X1 U9757 ( .C1(n8063), .C2(n9355), .A(n8804), .B(n8062), .ZN(P2_U3272) );
  NAND2_X1 U9758 ( .A1(n8065), .A2(n8064), .ZN(n8067) );
  OAI211_X1 U9759 ( .C1(n8068), .C2(n9952), .A(n8067), .B(n8066), .ZN(P1_U3332) );
  XNOR2_X1 U9760 ( .A(n8126), .B(n8125), .ZN(n10207) );
  NAND2_X1 U9761 ( .A1(n8073), .A2(n8072), .ZN(n8075) );
  NAND2_X1 U9762 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  NAND3_X1 U9763 ( .A1(n8076), .A2(n8117), .A3(n10092), .ZN(n8079) );
  OAI22_X1 U9764 ( .A1(n8428), .A2(n9991), .B1(n9504), .B2(n9989), .ZN(n8077)
         );
  INV_X1 U9765 ( .A(n8077), .ZN(n8078) );
  NAND2_X1 U9766 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  AOI21_X1 U9767 ( .B1(n10207), .B2(n8081), .A(n8080), .ZN(n10209) );
  OAI21_X1 U9768 ( .B1(n8082), .B2(n10204), .A(n10099), .ZN(n8083) );
  OR2_X1 U9769 ( .A1(n8127), .A2(n8083), .ZN(n10203) );
  AOI22_X1 U9770 ( .A1(n10121), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8425), .B2(
        n10096), .ZN(n8085) );
  NAND2_X1 U9771 ( .A1(n8431), .A2(n10094), .ZN(n8084) );
  OAI211_X1 U9772 ( .C1(n10203), .C2(n9847), .A(n8085), .B(n8084), .ZN(n8086)
         );
  AOI21_X1 U9773 ( .B1(n10207), .B2(n8087), .A(n8086), .ZN(n8088) );
  OAI21_X1 U9774 ( .B1(n10209), .B2(n10121), .A(n8088), .ZN(P1_U3282) );
  OAI21_X1 U9775 ( .B1(n4603), .B2(n5352), .A(n8089), .ZN(n8100) );
  XNOR2_X1 U9776 ( .A(n8090), .B(n8780), .ZN(n8091) );
  OAI222_X1 U9777 ( .A1(n10346), .A2(n8409), .B1(n10348), .B2(n8168), .C1(
        n9187), .C2(n8091), .ZN(n8097) );
  NAND2_X1 U9778 ( .A1(n8097), .A2(n9211), .ZN(n8094) );
  OAI22_X1 U9779 ( .A1(n10357), .A2(n8149), .B1(n8172), .B2(n10343), .ZN(n8092) );
  AOI21_X1 U9780 ( .B1(n8669), .B2(n9226), .A(n8092), .ZN(n8093) );
  OAI211_X1 U9781 ( .C1(n8100), .C2(n9229), .A(n8094), .B(n8093), .ZN(P2_U3221) );
  INV_X1 U9782 ( .A(n10414), .ZN(n10396) );
  NOR2_X1 U9783 ( .A1(n10423), .A2(n10396), .ZN(n9318) );
  INV_X1 U9784 ( .A(n9318), .ZN(n9342) );
  NAND2_X1 U9785 ( .A1(n8097), .A2(n10421), .ZN(n8096) );
  AOI22_X1 U9786 ( .A1(n8669), .A2(n9338), .B1(n10423), .B2(
        P2_REG0_REG_12__SCAN_IN), .ZN(n8095) );
  OAI211_X1 U9787 ( .C1(n8100), .C2(n9342), .A(n8096), .B(n8095), .ZN(P2_U3426) );
  AND2_X1 U9788 ( .A1(n10440), .A2(n10414), .ZN(n9253) );
  INV_X1 U9789 ( .A(n9253), .ZN(n9273) );
  NAND2_X1 U9790 ( .A1(n8097), .A2(n10440), .ZN(n8099) );
  AOI22_X1 U9791 ( .A1(n8669), .A2(n9270), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n10437), .ZN(n8098) );
  OAI211_X1 U9792 ( .C1(n9273), .C2(n8100), .A(n8099), .B(n8098), .ZN(P2_U3471) );
  INV_X1 U9793 ( .A(n8258), .ZN(n8115) );
  INV_X1 U9794 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8101) );
  MUX2_X1 U9795 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n8101), .S(n8258), .Z(n8102)
         );
  INV_X1 U9796 ( .A(n8102), .ZN(n8105) );
  OAI21_X1 U9797 ( .B1(n8107), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8103), .ZN(
        n8104) );
  NOR2_X1 U9798 ( .A1(n8104), .A2(n8105), .ZN(n8257) );
  AOI211_X1 U9799 ( .C1(n8105), .C2(n8104), .A(n8257), .B(n10022), .ZN(n8111)
         );
  OAI21_X1 U9800 ( .B1(n8107), .B2(P1_REG1_REG_12__SCAN_IN), .A(n8106), .ZN(
        n8109) );
  INV_X1 U9801 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10245) );
  MUX2_X1 U9802 ( .A(n10245), .B(P1_REG1_REG_13__SCAN_IN), .S(n8258), .Z(n8108) );
  NOR2_X1 U9803 ( .A1(n8109), .A2(n8108), .ZN(n8254) );
  AOI211_X1 U9804 ( .C1(n8109), .C2(n8108), .A(n8254), .B(n9631), .ZN(n8110)
         );
  NOR2_X1 U9805 ( .A1(n8111), .A2(n8110), .ZN(n8114) );
  AND2_X1 U9806 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8112) );
  AOI21_X1 U9807 ( .B1(n10049), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n8112), .ZN(
        n8113) );
  OAI211_X1 U9808 ( .C1(n8115), .C2(n9629), .A(n8114), .B(n8113), .ZN(P1_U3256) );
  AND2_X1 U9809 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  OAI21_X1 U9810 ( .B1(n8119), .B2(n8118), .A(n8306), .ZN(n8122) );
  OR2_X1 U9811 ( .A1(n8123), .A2(n9991), .ZN(n8121) );
  OR2_X1 U9812 ( .A1(n8288), .A2(n9989), .ZN(n8120) );
  NAND2_X1 U9813 ( .A1(n8121), .A2(n8120), .ZN(n8437) );
  AOI21_X1 U9814 ( .B1(n8122), .B2(n10092), .A(n8437), .ZN(n10212) );
  INV_X1 U9815 ( .A(n8123), .ZN(n9505) );
  XNOR2_X1 U9816 ( .A(n8292), .B(n8291), .ZN(n10215) );
  NAND2_X1 U9817 ( .A1(n10215), .A2(n10104), .ZN(n8132) );
  OAI211_X1 U9818 ( .C1(n8127), .C2(n10213), .A(n10099), .B(n8314), .ZN(n10211) );
  INV_X1 U9819 ( .A(n10211), .ZN(n8130) );
  AOI22_X1 U9820 ( .A1(n10121), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8436), .B2(
        n10096), .ZN(n8128) );
  OAI21_X1 U9821 ( .B1(n10213), .B2(n9815), .A(n8128), .ZN(n8129) );
  AOI21_X1 U9822 ( .B1(n8130), .B2(n10103), .A(n8129), .ZN(n8131) );
  OAI211_X1 U9823 ( .C1(n10121), .C2(n10212), .A(n8132), .B(n8131), .ZN(
        P1_U3281) );
  NOR2_X1 U9824 ( .A1(n8147), .A2(n8133), .ZN(n8135) );
  NAND2_X1 U9825 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8197), .ZN(n8136) );
  OAI21_X1 U9826 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8197), .A(n8136), .ZN(
        n8137) );
  AOI21_X1 U9827 ( .B1(n4595), .B2(n8137), .A(n8194), .ZN(n8163) );
  AOI22_X1 U9828 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8197), .B1(n8157), .B2(
        n8149), .ZN(n8143) );
  NAND2_X1 U9829 ( .A1(n8139), .A2(n8138), .ZN(n8141) );
  NAND2_X1 U9830 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  NAND2_X1 U9831 ( .A1(n8143), .A2(n8142), .ZN(n8198) );
  OAI21_X1 U9832 ( .B1(n8143), .B2(n8142), .A(n8198), .ZN(n8161) );
  INV_X1 U9833 ( .A(n8144), .ZN(n8146) );
  MUX2_X1 U9834 ( .A(n8149), .B(n8148), .S(n8049), .Z(n8150) );
  NOR2_X1 U9835 ( .A1(n8150), .A2(n8157), .ZN(n8202) );
  NAND2_X1 U9836 ( .A1(n8150), .A2(n8157), .ZN(n8203) );
  INV_X1 U9837 ( .A(n8203), .ZN(n8151) );
  NOR2_X1 U9838 ( .A1(n8202), .A2(n8151), .ZN(n8153) );
  NAND2_X1 U9839 ( .A1(n8204), .A2(n8153), .ZN(n8152) );
  OAI211_X1 U9840 ( .C1(n8204), .C2(n8153), .A(n10272), .B(n8152), .ZN(n8159)
         );
  NOR2_X1 U9841 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8154), .ZN(n8170) );
  NOR2_X1 U9842 ( .A1(n10321), .A2(n8155), .ZN(n8156) );
  AOI211_X1 U9843 ( .C1(n9045), .C2(n8157), .A(n8170), .B(n8156), .ZN(n8158)
         );
  NAND2_X1 U9844 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  AOI21_X1 U9845 ( .B1(n8161), .B2(n10308), .A(n8160), .ZN(n8162) );
  OAI21_X1 U9846 ( .B1(n8163), .B2(n10283), .A(n8162), .ZN(P2_U3194) );
  XNOR2_X1 U9847 ( .A(n8164), .B(n8838), .ZN(n8225) );
  XNOR2_X1 U9848 ( .A(n8669), .B(n8838), .ZN(n8343) );
  XNOR2_X1 U9849 ( .A(n8343), .B(n8668), .ZN(n8167) );
  XNOR2_X1 U9850 ( .A(n8344), .B(n8167), .ZN(n8175) );
  NOR2_X1 U9851 ( .A1(n8948), .A2(n8168), .ZN(n8169) );
  AOI211_X1 U9852 ( .C1(n8944), .C2(n8962), .A(n8170), .B(n8169), .ZN(n8171)
         );
  OAI21_X1 U9853 ( .B1(n8172), .B2(n8221), .A(n8171), .ZN(n8173) );
  AOI21_X1 U9854 ( .B1(n8669), .B2(n8951), .A(n8173), .ZN(n8174) );
  OAI21_X1 U9855 ( .B1(n8175), .B2(n8953), .A(n8174), .ZN(P2_U3164) );
  INV_X1 U9856 ( .A(n8176), .ZN(n8180) );
  OAI222_X1 U9857 ( .A1(n8178), .A2(P1_U3086), .B1(n9949), .B2(n8180), .C1(
        n8177), .C2(n9952), .ZN(P1_U3331) );
  OAI222_X1 U9858 ( .A1(n8181), .A2(P2_U3151), .B1(n9355), .B2(n8180), .C1(
        n8179), .C2(n8849), .ZN(P2_U3271) );
  INV_X1 U9859 ( .A(n8182), .ZN(n8183) );
  AOI21_X1 U9860 ( .B1(n8777), .B2(n8184), .A(n8183), .ZN(n8185) );
  OAI222_X1 U9861 ( .A1(n10346), .A2(n8512), .B1(n10348), .B2(n8668), .C1(
        n9187), .C2(n8185), .ZN(n8248) );
  INV_X1 U9862 ( .A(n5714), .ZN(n8357) );
  OAI22_X1 U9863 ( .A1(n8357), .A2(n10341), .B1(n8350), .B2(n10343), .ZN(n8186) );
  OAI21_X1 U9864 ( .B1(n8248), .B2(n8186), .A(n9211), .ZN(n8189) );
  XOR2_X1 U9865 ( .A(n8187), .B(n8777), .Z(n8245) );
  INV_X1 U9866 ( .A(n9229), .ZN(n10336) );
  NAND2_X1 U9867 ( .A1(n8245), .A2(n10336), .ZN(n8188) );
  OAI211_X1 U9868 ( .C1(n10357), .C2(n8190), .A(n8189), .B(n8188), .ZN(
        P2_U3220) );
  INV_X1 U9869 ( .A(n8191), .ZN(n8215) );
  AOI22_X1 U9870 ( .A1(n8192), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9352), .ZN(n8193) );
  OAI21_X1 U9871 ( .B1(n8215), .B2(n9355), .A(n8193), .ZN(P2_U3270) );
  AOI21_X1 U9872 ( .B1(n8196), .B2(n8195), .A(n8365), .ZN(n8213) );
  NAND2_X1 U9873 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8197), .ZN(n8199) );
  OAI21_X1 U9874 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8200), .A(n8370), .ZN(
        n8211) );
  NOR2_X1 U9875 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5362), .ZN(n8351) );
  NOR2_X1 U9876 ( .A1(n10312), .A2(n8374), .ZN(n8201) );
  AOI211_X1 U9877 ( .C1(n10248), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n8351), .B(
        n8201), .ZN(n8209) );
  MUX2_X1 U9878 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8049), .Z(n8375) );
  XNOR2_X1 U9879 ( .A(n8375), .B(n8364), .ZN(n8206) );
  AOI21_X1 U9880 ( .B1(n8204), .B2(n8203), .A(n8202), .ZN(n8205) );
  NAND2_X1 U9881 ( .A1(n8205), .A2(n8206), .ZN(n8376) );
  OAI21_X1 U9882 ( .B1(n8206), .B2(n8205), .A(n8376), .ZN(n8207) );
  NAND2_X1 U9883 ( .A1(n8207), .A2(n10272), .ZN(n8208) );
  NAND2_X1 U9884 ( .A1(n8209), .A2(n8208), .ZN(n8210) );
  AOI21_X1 U9885 ( .B1(n8211), .B2(n10308), .A(n8210), .ZN(n8212) );
  OAI21_X1 U9886 ( .B1(n8213), .B2(n10283), .A(n8212), .ZN(P2_U3195) );
  OAI222_X1 U9887 ( .A1(n8216), .A2(P1_U3086), .B1(n9949), .B2(n8215), .C1(
        n8214), .C2(n9952), .ZN(P1_U3330) );
  NOR2_X1 U9888 ( .A1(n8948), .A2(n8217), .ZN(n8218) );
  AOI211_X1 U9889 ( .C1(n8944), .C2(n8963), .A(n8219), .B(n8218), .ZN(n8220)
         );
  OAI21_X1 U9890 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8227) );
  AOI211_X1 U9891 ( .C1(n8225), .C2(n8224), .A(n8953), .B(n8223), .ZN(n8226)
         );
  AOI211_X1 U9892 ( .C1(n10417), .C2(n8951), .A(n8227), .B(n8226), .ZN(n8228)
         );
  INV_X1 U9893 ( .A(n8228), .ZN(P2_U3176) );
  INV_X1 U9894 ( .A(n8691), .ZN(n8229) );
  XNOR2_X1 U9895 ( .A(n8230), .B(n8781), .ZN(n8241) );
  INV_X1 U9896 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8233) );
  XNOR2_X1 U9897 ( .A(n8231), .B(n8781), .ZN(n8232) );
  AOI222_X1 U9898 ( .A1(n10350), .A2(n8232), .B1(n8959), .B2(n10328), .C1(
        n8961), .C2(n10326), .ZN(n8238) );
  MUX2_X1 U9899 ( .A(n8233), .B(n8238), .S(n10421), .Z(n8235) );
  NAND2_X1 U9900 ( .A1(n8508), .A2(n9338), .ZN(n8234) );
  OAI211_X1 U9901 ( .C1(n8241), .C2(n9342), .A(n8235), .B(n8234), .ZN(P2_U3435) );
  MUX2_X1 U9902 ( .A(n8986), .B(n8238), .S(n10357), .Z(n8237) );
  AOI22_X1 U9903 ( .A1(n8508), .A2(n9226), .B1(n9225), .B2(n8514), .ZN(n8236)
         );
  OAI211_X1 U9904 ( .C1(n8241), .C2(n9229), .A(n8237), .B(n8236), .ZN(P2_U3218) );
  MUX2_X1 U9905 ( .A(n8976), .B(n8238), .S(n10440), .Z(n8240) );
  NAND2_X1 U9906 ( .A1(n8508), .A2(n9270), .ZN(n8239) );
  OAI211_X1 U9907 ( .C1(n9273), .C2(n8241), .A(n8240), .B(n8239), .ZN(P2_U3474) );
  INV_X1 U9908 ( .A(n8242), .ZN(n8302) );
  AOI22_X1 U9909 ( .A1(n8243), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9352), .ZN(n8244) );
  OAI21_X1 U9910 ( .B1(n8302), .B2(n9355), .A(n8244), .ZN(P2_U3269) );
  MUX2_X1 U9911 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8248), .S(n10440), .Z(n8247) );
  INV_X1 U9912 ( .A(n8245), .ZN(n8249) );
  OAI22_X1 U9913 ( .A1(n8249), .A2(n9273), .B1(n8357), .B2(n9263), .ZN(n8246)
         );
  OR2_X1 U9914 ( .A1(n8247), .A2(n8246), .ZN(P2_U3472) );
  MUX2_X1 U9915 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8248), .S(n10421), .Z(n8251) );
  OAI22_X1 U9916 ( .A1(n8249), .A2(n9342), .B1(n8357), .B2(n9331), .ZN(n8250)
         );
  OR2_X1 U9917 ( .A1(n8251), .A2(n8250), .ZN(P2_U3429) );
  OR2_X1 U9918 ( .A1(n9553), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U9919 ( .A1(n9553), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U9920 ( .A1(n8253), .A2(n8252), .ZN(n9555) );
  AOI21_X1 U9921 ( .B1(n8258), .B2(P1_REG1_REG_13__SCAN_IN), .A(n8254), .ZN(
        n9556) );
  XOR2_X1 U9922 ( .A(n9555), .B(n9556), .Z(n8264) );
  AND2_X1 U9923 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8255) );
  AOI21_X1 U9924 ( .B1(n10049), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n8255), .ZN(
        n8256) );
  OAI21_X1 U9925 ( .B1(n9629), .B2(n9558), .A(n8256), .ZN(n8263) );
  INV_X1 U9926 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8259) );
  AOI22_X1 U9927 ( .A1(n9553), .A2(n8259), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n9558), .ZN(n8260) );
  AOI211_X1 U9928 ( .C1(n8261), .C2(n8260), .A(n9552), .B(n10022), .ZN(n8262)
         );
  AOI211_X1 U9929 ( .C1(n10053), .C2(n8264), .A(n8263), .B(n8262), .ZN(n8265)
         );
  INV_X1 U9930 ( .A(n8265), .ZN(P1_U3257) );
  INV_X1 U9931 ( .A(n8266), .ZN(n8681) );
  OR2_X1 U9932 ( .A1(n8680), .A2(n8681), .ZN(n8779) );
  XNOR2_X1 U9933 ( .A(n8267), .B(n8779), .ZN(n8268) );
  AOI222_X1 U9934 ( .A1(n10350), .A2(n8268), .B1(n8960), .B2(n10328), .C1(
        n8962), .C2(n10326), .ZN(n8278) );
  MUX2_X1 U9935 ( .A(n8269), .B(n8278), .S(n10440), .Z(n8274) );
  NAND2_X1 U9936 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  XNOR2_X1 U9937 ( .A(n8272), .B(n8779), .ZN(n8281) );
  AOI22_X1 U9938 ( .A1(n8281), .A2(n9253), .B1(n9270), .B2(n8402), .ZN(n8273)
         );
  NAND2_X1 U9939 ( .A1(n8274), .A2(n8273), .ZN(P2_U3473) );
  INV_X1 U9940 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8275) );
  MUX2_X1 U9941 ( .A(n8275), .B(n8278), .S(n10421), .Z(n8277) );
  AOI22_X1 U9942 ( .A1(n8281), .A2(n9318), .B1(n9338), .B2(n8402), .ZN(n8276)
         );
  NAND2_X1 U9943 ( .A1(n8277), .A2(n8276), .ZN(P2_U3432) );
  INV_X1 U9944 ( .A(n8402), .ZN(n8414) );
  NOR2_X1 U9945 ( .A1(n8414), .A2(n10341), .ZN(n8280) );
  INV_X1 U9946 ( .A(n8278), .ZN(n8279) );
  AOI211_X1 U9947 ( .C1(n9225), .C2(n8411), .A(n8280), .B(n8279), .ZN(n8283)
         );
  INV_X1 U9948 ( .A(n9211), .ZN(n10339) );
  AOI22_X1 U9949 ( .A1(n8281), .A2(n10336), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10339), .ZN(n8282) );
  OAI21_X1 U9950 ( .B1(n8283), .B2(n10339), .A(n8282), .ZN(P2_U3219) );
  NAND2_X1 U9951 ( .A1(n8284), .A2(n8285), .ZN(n8287) );
  NAND2_X1 U9952 ( .A1(n8287), .A2(n8293), .ZN(n8286) );
  OAI21_X1 U9953 ( .B1(n8293), .B2(n8287), .A(n8286), .ZN(n8295) );
  OAI22_X1 U9954 ( .A1(n9395), .A2(n9989), .B1(n8288), .B2(n9991), .ZN(n8395)
         );
  OAI22_X1 U9955 ( .A1(n8312), .A2(n8311), .B1(n8528), .B2(n9503), .ZN(n8326)
         );
  XNOR2_X1 U9956 ( .A(n8326), .B(n8293), .ZN(n9923) );
  NOR2_X1 U9957 ( .A1(n9923), .A2(n9859), .ZN(n8294) );
  AOI211_X1 U9958 ( .C1(n10092), .C2(n8295), .A(n8395), .B(n8294), .ZN(n9922)
         );
  AOI211_X1 U9959 ( .C1(n9920), .C2(n8315), .A(n9810), .B(n4602), .ZN(n9919)
         );
  AOI22_X1 U9960 ( .A1(n10121), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8394), .B2(
        n10096), .ZN(n8296) );
  OAI21_X1 U9961 ( .B1(n8324), .B2(n9815), .A(n8296), .ZN(n8299) );
  NOR2_X1 U9962 ( .A1(n9923), .A2(n8297), .ZN(n8298) );
  AOI211_X1 U9963 ( .C1(n9919), .C2(n10103), .A(n8299), .B(n8298), .ZN(n8300)
         );
  OAI21_X1 U9964 ( .B1(n9922), .B2(n10121), .A(n8300), .ZN(P1_U3279) );
  OAI222_X1 U9965 ( .A1(n8303), .A2(P1_U3086), .B1(n9949), .B2(n8302), .C1(
        n8301), .C2(n9952), .ZN(P1_U3329) );
  INV_X1 U9966 ( .A(n8311), .ZN(n8305) );
  NAND3_X1 U9967 ( .A1(n8306), .A2(n8305), .A3(n8304), .ZN(n8307) );
  NAND2_X1 U9968 ( .A1(n8284), .A2(n8307), .ZN(n8310) );
  NAND2_X1 U9969 ( .A1(n9502), .A2(n9834), .ZN(n8308) );
  OAI21_X1 U9970 ( .B1(n9504), .B2(n9991), .A(n8308), .ZN(n8309) );
  AOI21_X1 U9971 ( .B1(n8310), .B2(n10092), .A(n8309), .ZN(n10218) );
  XNOR2_X1 U9972 ( .A(n8312), .B(n8311), .ZN(n10223) );
  NAND2_X1 U9973 ( .A1(n10223), .A2(n10104), .ZN(n8320) );
  INV_X1 U9974 ( .A(n8313), .ZN(n8525) );
  OAI22_X1 U9975 ( .A1(n10118), .A2(n8101), .B1(n8525), .B2(n10108), .ZN(n8318) );
  INV_X1 U9976 ( .A(n8314), .ZN(n8316) );
  INV_X1 U9977 ( .A(n8528), .ZN(n10220) );
  OAI211_X1 U9978 ( .C1(n8316), .C2(n10220), .A(n10099), .B(n8315), .ZN(n10217) );
  NOR2_X1 U9979 ( .A1(n10217), .A2(n9847), .ZN(n8317) );
  AOI211_X1 U9980 ( .C1(n10094), .C2(n8528), .A(n8318), .B(n8317), .ZN(n8319)
         );
  OAI211_X1 U9981 ( .C1(n10121), .C2(n10218), .A(n8320), .B(n8319), .ZN(
        P1_U3280) );
  INV_X1 U9982 ( .A(n8321), .ZN(n8358) );
  AOI21_X1 U9983 ( .B1(n9352), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8322), .ZN(
        n8323) );
  OAI21_X1 U9984 ( .B1(n8358), .B2(n9355), .A(n8323), .ZN(P2_U3268) );
  NAND2_X1 U9985 ( .A1(n9920), .A2(n9502), .ZN(n8325) );
  AOI22_X1 U9986 ( .A1(n8326), .A2(n8325), .B1(n8324), .B2(n9489), .ZN(n8486)
         );
  XNOR2_X1 U9987 ( .A(n8486), .B(n8329), .ZN(n9918) );
  OAI21_X1 U9988 ( .B1(n4602), .B2(n8487), .A(n10099), .ZN(n8327) );
  NOR2_X1 U9989 ( .A1(n8327), .A2(n8494), .ZN(n9915) );
  INV_X1 U9990 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8328) );
  OAI22_X1 U9991 ( .A1(n8487), .A2(n9815), .B1(n10118), .B2(n8328), .ZN(n8334)
         );
  XNOR2_X1 U9992 ( .A(n8330), .B(n8329), .ZN(n8331) );
  OAI222_X1 U9993 ( .A1(n9989), .A2(n9486), .B1(n9991), .B2(n9489), .C1(n8331), 
        .C2(n10129), .ZN(n9914) );
  AOI21_X1 U9994 ( .B1(n9484), .B2(n10096), .A(n9914), .ZN(n8332) );
  NOR2_X1 U9995 ( .A1(n8332), .A2(n10121), .ZN(n8333) );
  AOI211_X1 U9996 ( .C1(n9915), .C2(n10103), .A(n8334), .B(n8333), .ZN(n8335)
         );
  OAI21_X1 U9997 ( .B1(n9918), .B2(n9829), .A(n8335), .ZN(P1_U3278) );
  INV_X1 U9998 ( .A(n8336), .ZN(n8783) );
  XNOR2_X1 U9999 ( .A(n8337), .B(n8783), .ZN(n8338) );
  AOI222_X1 U10000 ( .A1(n10350), .A2(n8338), .B1(n8958), .B2(n10328), .C1(
        n8960), .C2(n10326), .ZN(n9277) );
  OAI21_X1 U10001 ( .B1(n4541), .B2(n8783), .A(n4596), .ZN(n9275) );
  INV_X1 U10002 ( .A(n9274), .ZN(n8546) );
  AOI22_X1 U10003 ( .A1(n10339), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9225), 
        .B2(n8543), .ZN(n8339) );
  OAI21_X1 U10004 ( .B1(n8546), .B2(n10334), .A(n8339), .ZN(n8340) );
  AOI21_X1 U10005 ( .B1(n9275), .B2(n10336), .A(n8340), .ZN(n8341) );
  OAI21_X1 U10006 ( .B1(n9277), .B2(n10339), .A(n8341), .ZN(P2_U3217) );
  INV_X1 U10007 ( .A(n8951), .ZN(n8939) );
  XNOR2_X1 U10008 ( .A(n5714), .B(n4527), .ZN(n8342) );
  NOR2_X1 U10009 ( .A1(n8342), .A2(n8962), .ZN(n8401) );
  AOI21_X1 U10010 ( .B1(n8342), .B2(n8962), .A(n8401), .ZN(n8348) );
  INV_X1 U10011 ( .A(n8344), .ZN(n8346) );
  AOI21_X1 U10012 ( .B1(n8344), .B2(n8668), .A(n8343), .ZN(n8345) );
  AOI21_X1 U10013 ( .B1(n8963), .B2(n8346), .A(n8345), .ZN(n8347) );
  NAND2_X1 U10014 ( .A1(n8347), .A2(n8348), .ZN(n8405) );
  OAI21_X1 U10015 ( .B1(n8348), .B2(n8347), .A(n8405), .ZN(n8349) );
  NAND2_X1 U10016 ( .A1(n8349), .A2(n8928), .ZN(n8356) );
  INV_X1 U10017 ( .A(n8350), .ZN(n8354) );
  AOI21_X1 U10018 ( .B1(n8931), .B2(n8963), .A(n8351), .ZN(n8352) );
  OAI21_X1 U10019 ( .B1(n8512), .B2(n8933), .A(n8352), .ZN(n8353) );
  AOI21_X1 U10020 ( .B1(n8354), .B2(n8945), .A(n8353), .ZN(n8355) );
  OAI211_X1 U10021 ( .C1(n8357), .C2(n8939), .A(n8356), .B(n8355), .ZN(
        P2_U3174) );
  OAI222_X1 U10022 ( .A1(n9952), .A2(n8359), .B1(P1_U3086), .B2(n10028), .C1(
        n9949), .C2(n8358), .ZN(P1_U3328) );
  INV_X1 U10023 ( .A(n8360), .ZN(n8503) );
  AOI21_X1 U10024 ( .B1(n9352), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8361), .ZN(
        n8362) );
  OAI21_X1 U10025 ( .B1(n8503), .B2(n9355), .A(n8362), .ZN(P2_U3267) );
  NOR2_X1 U10026 ( .A1(n8364), .A2(n8363), .ZN(n8366) );
  NAND2_X1 U10027 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8985), .ZN(n8367) );
  OAI21_X1 U10028 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8985), .A(n8367), .ZN(
        n8368) );
  AOI21_X1 U10029 ( .B1(n4593), .B2(n8368), .A(n8974), .ZN(n8388) );
  NAND2_X1 U10030 ( .A1(n8373), .A2(n5382), .ZN(n8984) );
  OAI21_X1 U10031 ( .B1(n8373), .B2(n5382), .A(n8984), .ZN(n8372) );
  NAND2_X1 U10032 ( .A1(n8374), .A2(n8369), .ZN(n8371) );
  XOR2_X1 U10033 ( .A(n8372), .B(n8983), .Z(n8386) );
  MUX2_X1 U10034 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8049), .Z(n8977) );
  XNOR2_X1 U10035 ( .A(n8977), .B(n8373), .ZN(n8379) );
  OR2_X1 U10036 ( .A1(n8375), .A2(n8374), .ZN(n8377) );
  NAND2_X1 U10037 ( .A1(n8377), .A2(n8376), .ZN(n8378) );
  NAND2_X1 U10038 ( .A1(n8379), .A2(n8378), .ZN(n8978) );
  OAI21_X1 U10039 ( .B1(n8379), .B2(n8378), .A(n8978), .ZN(n8383) );
  NOR2_X1 U10040 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8380), .ZN(n8407) );
  NOR2_X1 U10041 ( .A1(n10321), .A2(n8381), .ZN(n8382) );
  AOI211_X1 U10042 ( .C1(n10272), .C2(n8383), .A(n8407), .B(n8382), .ZN(n8384)
         );
  OAI21_X1 U10043 ( .B1(n8985), .B2(n10312), .A(n8384), .ZN(n8385) );
  AOI21_X1 U10044 ( .B1(n8386), .B2(n10308), .A(n8385), .ZN(n8387) );
  OAI21_X1 U10045 ( .B1(n8388), .B2(n10283), .A(n8387), .ZN(P2_U3196) );
  INV_X1 U10046 ( .A(n8389), .ZN(n8393) );
  XNOR2_X1 U10047 ( .A(n8391), .B(n8390), .ZN(n8392) );
  XNOR2_X1 U10048 ( .A(n8393), .B(n8392), .ZN(n8400) );
  INV_X1 U10049 ( .A(n8394), .ZN(n8397) );
  AOI22_X1 U10050 ( .A1(n8395), .A2(n9996), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8396) );
  OAI21_X1 U10051 ( .B1(n8397), .B2(n10003), .A(n8396), .ZN(n8398) );
  AOI21_X1 U10052 ( .B1(n9920), .B2(n9492), .A(n8398), .ZN(n8399) );
  OAI21_X1 U10053 ( .B1(n8400), .B2(n9494), .A(n8399), .ZN(P1_U3215) );
  INV_X1 U10054 ( .A(n8401), .ZN(n8403) );
  XNOR2_X1 U10055 ( .A(n8402), .B(n4527), .ZN(n8505) );
  XNOR2_X1 U10056 ( .A(n8505), .B(n8961), .ZN(n8404) );
  AND3_X1 U10057 ( .A1(n8405), .A2(n8404), .A3(n8403), .ZN(n8406) );
  OAI21_X1 U10058 ( .B1(n8506), .B2(n8406), .A(n8928), .ZN(n8413) );
  AOI21_X1 U10059 ( .B1(n8944), .B2(n8960), .A(n8407), .ZN(n8408) );
  OAI21_X1 U10060 ( .B1(n8409), .B2(n8948), .A(n8408), .ZN(n8410) );
  AOI21_X1 U10061 ( .B1(n8411), .B2(n8945), .A(n8410), .ZN(n8412) );
  OAI211_X1 U10062 ( .C1(n8414), .C2(n8939), .A(n8413), .B(n8412), .ZN(
        P2_U3155) );
  NOR2_X1 U10063 ( .A1(n8415), .A2(n8416), .ZN(n8419) );
  AOI21_X1 U10064 ( .B1(n8415), .B2(n8416), .A(n8419), .ZN(n8458) );
  INV_X1 U10065 ( .A(n8417), .ZN(n8459) );
  NAND2_X1 U10066 ( .A1(n8458), .A2(n8459), .ZN(n8457) );
  INV_X1 U10067 ( .A(n8418), .ZN(n8420) );
  AOI21_X1 U10068 ( .B1(n8420), .B2(n8434), .A(n8419), .ZN(n8424) );
  NAND2_X1 U10069 ( .A1(n8421), .A2(n8422), .ZN(n8435) );
  INV_X1 U10070 ( .A(n8435), .ZN(n8423) );
  AOI22_X1 U10071 ( .A1(n8457), .A2(n8424), .B1(n8423), .B2(n8434), .ZN(n8433)
         );
  INV_X1 U10072 ( .A(n8425), .ZN(n8427) );
  OAI22_X1 U10073 ( .A1(n10003), .A2(n8427), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8426), .ZN(n8430) );
  INV_X1 U10074 ( .A(n9474), .ZN(n9488) );
  OAI22_X1 U10075 ( .A1(n8428), .A2(n9488), .B1(n9487), .B2(n9504), .ZN(n8429)
         );
  AOI211_X1 U10076 ( .C1(n8431), .C2(n9492), .A(n8430), .B(n8429), .ZN(n8432)
         );
  OAI21_X1 U10077 ( .B1(n8433), .B2(n9494), .A(n8432), .ZN(P1_U3236) );
  NAND2_X1 U10078 ( .A1(n8435), .A2(n8434), .ZN(n8519) );
  XOR2_X1 U10079 ( .A(n8518), .B(n8519), .Z(n8444) );
  INV_X1 U10080 ( .A(n8436), .ZN(n8440) );
  NAND2_X1 U10081 ( .A1(n8437), .A2(n9996), .ZN(n8439) );
  OAI211_X1 U10082 ( .C1(n10003), .C2(n8440), .A(n8439), .B(n8438), .ZN(n8441)
         );
  AOI21_X1 U10083 ( .B1(n8442), .B2(n9492), .A(n8441), .ZN(n8443) );
  OAI21_X1 U10084 ( .B1(n8444), .B2(n9494), .A(n8443), .ZN(P1_U3224) );
  XOR2_X1 U10085 ( .A(n8445), .B(n8696), .Z(n8456) );
  INV_X1 U10086 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8448) );
  XOR2_X1 U10087 ( .A(n8446), .B(n8696), .Z(n8447) );
  AOI222_X1 U10088 ( .A1(n10350), .A2(n8447), .B1(n8959), .B2(n10326), .C1(
        n8957), .C2(n10328), .ZN(n8453) );
  MUX2_X1 U10089 ( .A(n8448), .B(n8453), .S(n10421), .Z(n8450) );
  NAND2_X1 U10090 ( .A1(n8889), .A2(n9338), .ZN(n8449) );
  OAI211_X1 U10091 ( .C1(n8456), .C2(n9342), .A(n8450), .B(n8449), .ZN(
        P2_U3441) );
  INV_X1 U10092 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9037) );
  MUX2_X1 U10093 ( .A(n9037), .B(n8453), .S(n10357), .Z(n8452) );
  AOI22_X1 U10094 ( .A1(n8889), .A2(n9226), .B1(n9225), .B2(n8897), .ZN(n8451)
         );
  OAI211_X1 U10095 ( .C1(n8456), .C2(n9229), .A(n8452), .B(n8451), .ZN(
        P2_U3216) );
  MUX2_X1 U10096 ( .A(n9027), .B(n8453), .S(n10440), .Z(n8455) );
  NAND2_X1 U10097 ( .A1(n8889), .A2(n9270), .ZN(n8454) );
  OAI211_X1 U10098 ( .C1(n9273), .C2(n8456), .A(n8455), .B(n8454), .ZN(
        P2_U3476) );
  OAI21_X1 U10099 ( .B1(n8459), .B2(n8458), .A(n8457), .ZN(n8460) );
  NAND2_X1 U10100 ( .A1(n8460), .A2(n10000), .ZN(n8467) );
  INV_X1 U10101 ( .A(n8461), .ZN(n8462) );
  NOR2_X1 U10102 ( .A1(n10003), .A2(n8462), .ZN(n8463) );
  AOI211_X1 U10103 ( .C1(n9996), .C2(n8465), .A(n8464), .B(n8463), .ZN(n8466)
         );
  OAI211_X1 U10104 ( .C1(n10199), .C2(n9998), .A(n8467), .B(n8466), .ZN(
        P1_U3217) );
  NAND2_X1 U10105 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  INV_X1 U10106 ( .A(n8690), .ZN(n8701) );
  AND2_X1 U10107 ( .A1(n8701), .A2(n8699), .ZN(n8472) );
  XNOR2_X1 U10108 ( .A(n8470), .B(n8472), .ZN(n8484) );
  INV_X1 U10109 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8474) );
  XNOR2_X1 U10110 ( .A(n8471), .B(n8472), .ZN(n8473) );
  AOI222_X1 U10111 ( .A1(n10350), .A2(n8473), .B1(n9203), .B2(n10328), .C1(
        n8958), .C2(n10326), .ZN(n8480) );
  MUX2_X1 U10112 ( .A(n8474), .B(n8480), .S(n10357), .Z(n8476) );
  AOI22_X1 U10113 ( .A1(n8924), .A2(n9226), .B1(n9225), .B2(n8936), .ZN(n8475)
         );
  OAI211_X1 U10114 ( .C1(n8484), .C2(n9229), .A(n8476), .B(n8475), .ZN(
        P2_U3215) );
  MUX2_X1 U10115 ( .A(n8477), .B(n8480), .S(n10440), .Z(n8479) );
  NAND2_X1 U10116 ( .A1(n8924), .A2(n9270), .ZN(n8478) );
  OAI211_X1 U10117 ( .C1(n8484), .C2(n9273), .A(n8479), .B(n8478), .ZN(
        P2_U3477) );
  INV_X1 U10118 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8481) );
  MUX2_X1 U10119 ( .A(n8481), .B(n8480), .S(n10421), .Z(n8483) );
  NAND2_X1 U10120 ( .A1(n8924), .A2(n9338), .ZN(n8482) );
  OAI211_X1 U10121 ( .C1(n8484), .C2(n9342), .A(n8483), .B(n8482), .ZN(
        P2_U3444) );
  XNOR2_X1 U10122 ( .A(n8548), .B(n4850), .ZN(n9975) );
  INV_X1 U10123 ( .A(n9975), .ZN(n8500) );
  NAND2_X1 U10124 ( .A1(n8488), .A2(n8547), .ZN(n8489) );
  NAND2_X1 U10125 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  NAND2_X1 U10126 ( .A1(n8491), .A2(n10092), .ZN(n8493) );
  AOI22_X1 U10127 ( .A1(n9794), .A2(n9501), .B1(n9499), .B2(n9834), .ZN(n8492)
         );
  NAND2_X1 U10128 ( .A1(n8493), .A2(n8492), .ZN(n9974) );
  OAI211_X1 U10129 ( .C1(n8494), .C2(n9972), .A(n10099), .B(n8553), .ZN(n9971)
         );
  AOI22_X1 U10130 ( .A1(n10121), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10096), 
        .B2(n8495), .ZN(n8497) );
  NAND2_X1 U10131 ( .A1(n9398), .A2(n10094), .ZN(n8496) );
  OAI211_X1 U10132 ( .C1(n9971), .C2(n9847), .A(n8497), .B(n8496), .ZN(n8498)
         );
  AOI21_X1 U10133 ( .B1(n9974), .B2(n10118), .A(n8498), .ZN(n8499) );
  OAI21_X1 U10134 ( .B1(n8500), .B2(n9829), .A(n8499), .ZN(P1_U3277) );
  INV_X1 U10135 ( .A(n5825), .ZN(n9948) );
  AOI22_X1 U10136 ( .A1(n8501), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9352), .ZN(n8502) );
  OAI21_X1 U10137 ( .B1(n9948), .B2(n9355), .A(n8502), .ZN(P2_U3266) );
  OAI222_X1 U10138 ( .A1(n9952), .A2(n8504), .B1(P1_U3086), .B2(n6452), .C1(
        n9949), .C2(n8503), .ZN(P1_U3327) );
  INV_X1 U10139 ( .A(n8508), .ZN(n8517) );
  INV_X1 U10140 ( .A(n8505), .ZN(n8507) );
  AOI21_X1 U10141 ( .B1(n8512), .B2(n8507), .A(n8506), .ZN(n8510) );
  XNOR2_X1 U10142 ( .A(n8508), .B(n8838), .ZN(n8532) );
  XNOR2_X1 U10143 ( .A(n8532), .B(n8960), .ZN(n8509) );
  OAI211_X1 U10144 ( .C1(n8510), .C2(n8509), .A(n8537), .B(n8928), .ZN(n8516)
         );
  NAND2_X1 U10145 ( .A1(n8944), .A2(n8959), .ZN(n8511) );
  NAND2_X1 U10146 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8988) );
  OAI211_X1 U10147 ( .C1(n8512), .C2(n8948), .A(n8511), .B(n8988), .ZN(n8513)
         );
  AOI21_X1 U10148 ( .B1(n8514), .B2(n8945), .A(n8513), .ZN(n8515) );
  OAI211_X1 U10149 ( .C1(n8517), .C2(n8939), .A(n8516), .B(n8515), .ZN(
        P2_U3181) );
  NAND2_X1 U10150 ( .A1(n8519), .A2(n8518), .ZN(n8521) );
  NAND2_X1 U10151 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  XOR2_X1 U10152 ( .A(n8523), .B(n8522), .Z(n8530) );
  OAI22_X1 U10153 ( .A1(n10003), .A2(n8525), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8524), .ZN(n8527) );
  OAI22_X1 U10154 ( .A1(n9504), .A2(n9488), .B1(n9487), .B2(n9489), .ZN(n8526)
         );
  AOI211_X1 U10155 ( .C1(n8528), .C2(n9492), .A(n8527), .B(n8526), .ZN(n8529)
         );
  OAI21_X1 U10156 ( .B1(n8530), .B2(n9494), .A(n8529), .ZN(P1_U3234) );
  XNOR2_X1 U10157 ( .A(n9274), .B(n4527), .ZN(n8531) );
  NOR2_X1 U10158 ( .A1(n8531), .A2(n8959), .ZN(n8814) );
  AOI21_X1 U10159 ( .B1(n8531), .B2(n8959), .A(n8814), .ZN(n8535) );
  INV_X1 U10160 ( .A(n8532), .ZN(n8533) );
  NAND2_X1 U10161 ( .A1(n8533), .A2(n8960), .ZN(n8536) );
  INV_X1 U10162 ( .A(n8892), .ZN(n8539) );
  AOI21_X1 U10163 ( .B1(n8537), .B2(n8536), .A(n8535), .ZN(n8538) );
  OAI21_X1 U10164 ( .B1(n8539), .B2(n8538), .A(n8928), .ZN(n8545) );
  NAND2_X1 U10165 ( .A1(n8944), .A2(n8958), .ZN(n8540) );
  NAND2_X1 U10166 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9009) );
  OAI211_X1 U10167 ( .C1(n8541), .C2(n8948), .A(n8540), .B(n9009), .ZN(n8542)
         );
  AOI21_X1 U10168 ( .B1(n8543), .B2(n8945), .A(n8542), .ZN(n8544) );
  OAI211_X1 U10169 ( .C1(n8546), .C2(n8939), .A(n8545), .B(n8544), .ZN(
        P2_U3166) );
  XNOR2_X1 U10170 ( .A(n8558), .B(n5083), .ZN(n9913) );
  XNOR2_X1 U10171 ( .A(n8550), .B(n8549), .ZN(n8551) );
  OAI222_X1 U10172 ( .A1(n9989), .A2(n9837), .B1(n9991), .B2(n9486), .C1(n8551), .C2(n10129), .ZN(n9909) );
  INV_X1 U10173 ( .A(n9911), .ZN(n9412) );
  INV_X1 U10174 ( .A(n8552), .ZN(n8566) );
  AOI211_X1 U10175 ( .C1(n9911), .C2(n8553), .A(n9810), .B(n8566), .ZN(n9910)
         );
  NAND2_X1 U10176 ( .A1(n9910), .A2(n10103), .ZN(n8555) );
  AOI22_X1 U10177 ( .A1(n10121), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9409), 
        .B2(n10096), .ZN(n8554) );
  OAI211_X1 U10178 ( .C1(n9412), .C2(n9815), .A(n8555), .B(n8554), .ZN(n8556)
         );
  AOI21_X1 U10179 ( .B1(n9909), .B2(n10118), .A(n8556), .ZN(n8557) );
  OAI21_X1 U10180 ( .B1(n9913), .B2(n9829), .A(n8557), .ZN(P1_U3276) );
  XNOR2_X1 U10181 ( .A(n9644), .B(n8559), .ZN(n9969) );
  INV_X1 U10182 ( .A(n9969), .ZN(n8571) );
  INV_X1 U10183 ( .A(n8559), .ZN(n8560) );
  XNOR2_X1 U10184 ( .A(n8561), .B(n8560), .ZN(n8562) );
  NAND2_X1 U10185 ( .A1(n8562), .A2(n10092), .ZN(n8564) );
  AOI22_X1 U10186 ( .A1(n9794), .A2(n9499), .B1(n9648), .B2(n9834), .ZN(n8563)
         );
  NAND2_X1 U10187 ( .A1(n8564), .A2(n8563), .ZN(n9968) );
  INV_X1 U10188 ( .A(n9846), .ZN(n8565) );
  OAI211_X1 U10189 ( .C1(n9966), .C2(n8566), .A(n8565), .B(n10099), .ZN(n9965)
         );
  AOI22_X1 U10190 ( .A1(n10121), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9459), 
        .B2(n10096), .ZN(n8568) );
  NAND2_X1 U10191 ( .A1(n9645), .A2(n10094), .ZN(n8567) );
  OAI211_X1 U10192 ( .C1(n9965), .C2(n9847), .A(n8568), .B(n8567), .ZN(n8569)
         );
  AOI21_X1 U10193 ( .B1(n9968), .B2(n10118), .A(n8569), .ZN(n8570) );
  OAI21_X1 U10194 ( .B1(n8571), .B2(n9829), .A(n8570), .ZN(P1_U3275) );
  OAI21_X1 U10195 ( .B1(n8574), .B2(n8573), .A(n8572), .ZN(n8575) );
  NAND2_X1 U10196 ( .A1(n8575), .A2(n10000), .ZN(n8580) );
  OAI22_X1 U10197 ( .A1(n8577), .A2(n9991), .B1(n8576), .B2(n9989), .ZN(n10091) );
  AOI22_X1 U10198 ( .A1(n10091), .A2(n9996), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8578), .ZN(n8579) );
  OAI211_X1 U10199 ( .C1(n10143), .C2(n9998), .A(n8580), .B(n8579), .ZN(
        P1_U3237) );
  NAND2_X1 U10200 ( .A1(n8581), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8584) );
  AOI22_X1 U10201 ( .A1(n8928), .A2(n8765), .B1(n8582), .B2(n8951), .ZN(n8583)
         );
  OAI211_X1 U10202 ( .C1(n5692), .C2(n8933), .A(n8584), .B(n8583), .ZN(
        P2_U3172) );
  OR2_X2 U10203 ( .A1(n8585), .A2(n8587), .ZN(n9417) );
  INV_X1 U10204 ( .A(n9417), .ZN(n8586) );
  AOI21_X1 U10205 ( .B1(n8587), .B2(n8585), .A(n8586), .ZN(n8594) );
  OR2_X1 U10206 ( .A1(n9808), .A2(n9991), .ZN(n8589) );
  OR2_X1 U10207 ( .A1(n9747), .A2(n9989), .ZN(n8588) );
  AND2_X1 U10208 ( .A1(n8589), .A2(n8588), .ZN(n9892) );
  OAI22_X1 U10209 ( .A1(n9892), .A2(n9439), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8590), .ZN(n8592) );
  NOR2_X1 U10210 ( .A1(n9894), .A2(n9998), .ZN(n8591) );
  AOI211_X1 U10211 ( .C1(n9472), .C2(n9780), .A(n8592), .B(n8591), .ZN(n8593)
         );
  OAI21_X1 U10212 ( .B1(n8594), .B2(n9494), .A(n8593), .ZN(P1_U3216) );
  INV_X1 U10213 ( .A(n8791), .ZN(n8599) );
  NAND2_X1 U10214 ( .A1(n9351), .A2(n5421), .ZN(n8596) );
  NAND2_X1 U10215 ( .A1(n5539), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U10216 ( .A1(n9345), .A2(n5421), .ZN(n8598) );
  NAND2_X1 U10217 ( .A1(n5539), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8597) );
  NOR2_X1 U10218 ( .A1(n9278), .A2(n8601), .ZN(n8758) );
  INV_X1 U10219 ( .A(n8758), .ZN(n8605) );
  INV_X1 U10220 ( .A(n8955), .ZN(n8602) );
  NAND2_X1 U10221 ( .A1(n9231), .A2(n8602), .ZN(n8747) );
  NAND2_X1 U10222 ( .A1(n8747), .A2(n8603), .ZN(n8745) );
  INV_X1 U10223 ( .A(n8745), .ZN(n8604) );
  NAND2_X1 U10224 ( .A1(n8605), .A2(n8604), .ZN(n8794) );
  NAND2_X1 U10225 ( .A1(n9284), .A2(n8955), .ZN(n8761) );
  OAI22_X1 U10226 ( .A1(n8606), .A2(n8794), .B1(n9100), .B2(n8761), .ZN(n8798)
         );
  INV_X1 U10227 ( .A(n8607), .ZN(n8797) );
  MUX2_X1 U10228 ( .A(n8746), .B(n9290), .S(n8748), .Z(n8743) );
  INV_X1 U10229 ( .A(n8608), .ZN(n8611) );
  OAI21_X1 U10230 ( .B1(n8609), .B2(n8766), .A(n8615), .ZN(n8610) );
  NAND2_X1 U10231 ( .A1(n8612), .A2(n5790), .ZN(n8613) );
  OAI21_X1 U10232 ( .B1(n8614), .B2(n8801), .A(n8613), .ZN(n8616) );
  NAND2_X1 U10233 ( .A1(n8616), .A2(n8615), .ZN(n8618) );
  NAND2_X1 U10234 ( .A1(n8618), .A2(n8617), .ZN(n8624) );
  OR2_X1 U10235 ( .A1(n10347), .A2(n10369), .ZN(n8625) );
  NAND2_X1 U10236 ( .A1(n8625), .A2(n8619), .ZN(n8622) );
  NAND2_X1 U10237 ( .A1(n8620), .A2(n8649), .ZN(n8621) );
  MUX2_X1 U10238 ( .A(n8622), .B(n8621), .S(n8748), .Z(n8623) );
  INV_X1 U10239 ( .A(n8625), .ZN(n8627) );
  OAI211_X1 U10240 ( .C1(n8628), .C2(n8627), .A(n8651), .B(n8626), .ZN(n8632)
         );
  INV_X1 U10241 ( .A(n8645), .ZN(n8630) );
  NAND2_X1 U10242 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  NAND3_X1 U10243 ( .A1(n8632), .A2(n8652), .A3(n8631), .ZN(n8635) );
  INV_X1 U10244 ( .A(n8633), .ZN(n8634) );
  AOI21_X1 U10245 ( .B1(n8635), .B2(n8653), .A(n8634), .ZN(n8643) );
  AND2_X1 U10246 ( .A1(n8662), .A2(n8657), .ZN(n8638) );
  AND2_X1 U10247 ( .A1(n8639), .A2(n8636), .ZN(n8637) );
  MUX2_X1 U10248 ( .A(n8638), .B(n8637), .S(n8753), .Z(n8659) );
  INV_X1 U10249 ( .A(n8659), .ZN(n8642) );
  INV_X1 U10250 ( .A(n8639), .ZN(n8640) );
  NOR2_X1 U10251 ( .A1(n8664), .A2(n8640), .ZN(n8641) );
  NAND2_X1 U10252 ( .A1(n8665), .A2(n8661), .ZN(n8644) );
  OAI21_X1 U10253 ( .B1(n8647), .B2(n8646), .A(n8645), .ZN(n8648) );
  AOI21_X1 U10254 ( .B1(n8650), .B2(n8649), .A(n8648), .ZN(n8655) );
  INV_X1 U10255 ( .A(n8651), .ZN(n8654) );
  OAI211_X1 U10256 ( .C1(n8655), .C2(n8654), .A(n8653), .B(n8652), .ZN(n8658)
         );
  NAND3_X1 U10257 ( .A1(n8658), .A2(n8657), .A3(n8656), .ZN(n8660) );
  NAND2_X1 U10258 ( .A1(n8660), .A2(n8659), .ZN(n8663) );
  NAND2_X1 U10259 ( .A1(n8665), .A2(n8664), .ZN(n8666) );
  NAND2_X1 U10260 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  MUX2_X1 U10261 ( .A(n8671), .B(n8670), .S(n8748), .Z(n8672) );
  NAND2_X1 U10262 ( .A1(n8673), .A2(n8672), .ZN(n8678) );
  INV_X1 U10263 ( .A(n8674), .ZN(n8675) );
  MUX2_X1 U10264 ( .A(n8962), .B(n5714), .S(n8753), .Z(n8676) );
  INV_X1 U10265 ( .A(n8779), .ZN(n8679) );
  MUX2_X1 U10266 ( .A(n8681), .B(n8680), .S(n8748), .Z(n8682) );
  NOR2_X1 U10267 ( .A1(n8781), .A2(n8682), .ZN(n8683) );
  NAND2_X1 U10268 ( .A1(n8684), .A2(n8683), .ZN(n8693) );
  INV_X1 U10269 ( .A(n8685), .ZN(n8686) );
  NAND3_X1 U10270 ( .A1(n8693), .A2(n8686), .A3(n8695), .ZN(n8687) );
  INV_X1 U10271 ( .A(n8688), .ZN(n8689) );
  NOR2_X1 U10272 ( .A1(n8690), .A2(n8689), .ZN(n8784) );
  NAND3_X1 U10273 ( .A1(n8693), .A2(n8692), .A3(n8691), .ZN(n8694) );
  NAND2_X1 U10274 ( .A1(n5002), .A2(n8753), .ZN(n8697) );
  NAND2_X1 U10275 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  INV_X1 U10276 ( .A(n8699), .ZN(n8700) );
  NOR3_X1 U10277 ( .A1(n8703), .A2(n8700), .A3(n9216), .ZN(n8705) );
  NAND2_X1 U10278 ( .A1(n8706), .A2(n8701), .ZN(n8702) );
  NAND2_X1 U10279 ( .A1(n8710), .A2(n8706), .ZN(n8709) );
  NAND2_X1 U10280 ( .A1(n9199), .A2(n8707), .ZN(n8708) );
  MUX2_X1 U10281 ( .A(n8709), .B(n8708), .S(n8748), .Z(n8713) );
  INV_X1 U10282 ( .A(n8710), .ZN(n8711) );
  OAI21_X1 U10283 ( .B1(n8717), .B2(n8711), .A(n8748), .ZN(n8712) );
  AOI21_X1 U10284 ( .B1(n8716), .B2(n8714), .A(n8748), .ZN(n8715) );
  NAND2_X1 U10285 ( .A1(n8764), .A2(n8718), .ZN(n8721) );
  INV_X1 U10286 ( .A(n8719), .ZN(n8720) );
  MUX2_X1 U10287 ( .A(n8721), .B(n8720), .S(n8748), .Z(n8722) );
  INV_X1 U10288 ( .A(n8723), .ZN(n8724) );
  OAI21_X1 U10289 ( .B1(n8725), .B2(n8724), .A(n8763), .ZN(n8728) );
  INV_X1 U10290 ( .A(n9158), .ZN(n8726) );
  INV_X1 U10291 ( .A(n9118), .ZN(n8730) );
  OR2_X1 U10292 ( .A1(n8734), .A2(n8730), .ZN(n9132) );
  INV_X1 U10293 ( .A(n9132), .ZN(n9130) );
  MUX2_X1 U10294 ( .A(n8732), .B(n8731), .S(n8748), .Z(n8733) );
  INV_X1 U10295 ( .A(n8734), .ZN(n8735) );
  MUX2_X1 U10296 ( .A(n8735), .B(n9118), .S(n8748), .Z(n8736) );
  NAND3_X1 U10297 ( .A1(n8737), .A2(n8789), .A3(n8736), .ZN(n8741) );
  NAND2_X1 U10298 ( .A1(n9293), .A2(n8843), .ZN(n8739) );
  MUX2_X1 U10299 ( .A(n8739), .B(n8738), .S(n8748), .Z(n8740) );
  NAND3_X1 U10300 ( .A1(n5733), .A2(n8741), .A3(n8740), .ZN(n8744) );
  OAI21_X1 U10301 ( .B1(n8743), .B2(n8742), .A(n8744), .ZN(n8751) );
  NOR2_X1 U10302 ( .A1(n8744), .A2(n8743), .ZN(n8750) );
  AOI211_X1 U10303 ( .C1(n8746), .C2(n8751), .A(n8745), .B(n8750), .ZN(n8757)
         );
  INV_X1 U10304 ( .A(n8747), .ZN(n8749) );
  NOR2_X1 U10305 ( .A1(n8749), .A2(n8748), .ZN(n8756) );
  INV_X1 U10306 ( .A(n8750), .ZN(n8754) );
  NAND2_X1 U10307 ( .A1(n8751), .A2(n9290), .ZN(n8752) );
  NAND4_X1 U10308 ( .A1(n8754), .A2(n8753), .A3(n8752), .A4(n8791), .ZN(n8755)
         );
  OAI21_X1 U10309 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n8760) );
  INV_X1 U10310 ( .A(n8761), .ZN(n8793) );
  NAND2_X1 U10311 ( .A1(n8763), .A2(n8762), .ZN(n9161) );
  INV_X1 U10312 ( .A(n9177), .ZN(n9175) );
  INV_X1 U10313 ( .A(n9199), .ZN(n9198) );
  NOR4_X1 U10314 ( .A1(n8767), .A2(n8766), .A3(n10344), .A4(n8765), .ZN(n8770)
         );
  NAND4_X1 U10315 ( .A1(n8770), .A2(n10332), .A3(n8769), .A4(n8768), .ZN(n8772) );
  NOR4_X1 U10316 ( .A1(n4984), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n8774)
         );
  NAND4_X1 U10317 ( .A1(n8777), .A2(n8776), .A3(n8775), .A4(n8774), .ZN(n8778)
         );
  NOR4_X1 U10318 ( .A1(n8781), .A2(n8780), .A3(n8779), .A4(n8778), .ZN(n8782)
         );
  NAND4_X1 U10319 ( .A1(n8785), .A2(n8784), .A3(n8783), .A4(n8782), .ZN(n8786)
         );
  NOR3_X1 U10320 ( .A1(n9198), .A2(n9216), .A3(n8786), .ZN(n8787) );
  NAND4_X1 U10321 ( .A1(n9165), .A2(n9175), .A3(n9189), .A4(n8787), .ZN(n8788)
         );
  NOR4_X1 U10322 ( .A1(n9132), .A2(n9147), .A3(n9161), .A4(n8788), .ZN(n8790)
         );
  NAND4_X1 U10323 ( .A1(n8791), .A2(n8790), .A3(n9104), .A4(n8789), .ZN(n8792)
         );
  NOR3_X1 U10324 ( .A1(n8794), .A2(n8793), .A3(n8792), .ZN(n8795) );
  OAI22_X1 U10325 ( .A1(n8795), .A2(n6942), .B1(n9100), .B2(n9097), .ZN(n8796)
         );
  NOR3_X1 U10326 ( .A1(n8800), .A2(n8799), .A3(n5680), .ZN(n8803) );
  OAI21_X1 U10327 ( .B1(n8804), .B2(n8801), .A(P2_B_REG_SCAN_IN), .ZN(n8802)
         );
  OAI22_X1 U10328 ( .A1(n8805), .A2(n8804), .B1(n8803), .B2(n8802), .ZN(
        P2_U3296) );
  NAND2_X1 U10329 ( .A1(n8806), .A2(n9211), .ZN(n8811) );
  NOR2_X1 U10330 ( .A1(n8807), .A2(n10343), .ZN(n9098) );
  NOR2_X1 U10331 ( .A1(n8808), .A2(n10334), .ZN(n8809) );
  AOI211_X1 U10332 ( .C1(n10339), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9098), .B(
        n8809), .ZN(n8810) );
  OAI211_X1 U10333 ( .C1(n8813), .C2(n8812), .A(n8811), .B(n8810), .ZN(
        P2_U3204) );
  INV_X1 U10334 ( .A(n8814), .ZN(n8891) );
  XNOR2_X1 U10335 ( .A(n8889), .B(n8838), .ZN(n8816) );
  NAND2_X1 U10336 ( .A1(n8816), .A2(n8815), .ZN(n8819) );
  INV_X1 U10337 ( .A(n8816), .ZN(n8817) );
  NAND2_X1 U10338 ( .A1(n8817), .A2(n8958), .ZN(n8818) );
  NAND2_X1 U10339 ( .A1(n8819), .A2(n8818), .ZN(n8890) );
  INV_X1 U10340 ( .A(n8819), .ZN(n8926) );
  XNOR2_X1 U10341 ( .A(n8924), .B(n8838), .ZN(n8820) );
  XNOR2_X1 U10342 ( .A(n8820), .B(n8957), .ZN(n8925) );
  XNOR2_X1 U10343 ( .A(n9339), .B(n4527), .ZN(n8821) );
  NOR2_X1 U10344 ( .A1(n8821), .A2(n9203), .ZN(n8865) );
  NAND2_X1 U10345 ( .A1(n8821), .A2(n9203), .ZN(n8866) );
  XNOR2_X1 U10346 ( .A(n9334), .B(n8838), .ZN(n8822) );
  XNOR2_X1 U10347 ( .A(n8822), .B(n9219), .ZN(n8909) );
  INV_X1 U10348 ( .A(n8822), .ZN(n8823) );
  INV_X1 U10349 ( .A(n9219), .ZN(n8956) );
  XNOR2_X1 U10350 ( .A(n9191), .B(n8838), .ZN(n8824) );
  XNOR2_X1 U10351 ( .A(n8824), .B(n9204), .ZN(n8876) );
  XNOR2_X1 U10352 ( .A(n9324), .B(n8838), .ZN(n8826) );
  XNOR2_X1 U10353 ( .A(n8826), .B(n9168), .ZN(n8916) );
  NAND2_X1 U10354 ( .A1(n8917), .A2(n8916), .ZN(n8915) );
  XNOR2_X1 U10355 ( .A(n9317), .B(n4527), .ZN(n8828) );
  XNOR2_X1 U10356 ( .A(n9311), .B(n8838), .ZN(n8830) );
  XNOR2_X1 U10357 ( .A(n8830), .B(n9167), .ZN(n8902) );
  XNOR2_X1 U10358 ( .A(n9305), .B(n8838), .ZN(n8832) );
  XOR2_X1 U10359 ( .A(n9153), .B(n8832), .Z(n8883) );
  INV_X1 U10360 ( .A(n8832), .ZN(n8833) );
  XNOR2_X1 U10361 ( .A(n9299), .B(n4527), .ZN(n8942) );
  NOR2_X1 U10362 ( .A1(n8942), .A2(n9124), .ZN(n8835) );
  INV_X1 U10363 ( .A(n8942), .ZN(n8834) );
  XNOR2_X1 U10364 ( .A(n9293), .B(n8838), .ZN(n8836) );
  XNOR2_X1 U10365 ( .A(n8836), .B(n9134), .ZN(n8852) );
  INV_X1 U10366 ( .A(n8836), .ZN(n8837) );
  AOI22_X1 U10367 ( .A1(n8853), .A2(n8852), .B1(n8837), .B2(n9134), .ZN(n8840)
         );
  XOR2_X1 U10368 ( .A(n8838), .B(n9104), .Z(n8839) );
  XNOR2_X1 U10369 ( .A(n8840), .B(n8839), .ZN(n8846) );
  NAND2_X1 U10370 ( .A1(n9107), .A2(n8944), .ZN(n8842) );
  AOI22_X1 U10371 ( .A1(n9113), .A2(n8945), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8841) );
  OAI211_X1 U10372 ( .C1(n8843), .C2(n8948), .A(n8842), .B(n8841), .ZN(n8844)
         );
  AOI21_X1 U10373 ( .B1(n9114), .B2(n8951), .A(n8844), .ZN(n8845) );
  OAI21_X1 U10374 ( .B1(n8846), .B2(n8953), .A(n8845), .ZN(P2_U3160) );
  OAI222_X1 U10375 ( .A1(n9952), .A2(n8848), .B1(n9949), .B2(n8847), .C1(
        P1_U3086), .C2(n4507), .ZN(P1_U3336) );
  INV_X1 U10376 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8850) );
  OAI222_X1 U10377 ( .A1(n5790), .A2(P2_U3151), .B1(n9355), .B2(n8851), .C1(
        n8850), .C2(n8849), .ZN(P2_U3274) );
  XNOR2_X1 U10378 ( .A(n8853), .B(n8852), .ZN(n8858) );
  NAND2_X1 U10379 ( .A1(n9123), .A2(n8944), .ZN(n8855) );
  AOI22_X1 U10380 ( .A1(n9127), .A2(n8945), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8854) );
  OAI211_X1 U10381 ( .C1(n9143), .C2(n8948), .A(n8855), .B(n8854), .ZN(n8856)
         );
  AOI21_X1 U10382 ( .B1(n9293), .B2(n8951), .A(n8856), .ZN(n8857) );
  OAI21_X1 U10383 ( .B1(n8858), .B2(n8953), .A(n8857), .ZN(P2_U3154) );
  XNOR2_X1 U10384 ( .A(n8859), .B(n8919), .ZN(n8864) );
  AOI22_X1 U10385 ( .A1(n9168), .A2(n8931), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8861) );
  NAND2_X1 U10386 ( .A1(n9171), .A2(n8945), .ZN(n8860) );
  OAI211_X1 U10387 ( .C1(n9142), .C2(n8933), .A(n8861), .B(n8860), .ZN(n8862)
         );
  AOI21_X1 U10388 ( .B1(n9317), .B2(n8951), .A(n8862), .ZN(n8863) );
  OAI21_X1 U10389 ( .B1(n8864), .B2(n8953), .A(n8863), .ZN(P2_U3156) );
  INV_X1 U10390 ( .A(n8865), .ZN(n8867) );
  NAND2_X1 U10391 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  XNOR2_X1 U10392 ( .A(n8869), .B(n8868), .ZN(n8874) );
  NAND2_X1 U10393 ( .A1(n8931), .A2(n8957), .ZN(n8870) );
  NAND2_X1 U10394 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9091) );
  OAI211_X1 U10395 ( .C1(n9219), .C2(n8933), .A(n8870), .B(n9091), .ZN(n8871)
         );
  AOI21_X1 U10396 ( .B1(n9224), .B2(n8945), .A(n8871), .ZN(n8873) );
  NAND2_X1 U10397 ( .A1(n9339), .A2(n8951), .ZN(n8872) );
  OAI211_X1 U10398 ( .C1(n8874), .C2(n8953), .A(n8873), .B(n8872), .ZN(
        P2_U3159) );
  XOR2_X1 U10399 ( .A(n8876), .B(n8875), .Z(n8881) );
  AOI22_X1 U10400 ( .A1(n9168), .A2(n8944), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8878) );
  NAND2_X1 U10401 ( .A1(n8945), .A2(n9192), .ZN(n8877) );
  OAI211_X1 U10402 ( .C1(n9219), .C2(n8948), .A(n8878), .B(n8877), .ZN(n8879)
         );
  AOI21_X1 U10403 ( .B1(n9191), .B2(n8951), .A(n8879), .ZN(n8880) );
  OAI21_X1 U10404 ( .B1(n8881), .B2(n8953), .A(n8880), .ZN(P2_U3163) );
  XOR2_X1 U10405 ( .A(n8883), .B(n8882), .Z(n8888) );
  AOI22_X1 U10406 ( .A1(n9167), .A2(n8931), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8885) );
  NAND2_X1 U10407 ( .A1(n9145), .A2(n8945), .ZN(n8884) );
  OAI211_X1 U10408 ( .C1(n9143), .C2(n8933), .A(n8885), .B(n8884), .ZN(n8886)
         );
  AOI21_X1 U10409 ( .B1(n9305), .B2(n8951), .A(n8886), .ZN(n8887) );
  OAI21_X1 U10410 ( .B1(n8888), .B2(n8953), .A(n8887), .ZN(P2_U3165) );
  INV_X1 U10411 ( .A(n8889), .ZN(n8900) );
  AND3_X1 U10412 ( .A1(n8892), .A2(n8891), .A3(n8890), .ZN(n8893) );
  OAI21_X1 U10413 ( .B1(n8927), .B2(n8893), .A(n8928), .ZN(n8899) );
  NAND2_X1 U10414 ( .A1(n8944), .A2(n8957), .ZN(n8894) );
  NAND2_X1 U10415 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9039) );
  OAI211_X1 U10416 ( .C1(n8895), .C2(n8948), .A(n8894), .B(n9039), .ZN(n8896)
         );
  AOI21_X1 U10417 ( .B1(n8897), .B2(n8945), .A(n8896), .ZN(n8898) );
  OAI211_X1 U10418 ( .C1(n8900), .C2(n8939), .A(n8899), .B(n8898), .ZN(
        P2_U3168) );
  XOR2_X1 U10419 ( .A(n8902), .B(n8901), .Z(n8907) );
  AOI22_X1 U10420 ( .A1(n9179), .A2(n8931), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8904) );
  NAND2_X1 U10421 ( .A1(n9157), .A2(n8945), .ZN(n8903) );
  OAI211_X1 U10422 ( .C1(n8949), .C2(n8933), .A(n8904), .B(n8903), .ZN(n8905)
         );
  AOI21_X1 U10423 ( .B1(n9311), .B2(n8951), .A(n8905), .ZN(n8906) );
  OAI21_X1 U10424 ( .B1(n8907), .B2(n8953), .A(n8906), .ZN(P2_U3169) );
  XOR2_X1 U10425 ( .A(n8909), .B(n8908), .Z(n8914) );
  AOI22_X1 U10426 ( .A1(n9204), .A2(n8944), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8911) );
  NAND2_X1 U10427 ( .A1(n8945), .A2(n9207), .ZN(n8910) );
  OAI211_X1 U10428 ( .C1(n8934), .C2(n8948), .A(n8911), .B(n8910), .ZN(n8912)
         );
  AOI21_X1 U10429 ( .B1(n9334), .B2(n8951), .A(n8912), .ZN(n8913) );
  OAI21_X1 U10430 ( .B1(n8914), .B2(n8953), .A(n8913), .ZN(P2_U3173) );
  OAI211_X1 U10431 ( .C1(n8917), .C2(n8916), .A(n8915), .B(n8928), .ZN(n8922)
         );
  AOI22_X1 U10432 ( .A1(n9204), .A2(n8931), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8918) );
  OAI21_X1 U10433 ( .B1(n8919), .B2(n8933), .A(n8918), .ZN(n8920) );
  AOI21_X1 U10434 ( .B1(n9182), .B2(n8945), .A(n8920), .ZN(n8921) );
  OAI211_X1 U10435 ( .C1(n8923), .C2(n8939), .A(n8922), .B(n8921), .ZN(
        P2_U3175) );
  INV_X1 U10436 ( .A(n8924), .ZN(n8940) );
  NOR3_X1 U10437 ( .A1(n8927), .A2(n8926), .A3(n8925), .ZN(n8929) );
  OAI21_X1 U10438 ( .B1(n4594), .B2(n8929), .A(n8928), .ZN(n8938) );
  NOR2_X1 U10439 ( .A1(n8930), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9065) );
  AOI21_X1 U10440 ( .B1(n8931), .B2(n8958), .A(n9065), .ZN(n8932) );
  OAI21_X1 U10441 ( .B1(n8934), .B2(n8933), .A(n8932), .ZN(n8935) );
  AOI21_X1 U10442 ( .B1(n8936), .B2(n8945), .A(n8935), .ZN(n8937) );
  OAI211_X1 U10443 ( .C1(n8940), .C2(n8939), .A(n8938), .B(n8937), .ZN(
        P2_U3178) );
  XNOR2_X1 U10444 ( .A(n8942), .B(n9124), .ZN(n8943) );
  XNOR2_X1 U10445 ( .A(n8941), .B(n8943), .ZN(n8954) );
  NAND2_X1 U10446 ( .A1(n9134), .A2(n8944), .ZN(n8947) );
  AOI22_X1 U10447 ( .A1(n9137), .A2(n8945), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8946) );
  OAI211_X1 U10448 ( .C1(n8949), .C2(n8948), .A(n8947), .B(n8946), .ZN(n8950)
         );
  AOI21_X1 U10449 ( .B1(n9299), .B2(n8951), .A(n8950), .ZN(n8952) );
  OAI21_X1 U10450 ( .B1(n8954), .B2(n8953), .A(n8952), .ZN(P2_U3180) );
  MUX2_X1 U10451 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8955), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10452 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9107), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10453 ( .A(n9123), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8972), .Z(
        P2_U3519) );
  MUX2_X1 U10454 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9134), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10455 ( .A(n9124), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8972), .Z(
        P2_U3517) );
  MUX2_X1 U10456 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9153), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10457 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9167), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10458 ( .A(n9179), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8972), .Z(
        P2_U3514) );
  MUX2_X1 U10459 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9168), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10460 ( .A(n9204), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8972), .Z(
        P2_U3512) );
  MUX2_X1 U10461 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8956), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10462 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9203), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10463 ( .A(n8957), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8972), .Z(
        P2_U3509) );
  MUX2_X1 U10464 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8958), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10465 ( .A(n8959), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8972), .Z(
        P2_U3507) );
  MUX2_X1 U10466 ( .A(n8960), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8972), .Z(
        P2_U3506) );
  MUX2_X1 U10467 ( .A(n8961), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8972), .Z(
        P2_U3505) );
  MUX2_X1 U10468 ( .A(n8962), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8972), .Z(
        P2_U3504) );
  MUX2_X1 U10469 ( .A(n8963), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8972), .Z(
        P2_U3503) );
  MUX2_X1 U10470 ( .A(n8964), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8972), .Z(
        P2_U3502) );
  MUX2_X1 U10471 ( .A(n8965), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8972), .Z(
        P2_U3501) );
  MUX2_X1 U10472 ( .A(n8966), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8972), .Z(
        P2_U3500) );
  MUX2_X1 U10473 ( .A(n8967), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8972), .Z(
        P2_U3499) );
  MUX2_X1 U10474 ( .A(n8968), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8972), .Z(
        P2_U3498) );
  MUX2_X1 U10475 ( .A(n8969), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8972), .Z(
        P2_U3497) );
  MUX2_X1 U10476 ( .A(n8970), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8972), .Z(
        P2_U3496) );
  MUX2_X1 U10477 ( .A(n10329), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8972), .Z(
        P2_U3495) );
  MUX2_X1 U10478 ( .A(n8971), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8972), .Z(
        P2_U3494) );
  MUX2_X1 U10479 ( .A(n10327), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8972), .Z(
        P2_U3493) );
  MUX2_X1 U10480 ( .A(n6948), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8972), .Z(
        P2_U3492) );
  MUX2_X1 U10481 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8973), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U10482 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8985), .A(n8974), .ZN(
        n8996) );
  XOR2_X1 U10483 ( .A(n9002), .B(n8996), .Z(n8975) );
  NOR2_X1 U10484 ( .A1(n8975), .A2(n8976), .ZN(n8998) );
  AOI21_X1 U10485 ( .B1(n8976), .B2(n8975), .A(n8998), .ZN(n8995) );
  MUX2_X1 U10486 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8049), .Z(n9003) );
  XNOR2_X1 U10487 ( .A(n9003), .B(n9013), .ZN(n8981) );
  OR2_X1 U10488 ( .A1(n8977), .A2(n8985), .ZN(n8979) );
  NAND2_X1 U10489 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  NAND2_X1 U10490 ( .A1(n8981), .A2(n8980), .ZN(n9004) );
  OAI21_X1 U10491 ( .B1(n8981), .B2(n8980), .A(n9004), .ZN(n8992) );
  NOR2_X1 U10492 ( .A1(n10321), .A2(n8982), .ZN(n8991) );
  INV_X1 U10493 ( .A(n10308), .ZN(n9041) );
  AOI22_X1 U10494 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8985), .B1(n8984), .B2(
        n8983), .ZN(n9012) );
  AOI21_X1 U10495 ( .B1(n8987), .B2(n8986), .A(n9014), .ZN(n8989) );
  OAI21_X1 U10496 ( .B1(n9041), .B2(n8989), .A(n8988), .ZN(n8990) );
  AOI211_X1 U10497 ( .C1(n10272), .C2(n8992), .A(n8991), .B(n8990), .ZN(n8994)
         );
  NAND2_X1 U10498 ( .A1(n9045), .A2(n9013), .ZN(n8993) );
  OAI211_X1 U10499 ( .C1(n8995), .C2(n10283), .A(n8994), .B(n8993), .ZN(
        P2_U3197) );
  NOR2_X1 U10500 ( .A1(n9013), .A2(n8996), .ZN(n8997) );
  AOI22_X1 U10501 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n9021), .B1(n9036), .B2(
        n8999), .ZN(n9000) );
  AOI21_X1 U10502 ( .B1(n9001), .B2(n9000), .A(n9025), .ZN(n9023) );
  MUX2_X1 U10503 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8049), .Z(n9029) );
  XNOR2_X1 U10504 ( .A(n9029), .B(n9021), .ZN(n9007) );
  OR2_X1 U10505 ( .A1(n9003), .A2(n9002), .ZN(n9005) );
  NAND2_X1 U10506 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U10507 ( .A1(n9007), .A2(n9006), .ZN(n9030) );
  OAI21_X1 U10508 ( .B1(n9007), .B2(n9006), .A(n9030), .ZN(n9008) );
  NAND2_X1 U10509 ( .A1(n9008), .A2(n10272), .ZN(n9010) );
  OAI211_X1 U10510 ( .C1(n10321), .C2(n9011), .A(n9010), .B(n9009), .ZN(n9020)
         );
  NOR2_X1 U10511 ( .A1(n9013), .A2(n9012), .ZN(n9015) );
  MUX2_X1 U10512 ( .A(n5432), .B(P2_REG2_REG_16__SCAN_IN), .S(n9021), .Z(n9016) );
  INV_X1 U10513 ( .A(n9016), .ZN(n9017) );
  AOI21_X1 U10514 ( .B1(n4562), .B2(n9017), .A(n9035), .ZN(n9018) );
  NOR2_X1 U10515 ( .A1(n9018), .A2(n9041), .ZN(n9019) );
  AOI211_X1 U10516 ( .C1(n9045), .C2(n9021), .A(n9020), .B(n9019), .ZN(n9022)
         );
  OAI21_X1 U10517 ( .B1(n9023), .B2(n10283), .A(n9022), .ZN(P2_U3198) );
  NOR2_X1 U10518 ( .A1(n9027), .A2(n9026), .ZN(n9051) );
  AOI21_X1 U10519 ( .B1(n9027), .B2(n9026), .A(n9051), .ZN(n9048) );
  MUX2_X1 U10520 ( .A(n9037), .B(n9027), .S(n8049), .Z(n9055) );
  XNOR2_X1 U10521 ( .A(n9028), .B(n9055), .ZN(n9033) );
  OR2_X1 U10522 ( .A1(n9029), .A2(n9036), .ZN(n9031) );
  NAND2_X1 U10523 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  OAI21_X1 U10524 ( .B1(n9033), .B2(n9032), .A(n9054), .ZN(n9044) );
  NOR2_X1 U10525 ( .A1(n10321), .A2(n9034), .ZN(n9043) );
  AOI21_X1 U10526 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9036), .A(n9035), .ZN(
        n9066) );
  XNOR2_X1 U10527 ( .A(n9067), .B(n9066), .ZN(n9038) );
  AOI21_X1 U10528 ( .B1(n9038), .B2(n9037), .A(n9068), .ZN(n9040) );
  OAI21_X1 U10529 ( .B1(n9041), .B2(n9040), .A(n9039), .ZN(n9042) );
  AOI211_X1 U10530 ( .C1(n10272), .C2(n9044), .A(n9043), .B(n9042), .ZN(n9047)
         );
  NAND2_X1 U10531 ( .A1(n9045), .A2(n9067), .ZN(n9046) );
  OAI211_X1 U10532 ( .C1(n9048), .C2(n10283), .A(n9047), .B(n9046), .ZN(
        P2_U3199) );
  NOR2_X1 U10533 ( .A1(n9067), .A2(n9049), .ZN(n9050) );
  NAND2_X1 U10534 ( .A1(n9083), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9076) );
  OAI21_X1 U10535 ( .B1(n9083), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9076), .ZN(
        n9052) );
  AOI21_X1 U10536 ( .B1(n9053), .B2(n9052), .A(n9078), .ZN(n9075) );
  MUX2_X1 U10537 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8049), .Z(n9057) );
  AND2_X1 U10538 ( .A1(n9056), .A2(n9057), .ZN(n9084) );
  INV_X1 U10539 ( .A(n9057), .ZN(n9058) );
  NAND2_X1 U10540 ( .A1(n9059), .A2(n9058), .ZN(n9082) );
  INV_X1 U10541 ( .A(n9082), .ZN(n9060) );
  NAND2_X1 U10542 ( .A1(n9061), .A2(P2_U3893), .ZN(n9062) );
  NAND2_X1 U10543 ( .A1(n10312), .A2(n9062), .ZN(n9064) );
  NOR2_X1 U10544 ( .A1(n9067), .A2(n9066), .ZN(n9069) );
  NOR2_X1 U10545 ( .A1(n9069), .A2(n9068), .ZN(n9071) );
  NAND2_X1 U10546 ( .A1(n9083), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9080) );
  OAI21_X1 U10547 ( .B1(n9083), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9080), .ZN(
        n9070) );
  AND2_X1 U10548 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  OAI21_X1 U10549 ( .B1(n9081), .B2(n9072), .A(n10308), .ZN(n9073) );
  OAI211_X1 U10550 ( .C1(n9075), .C2(n10283), .A(n9074), .B(n9073), .ZN(
        P2_U3200) );
  INV_X1 U10551 ( .A(n9076), .ZN(n9077) );
  XNOR2_X1 U10552 ( .A(n9079), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9085) );
  MUX2_X1 U10553 ( .A(n9223), .B(P2_REG2_REG_19__SCAN_IN), .S(n9093), .Z(n9087) );
  OAI21_X1 U10554 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n9089) );
  INV_X1 U10555 ( .A(n9085), .ZN(n9086) );
  MUX2_X1 U10556 ( .A(n9087), .B(n9086), .S(n8049), .Z(n9088) );
  XNOR2_X1 U10557 ( .A(n9089), .B(n9088), .ZN(n9090) );
  NAND2_X1 U10558 ( .A1(n10248), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9092) );
  OAI211_X1 U10559 ( .C1(n10312), .C2(n9093), .A(n9092), .B(n9091), .ZN(n9094)
         );
  AOI21_X1 U10560 ( .B1(n9279), .B2(n9211), .A(n9098), .ZN(n9102) );
  NAND2_X1 U10561 ( .A1(n10339), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9099) );
  OAI211_X1 U10562 ( .C1(n9100), .C2(n10334), .A(n9102), .B(n9099), .ZN(
        P2_U3202) );
  NAND2_X1 U10563 ( .A1(n10339), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9101) );
  OAI211_X1 U10564 ( .C1(n9284), .C2(n10334), .A(n9102), .B(n9101), .ZN(
        P2_U3203) );
  INV_X1 U10565 ( .A(n9287), .ZN(n9117) );
  INV_X1 U10566 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9112) );
  INV_X1 U10567 ( .A(n9104), .ZN(n9105) );
  XNOR2_X1 U10568 ( .A(n9106), .B(n9105), .ZN(n9111) );
  AOI21_X1 U10569 ( .B1(n9111), .B2(n10350), .A(n9110), .ZN(n9285) );
  MUX2_X1 U10570 ( .A(n9112), .B(n9285), .S(n10357), .Z(n9116) );
  AOI22_X1 U10571 ( .A1(n9114), .A2(n9226), .B1(n9225), .B2(n9113), .ZN(n9115)
         );
  OAI211_X1 U10572 ( .C1(n9117), .C2(n9229), .A(n9116), .B(n9115), .ZN(
        P2_U3205) );
  NAND2_X1 U10573 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  XNOR2_X1 U10574 ( .A(n9120), .B(n9121), .ZN(n9296) );
  INV_X1 U10575 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9126) );
  XNOR2_X1 U10576 ( .A(n9122), .B(n9121), .ZN(n9125) );
  AOI222_X1 U10577 ( .A1(n10350), .A2(n9125), .B1(n9124), .B2(n10326), .C1(
        n9123), .C2(n10328), .ZN(n9291) );
  MUX2_X1 U10578 ( .A(n9126), .B(n9291), .S(n10357), .Z(n9129) );
  AOI22_X1 U10579 ( .A1(n9293), .A2(n9226), .B1(n9225), .B2(n9127), .ZN(n9128)
         );
  OAI211_X1 U10580 ( .C1(n9296), .C2(n9229), .A(n9129), .B(n9128), .ZN(
        P2_U3206) );
  XNOR2_X1 U10581 ( .A(n9131), .B(n9130), .ZN(n9302) );
  INV_X1 U10582 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9136) );
  XNOR2_X1 U10583 ( .A(n9133), .B(n9132), .ZN(n9135) );
  AOI222_X1 U10584 ( .A1(n10350), .A2(n9135), .B1(n9153), .B2(n10326), .C1(
        n9134), .C2(n10328), .ZN(n9297) );
  MUX2_X1 U10585 ( .A(n9136), .B(n9297), .S(n10357), .Z(n9139) );
  AOI22_X1 U10586 ( .A1(n9299), .A2(n9226), .B1(n9225), .B2(n9137), .ZN(n9138)
         );
  OAI211_X1 U10587 ( .C1(n9302), .C2(n9229), .A(n9139), .B(n9138), .ZN(
        P2_U3207) );
  XNOR2_X1 U10588 ( .A(n9140), .B(n9147), .ZN(n9141) );
  OAI222_X1 U10589 ( .A1(n10346), .A2(n9143), .B1(n10348), .B2(n9142), .C1(
        n9187), .C2(n9141), .ZN(n9245) );
  AOI21_X1 U10590 ( .B1(n9144), .B2(n9305), .A(n9245), .ZN(n9150) );
  AOI22_X1 U10591 ( .A1(n9145), .A2(n9225), .B1(n10339), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9149) );
  XNOR2_X1 U10592 ( .A(n9146), .B(n9147), .ZN(n9306) );
  NAND2_X1 U10593 ( .A1(n9306), .A2(n10336), .ZN(n9148) );
  OAI211_X1 U10594 ( .C1(n9150), .C2(n10339), .A(n9149), .B(n9148), .ZN(
        P2_U3208) );
  NOR2_X1 U10595 ( .A1(n9151), .A2(n10341), .ZN(n9156) );
  XOR2_X1 U10596 ( .A(n9161), .B(n9152), .Z(n9154) );
  AOI222_X1 U10597 ( .A1(n10350), .A2(n9154), .B1(n9179), .B2(n10326), .C1(
        n9153), .C2(n10328), .ZN(n9309) );
  INV_X1 U10598 ( .A(n9309), .ZN(n9155) );
  AOI211_X1 U10599 ( .C1(n9225), .C2(n9157), .A(n9156), .B(n9155), .ZN(n9163)
         );
  NAND2_X1 U10600 ( .A1(n9159), .A2(n9158), .ZN(n9160) );
  XOR2_X1 U10601 ( .A(n9161), .B(n9160), .Z(n9312) );
  AOI22_X1 U10602 ( .A1(n9312), .A2(n10336), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10339), .ZN(n9162) );
  OAI21_X1 U10603 ( .B1(n9163), .B2(n10339), .A(n9162), .ZN(P2_U3209) );
  XNOR2_X1 U10604 ( .A(n9164), .B(n9165), .ZN(n9319) );
  INV_X1 U10605 ( .A(n9319), .ZN(n9174) );
  INV_X1 U10606 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9170) );
  XNOR2_X1 U10607 ( .A(n9166), .B(n9165), .ZN(n9169) );
  AOI222_X1 U10608 ( .A1(n10350), .A2(n9169), .B1(n9168), .B2(n10326), .C1(
        n9167), .C2(n10328), .ZN(n9315) );
  MUX2_X1 U10609 ( .A(n9170), .B(n9315), .S(n10357), .Z(n9173) );
  AOI22_X1 U10610 ( .A1(n9317), .A2(n9226), .B1(n9225), .B2(n9171), .ZN(n9172)
         );
  OAI211_X1 U10611 ( .C1(n9174), .C2(n9229), .A(n9173), .B(n9172), .ZN(
        P2_U3210) );
  XNOR2_X1 U10612 ( .A(n9176), .B(n9175), .ZN(n9327) );
  INV_X1 U10613 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9181) );
  XNOR2_X1 U10614 ( .A(n9178), .B(n9177), .ZN(n9180) );
  AOI222_X1 U10615 ( .A1(n10350), .A2(n9180), .B1(n9179), .B2(n10328), .C1(
        n9204), .C2(n10326), .ZN(n9322) );
  MUX2_X1 U10616 ( .A(n9181), .B(n9322), .S(n10357), .Z(n9184) );
  AOI22_X1 U10617 ( .A1(n9324), .A2(n9226), .B1(n9225), .B2(n9182), .ZN(n9183)
         );
  OAI211_X1 U10618 ( .C1(n9327), .C2(n9229), .A(n9184), .B(n9183), .ZN(
        P2_U3211) );
  XOR2_X1 U10619 ( .A(n9189), .B(n9185), .Z(n9186) );
  OAI222_X1 U10620 ( .A1(n10346), .A2(n9188), .B1(n10348), .B2(n9219), .C1(
        n9187), .C2(n9186), .ZN(n9259) );
  INV_X1 U10621 ( .A(n9259), .ZN(n9196) );
  XNOR2_X1 U10622 ( .A(n9190), .B(n9189), .ZN(n9260) );
  AOI22_X1 U10623 ( .A1(n9225), .A2(n9192), .B1(n10339), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n9193) );
  OAI21_X1 U10624 ( .B1(n4828), .B2(n10334), .A(n9193), .ZN(n9194) );
  AOI21_X1 U10625 ( .B1(n9260), .B2(n10336), .A(n9194), .ZN(n9195) );
  OAI21_X1 U10626 ( .B1(n9196), .B2(n10339), .A(n9195), .ZN(P2_U3212) );
  XNOR2_X1 U10627 ( .A(n9197), .B(n9198), .ZN(n9264) );
  INV_X1 U10628 ( .A(n9264), .ZN(n9213) );
  AND2_X1 U10629 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  OAI21_X1 U10630 ( .B1(n9202), .B2(n9201), .A(n10350), .ZN(n9206) );
  AOI22_X1 U10631 ( .A1(n9204), .A2(n10328), .B1(n10326), .B2(n9203), .ZN(
        n9205) );
  NAND2_X1 U10632 ( .A1(n9206), .A2(n9205), .ZN(n9266) );
  AOI22_X1 U10633 ( .A1(n10339), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9207), 
        .B2(n9225), .ZN(n9208) );
  OAI21_X1 U10634 ( .B1(n9209), .B2(n10334), .A(n9208), .ZN(n9210) );
  AOI21_X1 U10635 ( .B1(n9266), .B2(n9211), .A(n9210), .ZN(n9212) );
  OAI21_X1 U10636 ( .B1(n9213), .B2(n9229), .A(n9212), .ZN(P2_U3213) );
  XOR2_X1 U10637 ( .A(n9214), .B(n9216), .Z(n9343) );
  OAI211_X1 U10638 ( .C1(n9217), .C2(n9216), .A(n9215), .B(n10350), .ZN(n9222)
         );
  OAI22_X1 U10639 ( .A1(n9219), .A2(n10346), .B1(n9218), .B2(n10348), .ZN(
        n9220) );
  INV_X1 U10640 ( .A(n9220), .ZN(n9221) );
  MUX2_X1 U10641 ( .A(n9337), .B(n9223), .S(n10339), .Z(n9228) );
  AOI22_X1 U10642 ( .A1(n9339), .A2(n9226), .B1(n9225), .B2(n9224), .ZN(n9227)
         );
  OAI211_X1 U10643 ( .C1(n9343), .C2(n9229), .A(n9228), .B(n9227), .ZN(
        P2_U3214) );
  NAND2_X1 U10644 ( .A1(n9278), .A2(n9270), .ZN(n9230) );
  NAND2_X1 U10645 ( .A1(n9279), .A2(n10440), .ZN(n9232) );
  OAI211_X1 U10646 ( .C1(n10440), .C2(n7423), .A(n9230), .B(n9232), .ZN(
        P2_U3490) );
  NAND2_X1 U10647 ( .A1(n9231), .A2(n9270), .ZN(n9233) );
  OAI211_X1 U10648 ( .C1(n10440), .C2(n5684), .A(n9233), .B(n9232), .ZN(
        P2_U3489) );
  NAND2_X1 U10649 ( .A1(n10437), .A2(n9234), .ZN(n9235) );
  NAND2_X1 U10650 ( .A1(n9287), .A2(n9253), .ZN(n9237) );
  OAI211_X1 U10651 ( .C1(n9290), .C2(n9263), .A(n9238), .B(n9237), .ZN(
        P2_U3487) );
  MUX2_X1 U10652 ( .A(n9239), .B(n9291), .S(n10440), .Z(n9241) );
  NAND2_X1 U10653 ( .A1(n9293), .A2(n9270), .ZN(n9240) );
  OAI211_X1 U10654 ( .C1(n9296), .C2(n9273), .A(n9241), .B(n9240), .ZN(
        P2_U3486) );
  MUX2_X1 U10655 ( .A(n9242), .B(n9297), .S(n10440), .Z(n9244) );
  NAND2_X1 U10656 ( .A1(n9299), .A2(n9270), .ZN(n9243) );
  OAI211_X1 U10657 ( .C1(n9302), .C2(n9273), .A(n9244), .B(n9243), .ZN(
        P2_U3485) );
  INV_X1 U10658 ( .A(n9245), .ZN(n9303) );
  MUX2_X1 U10659 ( .A(n9246), .B(n9303), .S(n10440), .Z(n9248) );
  AOI22_X1 U10660 ( .A1(n9306), .A2(n9253), .B1(n9270), .B2(n9305), .ZN(n9247)
         );
  NAND2_X1 U10661 ( .A1(n9248), .A2(n9247), .ZN(P2_U3484) );
  MUX2_X1 U10662 ( .A(n9249), .B(n9309), .S(n10440), .Z(n9251) );
  AOI22_X1 U10663 ( .A1(n9312), .A2(n9253), .B1(n9270), .B2(n9311), .ZN(n9250)
         );
  NAND2_X1 U10664 ( .A1(n9251), .A2(n9250), .ZN(P2_U3483) );
  MUX2_X1 U10665 ( .A(n9252), .B(n9315), .S(n10440), .Z(n9255) );
  AOI22_X1 U10666 ( .A1(n9319), .A2(n9253), .B1(n9270), .B2(n9317), .ZN(n9254)
         );
  NAND2_X1 U10667 ( .A1(n9255), .A2(n9254), .ZN(P2_U3482) );
  MUX2_X1 U10668 ( .A(n9256), .B(n9322), .S(n10440), .Z(n9258) );
  NAND2_X1 U10669 ( .A1(n9324), .A2(n9270), .ZN(n9257) );
  OAI211_X1 U10670 ( .C1(n9327), .C2(n9273), .A(n9258), .B(n9257), .ZN(
        P2_U3481) );
  AOI21_X1 U10671 ( .B1(n9260), .B2(n10414), .A(n9259), .ZN(n9328) );
  MUX2_X1 U10672 ( .A(n9261), .B(n9328), .S(n10440), .Z(n9262) );
  OAI21_X1 U10673 ( .B1(n4828), .B2(n9263), .A(n9262), .ZN(P2_U3480) );
  AND2_X1 U10674 ( .A1(n9264), .A2(n10414), .ZN(n9265) );
  MUX2_X1 U10675 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9332), .S(n10440), .Z(
        n9267) );
  AOI21_X1 U10676 ( .B1(n9270), .B2(n9334), .A(n9267), .ZN(n9268) );
  INV_X1 U10677 ( .A(n9268), .ZN(P2_U3479) );
  INV_X1 U10678 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9269) );
  MUX2_X1 U10679 ( .A(n9269), .B(n9337), .S(n10440), .Z(n9272) );
  NAND2_X1 U10680 ( .A1(n9339), .A2(n9270), .ZN(n9271) );
  OAI211_X1 U10681 ( .C1(n9273), .C2(n9343), .A(n9272), .B(n9271), .ZN(
        P2_U3478) );
  AOI22_X1 U10682 ( .A1(n9275), .A2(n10414), .B1(n10416), .B2(n9274), .ZN(
        n9276) );
  NAND2_X1 U10683 ( .A1(n9277), .A2(n9276), .ZN(n9344) );
  MUX2_X1 U10684 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9344), .S(n10440), .Z(
        P2_U3475) );
  INV_X1 U10685 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U10686 ( .A1(n9278), .A2(n9338), .ZN(n9280) );
  NAND2_X1 U10687 ( .A1(n9279), .A2(n10421), .ZN(n9282) );
  OAI211_X1 U10688 ( .C1(n9281), .C2(n10421), .A(n9280), .B(n9282), .ZN(
        P2_U3458) );
  NAND2_X1 U10689 ( .A1(n10423), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9283) );
  OAI211_X1 U10690 ( .C1(n9284), .C2(n9331), .A(n9283), .B(n9282), .ZN(
        P2_U3457) );
  INV_X1 U10691 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9286) );
  MUX2_X1 U10692 ( .A(n9286), .B(n9285), .S(n10421), .Z(n9289) );
  NAND2_X1 U10693 ( .A1(n9287), .A2(n9318), .ZN(n9288) );
  OAI211_X1 U10694 ( .C1(n9290), .C2(n9331), .A(n9289), .B(n9288), .ZN(
        P2_U3455) );
  INV_X1 U10695 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9292) );
  MUX2_X1 U10696 ( .A(n9292), .B(n9291), .S(n10421), .Z(n9295) );
  NAND2_X1 U10697 ( .A1(n9293), .A2(n9338), .ZN(n9294) );
  OAI211_X1 U10698 ( .C1(n9296), .C2(n9342), .A(n9295), .B(n9294), .ZN(
        P2_U3454) );
  INV_X1 U10699 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9298) );
  MUX2_X1 U10700 ( .A(n9298), .B(n9297), .S(n10421), .Z(n9301) );
  NAND2_X1 U10701 ( .A1(n9299), .A2(n9338), .ZN(n9300) );
  OAI211_X1 U10702 ( .C1(n9302), .C2(n9342), .A(n9301), .B(n9300), .ZN(
        P2_U3453) );
  INV_X1 U10703 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9304) );
  MUX2_X1 U10704 ( .A(n9304), .B(n9303), .S(n10421), .Z(n9308) );
  AOI22_X1 U10705 ( .A1(n9306), .A2(n9318), .B1(n9338), .B2(n9305), .ZN(n9307)
         );
  NAND2_X1 U10706 ( .A1(n9308), .A2(n9307), .ZN(P2_U3452) );
  INV_X1 U10707 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9310) );
  MUX2_X1 U10708 ( .A(n9310), .B(n9309), .S(n10421), .Z(n9314) );
  AOI22_X1 U10709 ( .A1(n9312), .A2(n9318), .B1(n9338), .B2(n9311), .ZN(n9313)
         );
  NAND2_X1 U10710 ( .A1(n9314), .A2(n9313), .ZN(P2_U3451) );
  INV_X1 U10711 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9316) );
  MUX2_X1 U10712 ( .A(n9316), .B(n9315), .S(n10421), .Z(n9321) );
  AOI22_X1 U10713 ( .A1(n9319), .A2(n9318), .B1(n9338), .B2(n9317), .ZN(n9320)
         );
  NAND2_X1 U10714 ( .A1(n9321), .A2(n9320), .ZN(P2_U3450) );
  INV_X1 U10715 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9323) );
  MUX2_X1 U10716 ( .A(n9323), .B(n9322), .S(n10421), .Z(n9326) );
  NAND2_X1 U10717 ( .A1(n9324), .A2(n9338), .ZN(n9325) );
  OAI211_X1 U10718 ( .C1(n9327), .C2(n9342), .A(n9326), .B(n9325), .ZN(
        P2_U3449) );
  INV_X1 U10719 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9329) );
  MUX2_X1 U10720 ( .A(n9329), .B(n9328), .S(n10421), .Z(n9330) );
  OAI21_X1 U10721 ( .B1(n4828), .B2(n9331), .A(n9330), .ZN(P2_U3448) );
  MUX2_X1 U10722 ( .A(n9332), .B(P2_REG0_REG_20__SCAN_IN), .S(n10423), .Z(
        n9333) );
  AOI21_X1 U10723 ( .B1(n9338), .B2(n9334), .A(n9333), .ZN(n9335) );
  INV_X1 U10724 ( .A(n9335), .ZN(P2_U3447) );
  INV_X1 U10725 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9336) );
  MUX2_X1 U10726 ( .A(n9337), .B(n9336), .S(n10423), .Z(n9341) );
  NAND2_X1 U10727 ( .A1(n9339), .A2(n9338), .ZN(n9340) );
  OAI211_X1 U10728 ( .C1(n9343), .C2(n9342), .A(n9341), .B(n9340), .ZN(
        P2_U3446) );
  MUX2_X1 U10729 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9344), .S(n10421), .Z(
        P2_U3438) );
  INV_X1 U10730 ( .A(n9345), .ZN(n9943) );
  NOR4_X1 U10731 ( .A1(n9348), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9346), .ZN(n9349) );
  AOI21_X1 U10732 ( .B1(n9352), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9349), .ZN(
        n9350) );
  OAI21_X1 U10733 ( .B1(n9943), .B2(n9355), .A(n9350), .ZN(P2_U3264) );
  INV_X1 U10734 ( .A(n9351), .ZN(n9947) );
  AOI22_X1 U10735 ( .A1(n9353), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9352), .ZN(n9354) );
  OAI21_X1 U10736 ( .B1(n9947), .B2(n9355), .A(n9354), .ZN(P2_U3265) );
  MUX2_X1 U10737 ( .A(n9356), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10738 ( .B1(n9469), .B2(n9358), .A(n9357), .ZN(n9360) );
  OAI21_X1 U10739 ( .B1(n9360), .B2(n9359), .A(n10000), .ZN(n9364) );
  AOI22_X1 U10740 ( .A1(n9472), .A2(n9723), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9363) );
  INV_X1 U10741 ( .A(n9748), .ZN(n9498) );
  INV_X1 U10742 ( .A(n9721), .ZN(n9668) );
  AOI22_X1 U10743 ( .A1(n9474), .A2(n9498), .B1(n9473), .B2(n9668), .ZN(n9362)
         );
  NAND2_X1 U10744 ( .A1(n9874), .A2(n9492), .ZN(n9361) );
  NAND4_X1 U10745 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(
        P1_U3214) );
  XOR2_X1 U10746 ( .A(n9366), .B(n9365), .Z(n9372) );
  INV_X1 U10747 ( .A(n9367), .ZN(n9842) );
  OAI22_X1 U10748 ( .A1(n10003), .A2(n9842), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9368), .ZN(n9370) );
  OAI22_X1 U10749 ( .A1(n9837), .A2(n9488), .B1(n9487), .B2(n9807), .ZN(n9369)
         );
  AOI211_X1 U10750 ( .C1(n9850), .C2(n9492), .A(n9370), .B(n9369), .ZN(n9371)
         );
  OAI21_X1 U10751 ( .B1(n9372), .B2(n9494), .A(n9371), .ZN(P1_U3219) );
  XNOR2_X1 U10752 ( .A(n9373), .B(n9374), .ZN(n9379) );
  INV_X1 U10753 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9375) );
  OAI22_X1 U10754 ( .A1(n10003), .A2(n9811), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9375), .ZN(n9377) );
  OAI22_X1 U10755 ( .A1(n9807), .A2(n9488), .B1(n9487), .B2(n9808), .ZN(n9376)
         );
  AOI211_X1 U10756 ( .C1(n9906), .C2(n9492), .A(n9377), .B(n9376), .ZN(n9378)
         );
  OAI21_X1 U10757 ( .B1(n9379), .B2(n9494), .A(n9378), .ZN(P1_U3223) );
  NAND2_X1 U10758 ( .A1(n9414), .A2(n9381), .ZN(n9382) );
  OAI21_X1 U10759 ( .B1(n9383), .B2(n9382), .A(n9468), .ZN(n9384) );
  NAND2_X1 U10760 ( .A1(n9384), .A2(n10000), .ZN(n9388) );
  AOI22_X1 U10761 ( .A1(n9472), .A2(n9750), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9387) );
  INV_X1 U10762 ( .A(n9747), .ZN(n9658) );
  AOI22_X1 U10763 ( .A1(n9474), .A2(n9658), .B1(n9473), .B2(n9498), .ZN(n9386)
         );
  NAND2_X1 U10764 ( .A1(n9884), .A2(n9492), .ZN(n9385) );
  NAND4_X1 U10765 ( .A1(n9388), .A2(n9387), .A3(n9386), .A4(n9385), .ZN(
        P1_U3225) );
  NAND2_X1 U10766 ( .A1(n9391), .A2(n9390), .ZN(n9392) );
  XNOR2_X1 U10767 ( .A(n9389), .B(n9392), .ZN(n9400) );
  INV_X1 U10768 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9393) );
  OAI22_X1 U10769 ( .A1(n10003), .A2(n9394), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9393), .ZN(n9397) );
  OAI22_X1 U10770 ( .A1(n9395), .A2(n9488), .B1(n9487), .B2(n9462), .ZN(n9396)
         );
  AOI211_X1 U10771 ( .C1(n9398), .C2(n9492), .A(n9397), .B(n9396), .ZN(n9399)
         );
  OAI21_X1 U10772 ( .B1(n9400), .B2(n9494), .A(n9399), .ZN(P1_U3226) );
  INV_X1 U10773 ( .A(n9404), .ZN(n9401) );
  NOR2_X1 U10774 ( .A1(n9402), .A2(n9401), .ZN(n9407) );
  AOI21_X1 U10775 ( .B1(n9405), .B2(n9404), .A(n9403), .ZN(n9406) );
  OAI21_X1 U10776 ( .B1(n9407), .B2(n9406), .A(n10000), .ZN(n9411) );
  AND2_X1 U10777 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9601) );
  OAI22_X1 U10778 ( .A1(n9486), .A2(n9488), .B1(n9487), .B2(n9837), .ZN(n9408)
         );
  AOI211_X1 U10779 ( .C1(n9472), .C2(n9409), .A(n9601), .B(n9408), .ZN(n9410)
         );
  OAI211_X1 U10780 ( .C1(n9412), .C2(n9998), .A(n9411), .B(n9410), .ZN(
        P1_U3228) );
  AND2_X1 U10781 ( .A1(n9414), .A2(n9413), .ZN(n9419) );
  NAND3_X1 U10782 ( .A1(n9417), .A2(n9416), .A3(n9415), .ZN(n9418) );
  AOI21_X1 U10783 ( .B1(n9419), .B2(n9418), .A(n9494), .ZN(n9423) );
  AOI22_X1 U10784 ( .A1(n9472), .A2(n9767), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9421) );
  AOI22_X1 U10785 ( .A1(n9474), .A2(n9796), .B1(n9473), .B2(n9661), .ZN(n9420)
         );
  OAI211_X1 U10786 ( .C1(n9770), .C2(n9998), .A(n9421), .B(n9420), .ZN(n9422)
         );
  OR2_X1 U10787 ( .A1(n9423), .A2(n9422), .ZN(P1_U3229) );
  AND2_X1 U10788 ( .A1(n9986), .A2(n9424), .ZN(n9427) );
  OAI211_X1 U10789 ( .C1(n9427), .C2(n9426), .A(n10000), .B(n9425), .ZN(n9434)
         );
  AOI21_X1 U10790 ( .B1(n9472), .B2(n9429), .A(n9428), .ZN(n9433) );
  AOI22_X1 U10791 ( .A1(n9474), .A2(n9508), .B1(n9473), .B2(n9506), .ZN(n9432)
         );
  NAND2_X1 U10792 ( .A1(n9492), .A2(n9430), .ZN(n9431) );
  NAND4_X1 U10793 ( .A1(n9434), .A2(n9433), .A3(n9432), .A4(n9431), .ZN(
        P1_U3231) );
  XNOR2_X1 U10794 ( .A(n9437), .B(n9436), .ZN(n9438) );
  XNOR2_X1 U10795 ( .A(n9435), .B(n9438), .ZN(n9444) );
  AOI22_X1 U10796 ( .A1(n9795), .A2(n9834), .B1(n9794), .B2(n9648), .ZN(n9820)
         );
  NOR2_X1 U10797 ( .A1(n9820), .A2(n9439), .ZN(n9442) );
  OAI22_X1 U10798 ( .A1(n10003), .A2(n9822), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9440), .ZN(n9441) );
  AOI211_X1 U10799 ( .C1(n9824), .C2(n9492), .A(n9442), .B(n9441), .ZN(n9443)
         );
  OAI21_X1 U10800 ( .B1(n9444), .B2(n9494), .A(n9443), .ZN(P1_U3233) );
  XNOR2_X1 U10801 ( .A(n9446), .B(n9445), .ZN(n9447) );
  XNOR2_X1 U10802 ( .A(n9448), .B(n9447), .ZN(n9454) );
  INV_X1 U10803 ( .A(n9788), .ZN(n9450) );
  OAI22_X1 U10804 ( .A1(n10003), .A2(n9450), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9449), .ZN(n9452) );
  OAI22_X1 U10805 ( .A1(n9653), .A2(n9488), .B1(n9487), .B2(n9762), .ZN(n9451)
         );
  AOI211_X1 U10806 ( .C1(n9900), .C2(n9492), .A(n9452), .B(n9451), .ZN(n9453)
         );
  OAI21_X1 U10807 ( .B1(n9454), .B2(n9494), .A(n9453), .ZN(P1_U3235) );
  NAND2_X1 U10808 ( .A1(n9456), .A2(n9455), .ZN(n9457) );
  XOR2_X1 U10809 ( .A(n9458), .B(n9457), .Z(n9466) );
  INV_X1 U10810 ( .A(n9459), .ZN(n9461) );
  INV_X1 U10811 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9460) );
  OAI22_X1 U10812 ( .A1(n10003), .A2(n9461), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9460), .ZN(n9464) );
  OAI22_X1 U10813 ( .A1(n9462), .A2(n9488), .B1(n9487), .B2(n9649), .ZN(n9463)
         );
  AOI211_X1 U10814 ( .C1(n9645), .C2(n9492), .A(n9464), .B(n9463), .ZN(n9465)
         );
  OAI21_X1 U10815 ( .B1(n9466), .B2(n9494), .A(n9465), .ZN(P1_U3238) );
  AND2_X1 U10816 ( .A1(n9468), .A2(n9467), .ZN(n9471) );
  OAI211_X1 U10817 ( .C1(n9471), .C2(n9470), .A(n10000), .B(n9469), .ZN(n9478)
         );
  AOI22_X1 U10818 ( .A1(n9472), .A2(n9736), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9477) );
  INV_X1 U10819 ( .A(n9732), .ZN(n9497) );
  AOI22_X1 U10820 ( .A1(n9474), .A2(n9661), .B1(n9473), .B2(n9497), .ZN(n9476)
         );
  NAND2_X1 U10821 ( .A1(n9879), .A2(n9492), .ZN(n9475) );
  NAND4_X1 U10822 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), .ZN(
        P1_U3240) );
  INV_X1 U10823 ( .A(n9479), .ZN(n9483) );
  XNOR2_X1 U10824 ( .A(n9481), .B(n9480), .ZN(n9482) );
  XNOR2_X1 U10825 ( .A(n9483), .B(n9482), .ZN(n9495) );
  INV_X1 U10826 ( .A(n9484), .ZN(n9485) );
  OAI22_X1 U10827 ( .A1(n10003), .A2(n9485), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9561), .ZN(n9491) );
  OAI22_X1 U10828 ( .A1(n9489), .A2(n9488), .B1(n9487), .B2(n9486), .ZN(n9490)
         );
  AOI211_X1 U10829 ( .C1(n9916), .C2(n9492), .A(n9491), .B(n9490), .ZN(n9493)
         );
  OAI21_X1 U10830 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(P1_U3241) );
  MUX2_X1 U10831 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n4957), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10832 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9496), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10833 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9668), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10834 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9497), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10835 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9498), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10836 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9661), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10837 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9658), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10838 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9796), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10839 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9654), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10840 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9795), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10841 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9835), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10842 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9648), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10843 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9646), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10844 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9499), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10845 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9500), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10846 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9501), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10847 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9502), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10848 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9503), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10849 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8289), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10850 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9505), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10851 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9506), .S(P1_U3973), .Z(
        P1_U3564) );
  INV_X1 U10852 ( .A(n9990), .ZN(n9507) );
  MUX2_X1 U10853 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9507), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10854 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9508), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10855 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9509), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10856 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n6034), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10857 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9510), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10858 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9511), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10859 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9512), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10860 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9513), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10861 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5981), .S(P1_U3973), .Z(
        P1_U3555) );
  NOR2_X1 U10862 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9514), .ZN(n9517) );
  NOR2_X1 U10863 ( .A1(n9629), .A2(n9515), .ZN(n9516) );
  AOI211_X1 U10864 ( .C1(n10049), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9517), .B(
        n9516), .ZN(n9527) );
  AOI211_X1 U10865 ( .C1(n9520), .C2(n9519), .A(n9518), .B(n10022), .ZN(n9521)
         );
  INV_X1 U10866 ( .A(n9521), .ZN(n9526) );
  OAI211_X1 U10867 ( .C1(n9524), .C2(n9523), .A(n10053), .B(n9522), .ZN(n9525)
         );
  NAND3_X1 U10868 ( .A1(n9527), .A2(n9526), .A3(n9525), .ZN(P1_U3246) );
  OAI211_X1 U10869 ( .C1(n9530), .C2(n9529), .A(n10043), .B(n9528), .ZN(n9539)
         );
  OAI211_X1 U10870 ( .C1(n9533), .C2(n9532), .A(n10053), .B(n9531), .ZN(n9538)
         );
  AND2_X1 U10871 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9534) );
  AOI21_X1 U10872 ( .B1(n10049), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9534), .ZN(
        n9537) );
  NAND2_X1 U10873 ( .A1(n10051), .A2(n9535), .ZN(n9536) );
  NAND4_X1 U10874 ( .A1(n9539), .A2(n9538), .A3(n9537), .A4(n9536), .ZN(
        P1_U3248) );
  AOI211_X1 U10875 ( .C1(n9542), .C2(n9541), .A(n9540), .B(n10022), .ZN(n9543)
         );
  INV_X1 U10876 ( .A(n9543), .ZN(n9551) );
  AND2_X1 U10877 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9995) );
  AOI21_X1 U10878 ( .B1(n10049), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9995), .ZN(
        n9550) );
  NAND2_X1 U10879 ( .A1(n10051), .A2(n9544), .ZN(n9549) );
  OAI211_X1 U10880 ( .C1(n9547), .C2(n9546), .A(n10053), .B(n9545), .ZN(n9548)
         );
  NAND4_X1 U10881 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(
        P1_U3251) );
  NOR2_X1 U10882 ( .A1(n8328), .A2(n9554), .ZN(n9576) );
  AOI211_X1 U10883 ( .C1(n9554), .C2(n8328), .A(n9576), .B(n10022), .ZN(n9566)
         );
  INV_X1 U10884 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9559) );
  OR2_X1 U10885 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  OAI21_X1 U10886 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9567) );
  XNOR2_X1 U10887 ( .A(n9574), .B(n9567), .ZN(n9560) );
  NAND2_X1 U10888 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9560), .ZN(n9569) );
  OAI211_X1 U10889 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9560), .A(n10053), .B(
        n9569), .ZN(n9564) );
  NOR2_X1 U10890 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9561), .ZN(n9562) );
  AOI21_X1 U10891 ( .B1(n10049), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9562), .ZN(
        n9563) );
  OAI211_X1 U10892 ( .C1(n9629), .C2(n9574), .A(n9564), .B(n9563), .ZN(n9565)
         );
  OR2_X1 U10893 ( .A1(n9566), .A2(n9565), .ZN(P1_U3258) );
  NAND2_X1 U10894 ( .A1(n9568), .A2(n9567), .ZN(n9570) );
  NAND2_X1 U10895 ( .A1(n9570), .A2(n9569), .ZN(n9573) );
  INV_X1 U10896 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9976) );
  NOR2_X1 U10897 ( .A1(n9589), .A2(n9976), .ZN(n9571) );
  AOI21_X1 U10898 ( .B1(n9589), .B2(n9976), .A(n9571), .ZN(n9572) );
  NOR2_X1 U10899 ( .A1(n9572), .A2(n9573), .ZN(n9594) );
  AOI21_X1 U10900 ( .B1(n9573), .B2(n9572), .A(n9594), .ZN(n9586) );
  NOR2_X1 U10901 ( .A1(n9575), .A2(n9574), .ZN(n9577) );
  NAND2_X1 U10902 ( .A1(n9589), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9578) );
  OAI21_X1 U10903 ( .B1(n9589), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9578), .ZN(
        n9579) );
  NOR2_X1 U10904 ( .A1(n9580), .A2(n9579), .ZN(n9588) );
  AOI211_X1 U10905 ( .C1(n9580), .C2(n9579), .A(n9588), .B(n10022), .ZN(n9581)
         );
  INV_X1 U10906 ( .A(n9581), .ZN(n9585) );
  AND2_X1 U10907 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9583) );
  NOR2_X1 U10908 ( .A1(n9629), .A2(n9595), .ZN(n9582) );
  AOI211_X1 U10909 ( .C1(n10049), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9583), .B(
        n9582), .ZN(n9584) );
  OAI211_X1 U10910 ( .C1(n9586), .C2(n9631), .A(n9585), .B(n9584), .ZN(
        P1_U3259) );
  INV_X1 U10911 ( .A(n9605), .ZN(n9604) );
  OR2_X1 U10912 ( .A1(n9605), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U10913 ( .A1(n9605), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9587) );
  AOI21_X1 U10914 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9589), .A(n9588), .ZN(
        n9590) );
  OAI21_X1 U10915 ( .B1(n4611), .B2(n9590), .A(n9612), .ZN(n9600) );
  INV_X1 U10916 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9591) );
  OR2_X1 U10917 ( .A1(n9605), .A2(n9591), .ZN(n9593) );
  NAND2_X1 U10918 ( .A1(n9605), .A2(n9591), .ZN(n9592) );
  NAND2_X1 U10919 ( .A1(n9593), .A2(n9592), .ZN(n9598) );
  AOI21_X1 U10920 ( .B1(n9595), .B2(n9976), .A(n9594), .ZN(n9596) );
  INV_X1 U10921 ( .A(n9596), .ZN(n9597) );
  NAND2_X1 U10922 ( .A1(n9598), .A2(n9597), .ZN(n9607) );
  OAI21_X1 U10923 ( .B1(n9598), .B2(n9597), .A(n9607), .ZN(n9599) );
  AOI22_X1 U10924 ( .A1(n10043), .A2(n9600), .B1(n10053), .B2(n9599), .ZN(
        n9603) );
  AOI21_X1 U10925 ( .B1(n10049), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9601), .ZN(
        n9602) );
  OAI211_X1 U10926 ( .C1(n9604), .C2(n9629), .A(n9603), .B(n9602), .ZN(
        P1_U3260) );
  OR2_X1 U10927 ( .A1(n9605), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9606) );
  AND2_X1 U10928 ( .A1(n9607), .A2(n9606), .ZN(n9610) );
  NAND2_X1 U10929 ( .A1(n9622), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9626) );
  OAI21_X1 U10930 ( .B1(n9622), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9626), .ZN(
        n9608) );
  INV_X1 U10931 ( .A(n9608), .ZN(n9609) );
  NAND2_X1 U10932 ( .A1(n9610), .A2(n9609), .ZN(n9627) );
  OAI211_X1 U10933 ( .C1(n9610), .C2(n9609), .A(n10053), .B(n9627), .ZN(n9621)
         );
  INV_X1 U10934 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U10935 ( .A1(n9622), .A2(n9614), .ZN(n9613) );
  OAI21_X1 U10936 ( .B1(n9622), .B2(n9614), .A(n9613), .ZN(n9615) );
  OAI211_X1 U10937 ( .C1(n9616), .C2(n9615), .A(n10043), .B(n9624), .ZN(n9620)
         );
  AND2_X1 U10938 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9617) );
  AOI21_X1 U10939 ( .B1(n10049), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9617), .ZN(
        n9619) );
  NAND2_X1 U10940 ( .A1(n10051), .A2(n9622), .ZN(n9618) );
  NAND4_X1 U10941 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(
        P1_U3261) );
  NAND2_X1 U10942 ( .A1(n9622), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U10943 ( .A1(n9624), .A2(n9623), .ZN(n9625) );
  INV_X1 U10944 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U10945 ( .A1(n9627), .A2(n9626), .ZN(n9628) );
  XNOR2_X1 U10946 ( .A(n9628), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U10947 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9632) );
  OAI211_X1 U10948 ( .C1(n9635), .C2(n9634), .A(n9633), .B(n9632), .ZN(
        P1_U3262) );
  NOR2_X1 U10949 ( .A1(n9855), .A2(n10121), .ZN(n9642) );
  NOR2_X1 U10950 ( .A1(n9636), .A2(n9815), .ZN(n9637) );
  AOI211_X1 U10951 ( .C1(n10121), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9642), .B(
        n9637), .ZN(n9638) );
  OAI21_X1 U10952 ( .B1(n9639), .B2(n9847), .A(n9638), .ZN(P1_U3263) );
  OAI211_X1 U10953 ( .C1(n4743), .C2(n9691), .A(n10099), .B(n9640), .ZN(n9856)
         );
  NOR2_X1 U10954 ( .A1(n4743), .A2(n9815), .ZN(n9641) );
  AOI211_X1 U10955 ( .C1(n10121), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9642), .B(
        n9641), .ZN(n9643) );
  OAI21_X1 U10956 ( .B1(n9847), .B2(n9856), .A(n9643), .ZN(P1_U3264) );
  AOI21_X1 U10957 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9647) );
  OAI21_X1 U10958 ( .B1(n9648), .B2(n9850), .A(n9841), .ZN(n9650) );
  NAND2_X1 U10959 ( .A1(n9650), .A2(n5095), .ZN(n9818) );
  NAND2_X1 U10960 ( .A1(n9651), .A2(n9653), .ZN(n9652) );
  NAND2_X1 U10961 ( .A1(n9790), .A2(n9808), .ZN(n9656) );
  NAND2_X1 U10962 ( .A1(n9774), .A2(n9796), .ZN(n9657) );
  NAND2_X1 U10963 ( .A1(n9770), .A2(n9747), .ZN(n9660) );
  AOI21_X1 U10964 ( .B1(n9756), .B2(n9660), .A(n9659), .ZN(n9742) );
  NAND2_X1 U10965 ( .A1(n9884), .A2(n9661), .ZN(n9663) );
  NOR2_X1 U10966 ( .A1(n9884), .A2(n9661), .ZN(n9662) );
  NAND2_X1 U10967 ( .A1(n9739), .A2(n9748), .ZN(n9665) );
  NOR2_X1 U10968 ( .A1(n9739), .A2(n9748), .ZN(n9664) );
  INV_X1 U10969 ( .A(n9699), .ZN(n9667) );
  INV_X1 U10970 ( .A(n9702), .ZN(n9666) );
  NAND2_X1 U10971 ( .A1(n9667), .A2(n9666), .ZN(n9701) );
  NAND2_X1 U10972 ( .A1(n9870), .A2(n9668), .ZN(n9669) );
  NAND2_X1 U10973 ( .A1(n9701), .A2(n9669), .ZN(n9671) );
  XNOR2_X1 U10974 ( .A(n9671), .B(n9670), .ZN(n9860) );
  INV_X1 U10975 ( .A(n9860), .ZN(n9698) );
  INV_X1 U10976 ( .A(n9680), .ZN(n9681) );
  AOI21_X1 U10977 ( .B1(n9703), .B2(n9683), .A(n9682), .ZN(n9685) );
  XNOR2_X1 U10978 ( .A(n9685), .B(n9684), .ZN(n9690) );
  INV_X1 U10979 ( .A(n9688), .ZN(n9689) );
  OAI21_X1 U10980 ( .B1(n9690), .B2(n10129), .A(n9689), .ZN(n9864) );
  INV_X1 U10981 ( .A(n9861), .ZN(n9695) );
  AOI211_X1 U10982 ( .C1(n9861), .C2(n9706), .A(n9810), .B(n9691), .ZN(n9863)
         );
  NAND2_X1 U10983 ( .A1(n9863), .A2(n10103), .ZN(n9694) );
  AOI22_X1 U10984 ( .A1(n10121), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9692), 
        .B2(n10096), .ZN(n9693) );
  OAI211_X1 U10985 ( .C1(n9695), .C2(n9815), .A(n9694), .B(n9693), .ZN(n9696)
         );
  AOI21_X1 U10986 ( .B1(n9864), .B2(n10118), .A(n9696), .ZN(n9697) );
  OAI21_X1 U10987 ( .B1(n9698), .B2(n9829), .A(n9697), .ZN(P1_U3356) );
  NAND2_X1 U10988 ( .A1(n9699), .A2(n9702), .ZN(n9700) );
  INV_X1 U10989 ( .A(n9867), .ZN(n9715) );
  AOI22_X1 U10990 ( .A1(n9870), .A2(n10094), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10121), .ZN(n9714) );
  XNOR2_X1 U10991 ( .A(n9703), .B(n9702), .ZN(n9705) );
  INV_X1 U10992 ( .A(n9722), .ZN(n9708) );
  INV_X1 U10993 ( .A(n9706), .ZN(n9707) );
  AOI211_X1 U10994 ( .C1(n9870), .C2(n9708), .A(n9810), .B(n9707), .ZN(n9869)
         );
  INV_X1 U10995 ( .A(n9869), .ZN(n9711) );
  INV_X1 U10996 ( .A(n9709), .ZN(n9710) );
  OAI22_X1 U10997 ( .A1(n9711), .A2(n6504), .B1(n9710), .B2(n10108), .ZN(n9712) );
  OAI21_X1 U10998 ( .B1(n9868), .B2(n9712), .A(n10118), .ZN(n9713) );
  OAI211_X1 U10999 ( .C1(n9715), .C2(n9829), .A(n9714), .B(n9713), .ZN(
        P1_U3265) );
  XOR2_X1 U11000 ( .A(n9718), .B(n9716), .Z(n9876) );
  AOI21_X1 U11001 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9720) );
  OAI222_X1 U11002 ( .A1(n9989), .A2(n9721), .B1(n9991), .B2(n9748), .C1(
        n10129), .C2(n9720), .ZN(n9872) );
  AOI211_X1 U11003 ( .C1(n9874), .C2(n9733), .A(n9810), .B(n9722), .ZN(n9873)
         );
  NAND2_X1 U11004 ( .A1(n9873), .A2(n10103), .ZN(n9725) );
  AOI22_X1 U11005 ( .A1(n10121), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9723), 
        .B2(n10096), .ZN(n9724) );
  OAI211_X1 U11006 ( .C1(n4866), .C2(n9815), .A(n9725), .B(n9724), .ZN(n9726)
         );
  AOI21_X1 U11007 ( .B1(n9872), .B2(n10118), .A(n9726), .ZN(n9727) );
  OAI21_X1 U11008 ( .B1(n9876), .B2(n9829), .A(n9727), .ZN(P1_U3266) );
  XNOR2_X1 U11009 ( .A(n9728), .B(n9729), .ZN(n9881) );
  AOI21_X1 U11010 ( .B1(n9730), .B2(n9729), .A(n4566), .ZN(n9731) );
  OAI222_X1 U11011 ( .A1(n9989), .A2(n9732), .B1(n9991), .B2(n9763), .C1(
        n10129), .C2(n9731), .ZN(n9877) );
  INV_X1 U11012 ( .A(n9749), .ZN(n9735) );
  INV_X1 U11013 ( .A(n9733), .ZN(n9734) );
  AOI211_X1 U11014 ( .C1(n9879), .C2(n9735), .A(n9810), .B(n9734), .ZN(n9878)
         );
  NAND2_X1 U11015 ( .A1(n9878), .A2(n10103), .ZN(n9738) );
  AOI22_X1 U11016 ( .A1(n10121), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9736), 
        .B2(n10096), .ZN(n9737) );
  OAI211_X1 U11017 ( .C1(n9739), .C2(n9815), .A(n9738), .B(n9737), .ZN(n9740)
         );
  AOI21_X1 U11018 ( .B1(n9877), .B2(n10118), .A(n9740), .ZN(n9741) );
  OAI21_X1 U11019 ( .B1(n9881), .B2(n9829), .A(n9741), .ZN(P1_U3267) );
  XOR2_X1 U11020 ( .A(n9745), .B(n9742), .Z(n9886) );
  AOI21_X1 U11021 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9746) );
  OAI222_X1 U11022 ( .A1(n9989), .A2(n9748), .B1(n9991), .B2(n9747), .C1(
        n10129), .C2(n9746), .ZN(n9882) );
  INV_X1 U11023 ( .A(n9884), .ZN(n9753) );
  AOI211_X1 U11024 ( .C1(n9884), .C2(n9764), .A(n9810), .B(n9749), .ZN(n9883)
         );
  NAND2_X1 U11025 ( .A1(n9883), .A2(n10103), .ZN(n9752) );
  AOI22_X1 U11026 ( .A1(n10121), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9750), 
        .B2(n10096), .ZN(n9751) );
  OAI211_X1 U11027 ( .C1(n9753), .C2(n9815), .A(n9752), .B(n9751), .ZN(n9754)
         );
  AOI21_X1 U11028 ( .B1(n9882), .B2(n10118), .A(n9754), .ZN(n9755) );
  OAI21_X1 U11029 ( .B1(n9886), .B2(n9829), .A(n9755), .ZN(P1_U3268) );
  XOR2_X1 U11030 ( .A(n9756), .B(n9760), .Z(n9891) );
  NAND2_X1 U11031 ( .A1(n9757), .A2(n9758), .ZN(n9759) );
  XOR2_X1 U11032 ( .A(n9760), .B(n9759), .Z(n9761) );
  OAI222_X1 U11033 ( .A1(n9989), .A2(n9763), .B1(n9991), .B2(n9762), .C1(n9761), .C2(n10129), .ZN(n9887) );
  INV_X1 U11034 ( .A(n9778), .ZN(n9766) );
  INV_X1 U11035 ( .A(n9764), .ZN(n9765) );
  AOI211_X1 U11036 ( .C1(n9889), .C2(n9766), .A(n9810), .B(n9765), .ZN(n9888)
         );
  NAND2_X1 U11037 ( .A1(n9888), .A2(n10103), .ZN(n9769) );
  AOI22_X1 U11038 ( .A1(n10121), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9767), 
        .B2(n10096), .ZN(n9768) );
  OAI211_X1 U11039 ( .C1(n9770), .C2(n9815), .A(n9769), .B(n9768), .ZN(n9771)
         );
  AOI21_X1 U11040 ( .B1(n9887), .B2(n10118), .A(n9771), .ZN(n9772) );
  OAI21_X1 U11041 ( .B1(n9891), .B2(n9829), .A(n9772), .ZN(P1_U3269) );
  XOR2_X1 U11042 ( .A(n9773), .B(n9775), .Z(n9897) );
  INV_X1 U11043 ( .A(n9897), .ZN(n9785) );
  AOI22_X1 U11044 ( .A1(n9774), .A2(n10094), .B1(n10121), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9784) );
  OR2_X1 U11045 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  AOI21_X1 U11046 ( .B1(n9757), .B2(n9777), .A(n10129), .ZN(n9896) );
  OAI21_X1 U11047 ( .B1(n9787), .B2(n9894), .A(n10099), .ZN(n9779) );
  OR2_X1 U11048 ( .A1(n9779), .A2(n9778), .ZN(n9893) );
  NAND2_X1 U11049 ( .A1(n10096), .A2(n9780), .ZN(n9781) );
  OAI211_X1 U11050 ( .C1(n9893), .C2(n6504), .A(n9892), .B(n9781), .ZN(n9782)
         );
  OAI21_X1 U11051 ( .B1(n9896), .B2(n9782), .A(n10118), .ZN(n9783) );
  OAI211_X1 U11052 ( .C1(n9785), .C2(n9829), .A(n9784), .B(n9783), .ZN(
        P1_U3270) );
  XOR2_X1 U11053 ( .A(n9786), .B(n9792), .Z(n9903) );
  AOI211_X1 U11054 ( .C1(n9900), .C2(n9809), .A(n9810), .B(n9787), .ZN(n9899)
         );
  AOI22_X1 U11055 ( .A1(n10121), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9788), 
        .B2(n10096), .ZN(n9789) );
  OAI21_X1 U11056 ( .B1(n9790), .B2(n9815), .A(n9789), .ZN(n9799) );
  OAI21_X1 U11057 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9797) );
  AOI222_X1 U11058 ( .A1(n10092), .A2(n9797), .B1(n9796), .B2(n9834), .C1(
        n9795), .C2(n9794), .ZN(n9902) );
  NOR2_X1 U11059 ( .A1(n9902), .A2(n10121), .ZN(n9798) );
  AOI211_X1 U11060 ( .C1(n9899), .C2(n10103), .A(n9799), .B(n9798), .ZN(n9800)
         );
  OAI21_X1 U11061 ( .B1(n9903), .B2(n9829), .A(n9800), .ZN(P1_U3271) );
  XNOR2_X1 U11062 ( .A(n9801), .B(n9805), .ZN(n9908) );
  INV_X1 U11063 ( .A(n9802), .ZN(n9803) );
  AOI21_X1 U11064 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9806) );
  OAI222_X1 U11065 ( .A1(n9989), .A2(n9808), .B1(n9991), .B2(n9807), .C1(
        n10129), .C2(n9806), .ZN(n9904) );
  AOI211_X1 U11066 ( .C1(n9906), .C2(n4540), .A(n9810), .B(n4857), .ZN(n9905)
         );
  NAND2_X1 U11067 ( .A1(n9905), .A2(n10103), .ZN(n9814) );
  INV_X1 U11068 ( .A(n9811), .ZN(n9812) );
  AOI22_X1 U11069 ( .A1(n10121), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9812), 
        .B2(n10096), .ZN(n9813) );
  OAI211_X1 U11070 ( .C1(n9651), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9816)
         );
  AOI21_X1 U11071 ( .B1(n9904), .B2(n10118), .A(n9816), .ZN(n9817) );
  OAI21_X1 U11072 ( .B1(n9908), .B2(n9829), .A(n9817), .ZN(P1_U3272) );
  XOR2_X1 U11073 ( .A(n9818), .B(n9819), .Z(n9958) );
  INV_X1 U11074 ( .A(n9958), .ZN(n9830) );
  XNOR2_X1 U11075 ( .A(n9672), .B(n9819), .ZN(n9821) );
  OAI21_X1 U11076 ( .B1(n9821), .B2(n10129), .A(n9820), .ZN(n9957) );
  OAI211_X1 U11077 ( .C1(n9844), .C2(n9955), .A(n10099), .B(n4540), .ZN(n9954)
         );
  INV_X1 U11078 ( .A(n9822), .ZN(n9823) );
  AOI22_X1 U11079 ( .A1(n10121), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9823), 
        .B2(n10096), .ZN(n9826) );
  NAND2_X1 U11080 ( .A1(n9824), .A2(n10094), .ZN(n9825) );
  OAI211_X1 U11081 ( .C1(n9954), .C2(n9847), .A(n9826), .B(n9825), .ZN(n9827)
         );
  AOI21_X1 U11082 ( .B1(n9957), .B2(n10118), .A(n9827), .ZN(n9828) );
  OAI21_X1 U11083 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(P1_U3273) );
  NAND2_X1 U11084 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  XNOR2_X1 U11085 ( .A(n9833), .B(n9840), .ZN(n9839) );
  NAND2_X1 U11086 ( .A1(n9835), .A2(n9834), .ZN(n9836) );
  OAI21_X1 U11087 ( .B1(n9837), .B2(n9991), .A(n9836), .ZN(n9838) );
  AOI21_X1 U11088 ( .B1(n9839), .B2(n10092), .A(n9838), .ZN(n9960) );
  XOR2_X1 U11089 ( .A(n9841), .B(n9840), .Z(n9963) );
  NAND2_X1 U11090 ( .A1(n9963), .A2(n10104), .ZN(n9852) );
  OAI22_X1 U11091 ( .A1(n10118), .A2(n9843), .B1(n9842), .B2(n10108), .ZN(
        n9849) );
  INV_X1 U11092 ( .A(n9844), .ZN(n9845) );
  OAI211_X1 U11093 ( .C1(n9961), .C2(n9846), .A(n9845), .B(n10099), .ZN(n9959)
         );
  NOR2_X1 U11094 ( .A1(n9959), .A2(n9847), .ZN(n9848) );
  AOI211_X1 U11095 ( .C1(n10094), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9851)
         );
  OAI211_X1 U11096 ( .C1(n10121), .C2(n9960), .A(n9852), .B(n9851), .ZN(
        P1_U3274) );
  AND2_X2 U11097 ( .A1(n9853), .A2(n9940), .ZN(n10247) );
  MUX2_X1 U11098 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9854), .S(n10247), .Z(
        P1_U3553) );
  OAI211_X1 U11099 ( .C1(n4743), .C2(n10219), .A(n9856), .B(n9855), .ZN(n9924)
         );
  MUX2_X1 U11100 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9924), .S(n10247), .Z(
        P1_U3552) );
  OR2_X1 U11101 ( .A1(n9858), .A2(n9857), .ZN(n10134) );
  NAND2_X1 U11102 ( .A1(n9860), .A2(n10222), .ZN(n9866) );
  NAND2_X1 U11103 ( .A1(n9866), .A2(n9865), .ZN(n9925) );
  MUX2_X1 U11104 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9925), .S(n10247), .Z(
        P1_U3551) );
  NAND2_X1 U11105 ( .A1(n9867), .A2(n10222), .ZN(n9871) );
  INV_X1 U11106 ( .A(n10222), .ZN(n10162) );
  AOI211_X1 U11107 ( .C1(n10158), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9875)
         );
  OAI21_X1 U11108 ( .B1(n9876), .B2(n10162), .A(n9875), .ZN(n9927) );
  MUX2_X1 U11109 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9927), .S(n10247), .Z(
        P1_U3549) );
  AOI211_X1 U11110 ( .C1(n10158), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9880)
         );
  OAI21_X1 U11111 ( .B1(n9881), .B2(n10162), .A(n9880), .ZN(n9928) );
  MUX2_X1 U11112 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9928), .S(n10247), .Z(
        P1_U3548) );
  AOI211_X1 U11113 ( .C1(n10158), .C2(n9884), .A(n9883), .B(n9882), .ZN(n9885)
         );
  OAI21_X1 U11114 ( .B1(n9886), .B2(n10162), .A(n9885), .ZN(n9929) );
  MUX2_X1 U11115 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9929), .S(n10247), .Z(
        P1_U3547) );
  AOI211_X1 U11116 ( .C1(n10158), .C2(n9889), .A(n9888), .B(n9887), .ZN(n9890)
         );
  OAI21_X1 U11117 ( .B1(n9891), .B2(n10162), .A(n9890), .ZN(n9930) );
  MUX2_X1 U11118 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9930), .S(n10247), .Z(
        P1_U3546) );
  OAI211_X1 U11119 ( .C1(n9894), .C2(n10219), .A(n9893), .B(n9892), .ZN(n9895)
         );
  AOI211_X1 U11120 ( .C1(n9897), .C2(n10222), .A(n9896), .B(n9895), .ZN(n9898)
         );
  INV_X1 U11121 ( .A(n9898), .ZN(n9931) );
  MUX2_X1 U11122 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9931), .S(n10247), .Z(
        P1_U3545) );
  AOI21_X1 U11123 ( .B1(n10158), .B2(n9900), .A(n9899), .ZN(n9901) );
  OAI211_X1 U11124 ( .C1(n9903), .C2(n10162), .A(n9902), .B(n9901), .ZN(n9932)
         );
  MUX2_X1 U11125 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9932), .S(n10247), .Z(
        P1_U3544) );
  AOI211_X1 U11126 ( .C1(n10158), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9907)
         );
  OAI21_X1 U11127 ( .B1(n9908), .B2(n10162), .A(n9907), .ZN(n9933) );
  MUX2_X1 U11128 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9933), .S(n10247), .Z(
        P1_U3543) );
  AOI211_X1 U11129 ( .C1(n10158), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9912)
         );
  OAI21_X1 U11130 ( .B1(n9913), .B2(n10162), .A(n9912), .ZN(n9934) );
  MUX2_X1 U11131 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9934), .S(n10247), .Z(
        P1_U3539) );
  AOI211_X1 U11132 ( .C1(n10158), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9917)
         );
  OAI21_X1 U11133 ( .B1(n9918), .B2(n10162), .A(n9917), .ZN(n9935) );
  MUX2_X1 U11134 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9935), .S(n10247), .Z(
        P1_U3537) );
  AOI21_X1 U11135 ( .B1(n10158), .B2(n9920), .A(n9919), .ZN(n9921) );
  OAI211_X1 U11136 ( .C1(n9923), .C2(n10134), .A(n9922), .B(n9921), .ZN(n9936)
         );
  MUX2_X1 U11137 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9936), .S(n10247), .Z(
        P1_U3536) );
  MUX2_X1 U11138 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9924), .S(n10226), .Z(
        P1_U3520) );
  MUX2_X1 U11139 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9925), .S(n10226), .Z(
        P1_U3519) );
  MUX2_X1 U11140 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9926), .S(n10226), .Z(
        P1_U3518) );
  MUX2_X1 U11141 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9927), .S(n10226), .Z(
        P1_U3517) );
  MUX2_X1 U11142 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9928), .S(n10226), .Z(
        P1_U3516) );
  MUX2_X1 U11143 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9929), .S(n10226), .Z(
        P1_U3515) );
  MUX2_X1 U11144 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9930), .S(n10226), .Z(
        P1_U3514) );
  MUX2_X1 U11145 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9931), .S(n10226), .Z(
        P1_U3513) );
  MUX2_X1 U11146 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9932), .S(n10226), .Z(
        P1_U3512) );
  MUX2_X1 U11147 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9933), .S(n10226), .Z(
        P1_U3511) );
  MUX2_X1 U11148 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9934), .S(n10226), .Z(
        P1_U3504) );
  MUX2_X1 U11149 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9935), .S(n10226), .Z(
        P1_U3498) );
  MUX2_X1 U11150 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9936), .S(n10226), .Z(
        P1_U3495) );
  NOR2_X1 U11151 ( .A1(n9939), .A2(n9937), .ZN(n10127) );
  MUX2_X1 U11152 ( .A(P1_D_REG_1__SCAN_IN), .B(n9938), .S(n10127), .Z(P1_U3440) );
  MUX2_X1 U11153 ( .A(n9940), .B(P1_D_REG_0__SCAN_IN), .S(n9939), .Z(P1_U3439)
         );
  NOR4_X1 U11154 ( .A1(n5832), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5815), .A4(
        P1_U3086), .ZN(n9941) );
  AOI21_X1 U11155 ( .B1(n9945), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9941), .ZN(
        n9942) );
  OAI21_X1 U11156 ( .B1(n9943), .B2(n9949), .A(n9942), .ZN(P1_U3324) );
  AOI22_X1 U11157 ( .A1(n9944), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9945), .ZN(n9946) );
  OAI21_X1 U11158 ( .B1(n9947), .B2(n9949), .A(n9946), .ZN(P1_U3325) );
  OAI222_X1 U11159 ( .A1(n9952), .A2(n9951), .B1(P1_U3086), .B2(n9950), .C1(
        n9949), .C2(n9948), .ZN(P1_U3326) );
  MUX2_X1 U11160 ( .A(n9953), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U11161 ( .B1(n9955), .B2(n10219), .A(n9954), .ZN(n9956) );
  AOI211_X1 U11162 ( .C1(n9958), .C2(n10222), .A(n9957), .B(n9956), .ZN(n9978)
         );
  AOI22_X1 U11163 ( .A1(n10247), .A2(n9978), .B1(n6184), .B2(n10244), .ZN(
        P1_U3542) );
  OAI211_X1 U11164 ( .C1(n9961), .C2(n10219), .A(n9960), .B(n9959), .ZN(n9962)
         );
  AOI21_X1 U11165 ( .B1(n9963), .B2(n10222), .A(n9962), .ZN(n9980) );
  INV_X1 U11166 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11167 ( .A1(n10247), .A2(n9980), .B1(n9964), .B2(n10244), .ZN(
        P1_U3541) );
  OAI21_X1 U11168 ( .B1(n9966), .B2(n10219), .A(n9965), .ZN(n9967) );
  AOI211_X1 U11169 ( .C1(n9969), .C2(n10222), .A(n9968), .B(n9967), .ZN(n9982)
         );
  INV_X1 U11170 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11171 ( .A1(n10247), .A2(n9982), .B1(n9970), .B2(n10244), .ZN(
        P1_U3540) );
  OAI21_X1 U11172 ( .B1(n9972), .B2(n10219), .A(n9971), .ZN(n9973) );
  AOI211_X1 U11173 ( .C1(n9975), .C2(n10222), .A(n9974), .B(n9973), .ZN(n9984)
         );
  AOI22_X1 U11174 ( .A1(n10247), .A2(n9984), .B1(n9976), .B2(n10244), .ZN(
        P1_U3538) );
  INV_X1 U11175 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11176 ( .A1(n10226), .A2(n9978), .B1(n9977), .B2(n10224), .ZN(
        P1_U3510) );
  INV_X1 U11177 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11178 ( .A1(n10226), .A2(n9980), .B1(n9979), .B2(n10224), .ZN(
        P1_U3509) );
  INV_X1 U11179 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11180 ( .A1(n10226), .A2(n9982), .B1(n9981), .B2(n10224), .ZN(
        P1_U3507) );
  INV_X1 U11181 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U11182 ( .A1(n10226), .A2(n9984), .B1(n9983), .B2(n10224), .ZN(
        P1_U3501) );
  XOR2_X1 U11183 ( .A(n9985), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U11184 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11185 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n10001) );
  OR2_X1 U11186 ( .A1(n9990), .A2(n9989), .ZN(n9994) );
  OR2_X1 U11187 ( .A1(n9992), .A2(n9991), .ZN(n9993) );
  NAND2_X1 U11188 ( .A1(n9994), .A2(n9993), .ZN(n10063) );
  AOI21_X1 U11189 ( .B1(n10063), .B2(n9996), .A(n9995), .ZN(n9997) );
  OAI21_X1 U11190 ( .B1(n10187), .B2(n9998), .A(n9997), .ZN(n9999) );
  AOI21_X1 U11191 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(n10002) );
  OAI21_X1 U11192 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(P1_U3221) );
  INV_X1 U11193 ( .A(n10028), .ZN(n10005) );
  AOI21_X1 U11194 ( .B1(n10005), .B2(n10120), .A(n6452), .ZN(n10034) );
  OAI21_X1 U11195 ( .B1(n10005), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10034), .ZN(
        n10006) );
  XOR2_X1 U11196 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10006), .Z(n10009) );
  AOI22_X1 U11197 ( .A1(n10049), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10007) );
  OAI21_X1 U11198 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(P1_U3243) );
  AOI22_X1 U11199 ( .A1(n10049), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10021) );
  AOI211_X1 U11200 ( .C1(n10012), .C2(n10011), .A(n10010), .B(n10022), .ZN(
        n10013) );
  AOI21_X1 U11201 ( .B1(n10051), .B2(n10014), .A(n10013), .ZN(n10020) );
  NOR2_X1 U11202 ( .A1(n10015), .A2(n10227), .ZN(n10018) );
  OAI211_X1 U11203 ( .C1(n10018), .C2(n10017), .A(n10053), .B(n10016), .ZN(
        n10019) );
  NAND3_X1 U11204 ( .A1(n10021), .A2(n10020), .A3(n10019), .ZN(P1_U3244) );
  AOI22_X1 U11205 ( .A1(n10049), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10040) );
  AOI211_X1 U11206 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10026) );
  AOI21_X1 U11207 ( .B1(n10051), .B2(n10027), .A(n10026), .ZN(n10039) );
  MUX2_X1 U11208 ( .A(n10030), .B(n10029), .S(n10028), .Z(n10032) );
  NAND2_X1 U11209 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  OAI211_X1 U11210 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10034), .A(n10033), .B(
        P1_U3973), .ZN(n10058) );
  OAI211_X1 U11211 ( .C1(n10037), .C2(n10036), .A(n10053), .B(n10035), .ZN(
        n10038) );
  NAND4_X1 U11212 ( .A1(n10040), .A2(n10039), .A3(n10058), .A4(n10038), .ZN(
        P1_U3245) );
  NOR2_X1 U11213 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10041), .ZN(n10048) );
  OAI211_X1 U11214 ( .C1(n10045), .C2(n10044), .A(n10043), .B(n10042), .ZN(
        n10046) );
  INV_X1 U11215 ( .A(n10046), .ZN(n10047) );
  AOI211_X1 U11216 ( .C1(n10049), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10048), .B(
        n10047), .ZN(n10059) );
  NAND2_X1 U11217 ( .A1(n10051), .A2(n10050), .ZN(n10057) );
  OAI211_X1 U11218 ( .C1(n10055), .C2(n10054), .A(n10053), .B(n10052), .ZN(
        n10056) );
  NAND4_X1 U11219 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        P1_U3247) );
  NOR2_X1 U11220 ( .A1(n10060), .A2(n10129), .ZN(n10065) );
  OAI21_X1 U11221 ( .B1(n10062), .B2(n10061), .A(n10071), .ZN(n10064) );
  AOI21_X1 U11222 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(n10186) );
  AOI222_X1 U11223 ( .A1(n10067), .A2(n10094), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n10121), .C1(n10096), .C2(n10066), .ZN(n10078) );
  NAND2_X1 U11224 ( .A1(n8012), .A2(n10068), .ZN(n10070) );
  NAND2_X1 U11225 ( .A1(n10070), .A2(n10069), .ZN(n10072) );
  XNOR2_X1 U11226 ( .A(n10072), .B(n10071), .ZN(n10189) );
  INV_X1 U11227 ( .A(n10073), .ZN(n10075) );
  OAI211_X1 U11228 ( .C1(n10075), .C2(n10187), .A(n10099), .B(n10074), .ZN(
        n10185) );
  INV_X1 U11229 ( .A(n10185), .ZN(n10076) );
  AOI22_X1 U11230 ( .A1(n10189), .A2(n10104), .B1(n10103), .B2(n10076), .ZN(
        n10077) );
  OAI211_X1 U11231 ( .C1(n10121), .C2(n10186), .A(n10078), .B(n10077), .ZN(
        P1_U3285) );
  XOR2_X1 U11232 ( .A(n10084), .B(n10079), .Z(n10081) );
  AOI21_X1 U11233 ( .B1(n10081), .B2(n10092), .A(n10080), .ZN(n10173) );
  AOI222_X1 U11234 ( .A1(n10083), .A2(n10094), .B1(n10082), .B2(n10096), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(n10121), .ZN(n10089) );
  XNOR2_X1 U11235 ( .A(n8012), .B(n10084), .ZN(n10176) );
  OAI211_X1 U11236 ( .C1(n10086), .C2(n10174), .A(n10099), .B(n10085), .ZN(
        n10172) );
  INV_X1 U11237 ( .A(n10172), .ZN(n10087) );
  AOI22_X1 U11238 ( .A1(n10176), .A2(n10104), .B1(n10103), .B2(n10087), .ZN(
        n10088) );
  OAI211_X1 U11239 ( .C1(n10121), .C2(n10173), .A(n10089), .B(n10088), .ZN(
        P1_U3287) );
  XOR2_X1 U11240 ( .A(n10090), .B(n10098), .Z(n10093) );
  AOI21_X1 U11241 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10144) );
  AOI222_X1 U11242 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n10121), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10096), .C1(n10095), .C2(n10094), .ZN(
        n10106) );
  XNOR2_X1 U11243 ( .A(n10098), .B(n10097), .ZN(n10147) );
  OAI211_X1 U11244 ( .C1(n10101), .C2(n10143), .A(n10100), .B(n10099), .ZN(
        n10142) );
  INV_X1 U11245 ( .A(n10142), .ZN(n10102) );
  AOI22_X1 U11246 ( .A1(n10147), .A2(n10104), .B1(n10103), .B2(n10102), .ZN(
        n10105) );
  OAI211_X1 U11247 ( .C1(n10121), .C2(n10144), .A(n10106), .B(n10105), .ZN(
        P1_U3291) );
  INV_X1 U11248 ( .A(n10128), .ZN(n10116) );
  NOR2_X1 U11249 ( .A1(n10111), .A2(n10107), .ZN(n10130) );
  INV_X1 U11250 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10109) );
  OAI22_X1 U11251 ( .A1(n10111), .A2(n10110), .B1(n10109), .B2(n10108), .ZN(
        n10112) );
  AOI211_X1 U11252 ( .C1(n10130), .C2(n4507), .A(n10112), .B(n10131), .ZN(
        n10114) );
  INV_X1 U11253 ( .A(n10114), .ZN(n10115) );
  AOI21_X1 U11254 ( .B1(n10117), .B2(n10116), .A(n10115), .ZN(n10119) );
  AOI22_X1 U11255 ( .A1(n10121), .A2(n10120), .B1(n10119), .B2(n10118), .ZN(
        P1_U3293) );
  AND2_X1 U11256 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10122), .ZN(P1_U3294) );
  AND2_X1 U11257 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10122), .ZN(P1_U3295) );
  AND2_X1 U11258 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10122), .ZN(P1_U3296) );
  AND2_X1 U11259 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10122), .ZN(P1_U3297) );
  AND2_X1 U11260 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10122), .ZN(P1_U3298) );
  AND2_X1 U11261 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10122), .ZN(P1_U3299) );
  AND2_X1 U11262 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10122), .ZN(P1_U3300) );
  AND2_X1 U11263 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10122), .ZN(P1_U3301) );
  AND2_X1 U11264 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10122), .ZN(P1_U3302) );
  AND2_X1 U11265 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10122), .ZN(P1_U3303) );
  AND2_X1 U11266 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10122), .ZN(P1_U3304) );
  AND2_X1 U11267 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10122), .ZN(P1_U3305) );
  AND2_X1 U11268 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10122), .ZN(P1_U3306) );
  AND2_X1 U11269 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10122), .ZN(P1_U3307) );
  AND2_X1 U11270 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10122), .ZN(P1_U3308) );
  AND2_X1 U11271 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10122), .ZN(P1_U3309) );
  AND2_X1 U11272 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10122), .ZN(P1_U3310) );
  AND2_X1 U11273 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10122), .ZN(P1_U3311) );
  AND2_X1 U11274 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10122), .ZN(P1_U3312) );
  AND2_X1 U11275 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10122), .ZN(P1_U3313) );
  AND2_X1 U11276 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10122), .ZN(P1_U3314) );
  AND2_X1 U11277 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10122), .ZN(P1_U3315) );
  AND2_X1 U11278 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10122), .ZN(P1_U3316) );
  AND2_X1 U11279 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10122), .ZN(P1_U3317) );
  AND2_X1 U11280 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10122), .ZN(P1_U3318) );
  AND2_X1 U11281 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10122), .ZN(P1_U3319) );
  NOR2_X1 U11282 ( .A1(n10127), .A2(n10123), .ZN(P1_U3320) );
  NOR2_X1 U11283 ( .A1(n10127), .A2(n10124), .ZN(P1_U3321) );
  NOR2_X1 U11284 ( .A1(n10127), .A2(n10125), .ZN(P1_U3322) );
  NOR2_X1 U11285 ( .A1(n10127), .A2(n10126), .ZN(P1_U3323) );
  AOI21_X1 U11286 ( .B1(n10162), .B2(n10129), .A(n10128), .ZN(n10132) );
  NOR3_X1 U11287 ( .A1(n10132), .A2(n10131), .A3(n10130), .ZN(n10228) );
  INV_X1 U11288 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11289 ( .A1(n10226), .A2(n10228), .B1(n10133), .B2(n10224), .ZN(
        P1_U3453) );
  INV_X1 U11290 ( .A(n10134), .ZN(n10206) );
  INV_X1 U11291 ( .A(n10135), .ZN(n10140) );
  OAI21_X1 U11292 ( .B1(n10137), .B2(n10219), .A(n10136), .ZN(n10139) );
  AOI211_X1 U11293 ( .C1(n10206), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        n10230) );
  INV_X1 U11294 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U11295 ( .A1(n10226), .A2(n10230), .B1(n10141), .B2(n10224), .ZN(
        P1_U3456) );
  OAI21_X1 U11296 ( .B1(n10143), .B2(n10219), .A(n10142), .ZN(n10146) );
  INV_X1 U11297 ( .A(n10144), .ZN(n10145) );
  AOI211_X1 U11298 ( .C1(n10222), .C2(n10147), .A(n10146), .B(n10145), .ZN(
        n10231) );
  INV_X1 U11299 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U11300 ( .A1(n10226), .A2(n10231), .B1(n10148), .B2(n10224), .ZN(
        P1_U3459) );
  OAI21_X1 U11301 ( .B1(n10150), .B2(n10219), .A(n10149), .ZN(n10151) );
  AOI21_X1 U11302 ( .B1(n10152), .B2(n10222), .A(n10151), .ZN(n10153) );
  AND2_X1 U11303 ( .A1(n10154), .A2(n10153), .ZN(n10232) );
  INV_X1 U11304 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11305 ( .A1(n10226), .A2(n10232), .B1(n10155), .B2(n10224), .ZN(
        P1_U3462) );
  AOI21_X1 U11306 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10159) );
  OAI211_X1 U11307 ( .C1(n10162), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        n10163) );
  INV_X1 U11308 ( .A(n10163), .ZN(n10233) );
  INV_X1 U11309 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U11310 ( .A1(n10226), .A2(n10233), .B1(n10164), .B2(n10224), .ZN(
        P1_U3465) );
  OAI21_X1 U11311 ( .B1(n10166), .B2(n10219), .A(n10165), .ZN(n10167) );
  AOI21_X1 U11312 ( .B1(n10168), .B2(n10222), .A(n10167), .ZN(n10169) );
  AND2_X1 U11313 ( .A1(n10170), .A2(n10169), .ZN(n10234) );
  INV_X1 U11314 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U11315 ( .A1(n10226), .A2(n10234), .B1(n10171), .B2(n10224), .ZN(
        P1_U3468) );
  OAI211_X1 U11316 ( .C1(n10174), .C2(n10219), .A(n10173), .B(n10172), .ZN(
        n10175) );
  AOI21_X1 U11317 ( .B1(n10222), .B2(n10176), .A(n10175), .ZN(n10236) );
  INV_X1 U11318 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U11319 ( .A1(n10226), .A2(n10236), .B1(n10177), .B2(n10224), .ZN(
        P1_U3471) );
  OAI21_X1 U11320 ( .B1(n10179), .B2(n10219), .A(n10178), .ZN(n10180) );
  AOI21_X1 U11321 ( .B1(n10181), .B2(n10206), .A(n10180), .ZN(n10182) );
  AND2_X1 U11322 ( .A1(n10183), .A2(n10182), .ZN(n10237) );
  INV_X1 U11323 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U11324 ( .A1(n10226), .A2(n10237), .B1(n10184), .B2(n10224), .ZN(
        P1_U3474) );
  OAI211_X1 U11325 ( .C1(n10187), .C2(n10219), .A(n10186), .B(n10185), .ZN(
        n10188) );
  AOI21_X1 U11326 ( .B1(n10222), .B2(n10189), .A(n10188), .ZN(n10238) );
  INV_X1 U11327 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U11328 ( .A1(n10226), .A2(n10238), .B1(n10190), .B2(n10224), .ZN(
        P1_U3477) );
  OAI211_X1 U11329 ( .C1(n10193), .C2(n10219), .A(n10192), .B(n10191), .ZN(
        n10194) );
  AOI21_X1 U11330 ( .B1(n10222), .B2(n10195), .A(n10194), .ZN(n10239) );
  INV_X1 U11331 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U11332 ( .A1(n10226), .A2(n10239), .B1(n10196), .B2(n10224), .ZN(
        P1_U3480) );
  OAI211_X1 U11333 ( .C1(n10199), .C2(n10219), .A(n10198), .B(n10197), .ZN(
        n10200) );
  AOI21_X1 U11334 ( .B1(n10201), .B2(n10222), .A(n10200), .ZN(n10240) );
  INV_X1 U11335 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U11336 ( .A1(n10226), .A2(n10240), .B1(n10202), .B2(n10224), .ZN(
        P1_U3483) );
  OAI21_X1 U11337 ( .B1(n10204), .B2(n10219), .A(n10203), .ZN(n10205) );
  AOI21_X1 U11338 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10208) );
  AND2_X1 U11339 ( .A1(n10209), .A2(n10208), .ZN(n10241) );
  INV_X1 U11340 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U11341 ( .A1(n10226), .A2(n10241), .B1(n10210), .B2(n10224), .ZN(
        P1_U3486) );
  OAI211_X1 U11342 ( .C1(n10213), .C2(n10219), .A(n10212), .B(n10211), .ZN(
        n10214) );
  AOI21_X1 U11343 ( .B1(n10215), .B2(n10222), .A(n10214), .ZN(n10243) );
  INV_X1 U11344 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11345 ( .A1(n10226), .A2(n10243), .B1(n10216), .B2(n10224), .ZN(
        P1_U3489) );
  OAI211_X1 U11346 ( .C1(n10220), .C2(n10219), .A(n10218), .B(n10217), .ZN(
        n10221) );
  AOI21_X1 U11347 ( .B1(n10223), .B2(n10222), .A(n10221), .ZN(n10246) );
  INV_X1 U11348 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U11349 ( .A1(n10226), .A2(n10246), .B1(n10225), .B2(n10224), .ZN(
        P1_U3492) );
  AOI22_X1 U11350 ( .A1(n10247), .A2(n10228), .B1(n10227), .B2(n10244), .ZN(
        P1_U3522) );
  AOI22_X1 U11351 ( .A1(n10247), .A2(n10230), .B1(n10229), .B2(n10244), .ZN(
        P1_U3523) );
  AOI22_X1 U11352 ( .A1(n10247), .A2(n10231), .B1(n6803), .B2(n10244), .ZN(
        P1_U3524) );
  AOI22_X1 U11353 ( .A1(n10247), .A2(n10232), .B1(n6802), .B2(n10244), .ZN(
        P1_U3525) );
  AOI22_X1 U11354 ( .A1(n10247), .A2(n10233), .B1(n6800), .B2(n10244), .ZN(
        P1_U3526) );
  AOI22_X1 U11355 ( .A1(n10247), .A2(n10234), .B1(n6808), .B2(n10244), .ZN(
        P1_U3527) );
  AOI22_X1 U11356 ( .A1(n10247), .A2(n10236), .B1(n10235), .B2(n10244), .ZN(
        P1_U3528) );
  AOI22_X1 U11357 ( .A1(n10247), .A2(n10237), .B1(n7053), .B2(n10244), .ZN(
        P1_U3529) );
  AOI22_X1 U11358 ( .A1(n10247), .A2(n10238), .B1(n7050), .B2(n10244), .ZN(
        P1_U3530) );
  AOI22_X1 U11359 ( .A1(n10247), .A2(n10239), .B1(n7055), .B2(n10244), .ZN(
        P1_U3531) );
  AOI22_X1 U11360 ( .A1(n10247), .A2(n10240), .B1(n7298), .B2(n10244), .ZN(
        P1_U3532) );
  AOI22_X1 U11361 ( .A1(n10247), .A2(n10241), .B1(n7355), .B2(n10244), .ZN(
        P1_U3533) );
  AOI22_X1 U11362 ( .A1(n10247), .A2(n10243), .B1(n10242), .B2(n10244), .ZN(
        P1_U3534) );
  AOI22_X1 U11363 ( .A1(n10247), .A2(n10246), .B1(n10245), .B2(n10244), .ZN(
        P1_U3535) );
  AOI22_X1 U11364 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n10248), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10254) );
  OAI21_X1 U11365 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10250), .A(n10249), .ZN(
        n10251) );
  OAI21_X1 U11366 ( .B1(n10252), .B2(n10272), .A(n10251), .ZN(n10253) );
  OAI211_X1 U11367 ( .C1(n10312), .C2(n10255), .A(n10254), .B(n10253), .ZN(
        P2_U3182) );
  OR2_X1 U11368 ( .A1(n10312), .A2(n10256), .ZN(n10269) );
  OAI21_X1 U11369 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10260) );
  INV_X1 U11370 ( .A(n10260), .ZN(n10261) );
  OR2_X1 U11371 ( .A1(n10283), .A2(n10261), .ZN(n10268) );
  OAI21_X1 U11372 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(n10265) );
  NAND2_X1 U11373 ( .A1(n10308), .A2(n10265), .ZN(n10267) );
  NAND2_X1 U11374 ( .A1(P2_U3151), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10266) );
  AND4_X1 U11375 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10275) );
  XOR2_X1 U11376 ( .A(n10271), .B(n10270), .Z(n10273) );
  NAND2_X1 U11377 ( .A1(n10273), .A2(n10272), .ZN(n10274) );
  OAI211_X1 U11378 ( .C1(n10276), .C2(n10321), .A(n10275), .B(n10274), .ZN(
        P2_U3184) );
  XNOR2_X1 U11379 ( .A(n10277), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n10279) );
  AOI21_X1 U11380 ( .B1(n10308), .B2(n10279), .A(n10278), .ZN(n10285) );
  AND2_X1 U11381 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  OR2_X1 U11382 ( .A1(n10283), .A2(n10282), .ZN(n10284) );
  OAI211_X1 U11383 ( .C1(n10312), .C2(n10286), .A(n10285), .B(n10284), .ZN(
        n10287) );
  INV_X1 U11384 ( .A(n10287), .ZN(n10293) );
  AOI21_X1 U11385 ( .B1(n10290), .B2(n10289), .A(n10288), .ZN(n10291) );
  OR2_X1 U11386 ( .A1(n10291), .A2(n10317), .ZN(n10292) );
  OAI211_X1 U11387 ( .C1(n10294), .C2(n10321), .A(n10293), .B(n10292), .ZN(
        P2_U3185) );
  INV_X1 U11388 ( .A(n10295), .ZN(n10300) );
  NAND3_X1 U11389 ( .A1(n10298), .A2(n10297), .A3(n10296), .ZN(n10299) );
  NAND2_X1 U11390 ( .A1(n10300), .A2(n10299), .ZN(n10302) );
  AOI21_X1 U11391 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(n10310) );
  OAI21_X1 U11392 ( .B1(n10306), .B2(n10305), .A(n10304), .ZN(n10307) );
  NAND2_X1 U11393 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  OAI211_X1 U11394 ( .C1(n10312), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        n10313) );
  INV_X1 U11395 ( .A(n10313), .ZN(n10320) );
  AOI21_X1 U11396 ( .B1(n10316), .B2(n10315), .A(n10314), .ZN(n10318) );
  OR2_X1 U11397 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  OAI211_X1 U11398 ( .C1(n10322), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        P2_U3188) );
  NAND2_X1 U11399 ( .A1(n10324), .A2(n10323), .ZN(n10325) );
  XOR2_X1 U11400 ( .A(n10332), .B(n10325), .Z(n10330) );
  AOI222_X1 U11401 ( .A1(n10350), .A2(n10330), .B1(n10329), .B2(n10328), .C1(
        n10327), .C2(n10326), .ZN(n10372) );
  INV_X1 U11402 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10338) );
  XNOR2_X1 U11403 ( .A(n10331), .B(n10332), .ZN(n10370) );
  OAI22_X1 U11404 ( .A1(n10334), .A2(n10333), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n10343), .ZN(n10335) );
  AOI21_X1 U11405 ( .B1(n10370), .B2(n10336), .A(n10335), .ZN(n10337) );
  OAI221_X1 U11406 ( .B1(n10339), .B2(n10372), .C1(n10357), .C2(n10338), .A(
        n10337), .ZN(P2_U3230) );
  XNOR2_X1 U11407 ( .A(n10340), .B(n10344), .ZN(n10366) );
  INV_X1 U11408 ( .A(n10366), .ZN(n10355) );
  OAI22_X1 U11409 ( .A1(n10343), .A2(n10342), .B1(n10365), .B2(n10341), .ZN(
        n10354) );
  XNOR2_X1 U11410 ( .A(n10345), .B(n10344), .ZN(n10351) );
  OAI22_X1 U11411 ( .A1(n5692), .A2(n10348), .B1(n10347), .B2(n10346), .ZN(
        n10349) );
  AOI21_X1 U11412 ( .B1(n10351), .B2(n10350), .A(n10349), .ZN(n10352) );
  OAI21_X1 U11413 ( .B1(n10366), .B2(n10353), .A(n10352), .ZN(n10368) );
  AOI211_X1 U11414 ( .C1(n10356), .C2(n10355), .A(n10354), .B(n10368), .ZN(
        n10358) );
  AOI22_X1 U11415 ( .A1(n10339), .A2(n6904), .B1(n10358), .B2(n10357), .ZN(
        P2_U3231) );
  INV_X1 U11416 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10364) );
  INV_X1 U11417 ( .A(n10359), .ZN(n10363) );
  OAI22_X1 U11418 ( .A1(n10361), .A2(n10396), .B1(n10360), .B2(n10390), .ZN(
        n10362) );
  NOR2_X1 U11419 ( .A1(n10363), .A2(n10362), .ZN(n10424) );
  AOI22_X1 U11420 ( .A1(n10423), .A2(n10364), .B1(n10424), .B2(n10421), .ZN(
        P2_U3393) );
  OAI22_X1 U11421 ( .A1(n10366), .A2(n5741), .B1(n10365), .B2(n10390), .ZN(
        n10367) );
  NOR2_X1 U11422 ( .A1(n10368), .A2(n10367), .ZN(n10426) );
  AOI22_X1 U11423 ( .A1(n10423), .A2(n5152), .B1(n10426), .B2(n10421), .ZN(
        P2_U3396) );
  AOI22_X1 U11424 ( .A1(n10370), .A2(n10414), .B1(n10416), .B2(n10369), .ZN(
        n10371) );
  AND2_X1 U11425 ( .A1(n10372), .A2(n10371), .ZN(n10427) );
  AOI22_X1 U11426 ( .A1(n10423), .A2(n5168), .B1(n10427), .B2(n10421), .ZN(
        P2_U3399) );
  INV_X1 U11427 ( .A(n10373), .ZN(n10377) );
  OAI21_X1 U11428 ( .B1(n10375), .B2(n10390), .A(n10374), .ZN(n10376) );
  AOI21_X1 U11429 ( .B1(n10414), .B2(n10377), .A(n10376), .ZN(n10428) );
  AOI22_X1 U11430 ( .A1(n10423), .A2(n5184), .B1(n10428), .B2(n10421), .ZN(
        P2_U3402) );
  INV_X1 U11431 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10383) );
  INV_X1 U11432 ( .A(n10378), .ZN(n10382) );
  NOR2_X1 U11433 ( .A1(n10379), .A2(n10390), .ZN(n10381) );
  AOI211_X1 U11434 ( .C1(n10404), .C2(n10382), .A(n10381), .B(n10380), .ZN(
        n10430) );
  AOI22_X1 U11435 ( .A1(n10423), .A2(n10383), .B1(n10430), .B2(n10421), .ZN(
        P2_U3405) );
  INV_X1 U11436 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10389) );
  INV_X1 U11437 ( .A(n10384), .ZN(n10388) );
  OAI21_X1 U11438 ( .B1(n10386), .B2(n10390), .A(n10385), .ZN(n10387) );
  AOI21_X1 U11439 ( .B1(n10414), .B2(n10388), .A(n10387), .ZN(n10431) );
  AOI22_X1 U11440 ( .A1(n10423), .A2(n10389), .B1(n10431), .B2(n10421), .ZN(
        P2_U3408) );
  INV_X1 U11441 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10395) );
  OAI22_X1 U11442 ( .A1(n10392), .A2(n5741), .B1(n10391), .B2(n10390), .ZN(
        n10393) );
  NOR2_X1 U11443 ( .A1(n10394), .A2(n10393), .ZN(n10432) );
  AOI22_X1 U11444 ( .A1(n10423), .A2(n10395), .B1(n10432), .B2(n10421), .ZN(
        P2_U3411) );
  INV_X1 U11445 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10401) );
  NOR2_X1 U11446 ( .A1(n10397), .A2(n10396), .ZN(n10399) );
  AOI211_X1 U11447 ( .C1(n10416), .C2(n10400), .A(n10399), .B(n10398), .ZN(
        n10433) );
  AOI22_X1 U11448 ( .A1(n10423), .A2(n10401), .B1(n10433), .B2(n10421), .ZN(
        P2_U3414) );
  INV_X1 U11449 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10408) );
  INV_X1 U11450 ( .A(n10402), .ZN(n10405) );
  AOI22_X1 U11451 ( .A1(n10405), .A2(n10404), .B1(n10416), .B2(n10403), .ZN(
        n10406) );
  AND2_X1 U11452 ( .A1(n10407), .A2(n10406), .ZN(n10435) );
  AOI22_X1 U11453 ( .A1(n10423), .A2(n10408), .B1(n10435), .B2(n10421), .ZN(
        P2_U3417) );
  INV_X1 U11454 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10413) );
  NOR2_X1 U11455 ( .A1(n10409), .A2(n5741), .ZN(n10411) );
  AOI211_X1 U11456 ( .C1(n10416), .C2(n10412), .A(n10411), .B(n10410), .ZN(
        n10436) );
  AOI22_X1 U11457 ( .A1(n10423), .A2(n10413), .B1(n10436), .B2(n10421), .ZN(
        P2_U3420) );
  INV_X1 U11458 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10422) );
  AND2_X1 U11459 ( .A1(n10415), .A2(n10414), .ZN(n10419) );
  AND2_X1 U11460 ( .A1(n10417), .A2(n10416), .ZN(n10418) );
  NOR3_X1 U11461 ( .A1(n10420), .A2(n10419), .A3(n10418), .ZN(n10439) );
  AOI22_X1 U11462 ( .A1(n10423), .A2(n10422), .B1(n10439), .B2(n10421), .ZN(
        P2_U3423) );
  AOI22_X1 U11463 ( .A1(n10440), .A2(n10424), .B1(n5131), .B2(n10437), .ZN(
        P2_U3460) );
  INV_X1 U11464 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U11465 ( .A1(n10440), .A2(n10426), .B1(n10425), .B2(n10437), .ZN(
        P2_U3461) );
  AOI22_X1 U11466 ( .A1(n10440), .A2(n10427), .B1(n5167), .B2(n10437), .ZN(
        P2_U3462) );
  AOI22_X1 U11467 ( .A1(n10440), .A2(n10428), .B1(n7020), .B2(n10437), .ZN(
        P2_U3463) );
  AOI22_X1 U11468 ( .A1(n10440), .A2(n10430), .B1(n10429), .B2(n10437), .ZN(
        P2_U3464) );
  AOI22_X1 U11469 ( .A1(n10440), .A2(n10431), .B1(n7024), .B2(n10437), .ZN(
        P2_U3465) );
  AOI22_X1 U11470 ( .A1(n10440), .A2(n10432), .B1(n7015), .B2(n10437), .ZN(
        P2_U3466) );
  AOI22_X1 U11471 ( .A1(n10440), .A2(n10433), .B1(n5269), .B2(n10437), .ZN(
        P2_U3467) );
  AOI22_X1 U11472 ( .A1(n10440), .A2(n10435), .B1(n10434), .B2(n10437), .ZN(
        P2_U3468) );
  AOI22_X1 U11473 ( .A1(n10440), .A2(n10436), .B1(n7476), .B2(n10437), .ZN(
        P2_U3469) );
  AOI22_X1 U11474 ( .A1(n10440), .A2(n10439), .B1(n10438), .B2(n10437), .ZN(
        P2_U3470) );
  NOR2_X1 U11475 ( .A1(n10442), .A2(n10441), .ZN(n10443) );
  XOR2_X1 U11476 ( .A(n10443), .B(P2_ADDR_REG_1__SCAN_IN), .Z(ADD_1068_U5) );
  XOR2_X1 U11477 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11478 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10445), .A(n10444), 
        .ZN(n10447) );
  XOR2_X1 U11479 ( .A(n10447), .B(n10446), .Z(ADD_1068_U55) );
  XNOR2_X1 U11480 ( .A(n10449), .B(n10448), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11481 ( .A(n10451), .B(n10450), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11482 ( .A(n10453), .B(n10452), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11483 ( .A(n10455), .B(n10454), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11484 ( .A(n10457), .B(n10456), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11485 ( .A(n10459), .B(n10458), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11486 ( .A(n10461), .B(n10460), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11487 ( .A(n10463), .B(n10462), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11488 ( .A(n10465), .B(n10464), .ZN(ADD_1068_U47) );
  XOR2_X1 U11489 ( .A(n10467), .B(n10466), .Z(ADD_1068_U54) );
  XNOR2_X1 U11490 ( .A(n10469), .B(n10468), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11491 ( .A(n10471), .B(n10470), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11492 ( .A(n10473), .B(n10472), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11493 ( .A(n10475), .B(n10474), .ZN(ADD_1068_U50) );
  XOR2_X1 U11494 ( .A(n10477), .B(n10476), .Z(ADD_1068_U53) );
  XNOR2_X1 U11495 ( .A(n10479), .B(n10478), .ZN(ADD_1068_U52) );
  NAND2_X1 U8141 ( .A1(n9986), .A2(n6565), .ZN(n9425) );
  CLKBUF_X2 U5018 ( .A(n6097), .Z(n6191) );
  NAND2_X1 U6391 ( .A1(n9353), .A2(n8501), .ZN(n5209) );
endmodule

