

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506;

  NAND2_X1 U4784 ( .A1(n9934), .A2(n9939), .ZN(n9935) );
  OR2_X1 U4785 ( .A1(n9425), .A2(n8800), .ZN(n6003) );
  NAND2_X1 U4786 ( .A1(n8506), .A2(n8503), .ZN(n8595) );
  CLKBUF_X2 U4787 ( .A(n9136), .Z(n4279) );
  CLKBUF_X2 U4788 ( .A(n4470), .Z(n4282) );
  INV_X2 U4790 ( .A(n6647), .ZN(n6618) );
  NAND2_X1 U4791 ( .A1(n5263), .A2(n5262), .ZN(n9136) );
  NAND2_X1 U4792 ( .A1(n5008), .A2(n5007), .ZN(n5263) );
  NAND2_X1 U4793 ( .A1(n7096), .A2(n5142), .ZN(n5328) );
  CLKBUF_X2 U4794 ( .A(n5175), .Z(n4280) );
  MUX2_X1 U4795 ( .A(n8476), .B(n8475), .S(n4285), .Z(n8483) );
  NAND2_X1 U4796 ( .A1(n8225), .A2(n6040), .ZN(n6153) );
  NOR2_X1 U4797 ( .A1(n8603), .A2(n7723), .ZN(n6351) );
  INV_X1 U4798 ( .A(n7795), .ZN(n4912) );
  INV_X2 U4799 ( .A(n7020), .ZN(n7035) );
  NAND2_X1 U4800 ( .A1(n8429), .A2(n10249), .ZN(n6306) );
  NAND2_X2 U4802 ( .A1(n7120), .A2(n9136), .ZN(n6739) );
  NOR2_X1 U4803 ( .A1(n10258), .A2(n10263), .ZN(n4915) );
  INV_X1 U4804 ( .A(n7169), .ZN(n6643) );
  INV_X1 U4805 ( .A(n10246), .ZN(n6251) );
  AND2_X1 U4806 ( .A1(n6402), .A2(n6401), .ZN(n8512) );
  AOI21_X1 U4807 ( .B1(n8965), .B2(n8963), .A(n8964), .ZN(n8967) );
  NAND2_X1 U4808 ( .A1(n6048), .A2(n5962), .ZN(n6752) );
  NAND2_X1 U4809 ( .A1(n5596), .A2(n5595), .ZN(n9281) );
  NAND2_X1 U4810 ( .A1(n5718), .A2(n5717), .ZN(n9419) );
  INV_X1 U4811 ( .A(n8188), .ZN(n10209) );
  NAND2_X1 U4812 ( .A1(n8534), .A2(n8537), .ZN(n10028) );
  NAND2_X1 U4813 ( .A1(n8480), .A2(n8471), .ZN(n8603) );
  INV_X1 U4814 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4803) );
  INV_X1 U4815 ( .A(n9484), .ZN(n9338) );
  AND3_X1 U4816 ( .A1(n5333), .A2(n5332), .A3(n5331), .ZN(n7748) );
  INV_X1 U4817 ( .A(n7455), .ZN(n9741) );
  NAND2_X1 U4818 ( .A1(n6633), .A2(n6725), .ZN(n8591) );
  XNOR2_X1 U4819 ( .A(n6637), .B(n6636), .ZN(n8600) );
  CLKBUF_X2 U4820 ( .A(n10365), .Z(n4278) );
  NAND2_X1 U4821 ( .A1(n6339), .A2(n4434), .ZN(n10365) );
  INV_X2 U4822 ( .A(n9737), .ZN(n7676) );
  INV_X2 U4823 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5382) );
  INV_X1 U4824 ( .A(n7730), .ZN(n7845) );
  NOR2_X2 U4825 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5134) );
  AOI21_X2 U4826 ( .B1(n7810), .B2(n7826), .A(n8251), .ZN(n7811) );
  NAND2_X2 U4827 ( .A1(n8445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6247) );
  BUF_X4 U4828 ( .A(n5175), .Z(n4281) );
  NAND2_X1 U4829 ( .A1(n4808), .A2(n4809), .ZN(n5175) );
  AOI211_X2 U4830 ( .C1(n10135), .C2(n10195), .A(n10134), .B(n10133), .ZN(
        n10219) );
  MUX2_X1 U4831 ( .A(n9350), .B(n9417), .S(n10448), .Z(n9352) );
  MUX2_X1 U4832 ( .A(n9418), .B(n9417), .S(n10440), .Z(n9422) );
  INV_X1 U4833 ( .A(n5335), .ZN(n4470) );
  XNOR2_X2 U4834 ( .A(n4492), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7208) );
  NAND3_X1 U4835 ( .A1(n4912), .A2(n7076), .A3(n4911), .ZN(n4283) );
  NAND3_X1 U4836 ( .A1(n4912), .A2(n7076), .A3(n4911), .ZN(n4284) );
  NAND3_X2 U4837 ( .A1(n4912), .A2(n7076), .A3(n4911), .ZN(n7020) );
  NAND2_X1 U4838 ( .A1(n6959), .A2(n4922), .ZN(n4921) );
  AOI21_X1 U4839 ( .B1(n5083), .B2(n4663), .A(n4662), .ZN(n4661) );
  NAND2_X1 U4840 ( .A1(n6571), .A2(n6570), .ZN(n9921) );
  AND2_X1 U4841 ( .A1(n5720), .A2(n5719), .ZN(n9148) );
  AND2_X1 U4842 ( .A1(n4368), .A2(n5897), .ZN(n9329) );
  AOI21_X1 U4843 ( .B1(n5098), .B2(n4344), .A(n5096), .ZN(n5095) );
  NAND2_X1 U4844 ( .A1(n5581), .A2(n5580), .ZN(n9393) );
  AND2_X1 U4845 ( .A1(n4396), .A2(n7712), .ZN(n8113) );
  AND2_X1 U4846 ( .A1(n5498), .A2(n5497), .ZN(n8790) );
  INV_X2 U4847 ( .A(n6147), .ZN(n6148) );
  AND2_X1 U4848 ( .A1(n5306), .A2(n4849), .ZN(n10427) );
  OR2_X1 U4849 ( .A1(n8923), .A2(n7583), .ZN(n5352) );
  NOR2_X1 U4850 ( .A1(n9745), .A2(n10381), .ZN(n8598) );
  OR2_X1 U4851 ( .A1(n8923), .A2(n10414), .ZN(n5856) );
  INV_X1 U4852 ( .A(n9743), .ZN(n7478) );
  INV_X4 U4853 ( .A(n7004), .ZN(n6849) );
  INV_X1 U4854 ( .A(n8921), .ZN(n8037) );
  INV_X1 U4855 ( .A(n6851), .ZN(n6834) );
  INV_X2 U4856 ( .A(n8582), .ZN(n4285) );
  INV_X1 U4857 ( .A(n8420), .ZN(n6592) );
  INV_X2 U4858 ( .A(n7082), .ZN(n6152) );
  INV_X1 U4859 ( .A(n6739), .ZN(n7084) );
  INV_X2 U4860 ( .A(n6306), .ZN(n7155) );
  NAND2_X2 U4861 ( .A1(n4915), .A2(n6728), .ZN(n7076) );
  OAI211_X2 U4862 ( .C1(n6502), .C2(n6501), .A(n6500), .B(n6499), .ZN(n8590)
         );
  INV_X1 U4863 ( .A(n8395), .ZN(n6252) );
  AND2_X1 U4864 ( .A1(n5329), .A2(n5366), .ZN(n7329) );
  INV_X2 U4865 ( .A(n4280), .ZN(n5184) );
  NAND2_X1 U4866 ( .A1(n4603), .A2(n6043), .ZN(n6052) );
  NAND2_X1 U4867 ( .A1(n4378), .A2(n4442), .ZN(n4535) );
  OAI21_X1 U4868 ( .B1(n6205), .B2(n9293), .A(n6204), .ZN(n9167) );
  NAND2_X1 U4869 ( .A1(n4831), .A2(n4340), .ZN(n8592) );
  AND2_X1 U4870 ( .A1(n4926), .A2(n4924), .ZN(n8718) );
  NAND2_X1 U4871 ( .A1(n9702), .A2(n7029), .ZN(n7041) );
  OR2_X1 U4872 ( .A1(n4666), .A2(n4664), .ZN(n10223) );
  INV_X1 U4873 ( .A(n6166), .ZN(n7075) );
  AOI21_X1 U4874 ( .B1(n4490), .B2(n10087), .A(n4488), .ZN(n10131) );
  NAND2_X1 U4875 ( .A1(n9903), .A2(n9905), .ZN(n9904) );
  OAI22_X1 U4876 ( .A1(n6207), .A2(n4520), .B1(n4521), .B2(n5108), .ZN(n6738)
         );
  OAI21_X1 U4877 ( .B1(n4479), .B2(n4478), .A(n4476), .ZN(n4701) );
  AND2_X1 U4878 ( .A1(n9114), .A2(n4572), .ZN(n9076) );
  AND2_X1 U4879 ( .A1(n6992), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U4880 ( .A1(n9552), .A2(n6950), .ZN(n6959) );
  NAND2_X1 U4881 ( .A1(n5995), .A2(n5994), .ZN(n9410) );
  NAND2_X1 U4882 ( .A1(n5809), .A2(n5808), .ZN(n6206) );
  NAND2_X1 U4883 ( .A1(n8422), .A2(n8421), .ZN(n8731) );
  AND2_X1 U4884 ( .A1(n6569), .A2(n4789), .ZN(n4788) );
  AND2_X1 U4885 ( .A1(n8705), .A2(n8555), .ZN(n8624) );
  NAND2_X1 U4886 ( .A1(n8417), .A2(n8416), .ZN(n10216) );
  AND2_X1 U4887 ( .A1(n5954), .A2(n5953), .ZN(n9416) );
  NOR2_X1 U4888 ( .A1(n5044), .A2(n5040), .ZN(n4599) );
  OR2_X1 U4889 ( .A1(n10127), .A2(n8559), .ZN(n8705) );
  NAND2_X1 U4890 ( .A1(n8805), .A2(n6114), .ZN(n8804) );
  OR2_X1 U4891 ( .A1(n6769), .A2(n6187), .ZN(n6048) );
  OR3_X1 U4892 ( .A1(n5979), .A2(n5982), .A3(n5978), .ZN(n5989) );
  NAND2_X1 U4893 ( .A1(n8645), .A2(n8632), .ZN(n9940) );
  NAND2_X1 U4894 ( .A1(n5702), .A2(n5701), .ZN(n6218) );
  AND2_X1 U4895 ( .A1(n5045), .A2(n5047), .ZN(n5044) );
  NOR2_X1 U4896 ( .A1(n6008), .A2(n5006), .ZN(n5005) );
  NAND2_X1 U4897 ( .A1(n6581), .A2(n6580), .ZN(n10129) );
  INV_X1 U4898 ( .A(n9190), .ZN(n9437) );
  OR2_X1 U4899 ( .A1(n9431), .A2(n8890), .ZN(n5931) );
  NAND2_X1 U4900 ( .A1(n5981), .A2(n5991), .ZN(n5979) );
  XNOR2_X1 U4901 ( .A(n5700), .B(n5712), .ZN(n9493) );
  OR2_X1 U4902 ( .A1(n5942), .A2(n5941), .ZN(n5981) );
  NAND2_X1 U4903 ( .A1(n6559), .A2(n6558), .ZN(n10139) );
  NAND2_X1 U4904 ( .A1(n5665), .A2(n5664), .ZN(n9431) );
  AND2_X1 U4905 ( .A1(n5265), .A2(n5264), .ZN(n9190) );
  NOR2_X1 U4906 ( .A1(n4772), .A2(n4496), .ZN(n4495) );
  AND2_X1 U4907 ( .A1(n5715), .A2(n5713), .ZN(n5700) );
  XNOR2_X1 U4908 ( .A(n5944), .B(n5943), .ZN(n8428) );
  NAND2_X1 U4909 ( .A1(n8238), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8347) );
  OAI222_X1 U4910 ( .A1(n10417), .A2(n10416), .B1(n10415), .B2(n10414), .C1(
        n10413), .C2(n10412), .ZN(n10418) );
  NAND2_X1 U4911 ( .A1(n5640), .A2(n5639), .ZN(n9370) );
  NAND2_X1 U4912 ( .A1(n6537), .A2(n6536), .ZN(n10151) );
  XNOR2_X1 U4913 ( .A(n5676), .B(n5675), .ZN(n8450) );
  XNOR2_X1 U4914 ( .A(n5260), .B(n5655), .ZN(n9501) );
  XNOR2_X1 U4915 ( .A(n5276), .B(n5275), .ZN(n8374) );
  AND2_X1 U4916 ( .A1(n5255), .A2(n5654), .ZN(n5260) );
  INV_X1 U4917 ( .A(n5089), .ZN(n5088) );
  AND2_X1 U4918 ( .A1(n5095), .A2(n6412), .ZN(n4545) );
  NAND2_X1 U4919 ( .A1(n5631), .A2(n5630), .ZN(n9454) );
  NAND2_X1 U4920 ( .A1(n6526), .A2(n6525), .ZN(n10231) );
  OR2_X1 U4921 ( .A1(n9270), .A2(n9247), .ZN(n9232) );
  AND2_X1 U4922 ( .A1(n9288), .A2(n4839), .ZN(n4471) );
  OR2_X1 U4923 ( .A1(n8002), .A2(n8594), .ZN(n4547) );
  OAI21_X1 U4924 ( .B1(n8278), .B2(n5064), .A(n6671), .ZN(n5063) );
  INV_X1 U4925 ( .A(n9288), .ZN(n4838) );
  AND2_X1 U4926 ( .A1(n5899), .A2(n5906), .ZN(n9318) );
  AOI21_X1 U4927 ( .B1(n9537), .B2(n9538), .A(n6887), .ZN(n6888) );
  OR2_X1 U4928 ( .A1(n9477), .A2(n6108), .ZN(n5899) );
  NAND2_X1 U4929 ( .A1(n4441), .A2(n4440), .ZN(n8094) );
  NAND2_X1 U4930 ( .A1(n5609), .A2(n5608), .ZN(n9270) );
  NAND2_X1 U4931 ( .A1(n6504), .A2(n6503), .ZN(n10168) );
  INV_X1 U4932 ( .A(n9291), .ZN(n9288) );
  NAND2_X1 U4933 ( .A1(n5514), .A2(n5513), .ZN(n9477) );
  AOI21_X1 U4934 ( .B1(n8200), .B2(n5491), .A(n4377), .ZN(n5038) );
  NAND2_X1 U4935 ( .A1(n7448), .A2(n7443), .ZN(n7464) );
  INV_X1 U4936 ( .A(n8093), .ZN(n4441) );
  INV_X1 U4937 ( .A(n8362), .ZN(n10198) );
  OR2_X1 U4938 ( .A1(n7668), .A2(n5992), .ZN(n5596) );
  INV_X1 U4939 ( .A(n8512), .ZN(n10204) );
  INV_X1 U4940 ( .A(n8283), .ZN(n9666) );
  AND2_X1 U4941 ( .A1(n5028), .A2(n5027), .ZN(n7448) );
  NAND2_X1 U4942 ( .A1(n5547), .A2(n5546), .ZN(n9484) );
  NAND2_X1 U4943 ( .A1(n6449), .A2(n6448), .ZN(n10190) );
  INV_X1 U4944 ( .A(n8790), .ZN(n8311) );
  OR2_X1 U4945 ( .A1(n7545), .A2(n7546), .ZN(n7543) );
  AND2_X1 U4946 ( .A1(n6435), .A2(n6434), .ZN(n8362) );
  OR2_X1 U4947 ( .A1(n7400), .A2(n5992), .ZN(n5547) );
  AOI21_X1 U4948 ( .B1(n4978), .B2(n4976), .A(n4303), .ZN(n4975) );
  NAND2_X1 U4949 ( .A1(n6468), .A2(n6467), .ZN(n10178) );
  AND2_X1 U4950 ( .A1(n7696), .A2(n6079), .ZN(n4978) );
  AND2_X1 U4951 ( .A1(n8505), .A2(n8508), .ZN(n8596) );
  NAND2_X1 U4952 ( .A1(n6458), .A2(n6457), .ZN(n10186) );
  NAND2_X1 U4953 ( .A1(n5570), .A2(n5569), .ZN(n9471) );
  NAND2_X1 U4954 ( .A1(n5460), .A2(n5459), .ZN(n8215) );
  NAND2_X1 U4955 ( .A1(n6374), .A2(n6373), .ZN(n10102) );
  NOR2_X1 U4956 ( .A1(n7718), .A2(n7730), .ZN(n7721) );
  NAND2_X2 U4957 ( .A1(n7625), .A2(n10417), .ZN(n10421) );
  NOR2_X1 U4958 ( .A1(n7513), .A2(n7809), .ZN(n7514) );
  OR2_X1 U4959 ( .A1(n7814), .A2(n4574), .ZN(n4757) );
  NAND2_X1 U4960 ( .A1(n7444), .A2(n5844), .ZN(n5849) );
  NAND2_X1 U4961 ( .A1(n5314), .A2(n7379), .ZN(n7444) );
  NAND2_X1 U4962 ( .A1(n8604), .A2(n8598), .ZN(n7477) );
  INV_X1 U4963 ( .A(n10427), .ZN(n7379) );
  NAND2_X1 U4964 ( .A1(n6067), .A2(n10427), .ZN(n5844) );
  NAND2_X1 U4965 ( .A1(n5437), .A2(n5436), .ZN(n8269) );
  NAND2_X1 U4966 ( .A1(n5856), .A2(n5862), .ZN(n6015) );
  NAND2_X1 U4967 ( .A1(n4514), .A2(n4512), .ZN(n7634) );
  INV_X1 U4968 ( .A(n8466), .ZN(n4286) );
  NAND2_X2 U4969 ( .A1(n7794), .A2(n10379), .ZN(n10386) );
  INV_X1 U4970 ( .A(n8016), .ZN(n7500) );
  XNOR2_X1 U4971 ( .A(n5448), .B(n5447), .ZN(n7174) );
  NAND2_X1 U4972 ( .A1(n4371), .A2(n6303), .ZN(n9745) );
  NAND2_X1 U4973 ( .A1(n7150), .A2(n6592), .ZN(n4502) );
  INV_X1 U4974 ( .A(n10414), .ZN(n7583) );
  NAND2_X1 U4975 ( .A1(n5312), .A2(n10422), .ZN(n5850) );
  INV_X1 U4976 ( .A(n5861), .ZN(n4287) );
  XNOR2_X1 U4977 ( .A(n5379), .B(n5378), .ZN(n7150) );
  AND4_X1 U4978 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n8232)
         );
  NAND4_X1 U4979 ( .A1(n6325), .A2(n6324), .A3(n6323), .A4(n6322), .ZN(n9743)
         );
  AND2_X1 U4980 ( .A1(n6309), .A2(n6308), .ZN(n6656) );
  INV_X1 U4981 ( .A(n5291), .ZN(n10422) );
  NAND2_X4 U4982 ( .A1(n4283), .A2(n7004), .ZN(n6821) );
  AND4_X1 U4983 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n7455)
         );
  AND2_X1 U4984 ( .A1(n6310), .A2(n6311), .ZN(n6655) );
  NAND3_X1 U4985 ( .A1(n5290), .A2(n5024), .A3(n5023), .ZN(n5291) );
  AND2_X1 U4986 ( .A1(n4794), .A2(n4403), .ZN(n4798) );
  NAND2_X1 U4987 ( .A1(n4722), .A2(n5195), .ZN(n5421) );
  XNOR2_X1 U4988 ( .A(n5304), .B(n5303), .ZN(n7132) );
  XNOR2_X1 U4989 ( .A(n5347), .B(n5346), .ZN(n7138) );
  NAND4_X1 U4990 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n8922)
         );
  NAND4_X1 U4991 ( .A1(n5404), .A2(n5403), .A3(n5402), .A4(n5401), .ZN(n8921)
         );
  NAND4_X1 U4992 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n8923)
         );
  NAND2_X1 U4993 ( .A1(n5754), .A2(n5756), .ZN(n5757) );
  NAND2_X1 U4994 ( .A1(n8588), .A2(n8590), .ZN(n4454) );
  NAND3_X1 U4995 ( .A1(n5310), .A2(n5311), .A3(n5309), .ZN(n6067) );
  NAND2_X2 U4996 ( .A1(n4697), .A2(n7076), .ZN(n6851) );
  INV_X1 U4997 ( .A(n8591), .ZN(n8588) );
  NAND4_X2 U4998 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n5312)
         );
  CLKBUF_X3 U4999 ( .A(n7084), .Z(n4289) );
  NAND2_X1 U5000 ( .A1(n4325), .A2(n5183), .ZN(n4724) );
  AND2_X2 U5001 ( .A1(n8395), .A2(n10246), .ZN(n6270) );
  NAND2_X2 U5002 ( .A1(n10246), .A2(n6252), .ZN(n7169) );
  AND2_X1 U5003 ( .A1(n6706), .A2(n6237), .ZN(n6728) );
  AND2_X4 U5004 ( .A1(n6739), .A2(n4281), .ZN(n5365) );
  CLKBUF_X1 U5005 ( .A(n5388), .Z(n5996) );
  AND2_X1 U5006 ( .A1(n4914), .A2(n4913), .ZN(n7795) );
  NAND2_X1 U5007 ( .A1(n4538), .A2(n4448), .ZN(n10249) );
  AND2_X1 U5008 ( .A1(n4357), .A2(n5449), .ZN(n4577) );
  NAND3_X1 U5009 ( .A1(n5174), .A2(n5173), .A3(n5301), .ZN(n5325) );
  XNOR2_X1 U5010 ( .A(n6708), .B(n6707), .ZN(n10258) );
  OR2_X1 U5011 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  NAND2_X1 U5012 ( .A1(n6632), .A2(n6631), .ZN(n6725) );
  NAND2_X1 U5013 ( .A1(n4669), .A2(n4672), .ZN(n10246) );
  NAND2_X1 U5014 ( .A1(n4536), .A2(n4450), .ZN(n8429) );
  NOR2_X1 U5015 ( .A1(n5753), .A2(n4324), .ZN(n5756) );
  NAND2_X1 U5016 ( .A1(n6630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6632) );
  OR2_X1 U5017 ( .A1(n6249), .A2(n6246), .ZN(n4672) );
  OAI22_X1 U5018 ( .A1(n4519), .A2(n4515), .B1(n9136), .B2(n4281), .ZN(n5380)
         );
  INV_X1 U5019 ( .A(n6650), .ZN(n8665) );
  XNOR2_X1 U5020 ( .A(n6638), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6650) );
  XNOR2_X1 U5021 ( .A(n5607), .B(n4984), .ZN(n9130) );
  OR2_X1 U5022 ( .A1(n6635), .A2(n6634), .ZN(n6637) );
  NAND2_X1 U5023 ( .A1(n6237), .A2(n4332), .ZN(n4538) );
  NAND2_X1 U5024 ( .A1(n8431), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U5025 ( .A1(n5080), .A2(n4301), .ZN(n8445) );
  NOR2_X1 U5026 ( .A1(n4453), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U5027 ( .A1(n4482), .A2(n6304), .ZN(n5284) );
  AND2_X2 U5028 ( .A1(n6234), .A2(n6432), .ZN(n5080) );
  OR2_X1 U5029 ( .A1(n5426), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5438) );
  NOR2_X1 U5030 ( .A1(n4288), .A2(n5593), .ZN(n4979) );
  CLKBUF_X3 U5031 ( .A(n5184), .Z(n6238) );
  INV_X4 U5032 ( .A(n4281), .ZN(n7131) );
  NAND2_X1 U5033 ( .A1(n4982), .A2(n5105), .ZN(n4981) );
  NOR2_X1 U5034 ( .A1(n4983), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U5035 ( .A1(n4803), .A2(n4804), .ZN(n4802) );
  AND3_X1 U5036 ( .A1(n6446), .A2(n6223), .A3(n6466), .ZN(n5053) );
  INV_X1 U5037 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6223) );
  NOR2_X1 U5038 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6228) );
  INV_X1 U5039 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6241) );
  NOR2_X1 U5040 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6229) );
  NOR2_X1 U5041 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6233) );
  NOR2_X1 U5042 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6240) );
  INV_X1 U5043 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5384) );
  INV_X1 U5044 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5367) );
  INV_X1 U5045 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5732) );
  NOR2_X1 U5046 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5136) );
  NOR2_X1 U5047 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5135) );
  INV_X4 U5048 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  OR2_X1 U5049 ( .A1(n4981), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4288) );
  OR2_X1 U5050 ( .A1(n5593), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4550) );
  XNOR2_X1 U5051 ( .A(n5749), .B(n5748), .ZN(n5758) );
  NAND2_X2 U5052 ( .A1(n5850), .A2(n5848), .ZN(n5293) );
  NAND2_X1 U5053 ( .A1(n6779), .A2(n8626), .ZN(n9874) );
  OAI22_X1 U5054 ( .A1(n10001), .A2(n6679), .B1(n10021), .B2(n10004), .ZN(
        n9978) );
  NAND2_X1 U5055 ( .A1(n7552), .A2(n5371), .ZN(n5373) );
  AOI21_X1 U5056 ( .B1(n8374), .B2(n5365), .A(n5113), .ZN(n6137) );
  OR2_X1 U5057 ( .A1(n6010), .A2(n6009), .ZN(n9282) );
  OAI222_X1 U5058 ( .A1(n10259), .A2(n7669), .B1(n10262), .B2(n7668), .C1(
        n10342), .C2(P1_U3086), .ZN(P1_U3337) );
  NAND2_X2 U5059 ( .A1(n5292), .A2(n5291), .ZN(n5848) );
  NAND2_X2 U5060 ( .A1(n4518), .A2(n4516), .ZN(n7120) );
  INV_X1 U5061 ( .A(n5849), .ZN(n7433) );
  OR2_X1 U5062 ( .A1(n4293), .A2(n5153), .ZN(n5154) );
  NAND2_X1 U5063 ( .A1(n5166), .A2(n5165), .ZN(n5282) );
  OR2_X1 U5064 ( .A1(n9393), .A2(n8812), .ZN(n5912) );
  OAI21_X1 U5065 ( .B1(n6238), .B2(n4580), .A(n4579), .ZN(n5197) );
  OR2_X1 U5066 ( .A1(n5472), .A2(n5471), .ZN(n4947) );
  NOR2_X2 U5067 ( .A1(n5643), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4763) );
  OR2_X2 U5068 ( .A1(n5641), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5643) );
  NOR2_X1 U5069 ( .A1(n5421), .A2(n4793), .ZN(n4792) );
  OR2_X1 U5070 ( .A1(n9281), .A2(n9297), .ZN(n9231) );
  NAND2_X2 U5071 ( .A1(n5373), .A2(n5372), .ZN(n7637) );
  NAND2_X2 U5072 ( .A1(n5912), .A2(n5799), .ZN(n9291) );
  XNOR2_X2 U5073 ( .A(n6247), .B(n8438), .ZN(n8395) );
  NAND2_X1 U5074 ( .A1(n5343), .A2(n5342), .ZN(n5347) );
  OR2_X2 U5075 ( .A1(n8269), .A2(n8164), .ZN(n5871) );
  NAND2_X1 U5076 ( .A1(n5506), .A2(n5505), .ZN(n8315) );
  OAI21_X2 U5077 ( .B1(n5757), .B2(P2_D_REG_0__SCAN_IN), .A(n7177), .ZN(n6062)
         );
  AOI21_X2 U5078 ( .B1(n5262), .B2(P2_IR_REG_31__SCAN_IN), .A(
        P2_IR_REG_28__SCAN_IN), .ZN(n4519) );
  NAND2_X2 U5079 ( .A1(n4795), .A2(n4798), .ZN(n5472) );
  NAND2_X1 U5080 ( .A1(n5588), .A2(n5233), .ZN(n5592) );
  AND2_X1 U5081 ( .A1(n5526), .A2(n5525), .ZN(n7338) );
  NAND2_X1 U5082 ( .A1(n5525), .A2(n5213), .ZN(n5537) );
  OR2_X2 U5083 ( .A1(n5334), .A2(n7748), .ZN(n5861) );
  INV_X2 U5084 ( .A(n5312), .ZN(n5292) );
  XNOR2_X2 U5085 ( .A(n5152), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5155) );
  AND2_X1 U5086 ( .A1(n6739), .A2(n4281), .ZN(n4290) );
  OAI21_X2 U5087 ( .B1(n8315), .B2(n5560), .A(n5559), .ZN(n9306) );
  INV_X1 U5088 ( .A(SI_16_), .ZN(n5222) );
  NAND2_X1 U5089 ( .A1(n5854), .A2(n7445), .ZN(n4467) );
  NOR2_X1 U5090 ( .A1(n7202), .A2(n4745), .ZN(n7204) );
  NOR2_X1 U5091 ( .A1(n7208), .A2(n10420), .ZN(n4745) );
  NAND2_X1 U5092 ( .A1(n9054), .A2(n9053), .ZN(n4633) );
  NAND2_X1 U5093 ( .A1(n9373), .A2(n9248), .ZN(n5051) );
  INV_X1 U5094 ( .A(n5889), .ZN(n5019) );
  NAND2_X1 U5095 ( .A1(n5150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5007) );
  OR2_X1 U5096 ( .A1(n5477), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U5097 ( .A1(n6688), .A2(n5077), .ZN(n5076) );
  NOR2_X1 U5098 ( .A1(n6690), .A2(n5078), .ZN(n5077) );
  INV_X1 U5099 ( .A(n6687), .ZN(n5078) );
  AND2_X1 U5100 ( .A1(n8588), .A2(n4914), .ZN(n7156) );
  AND2_X1 U5101 ( .A1(n8665), .A2(n8590), .ZN(n6802) );
  AOI21_X1 U5102 ( .B1(n4942), .B2(n4943), .A(n5523), .ZN(n4940) );
  NAND2_X1 U5103 ( .A1(n8201), .A2(n8200), .ZN(n8199) );
  NAND2_X1 U5104 ( .A1(n5039), .A2(n4598), .ZN(n4597) );
  NOR2_X1 U5105 ( .A1(n4599), .A2(n4359), .ZN(n4598) );
  NAND2_X1 U5106 ( .A1(n9245), .A2(n4345), .ZN(n5039) );
  AND2_X1 U5107 ( .A1(n6603), .A2(n6602), .ZN(n8559) );
  NAND2_X1 U5108 ( .A1(n7156), .A2(n8429), .ZN(n10045) );
  INV_X1 U5109 ( .A(n10085), .ZN(n10043) );
  NAND2_X1 U5110 ( .A1(n6306), .A2(n6238), .ZN(n8420) );
  NOR2_X1 U5111 ( .A1(n5853), .A2(n4287), .ZN(n4463) );
  AND2_X1 U5112 ( .A1(n9329), .A2(n4719), .ZN(n4718) );
  NOR2_X1 U5113 ( .A1(n4842), .A2(n5893), .ZN(n4719) );
  INV_X1 U5114 ( .A(n5894), .ZN(n4842) );
  INV_X1 U5115 ( .A(n5898), .ZN(n4717) );
  AND2_X1 U5116 ( .A1(n5899), .A2(n5908), .ZN(n4589) );
  NOR2_X1 U5117 ( .A1(n4837), .A2(n4471), .ZN(n4836) );
  NAND2_X1 U5118 ( .A1(n5905), .A2(n7082), .ZN(n4839) );
  AOI21_X1 U5119 ( .B1(n5917), .B2(n4346), .A(n4292), .ZN(n4841) );
  OAI21_X1 U5120 ( .B1(n8518), .B2(n8688), .A(n8528), .ZN(n8519) );
  NAND2_X1 U5121 ( .A1(n5334), .A2(n7748), .ZN(n5843) );
  NOR2_X1 U5122 ( .A1(n6752), .A2(n4366), .ZN(n4844) );
  NOR2_X1 U5123 ( .A1(n4352), .A2(n4846), .ZN(n4845) );
  NOR2_X1 U5124 ( .A1(n4333), .A2(n5042), .ZN(n5041) );
  INV_X1 U5125 ( .A(n5050), .ZN(n5042) );
  NOR2_X1 U5126 ( .A1(n5185), .A2(SI_5_), .ZN(n4727) );
  AND2_X1 U5127 ( .A1(n7223), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U5128 ( .A1(n7210), .A2(n7209), .ZN(n7212) );
  NAND2_X1 U5129 ( .A1(n4892), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4891) );
  INV_X1 U5130 ( .A(n9079), .ZN(n4627) );
  NOR2_X1 U5131 ( .A1(n5004), .A2(n5003), .ZN(n5002) );
  NAND2_X1 U5132 ( .A1(n9288), .A2(n5908), .ZN(n5004) );
  AND2_X1 U5133 ( .A1(n5530), .A2(n8739), .ZN(n5515) );
  INV_X1 U5134 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8766) );
  NOR2_X1 U5135 ( .A1(n6062), .A2(n6764), .ZN(n6151) );
  OR2_X1 U5136 ( .A1(n9454), .A2(n9248), .ZN(n5922) );
  NAND2_X1 U5137 ( .A1(n9313), .A2(n5906), .ZN(n5798) );
  NOR2_X1 U5138 ( .A1(n5148), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U5139 ( .A1(n6972), .A2(n6971), .ZN(n4684) );
  AND2_X1 U5140 ( .A1(n6803), .A2(n7076), .ZN(n4455) );
  INV_X1 U5141 ( .A(n9615), .ZN(n4907) );
  INV_X1 U5142 ( .A(n6925), .ZN(n4908) );
  INV_X1 U5143 ( .A(n4910), .ZN(n4909) );
  NAND2_X1 U5144 ( .A1(n4834), .A2(n9875), .ZN(n4833) );
  NAND2_X1 U5145 ( .A1(n4294), .A2(n4342), .ZN(n4929) );
  INV_X1 U5146 ( .A(n8662), .ZN(n4930) );
  NOR2_X1 U5147 ( .A1(n4900), .A2(n4899), .ZN(n4898) );
  OR2_X1 U5148 ( .A1(n9880), .A2(n10127), .ZN(n4900) );
  NAND2_X1 U5149 ( .A1(n6695), .A2(n9902), .ZN(n4899) );
  NAND2_X1 U5150 ( .A1(n4543), .A2(n8701), .ZN(n4542) );
  INV_X1 U5151 ( .A(n9905), .ZN(n4543) );
  INV_X1 U5152 ( .A(n8701), .ZN(n4544) );
  OR2_X1 U5153 ( .A1(n10129), .A2(n9916), .ZN(n8647) );
  AND2_X1 U5154 ( .A1(n5061), .A2(n4385), .ZN(n4773) );
  INV_X1 U5155 ( .A(n6670), .ZN(n5064) );
  AND2_X1 U5156 ( .A1(n7708), .A2(n4614), .ZN(n6665) );
  AND2_X1 U5157 ( .A1(n7707), .A2(n8045), .ZN(n4614) );
  OR2_X1 U5158 ( .A1(n9880), .A2(n7049), .ZN(n8654) );
  AND2_X1 U5159 ( .A1(n6579), .A2(n8632), .ZN(n5093) );
  NAND2_X1 U5160 ( .A1(n4788), .A2(n4791), .ZN(n4787) );
  NAND2_X1 U5161 ( .A1(n9969), .A2(n4788), .ZN(n4509) );
  AOI21_X1 U5162 ( .B1(n5070), .B2(n5069), .A(n4341), .ZN(n5068) );
  NAND2_X1 U5163 ( .A1(n5659), .A2(n4406), .ZN(n5694) );
  NOR2_X2 U5164 ( .A1(n4695), .A2(n6429), .ZN(n6432) );
  NOR2_X1 U5165 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6231) );
  NOR2_X1 U5166 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6232) );
  XNOR2_X1 U5167 ( .A(n5206), .B(SI_11_), .ZN(n5471) );
  NAND2_X1 U5168 ( .A1(n4802), .A2(n5162), .ZN(n4808) );
  NAND2_X1 U5169 ( .A1(n4698), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4809) );
  INV_X1 U5170 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5163) );
  INV_X1 U5171 ( .A(n4956), .ZN(n4569) );
  AOI21_X1 U5172 ( .B1(n8880), .B2(n4958), .A(n4957), .ZN(n4956) );
  NAND2_X1 U5173 ( .A1(n6129), .A2(n8773), .ZN(n8775) );
  OR2_X1 U5174 ( .A1(n5597), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5610) );
  AND2_X1 U5175 ( .A1(n6143), .A2(n8890), .ZN(n6144) );
  AND3_X1 U5176 ( .A1(n6062), .A2(n6157), .A3(n6764), .ZN(n6179) );
  INV_X1 U5177 ( .A(n4982), .ZN(n4980) );
  NAND2_X1 U5178 ( .A1(n9148), .A2(n5684), .ZN(n6001) );
  NAND2_X1 U5180 ( .A1(n4882), .A2(n7516), .ZN(n7814) );
  AND3_X1 U5181 ( .A1(n7529), .A2(n7814), .A3(P2_REG2_REG_7__SCAN_IN), .ZN(
        n8930) );
  AND2_X1 U5182 ( .A1(n8254), .A2(n8331), .ZN(n8255) );
  NAND2_X1 U5183 ( .A1(n8349), .A2(n8348), .ZN(n8988) );
  NAND2_X1 U5184 ( .A1(n9021), .A2(n4596), .ZN(n9023) );
  NAND2_X1 U5185 ( .A1(n9027), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4596) );
  INV_X1 U5186 ( .A(n9028), .ZN(n4635) );
  NAND2_X1 U5187 ( .A1(n5035), .A2(n5114), .ZN(n5034) );
  INV_X1 U5188 ( .A(n9273), .ZN(n5035) );
  AND2_X1 U5189 ( .A1(n5794), .A2(n5871), .ZN(n5009) );
  AND2_X1 U5190 ( .A1(n7080), .A2(n8446), .ZN(n6158) );
  INV_X1 U5191 ( .A(n9215), .ZN(n5045) );
  OR2_X1 U5192 ( .A1(n9370), .A2(n9206), .ZN(n5050) );
  NAND2_X1 U5193 ( .A1(n9462), .A2(n9227), .ZN(n5626) );
  INV_X1 U5194 ( .A(n9206), .ZN(n9226) );
  OR2_X1 U5195 ( .A1(n8835), .A2(n9227), .ZN(n9233) );
  INV_X1 U5196 ( .A(n5018), .ZN(n5017) );
  OAI21_X1 U5197 ( .B1(n5021), .B2(n4322), .A(n5797), .ZN(n5018) );
  AND2_X1 U5198 ( .A1(n6170), .A2(n7082), .ZN(n9331) );
  NAND2_X1 U5199 ( .A1(n8304), .A2(n8225), .ZN(n10434) );
  AND2_X1 U5200 ( .A1(n6154), .A2(n6049), .ZN(n9293) );
  NAND2_X1 U5201 ( .A1(n6802), .A2(n8591), .ZN(n4911) );
  NAND2_X1 U5202 ( .A1(n4503), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6572) );
  INV_X1 U5203 ( .A(n6803), .ZN(n4697) );
  AND2_X1 U5204 ( .A1(n4405), .A2(n6958), .ZN(n4922) );
  BUF_X1 U5205 ( .A(n6270), .Z(n7168) );
  BUF_X1 U5206 ( .A(n6617), .Z(n6529) );
  INV_X1 U5207 ( .A(n6270), .ZN(n6621) );
  NAND2_X2 U5208 ( .A1(n6252), .A2(n6251), .ZN(n6617) );
  INV_X1 U5209 ( .A(n8731), .ZN(n8581) );
  NAND2_X1 U5210 ( .A1(n9924), .A2(n4443), .ZN(n6792) );
  NOR2_X1 U5211 ( .A1(n9890), .A2(n4444), .ZN(n4443) );
  NAND2_X1 U5212 ( .A1(n9902), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U5213 ( .A1(n5073), .A2(n6693), .ZN(n6779) );
  OR2_X1 U5214 ( .A1(n5119), .A2(n6692), .ZN(n6693) );
  NAND2_X1 U5215 ( .A1(n5076), .A2(n5074), .ZN(n5073) );
  NAND2_X1 U5216 ( .A1(n9904), .A2(n8701), .ZN(n8402) );
  AND2_X1 U5217 ( .A1(n8647), .A2(n8701), .ZN(n9905) );
  NAND2_X1 U5218 ( .A1(n10011), .A2(n10163), .ZN(n10002) );
  NOR2_X1 U5219 ( .A1(n4343), .A2(n5057), .ZN(n5056) );
  INV_X1 U5220 ( .A(n8508), .ZN(n5096) );
  INV_X1 U5221 ( .A(n8503), .ZN(n5097) );
  AND2_X1 U5222 ( .A1(n7156), .A2(n7278), .ZN(n10085) );
  NAND2_X1 U5223 ( .A1(n4454), .A2(n8716), .ZN(n6651) );
  NAND2_X1 U5224 ( .A1(n6639), .A2(n8587), .ZN(n10087) );
  NAND2_X1 U5225 ( .A1(n4810), .A2(n6417), .ZN(n8283) );
  NAND2_X1 U5226 ( .A1(n7338), .A2(n6514), .ZN(n4810) );
  INV_X1 U5227 ( .A(n8429), .ZN(n7278) );
  AND2_X1 U5228 ( .A1(n7157), .A2(n6729), .ZN(n7162) );
  AND2_X1 U5229 ( .A1(n7076), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6729) );
  INV_X1 U5230 ( .A(n5080), .ZN(n6237) );
  XNOR2_X1 U5231 ( .A(n4529), .B(n5615), .ZN(n8102) );
  AOI21_X1 U5232 ( .B1(n4935), .B2(n5589), .A(n4313), .ZN(n4527) );
  INV_X1 U5233 ( .A(n4935), .ZN(n4528) );
  OR2_X1 U5234 ( .A1(n6371), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6385) );
  XNOR2_X1 U5235 ( .A(n4559), .B(n8831), .ZN(n4558) );
  AOI21_X1 U5236 ( .B1(n8828), .B2(n4557), .A(n4556), .ZN(n4559) );
  AND2_X1 U5237 ( .A1(n8827), .A2(n9193), .ZN(n4556) );
  NAND2_X1 U5238 ( .A1(n4595), .A2(n9054), .ZN(n4888) );
  INV_X1 U5239 ( .A(n9023), .ZN(n4595) );
  NAND2_X1 U5240 ( .A1(n8731), .A2(n8657), .ZN(n8627) );
  AND2_X1 U5241 ( .A1(n6791), .A2(n6790), .ZN(n9886) );
  AOI21_X1 U5242 ( .B1(n4465), .B2(n5866), .A(n5865), .ZN(n5867) );
  NAND2_X1 U5243 ( .A1(n4473), .A2(n4589), .ZN(n4472) );
  INV_X1 U5244 ( .A(n9318), .ZN(n4473) );
  OAI21_X1 U5245 ( .B1(n5895), .B2(n4304), .A(n4716), .ZN(n4475) );
  INV_X1 U5246 ( .A(n4589), .ZN(n4474) );
  NAND2_X1 U5247 ( .A1(n4836), .A2(n4838), .ZN(n4835) );
  INV_X1 U5248 ( .A(n5921), .ZN(n4702) );
  INV_X1 U5249 ( .A(n5922), .ZN(n4478) );
  NAND2_X1 U5250 ( .A1(n4826), .A2(n10051), .ZN(n8540) );
  AOI21_X1 U5251 ( .B1(n4335), .B2(n4285), .A(n4829), .ZN(n4828) );
  NOR2_X1 U5252 ( .A1(n4819), .A2(n4816), .ZN(n4815) );
  NOR2_X1 U5253 ( .A1(n8552), .A2(n4375), .ZN(n4816) );
  INV_X1 U5254 ( .A(n8553), .ZN(n4813) );
  NAND2_X1 U5255 ( .A1(n5419), .A2(n4336), .ZN(n5036) );
  OR2_X1 U5256 ( .A1(n9921), .A2(n9707), .ZN(n8635) );
  NOR2_X1 U5257 ( .A1(n6568), .A2(n9940), .ZN(n6569) );
  NAND2_X1 U5258 ( .A1(n9954), .A2(n4790), .ZN(n4789) );
  OAI21_X1 U5259 ( .B1(n7131), .B2(n4612), .A(n4611), .ZN(n5207) );
  NAND2_X1 U5260 ( .A1(n7131), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n4611) );
  NOR2_X1 U5261 ( .A1(n5206), .A2(SI_11_), .ZN(n4946) );
  NOR2_X1 U5262 ( .A1(n4727), .A2(n5196), .ZN(n4723) );
  NAND2_X1 U5263 ( .A1(n5374), .A2(n5377), .ZN(n5196) );
  NAND2_X1 U5264 ( .A1(n6238), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n4579) );
  OR2_X1 U5265 ( .A1(n4809), .A2(n4801), .ZN(n4807) );
  OAI21_X1 U5266 ( .B1(n4460), .B2(n4459), .A(n4457), .ZN(n5964) );
  INV_X1 U5267 ( .A(n4458), .ZN(n4457) );
  NAND2_X1 U5268 ( .A1(n4460), .A2(n4844), .ZN(n5966) );
  INV_X1 U5269 ( .A(n5262), .ZN(n4658) );
  INV_X1 U5270 ( .A(n8941), .ZN(n4864) );
  NAND2_X1 U5271 ( .A1(n8955), .A2(n4731), .ZN(n4730) );
  OR2_X1 U5272 ( .A1(n8253), .A2(n8242), .ZN(n4731) );
  NAND2_X1 U5273 ( .A1(n4881), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U5274 ( .A1(n4852), .A2(n4853), .ZN(n9033) );
  INV_X1 U5275 ( .A(n4855), .ZN(n4853) );
  OR2_X1 U5276 ( .A1(n8975), .A2(n4417), .ZN(n4852) );
  OAI21_X1 U5277 ( .B1(n4507), .B2(n4856), .A(n9032), .ZN(n4855) );
  INV_X1 U5278 ( .A(n9092), .ZN(n4738) );
  OAI21_X1 U5279 ( .B1(n6206), .B2(n4523), .A(n6044), .ZN(n4522) );
  INV_X1 U5280 ( .A(n6004), .ZN(n5932) );
  AND2_X1 U5281 ( .A1(n8766), .A2(n4769), .ZN(n4768) );
  INV_X1 U5282 ( .A(n5610), .ZN(n5131) );
  AND2_X1 U5283 ( .A1(n5858), .A2(n7634), .ZN(n5866) );
  NAND2_X1 U5284 ( .A1(n10422), .A2(n5292), .ZN(n7431) );
  NAND2_X1 U5285 ( .A1(n5293), .A2(n7503), .ZN(n7432) );
  OR2_X1 U5286 ( .A1(n9437), .A2(n8746), .ZN(n6006) );
  AND2_X1 U5287 ( .A1(n5051), .A2(n5626), .ZN(n5049) );
  AOI21_X1 U5288 ( .B1(n4999), .B2(n4997), .A(n4323), .ZN(n4623) );
  INV_X1 U5289 ( .A(n5002), .ZN(n4997) );
  AOI21_X1 U5290 ( .B1(n9259), .B2(n4298), .A(n4369), .ZN(n5030) );
  INV_X1 U5291 ( .A(n5114), .ZN(n5032) );
  AND2_X1 U5292 ( .A1(n8104), .A2(n9130), .ZN(n5814) );
  INV_X1 U5293 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5052) );
  INV_X1 U5294 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5773) );
  INV_X1 U5295 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U5296 ( .A1(n5732), .A2(n4984), .ZN(n4983) );
  NOR2_X1 U5297 ( .A1(n5565), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U5298 ( .A1(n9656), .A2(n6909), .ZN(n6912) );
  INV_X1 U5299 ( .A(n6377), .ZN(n4505) );
  NOR2_X1 U5300 ( .A1(n9573), .A2(n4683), .ZN(n4682) );
  INV_X1 U5301 ( .A(n6966), .ZN(n4683) );
  INV_X1 U5302 ( .A(n9614), .ZN(n4904) );
  AND2_X1 U5303 ( .A1(n4906), .A2(n4919), .ZN(n4686) );
  OR2_X1 U5304 ( .A1(n9890), .A2(n8562), .ZN(n8653) );
  OR2_X1 U5305 ( .A1(n6597), .A2(n6596), .ZN(n6607) );
  INV_X1 U5306 ( .A(n8696), .ZN(n5082) );
  NAND2_X1 U5307 ( .A1(n4508), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6540) );
  INV_X1 U5308 ( .A(n8537), .ZN(n4662) );
  INV_X1 U5309 ( .A(n6478), .ZN(n4663) );
  NAND2_X1 U5310 ( .A1(n4621), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U5311 ( .A1(n10071), .A2(n10072), .ZN(n10070) );
  INV_X1 U5312 ( .A(n8685), .ZN(n5090) );
  OAI21_X1 U5313 ( .B1(n6428), .B2(n5090), .A(n8529), .ZN(n5089) );
  OR2_X1 U5314 ( .A1(n6405), .A2(n6404), .ZN(n6420) );
  NAND2_X1 U5315 ( .A1(n4777), .A2(n8178), .ZN(n4576) );
  INV_X1 U5316 ( .A(n8151), .ZN(n4575) );
  AOI21_X1 U5317 ( .B1(n8151), .B2(n5066), .A(n4365), .ZN(n5065) );
  INV_X1 U5318 ( .A(n6666), .ZN(n5066) );
  INV_X1 U5319 ( .A(n4576), .ZN(n4480) );
  NAND2_X1 U5320 ( .A1(n4502), .A2(n4500), .ZN(n6663) );
  NOR2_X1 U5321 ( .A1(n8175), .A2(n4501), .ZN(n4500) );
  INV_X1 U5322 ( .A(n6277), .ZN(n4501) );
  NAND2_X1 U5323 ( .A1(n4435), .A2(n6661), .ZN(n7708) );
  NAND2_X1 U5324 ( .A1(n7478), .A2(n7500), .ZN(n8466) );
  OR2_X2 U5325 ( .A1(n9915), .A2(n10139), .ZN(n8632) );
  INV_X1 U5326 ( .A(n6681), .ZN(n5072) );
  INV_X1 U5327 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U5328 ( .A1(n5080), .A2(n5079), .ZN(n6248) );
  AND2_X1 U5329 ( .A1(n5829), .A2(n5699), .ZN(n5712) );
  AND2_X1 U5330 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  OR2_X1 U5331 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  INV_X1 U5332 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6704) );
  AOI21_X1 U5333 ( .B1(n4933), .B2(n4313), .A(n4415), .ZN(n4931) );
  XNOR2_X1 U5334 ( .A(n5226), .B(SI_17_), .ZN(n5576) );
  NAND2_X1 U5335 ( .A1(n4949), .A2(n4526), .ZN(n4525) );
  AOI21_X1 U5336 ( .B1(n4949), .B2(n4951), .A(n4374), .ZN(n4948) );
  INV_X1 U5337 ( .A(n4946), .ZN(n4944) );
  INV_X1 U5338 ( .A(n5405), .ZN(n4775) );
  NAND2_X1 U5339 ( .A1(n5325), .A2(n4581), .ZN(n5183) );
  AND2_X1 U5340 ( .A1(n5345), .A2(n5321), .ZN(n4581) );
  INV_X1 U5341 ( .A(n4727), .ZN(n4726) );
  INV_X1 U5342 ( .A(n4568), .ZN(n4567) );
  OAI21_X1 U5343 ( .B1(n4953), .B2(n4569), .A(n8763), .ZN(n4568) );
  INV_X1 U5344 ( .A(n8818), .ZN(n4954) );
  NAND2_X1 U5345 ( .A1(n8804), .A2(n8817), .ZN(n6118) );
  INV_X1 U5346 ( .A(n6146), .ZN(n4970) );
  INV_X1 U5347 ( .A(n4967), .ZN(n4966) );
  OAI21_X1 U5348 ( .B1(n8797), .B2(n6144), .A(n4968), .ZN(n4967) );
  INV_X1 U5349 ( .A(n8889), .ZN(n4968) );
  NAND2_X1 U5350 ( .A1(n4966), .A2(n6144), .ZN(n4964) );
  AND2_X1 U5351 ( .A1(n4971), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U5352 ( .A1(n4974), .A2(n4553), .ZN(n4552) );
  OAI21_X1 U5353 ( .B1(n8751), .B2(n8752), .A(n8868), .ZN(n6097) );
  NAND2_X1 U5354 ( .A1(n6118), .A2(n8818), .ZN(n8821) );
  NOR2_X1 U5355 ( .A1(n8899), .A2(n4961), .ZN(n4960) );
  INV_X1 U5356 ( .A(n6107), .ZN(n4961) );
  NAND2_X1 U5357 ( .A1(n4560), .A2(n8735), .ZN(n8736) );
  NAND2_X1 U5358 ( .A1(n8733), .A2(n8734), .ZN(n4560) );
  NAND2_X1 U5359 ( .A1(n6031), .A2(n4704), .ZN(n4703) );
  INV_X1 U5360 ( .A(n6041), .ZN(n6042) );
  NOR2_X1 U5361 ( .A1(n7082), .A2(n6040), .ZN(n4704) );
  AOI21_X1 U5362 ( .B1(n4996), .B2(n4339), .A(n4993), .ZN(n4992) );
  NAND2_X1 U5363 ( .A1(n4995), .A2(n4994), .ZN(n4993) );
  AND2_X1 U5364 ( .A1(n6001), .A2(n5737), .ZN(n6187) );
  AND2_X1 U5365 ( .A1(n5674), .A2(n5673), .ZN(n8890) );
  INV_X1 U5366 ( .A(n5958), .ZN(n5517) );
  NAND2_X1 U5367 ( .A1(n5354), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U5368 ( .A1(n5772), .A2(n5771), .ZN(n7080) );
  XNOR2_X1 U5369 ( .A(n7223), .B(n10444), .ZN(n7229) );
  NAND2_X1 U5370 ( .A1(n5305), .A2(n4493), .ZN(n5366) );
  NAND2_X1 U5371 ( .A1(n4740), .A2(n4739), .ZN(n7202) );
  OR2_X1 U5372 ( .A1(n7102), .A2(n7103), .ZN(n4739) );
  NAND2_X1 U5373 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  NAND2_X1 U5374 ( .A1(n4865), .A2(n7288), .ZN(n4866) );
  NAND2_X1 U5375 ( .A1(n7212), .A2(n7211), .ZN(n7304) );
  NAND3_X1 U5376 ( .A1(n4866), .A2(P2_REG1_REG_5__SCAN_IN), .A3(n7304), .ZN(
        n7306) );
  NAND2_X1 U5377 ( .A1(n7528), .A2(n7532), .ZN(n7529) );
  NAND2_X1 U5378 ( .A1(n4752), .A2(n4751), .ZN(n7528) );
  NAND2_X1 U5379 ( .A1(n4884), .A2(n7298), .ZN(n4751) );
  AOI21_X1 U5380 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7527), .A(n7511), .ZN(
        n7512) );
  OR2_X1 U5381 ( .A1(n4646), .A2(n8935), .ZN(n4639) );
  INV_X1 U5382 ( .A(n4647), .ZN(n4646) );
  OAI21_X1 U5383 ( .B1(n4648), .B2(n7523), .A(n8936), .ZN(n4647) );
  INV_X1 U5384 ( .A(n4648), .ZN(n4644) );
  NOR2_X1 U5385 ( .A1(n7512), .A2(n7532), .ZN(n7809) );
  NAND2_X1 U5386 ( .A1(n7514), .A2(n4328), .ZN(n4863) );
  NAND2_X1 U5387 ( .A1(n4758), .A2(n4755), .ZN(n4892) );
  AND2_X1 U5388 ( .A1(n4757), .A2(n4756), .ZN(n4755) );
  NOR2_X1 U5389 ( .A1(n4860), .A2(n4759), .ZN(n4756) );
  AND2_X1 U5390 ( .A1(n4506), .A2(n4863), .ZN(n7810) );
  INV_X1 U5391 ( .A(n4861), .ZN(n4506) );
  NAND2_X1 U5392 ( .A1(n7815), .A2(n4860), .ZN(n8951) );
  AND2_X1 U5393 ( .A1(n4757), .A2(n4760), .ZN(n4754) );
  OR2_X1 U5394 ( .A1(n4891), .A2(n4890), .ZN(n8953) );
  INV_X1 U5395 ( .A(n8951), .ZN(n4890) );
  AND2_X1 U5396 ( .A1(n4728), .A2(n8346), .ZN(n8238) );
  NAND2_X1 U5397 ( .A1(n4729), .A2(n8331), .ZN(n4728) );
  INV_X1 U5398 ( .A(n4730), .ZN(n4729) );
  NAND2_X1 U5399 ( .A1(n4730), .A2(n8241), .ZN(n8346) );
  NAND2_X1 U5400 ( .A1(n4872), .A2(n4873), .ZN(n8973) );
  AOI21_X1 U5401 ( .B1(n8335), .B2(n4875), .A(n4414), .ZN(n4873) );
  NAND2_X1 U5402 ( .A1(n8988), .A2(n4761), .ZN(n4881) );
  AND2_X1 U5403 ( .A1(n8980), .A2(n8987), .ZN(n4761) );
  NAND2_X1 U5404 ( .A1(n8989), .A2(n8999), .ZN(n9009) );
  NAND2_X1 U5405 ( .A1(n4878), .A2(n9009), .ZN(n9007) );
  INV_X1 U5406 ( .A(n4879), .ZN(n4878) );
  NAND2_X1 U5407 ( .A1(n4584), .A2(n9054), .ZN(n9035) );
  INV_X1 U5408 ( .A(n9033), .ZN(n4584) );
  NAND2_X1 U5409 ( .A1(n9062), .A2(n9061), .ZN(n4868) );
  NAND2_X1 U5410 ( .A1(n4416), .A2(n4633), .ZN(n4629) );
  NAND2_X1 U5411 ( .A1(n4632), .A2(n4634), .ZN(n4631) );
  INV_X1 U5412 ( .A(n9001), .ZN(n4632) );
  NAND2_X1 U5413 ( .A1(n4634), .A2(n4633), .ZN(n4630) );
  NAND2_X1 U5414 ( .A1(n5667), .A2(n5666), .ZN(n5682) );
  INV_X1 U5415 ( .A(n5668), .ZN(n5667) );
  NAND2_X1 U5416 ( .A1(n5048), .A2(n5051), .ZN(n5047) );
  INV_X1 U5417 ( .A(n9237), .ZN(n5048) );
  AND2_X1 U5418 ( .A1(n9259), .A2(n4319), .ZN(n5033) );
  NAND2_X1 U5419 ( .A1(n9290), .A2(n4838), .ZN(n4510) );
  AND2_X1 U5420 ( .A1(n4311), .A2(n4765), .ZN(n4764) );
  INV_X1 U5421 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4765) );
  AND4_X1 U5422 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n8784)
         );
  AND2_X1 U5423 ( .A1(n7760), .A2(n6012), .ZN(n5011) );
  NOR2_X1 U5424 ( .A1(n7082), .A2(n5779), .ZN(n6761) );
  NAND2_X1 U5425 ( .A1(n5760), .A2(n5759), .ZN(n6764) );
  OR2_X1 U5426 ( .A1(n5757), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U5427 ( .A1(n9172), .A2(n9331), .ZN(n5739) );
  NAND2_X1 U5428 ( .A1(n6207), .A2(n6206), .ZN(n9160) );
  AND2_X1 U5429 ( .A1(n6006), .A2(n6005), .ZN(n9198) );
  OR2_X1 U5430 ( .A1(n6008), .A2(n5804), .ZN(n9204) );
  NAND2_X1 U5431 ( .A1(n9245), .A2(n5049), .ZN(n5046) );
  INV_X1 U5432 ( .A(n9204), .ZN(n9201) );
  NAND2_X1 U5433 ( .A1(n7082), .A2(n6183), .ZN(n9298) );
  INV_X1 U5434 ( .A(n8812), .ZN(n9308) );
  AND2_X1 U5435 ( .A1(n5016), .A2(n5897), .ZN(n5015) );
  OAI21_X1 U5436 ( .B1(n5017), .B2(n5014), .A(n4368), .ZN(n5013) );
  INV_X1 U5437 ( .A(n5897), .ZN(n5014) );
  INV_X1 U5438 ( .A(n4322), .ZN(n5016) );
  AND4_X1 U5439 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n8873)
         );
  AND2_X1 U5440 ( .A1(n9314), .A2(n5896), .ZN(n8322) );
  INV_X1 U5441 ( .A(n8298), .ZN(n5021) );
  OR2_X1 U5442 ( .A1(n8194), .A2(n8200), .ZN(n8196) );
  INV_X1 U5443 ( .A(n9298), .ZN(n9333) );
  INV_X1 U5444 ( .A(n9293), .ZN(n9336) );
  NAND2_X1 U5445 ( .A1(n4516), .A2(n7131), .ZN(n4515) );
  NAND2_X1 U5446 ( .A1(n7082), .A2(n5814), .ZN(n6211) );
  AND2_X1 U5447 ( .A1(n6179), .A2(n6158), .ZN(n6215) );
  XNOR2_X1 U5448 ( .A(n5774), .B(n5773), .ZN(n7081) );
  OAI21_X1 U5449 ( .B1(n4316), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U5450 ( .A(n5496), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8986) );
  INV_X1 U5451 ( .A(n4606), .ZN(n5434) );
  NAND2_X1 U5452 ( .A1(n6835), .A2(n6836), .ZN(n6837) );
  NAND2_X1 U5453 ( .A1(n4619), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6584) );
  INV_X1 U5454 ( .A(n6572), .ZN(n4619) );
  NAND2_X1 U5455 ( .A1(n4678), .A2(n4681), .ZN(n4675) );
  INV_X1 U5456 ( .A(n6469), .ZN(n6470) );
  AOI21_X1 U5457 ( .B1(n6925), .B2(n6926), .A(n4360), .ZN(n4910) );
  INV_X1 U5458 ( .A(n6830), .ZN(n4916) );
  NAND2_X1 U5459 ( .A1(n9587), .A2(n4452), .ZN(n9685) );
  OR2_X1 U5460 ( .A1(n6895), .A2(n6894), .ZN(n4452) );
  NAND2_X1 U5461 ( .A1(n4833), .A2(n4832), .ZN(n4831) );
  AOI21_X1 U5462 ( .B1(n4925), .B2(n8664), .A(n8663), .ZN(n4924) );
  NAND2_X1 U5463 ( .A1(n4930), .A2(n4927), .ZN(n4926) );
  INV_X1 U5464 ( .A(n4929), .ZN(n4925) );
  AND3_X1 U5465 ( .A1(n6455), .A2(n6454), .A3(n6453), .ZN(n9519) );
  OR2_X1 U5466 ( .A1(n7169), .A2(n7188), .ZN(n6300) );
  NAND2_X1 U5467 ( .A1(n7367), .A2(n7368), .ZN(n4430) );
  NAND2_X1 U5468 ( .A1(n9816), .A2(n7275), .ZN(n7277) );
  OR2_X1 U5469 ( .A1(n7565), .A2(n7566), .ZN(n9836) );
  AND2_X1 U5470 ( .A1(n10283), .A2(n10282), .ZN(n10285) );
  AOI21_X1 U5471 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9851), .A(n10285), .ZN(
        n9839) );
  INV_X1 U5472 ( .A(n8419), .ZN(n9867) );
  NAND2_X1 U5473 ( .A1(n6616), .A2(n6615), .ZN(n9880) );
  NAND2_X1 U5474 ( .A1(n9941), .A2(n6686), .ZN(n6688) );
  AND2_X1 U5475 ( .A1(n6562), .A2(n6572), .ZN(n9937) );
  NAND2_X1 U5476 ( .A1(n9969), .A2(n8548), .ZN(n9945) );
  NAND2_X1 U5477 ( .A1(n6538), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6550) );
  INV_X1 U5478 ( .A(n6540), .ZN(n6538) );
  INV_X1 U5479 ( .A(n4503), .ZN(n6561) );
  NAND2_X1 U5480 ( .A1(n4486), .A2(n4487), .ZN(n6682) );
  INV_X1 U5481 ( .A(n9978), .ZN(n4486) );
  AND2_X1 U5482 ( .A1(n6524), .A2(n6523), .ZN(n9982) );
  NAND2_X1 U5483 ( .A1(n4447), .A2(n10016), .ZN(n4446) );
  INV_X1 U5484 ( .A(n4894), .ZN(n4447) );
  NOR2_X1 U5485 ( .A1(n10174), .A2(n10020), .ZN(n5057) );
  NOR2_X1 U5486 ( .A1(n6676), .A2(n5060), .ZN(n5059) );
  INV_X1 U5487 ( .A(n6674), .ZN(n5060) );
  NAND2_X1 U5488 ( .A1(n6469), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6487) );
  NOR2_X1 U5489 ( .A1(n10092), .A2(n4893), .ZN(n10054) );
  INV_X1 U5490 ( .A(n4895), .ZN(n4893) );
  NAND2_X1 U5491 ( .A1(n4498), .A2(n10063), .ZN(n4497) );
  INV_X1 U5492 ( .A(n4773), .ZN(n4772) );
  AOI21_X1 U5493 ( .B1(n5062), .B2(n5064), .A(n4362), .ZN(n5061) );
  AND2_X1 U5494 ( .A1(n8527), .A2(n8520), .ZN(n10083) );
  NAND2_X1 U5495 ( .A1(n8078), .A2(n6428), .ZN(n8273) );
  NAND2_X1 U5496 ( .A1(n8279), .A2(n8278), .ZN(n8277) );
  NAND2_X1 U5497 ( .A1(n8082), .A2(n8611), .ZN(n8081) );
  INV_X1 U5498 ( .A(n8596), .ZN(n8092) );
  OAI21_X1 U5499 ( .B1(n8110), .B2(n4485), .A(n4483), .ZN(n8091) );
  INV_X1 U5500 ( .A(n4484), .ZN(n4483) );
  OAI21_X1 U5501 ( .B1(n8595), .B2(n4485), .A(n8092), .ZN(n4484) );
  INV_X1 U5502 ( .A(n6667), .ZN(n4485) );
  NAND2_X1 U5503 ( .A1(n5099), .A2(n8597), .ZN(n8115) );
  OAI21_X1 U5504 ( .B1(n6665), .B2(n6664), .A(n4480), .ZN(n8172) );
  AND2_X1 U5505 ( .A1(n9742), .A2(n7605), .ZN(n7723) );
  INV_X1 U5506 ( .A(n10365), .ZN(n7605) );
  AND2_X1 U5507 ( .A1(n6355), .A2(n6354), .ZN(n7775) );
  NAND2_X1 U5508 ( .A1(n6592), .A2(n7136), .ZN(n6341) );
  NAND2_X1 U5509 ( .A1(n7155), .A2(n9760), .ZN(n6340) );
  INV_X1 U5510 ( .A(n10180), .ZN(n10397) );
  OAI211_X1 U5511 ( .C1(P1_B_REG_SCAN_IN), .C2(n10263), .A(n6728), .B(n6713), 
        .ZN(n7161) );
  INV_X1 U5512 ( .A(n8445), .ZN(n4671) );
  NAND2_X1 U5513 ( .A1(n5080), .A2(n7868), .ZN(n6236) );
  INV_X1 U5514 ( .A(n6248), .ZN(n4451) );
  INV_X1 U5515 ( .A(n6236), .ZN(n4449) );
  INV_X1 U5516 ( .A(n6702), .ZN(n4696) );
  OR2_X1 U5517 ( .A1(n7157), .A2(P1_U3086), .ZN(n8663) );
  XNOR2_X1 U5518 ( .A(n5606), .B(n5605), .ZN(n7837) );
  NAND2_X1 U5519 ( .A1(n5592), .A2(n5234), .ZN(n5606) );
  NAND2_X1 U5520 ( .A1(n5537), .A2(n5217), .ZN(n5540) );
  OAI21_X1 U5521 ( .B1(n4792), .B2(n4796), .A(n4942), .ZN(n5522) );
  XNOR2_X1 U5522 ( .A(n8828), .B(n8827), .ZN(n8829) );
  AND4_X1 U5523 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n8164)
         );
  AND2_X1 U5524 ( .A1(n5624), .A2(n5623), .ZN(n9227) );
  AND4_X1 U5525 ( .A1(n5536), .A2(n5535), .A3(n5534), .A4(n5533), .ZN(n8789)
         );
  INV_X1 U5526 ( .A(n8917), .ZN(n8751) );
  AOI21_X1 U5527 ( .B1(n9228), .B2(n5684), .A(n5636), .ZN(n9248) );
  AND2_X1 U5528 ( .A1(n5272), .A2(n5271), .ZN(n9214) );
  NAND2_X1 U5529 ( .A1(n6193), .A2(n10417), .ZN(n8896) );
  INV_X1 U5530 ( .A(n8890), .ZN(n9192) );
  INV_X1 U5531 ( .A(n9214), .ZN(n9193) );
  NAND2_X1 U5532 ( .A1(n5648), .A2(n5647), .ZN(n9206) );
  INV_X1 U5533 ( .A(n8873), .ZN(n8915) );
  INV_X1 U5534 ( .A(n8784), .ZN(n8916) );
  AOI21_X1 U5535 ( .B1(n7306), .B2(n7304), .A(n7305), .ZN(n7511) );
  NAND2_X1 U5536 ( .A1(n9026), .A2(n4634), .ZN(n9056) );
  INV_X1 U5537 ( .A(n4887), .ZN(n4886) );
  XNOR2_X1 U5538 ( .A(n4737), .B(n4420), .ZN(n4592) );
  NAND2_X1 U5539 ( .A1(n4733), .A2(n4732), .ZN(n4737) );
  AND2_X1 U5540 ( .A1(n4734), .A2(n9120), .ZN(n4732) );
  NAND2_X1 U5541 ( .A1(n4652), .A2(n9042), .ZN(n4651) );
  XNOR2_X1 U5542 ( .A(n4653), .B(n9138), .ZN(n4652) );
  INV_X1 U5543 ( .A(n9139), .ZN(n4653) );
  AOI21_X1 U5544 ( .B1(n9142), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9141), .ZN(
        n4654) );
  NOR2_X1 U5545 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  NOR2_X1 U5546 ( .A1(n8800), .A2(n9296), .ZN(n6203) );
  OR2_X1 U5547 ( .A1(n7625), .A2(n5812), .ZN(n9159) );
  NAND2_X1 U5548 ( .A1(n9404), .A2(n9394), .ZN(n9381) );
  NOR2_X1 U5549 ( .A1(n6759), .A2(n10428), .ZN(n6760) );
  INV_X1 U5550 ( .A(n6218), .ZN(n9356) );
  OR2_X1 U5551 ( .A1(n10441), .A2(n10434), .ZN(n9461) );
  AND4_X1 U5552 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(n9546)
         );
  NAND2_X1 U5553 ( .A1(n7406), .A2(n7407), .ZN(n4917) );
  XNOR2_X1 U5554 ( .A(n6837), .B(n6839), .ZN(n7453) );
  INV_X1 U5555 ( .A(n7041), .ZN(n9507) );
  INV_X1 U5556 ( .A(n9732), .ZN(n9583) );
  AND4_X1 U5557 ( .A1(n6383), .A2(n6382), .A3(n6381), .A4(n6380), .ZN(n9640)
         );
  NAND2_X1 U5558 ( .A1(n6516), .A2(n6515), .ZN(n10004) );
  AND2_X1 U5559 ( .A1(n7042), .A2(n7034), .ZN(n9672) );
  INV_X1 U5560 ( .A(n9709), .ZN(n9719) );
  AND2_X1 U5561 ( .A1(n7402), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9705) );
  INV_X1 U5562 ( .A(n9672), .ZN(n9724) );
  NAND2_X1 U5563 ( .A1(n7050), .A2(n7278), .ZN(n9717) );
  INV_X1 U5564 ( .A(n9712), .ZN(n9722) );
  INV_X1 U5565 ( .A(n9915), .ZN(n9950) );
  INV_X1 U5566 ( .A(n10046), .ZN(n10020) );
  INV_X1 U5567 ( .A(n10030), .ZN(n10074) );
  INV_X1 U5568 ( .A(n9519), .ZN(n10073) );
  NAND2_X1 U5569 ( .A1(n9790), .A2(n7271), .ZN(n9804) );
  NAND2_X1 U5570 ( .A1(n7420), .A2(n7419), .ZN(n9824) );
  OAI21_X1 U5571 ( .B1(n10349), .B2(n5162), .A(n9866), .ZN(n4618) );
  AOI21_X1 U5572 ( .B1(n8406), .B2(n10087), .A(n8405), .ZN(n8407) );
  XNOR2_X1 U5573 ( .A(n8400), .B(n4776), .ZN(n8414) );
  OAI21_X1 U5574 ( .B1(n9896), .B2(n8398), .A(n8399), .ZN(n4776) );
  INV_X1 U5575 ( .A(n4489), .ZN(n4488) );
  OAI21_X1 U5576 ( .B1(n9905), .B2(n9903), .A(n9904), .ZN(n4490) );
  AOI22_X1 U5577 ( .A1(n9906), .A2(n10377), .B1(n10085), .B2(n9932), .ZN(n4489) );
  NAND2_X1 U5578 ( .A1(n4668), .A2(n4667), .ZN(n4666) );
  AOI21_X1 U5579 ( .B1(n9932), .B2(n10377), .A(n4413), .ZN(n4667) );
  NAND2_X1 U5580 ( .A1(n9933), .A2(n10087), .ZN(n4668) );
  INV_X1 U5581 ( .A(n10369), .ZN(n10115) );
  NAND2_X1 U5582 ( .A1(n8190), .A2(n7841), .ZN(n10371) );
  AND2_X1 U5583 ( .A1(n10386), .A2(n7797), .ZN(n10366) );
  OR2_X1 U5584 ( .A1(n8433), .A2(n8420), .ZN(n8422) );
  AND3_X1 U5585 ( .A1(n4400), .A2(n6700), .A3(n4436), .ZN(n4442) );
  INV_X1 U5586 ( .A(n6699), .ZN(n4436) );
  NAND2_X1 U5587 ( .A1(n4504), .A2(n4355), .ZN(n6798) );
  AND2_X1 U5588 ( .A1(n6495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U5589 ( .A1(n6496), .A2(n6628), .ZN(n6500) );
  NAND2_X1 U5590 ( .A1(n4713), .A2(n6152), .ZN(n4712) );
  OAI21_X1 U5591 ( .B1(n4710), .B2(n4709), .A(n6152), .ZN(n4708) );
  NOR2_X1 U5592 ( .A1(n5876), .A2(n5872), .ZN(n4710) );
  OAI21_X1 U5593 ( .B1(n4707), .B2(n4706), .A(n7082), .ZN(n4705) );
  NAND2_X1 U5594 ( .A1(n5877), .A2(n5874), .ZN(n4706) );
  NOR2_X1 U5595 ( .A1(n5876), .A2(n5875), .ZN(n4707) );
  AND2_X1 U5596 ( .A1(n8486), .A2(n4285), .ZN(n4821) );
  INV_X1 U5597 ( .A(n5896), .ZN(n4843) );
  NAND2_X1 U5598 ( .A1(n4475), .A2(n9318), .ZN(n5907) );
  OAI21_X1 U5599 ( .B1(n4475), .B2(n4474), .A(n4353), .ZN(n4588) );
  INV_X1 U5600 ( .A(n4477), .ZN(n4476) );
  INV_X1 U5601 ( .A(n5924), .ZN(n4700) );
  NAND2_X1 U5602 ( .A1(n8532), .A2(n4327), .ZN(n4829) );
  INV_X1 U5603 ( .A(n8547), .ZN(n4817) );
  AND3_X1 U5604 ( .A1(n5936), .A2(n6006), .A3(n5805), .ZN(n5930) );
  NOR2_X1 U5605 ( .A1(n5931), .A2(n6152), .ZN(n4770) );
  NAND2_X1 U5606 ( .A1(n4814), .A2(n4812), .ZN(n8574) );
  INV_X1 U5607 ( .A(n8548), .ZN(n4790) );
  INV_X1 U5608 ( .A(n6684), .ZN(n5071) );
  INV_X1 U5609 ( .A(n9016), .ZN(n4856) );
  INV_X1 U5610 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5139) );
  INV_X1 U5611 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5140) );
  NAND4_X1 U5612 ( .A1(n5384), .A2(n5367), .A3(n5382), .A4(n5138), .ZN(n5565)
         );
  INV_X1 U5613 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5138) );
  INV_X1 U5614 ( .A(n5366), .ZN(n5567) );
  NOR2_X1 U5615 ( .A1(n6517), .A2(n9650), .ZN(n4508) );
  AND2_X1 U5616 ( .A1(n6278), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6266) );
  AND2_X1 U5617 ( .A1(n9739), .A2(n8009), .ZN(n8478) );
  INV_X1 U5618 ( .A(n7723), .ZN(n8467) );
  NOR2_X1 U5619 ( .A1(n4320), .A2(n5071), .ZN(n5069) );
  INV_X1 U5620 ( .A(n6685), .ZN(n5070) );
  NAND2_X1 U5621 ( .A1(n8113), .A2(n9551), .ZN(n8093) );
  OAI21_X2 U5622 ( .B1(n5659), .B2(n4939), .A(n4937), .ZN(n5833) );
  INV_X1 U5623 ( .A(n4938), .ZN(n4937) );
  OAI21_X1 U5624 ( .B1(n4406), .B2(n4939), .A(n5714), .ZN(n4938) );
  INV_X1 U5625 ( .A(n5693), .ZN(n4939) );
  INV_X1 U5626 ( .A(n4934), .ZN(n4933) );
  OAI21_X1 U5627 ( .B1(n4935), .B2(n4313), .A(n5615), .ZN(n4934) );
  INV_X1 U5628 ( .A(n5561), .ZN(n5223) );
  INV_X1 U5629 ( .A(n5218), .ZN(n4951) );
  INV_X1 U5630 ( .A(n5213), .ZN(n4526) );
  NAND2_X1 U5631 ( .A1(n6238), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n4601) );
  OAI21_X1 U5632 ( .B1(n6238), .B2(P1_DATAO_REG_10__SCAN_IN), .A(n4578), .ZN(
        n5203) );
  NAND2_X1 U5633 ( .A1(n6238), .A2(n5200), .ZN(n4578) );
  OAI21_X1 U5634 ( .B1(n4280), .B2(n4583), .A(n4582), .ZN(n5169) );
  NAND2_X1 U5635 ( .A1(n4280), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4582) );
  INV_X1 U5636 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4804) );
  INV_X1 U5637 ( .A(n8880), .ZN(n4959) );
  INV_X2 U5638 ( .A(n6147), .ZN(n6136) );
  NOR2_X1 U5639 ( .A1(n6085), .A2(n4554), .ZN(n4553) );
  AOI21_X1 U5640 ( .B1(n4974), .B2(n4972), .A(n4364), .ZN(n4971) );
  INV_X1 U5641 ( .A(n8158), .ZN(n4972) );
  INV_X1 U5642 ( .A(n8104), .ZN(n6040) );
  NAND2_X1 U5643 ( .A1(n9410), .A2(n6050), .ZN(n4995) );
  INV_X1 U5644 ( .A(n6049), .ZN(n4994) );
  NOR2_X1 U5645 ( .A1(n7296), .A2(n4883), .ZN(n4753) );
  NOR2_X1 U5646 ( .A1(n7298), .A2(n4750), .ZN(n4749) );
  OAI21_X1 U5647 ( .B1(n4649), .B2(n7520), .A(n7519), .ZN(n4648) );
  NAND2_X1 U5648 ( .A1(n4862), .A2(n4367), .ZN(n4861) );
  INV_X1 U5649 ( .A(n8928), .ZN(n4574) );
  NOR2_X1 U5650 ( .A1(n8339), .A2(n5481), .ZN(n4874) );
  OR2_X1 U5651 ( .A1(n8986), .A2(n8985), .ZN(n8987) );
  INV_X1 U5652 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4766) );
  INV_X1 U5653 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5130) );
  AND2_X1 U5654 ( .A1(n5129), .A2(n5128), .ZN(n5530) );
  INV_X1 U5655 ( .A(n5531), .ZN(n5129) );
  NOR2_X1 U5656 ( .A1(n5482), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4762) );
  AND2_X1 U5657 ( .A1(n5123), .A2(n5122), .ZN(n5389) );
  INV_X1 U5658 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5122) );
  OAI21_X1 U5659 ( .B1(n5293), .B2(n5847), .A(n5848), .ZN(n7430) );
  OR2_X1 U5660 ( .A1(n5757), .A2(n5770), .ZN(n6157) );
  NAND2_X1 U5661 ( .A1(n8800), .A2(n9425), .ZN(n6004) );
  INV_X1 U5662 ( .A(n5041), .ZN(n5040) );
  INV_X1 U5663 ( .A(n4999), .ZN(n4998) );
  NAND2_X1 U5664 ( .A1(n5036), .A2(n5432), .ZN(n7761) );
  INV_X1 U5665 ( .A(n5849), .ZN(n5029) );
  NAND2_X1 U5666 ( .A1(n5262), .A2(n4517), .ZN(n4516) );
  NOR2_X1 U5667 ( .A1(n5261), .A2(n5153), .ZN(n4517) );
  INV_X1 U5668 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U5669 ( .A1(n4606), .A2(n4605), .ZN(n5455) );
  INV_X1 U5670 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4605) );
  NOR2_X1 U5671 ( .A1(n5422), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5672 ( .A1(n5367), .A2(n5567), .ZN(n5381) );
  NOR2_X1 U5673 ( .A1(n6420), .A2(n6419), .ZN(n4620) );
  AND2_X1 U5674 ( .A1(n6266), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6253) );
  XNOR2_X1 U5675 ( .A(n6892), .B(n6849), .ZN(n6895) );
  INV_X1 U5676 ( .A(n8627), .ZN(n8712) );
  NOR2_X1 U5677 ( .A1(n8579), .A2(n8578), .ZN(n4832) );
  NOR2_X1 U5678 ( .A1(n9865), .A2(n8665), .ZN(n4928) );
  NOR2_X1 U5679 ( .A1(n6691), .A2(n5075), .ZN(n5074) );
  INV_X1 U5680 ( .A(n6689), .ZN(n5075) );
  NOR2_X1 U5681 ( .A1(n6550), .A2(n9529), .ZN(n4503) );
  INV_X1 U5682 ( .A(n4508), .ZN(n6527) );
  NAND2_X1 U5683 ( .A1(n10037), .A2(n4895), .ZN(n4894) );
  NOR2_X1 U5684 ( .A1(n6460), .A2(n6459), .ZN(n6469) );
  NOR2_X1 U5685 ( .A1(n6487), .A2(n6486), .ZN(n4621) );
  NOR2_X1 U5686 ( .A1(n4896), .A2(n10178), .ZN(n4895) );
  NAND2_X1 U5687 ( .A1(n10063), .A2(n6669), .ZN(n4496) );
  NAND2_X1 U5688 ( .A1(n6694), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U5689 ( .A1(n4620), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6451) );
  INV_X1 U5690 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6419) );
  INV_X1 U5691 ( .A(n4620), .ZN(n6437) );
  INV_X1 U5692 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U5693 ( .A1(n4505), .A2(n4356), .ZN(n6405) );
  AND3_X1 U5694 ( .A1(n6342), .A2(P1_REG3_REG_5__SCAN_IN), .A3(
        P1_REG3_REG_6__SCAN_IN), .ZN(n6278) );
  AND2_X1 U5695 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6342) );
  NOR2_X1 U5696 ( .A1(n6808), .A2(n9567), .ZN(n7483) );
  OAI21_X1 U5697 ( .B1(n9969), .B2(n4791), .A(n4788), .ZN(n5094) );
  NOR2_X2 U5698 ( .A1(n8094), .A2(n10204), .ZN(n8280) );
  NAND2_X1 U5699 ( .A1(n5833), .A2(n5829), .ZN(n5944) );
  AND2_X1 U5700 ( .A1(n5653), .A2(n5259), .ZN(n5655) );
  AND2_X1 U5701 ( .A1(n5273), .A2(n5274), .ZN(n5650) );
  NAND2_X1 U5702 ( .A1(n5242), .A2(n5241), .ZN(n4952) );
  NOR2_X1 U5703 ( .A1(n5605), .A2(n4936), .ZN(n4935) );
  INV_X1 U5704 ( .A(n5234), .ZN(n4936) );
  NAND2_X1 U5705 ( .A1(n6432), .A2(n4923), .ZN(n6626) );
  NOR2_X1 U5706 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4923) );
  AOI21_X1 U5707 ( .B1(n4945), .B2(n5471), .A(n4534), .ZN(n4942) );
  INV_X1 U5708 ( .A(n5208), .ZN(n4534) );
  INV_X1 U5709 ( .A(n4798), .ZN(n4793) );
  NAND2_X1 U5710 ( .A1(n4797), .A2(n4945), .ZN(n4796) );
  NAND2_X1 U5711 ( .A1(n4798), .A2(n4799), .ZN(n4797) );
  NAND2_X1 U5712 ( .A1(n4720), .A2(n4357), .ZN(n5448) );
  NAND2_X1 U5713 ( .A1(n5185), .A2(SI_5_), .ZN(n4725) );
  NAND2_X1 U5714 ( .A1(n7579), .A2(n7685), .ZN(n6077) );
  NAND2_X1 U5715 ( .A1(n4555), .A2(n6085), .ZN(n8030) );
  NAND2_X1 U5716 ( .A1(n5131), .A2(n8766), .ZN(n5618) );
  OR2_X1 U5717 ( .A1(n6063), .A2(n5292), .ZN(n6064) );
  XNOR2_X1 U5718 ( .A(n6137), .B(n6136), .ZN(n8827) );
  OR2_X1 U5719 ( .A1(n8827), .A2(n9193), .ZN(n4557) );
  NAND2_X1 U5720 ( .A1(n6086), .A2(n8158), .ZN(n8160) );
  NAND2_X1 U5721 ( .A1(n8030), .A2(n8157), .ZN(n6086) );
  NAND2_X1 U5722 ( .A1(n4566), .A2(n4564), .ZN(n6128) );
  AOI21_X1 U5723 ( .B1(n4567), .B2(n4569), .A(n4565), .ZN(n4564) );
  NAND2_X1 U5724 ( .A1(n6118), .A2(n4567), .ZN(n4566) );
  INV_X1 U5725 ( .A(n8904), .ZN(n8778) );
  XNOR2_X1 U5726 ( .A(n6148), .B(n10435), .ZN(n6080) );
  NAND2_X1 U5727 ( .A1(n6077), .A2(n7684), .ZN(n7687) );
  AND2_X1 U5728 ( .A1(n7080), .A2(n5776), .ZN(n6174) );
  AOI21_X1 U5729 ( .B1(n5968), .B2(n6152), .A(n5967), .ZN(n5974) );
  NAND2_X1 U5730 ( .A1(n9410), .A2(n9147), .ZN(n6051) );
  AND2_X1 U5731 ( .A1(n6051), .A2(n6053), .ZN(n4991) );
  NAND2_X1 U5732 ( .A1(n4470), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4468) );
  NOR2_X1 U5733 ( .A1(n7314), .A2(n7508), .ZN(n7313) );
  NAND2_X1 U5734 ( .A1(n4658), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4655) );
  OR2_X1 U5735 ( .A1(n5263), .A2(n10442), .ZN(n4656) );
  NOR2_X1 U5736 ( .A1(n7100), .A2(n7329), .ZN(n7101) );
  NAND2_X1 U5737 ( .A1(n4869), .A2(n7114), .ZN(n7332) );
  INV_X1 U5738 ( .A(n4870), .ZN(n4869) );
  INV_X1 U5739 ( .A(n4645), .ZN(n8937) );
  AOI21_X1 U5740 ( .B1(n7295), .B2(n7523), .A(n4648), .ZN(n4645) );
  NAND2_X1 U5741 ( .A1(n7809), .A2(n4864), .ZN(n4862) );
  AOI21_X1 U5742 ( .B1(n4291), .B2(n4643), .A(n4638), .ZN(n4637) );
  INV_X1 U5743 ( .A(n7830), .ZN(n4638) );
  NAND2_X1 U5744 ( .A1(n4880), .A2(n9008), .ZN(n9021) );
  NAND2_X1 U5745 ( .A1(n9002), .A2(n9001), .ZN(n9026) );
  NAND2_X1 U5746 ( .A1(n4626), .A2(n4625), .ZN(n9099) );
  AOI21_X1 U5747 ( .B1(n4312), .B2(n4630), .A(n4410), .ZN(n4625) );
  AND2_X1 U5748 ( .A1(n9097), .A2(n5111), .ZN(n4481) );
  NAND2_X1 U5749 ( .A1(n9069), .A2(n9082), .ZN(n9093) );
  NAND2_X1 U5750 ( .A1(n9070), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U5751 ( .A1(n4735), .A2(n4738), .ZN(n4734) );
  INV_X1 U5752 ( .A(n9093), .ZN(n4735) );
  AND2_X1 U5753 ( .A1(n4738), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U5754 ( .A1(n4524), .A2(n5810), .ZN(n4520) );
  INV_X1 U5755 ( .A(n4522), .ZN(n4521) );
  NAND2_X1 U5756 ( .A1(n5704), .A2(n5703), .ZN(n5721) );
  INV_X1 U5757 ( .A(n5705), .ZN(n5704) );
  NOR2_X1 U5758 ( .A1(n6201), .A2(n9298), .ZN(n6202) );
  NAND2_X1 U5759 ( .A1(n4763), .A2(n5132), .ZN(n5668) );
  INV_X1 U5760 ( .A(n4763), .ZN(n5267) );
  AND2_X1 U5761 ( .A1(n4768), .A2(n7862), .ZN(n4767) );
  NAND2_X1 U5762 ( .A1(n5131), .A2(n4768), .ZN(n5632) );
  NAND2_X1 U5763 ( .A1(n5031), .A2(n5030), .ZN(n9243) );
  NAND2_X1 U5764 ( .A1(n5798), .A2(n5002), .ZN(n5001) );
  INV_X1 U5765 ( .A(n9282), .ZN(n9274) );
  OAI21_X1 U5766 ( .B1(n9306), .B2(n6011), .A(n4350), .ZN(n9290) );
  NAND2_X1 U5767 ( .A1(n5515), .A2(n4311), .ZN(n5582) );
  NAND2_X1 U5768 ( .A1(n5515), .A2(n5130), .ZN(n5571) );
  NAND2_X1 U5769 ( .A1(n4762), .A2(n5127), .ZN(n5531) );
  INV_X1 U5770 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5127) );
  INV_X1 U5771 ( .A(n4762), .ZN(n5499) );
  OR2_X1 U5772 ( .A1(n5461), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U5773 ( .A1(n5126), .A2(n5125), .ZN(n5461) );
  INV_X1 U5774 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5125) );
  INV_X1 U5775 ( .A(n5438), .ZN(n5126) );
  NAND2_X1 U5776 ( .A1(n5389), .A2(n5124), .ZN(n5426) );
  INV_X1 U5777 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5124) );
  AOI21_X1 U5778 ( .B1(n7633), .B2(n5859), .A(n5792), .ZN(n7643) );
  AND2_X1 U5779 ( .A1(n7613), .A2(n5873), .ZN(n7648) );
  INV_X1 U5780 ( .A(SI_14_), .ZN(n7968) );
  NAND2_X1 U5781 ( .A1(n5856), .A2(n7461), .ZN(n7633) );
  NAND2_X1 U5782 ( .A1(n5120), .A2(n7549), .ZN(n5357) );
  NOR2_X1 U5783 ( .A1(n9147), .A2(n9146), .ZN(n9411) );
  AND2_X1 U5784 ( .A1(n6004), .A2(n6003), .ZN(n9170) );
  NOR2_X1 U5785 ( .A1(n9190), .A2(n8746), .ZN(n4511) );
  NAND2_X1 U5786 ( .A1(n5617), .A2(n5616), .ZN(n8835) );
  OR2_X1 U5787 ( .A1(n8315), .A2(n8316), .ZN(n9315) );
  INV_X1 U5788 ( .A(n7698), .ZN(n10435) );
  OR2_X1 U5789 ( .A1(n6154), .A2(n6153), .ZN(n6210) );
  AND2_X1 U5790 ( .A1(n6176), .A2(n6158), .ZN(n6213) );
  INV_X1 U5791 ( .A(n10426), .ZN(n10436) );
  INV_X1 U5792 ( .A(n5752), .ZN(n5753) );
  AND2_X1 U5793 ( .A1(n5731), .A2(n4316), .ZN(n5969) );
  AND2_X1 U5794 ( .A1(n5478), .A2(n4315), .ZN(n8331) );
  XNOR2_X1 U5795 ( .A(n5458), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U5796 ( .A1(n5409), .A2(n5384), .ZN(n5422) );
  NAND2_X1 U5797 ( .A1(n5366), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U5798 ( .A1(n4380), .A2(n4920), .ZN(n9514) );
  NAND2_X1 U5799 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  NAND2_X1 U5800 ( .A1(n4505), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U5801 ( .A1(n9594), .A2(n9595), .ZN(n9593) );
  NAND2_X1 U5802 ( .A1(n4620), .A2(n4491), .ZN(n6460) );
  NOR2_X1 U5803 ( .A1(n6450), .A2(n6436), .ZN(n4491) );
  INV_X1 U5804 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6459) );
  INV_X1 U5805 ( .A(n4684), .ZN(n4681) );
  NAND2_X1 U5806 ( .A1(n4680), .A2(n4684), .ZN(n4679) );
  INV_X1 U5807 ( .A(n4682), .ZN(n4680) );
  NAND2_X1 U5808 ( .A1(n6253), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6377) );
  INV_X1 U5809 ( .A(n7076), .ZN(n6807) );
  NOR2_X1 U5810 ( .A1(n9685), .A2(n6896), .ZN(n6897) );
  NAND2_X1 U5811 ( .A1(n4920), .A2(n4686), .ZN(n4685) );
  NAND2_X1 U5812 ( .A1(n9514), .A2(n6913), .ZN(n9603) );
  INV_X1 U5813 ( .A(n6802), .ZN(n8716) );
  AND2_X1 U5814 ( .A1(n6567), .A2(n6566), .ZN(n9915) );
  AND4_X1 U5815 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(n6364)
         );
  XNOR2_X1 U5816 ( .A(n9752), .B(n7799), .ZN(n9748) );
  NAND2_X1 U5817 ( .A1(n4616), .A2(n4615), .ZN(n7341) );
  INV_X1 U5818 ( .A(n7276), .ZN(n4615) );
  OR2_X1 U5819 ( .A1(n7349), .A2(n7350), .ZN(n7412) );
  NAND2_X1 U5820 ( .A1(n4428), .A2(n4427), .ZN(n7420) );
  INV_X1 U5821 ( .A(n7344), .ZN(n4427) );
  INV_X1 U5822 ( .A(n7343), .ZN(n4428) );
  NAND2_X1 U5823 ( .A1(n9822), .A2(n7422), .ZN(n7424) );
  OR2_X1 U5824 ( .A1(n7571), .A2(n7572), .ZN(n9850) );
  OR2_X1 U5825 ( .A1(n7424), .A2(n7423), .ZN(n7563) );
  AND2_X1 U5826 ( .A1(n10287), .A2(n10286), .ZN(n10289) );
  NAND2_X1 U5827 ( .A1(n9836), .A2(n9835), .ZN(n10283) );
  NOR2_X1 U5828 ( .A1(n10301), .A2(n9840), .ZN(n10311) );
  NAND2_X1 U5829 ( .A1(n8419), .A2(n8418), .ZN(n9868) );
  AND2_X1 U5830 ( .A1(n6624), .A2(n6623), .ZN(n7049) );
  NAND2_X1 U5831 ( .A1(n4317), .A2(n4544), .ZN(n4540) );
  NAND2_X1 U5832 ( .A1(n9903), .A2(n4317), .ZN(n4541) );
  AND2_X1 U5833 ( .A1(n6607), .A2(n6598), .ZN(n9509) );
  AND2_X1 U5834 ( .A1(n6614), .A2(n6613), .ZN(n8562) );
  OR2_X1 U5835 ( .A1(n9888), .A2(n6529), .ZN(n6614) );
  INV_X1 U5836 ( .A(n8624), .ZN(n8400) );
  NAND2_X1 U5837 ( .A1(n9924), .A2(n9902), .ZN(n9897) );
  NAND2_X1 U5838 ( .A1(n9945), .A2(n9954), .ZN(n9947) );
  AND2_X1 U5839 ( .A1(n6547), .A2(n6546), .ZN(n9983) );
  AND2_X1 U5840 ( .A1(n8640), .A2(n8543), .ZN(n9981) );
  NAND2_X1 U5841 ( .A1(n4384), .A2(n8461), .ZN(n5081) );
  NOR2_X2 U5842 ( .A1(n10002), .A2(n10231), .ZN(n9986) );
  NAND2_X1 U5843 ( .A1(n10018), .A2(n10019), .ZN(n10017) );
  NOR2_X1 U5844 ( .A1(n10092), .A2(n4894), .ZN(n10032) );
  INV_X1 U5845 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6486) );
  INV_X1 U5846 ( .A(n4621), .ZN(n6506) );
  AND2_X1 U5847 ( .A1(n6476), .A2(n6475), .ZN(n10030) );
  NAND2_X1 U5848 ( .A1(n4586), .A2(n6478), .ZN(n5085) );
  AND3_X1 U5849 ( .A1(n6464), .A2(n6463), .A3(n6462), .ZN(n10044) );
  CLKBUF_X1 U5850 ( .A(n10070), .Z(n4586) );
  NAND2_X1 U5851 ( .A1(n5088), .A2(n5090), .ZN(n5086) );
  NAND2_X1 U5852 ( .A1(n8091), .A2(n6668), .ZN(n8082) );
  NAND2_X1 U5853 ( .A1(n4547), .A2(n8677), .ZN(n8117) );
  NAND2_X1 U5854 ( .A1(n4779), .A2(n4351), .ZN(n8110) );
  NOR2_X1 U5855 ( .A1(n4576), .A2(n4575), .ZN(n4613) );
  NAND2_X1 U5856 ( .A1(n8110), .A2(n8595), .ZN(n8112) );
  AND2_X1 U5857 ( .A1(n7712), .A2(n4300), .ZN(n8184) );
  AND4_X1 U5858 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n8175)
         );
  AND2_X1 U5859 ( .A1(n8176), .A2(n6663), .ZN(n5115) );
  NAND2_X1 U5860 ( .A1(n7712), .A2(n4901), .ZN(n8185) );
  NAND2_X1 U5861 ( .A1(n7712), .A2(n8009), .ZN(n8054) );
  NAND2_X1 U5862 ( .A1(n6342), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U5863 ( .A1(n4438), .A2(n4348), .ZN(n7718) );
  NOR2_X1 U5864 ( .A1(n6808), .A2(n4439), .ZN(n4438) );
  NAND2_X1 U5865 ( .A1(n6328), .A2(n6340), .ZN(n4439) );
  NAND2_X1 U5866 ( .A1(n8466), .A2(n8668), .ZN(n8599) );
  NAND2_X1 U5867 ( .A1(n5067), .A2(n6684), .ZN(n9955) );
  NAND2_X1 U5868 ( .A1(n6682), .A2(n4320), .ZN(n5067) );
  AND3_X1 U5869 ( .A1(n6328), .A2(n6327), .A3(n6329), .ZN(n8016) );
  NAND2_X1 U5870 ( .A1(n7134), .A2(n7131), .ZN(n6313) );
  OAI211_X1 U5871 ( .C1(n5991), .C2(n5990), .A(n5989), .B(n5988), .ZN(n8433)
         );
  AND2_X1 U5872 ( .A1(n7868), .A2(n6235), .ZN(n5079) );
  INV_X1 U5873 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6235) );
  XNOR2_X1 U5874 ( .A(n5979), .B(n5952), .ZN(n8415) );
  NAND2_X1 U5875 ( .A1(n5694), .A2(n5693), .ZN(n5715) );
  XNOR2_X1 U5876 ( .A(n5681), .B(n5680), .ZN(n9498) );
  INV_X1 U5877 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6707) );
  INV_X1 U5878 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6631) );
  INV_X1 U5879 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6636) );
  NOR2_X1 U5880 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6628) );
  NOR2_X1 U5881 ( .A1(n5227), .A2(SI_17_), .ZN(n5228) );
  NAND2_X1 U5882 ( .A1(n6432), .A2(n6446), .ZN(n6465) );
  NAND2_X1 U5883 ( .A1(n5540), .A2(n5218), .ZN(n5509) );
  INV_X1 U5884 ( .A(n6432), .ZN(n6703) );
  NAND2_X1 U5885 ( .A1(n4945), .A2(n4947), .ZN(n5495) );
  NAND2_X1 U5886 ( .A1(n4947), .A2(n4944), .ZN(n5493) );
  NAND2_X1 U5887 ( .A1(n5408), .A2(n5375), .ZN(n5379) );
  OR2_X1 U5888 ( .A1(n6287), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U5889 ( .A1(n4724), .A2(n4726), .ZN(n5406) );
  NAND2_X1 U5890 ( .A1(n4963), .A2(n4962), .ZN(n7067) );
  AOI21_X1 U5891 ( .B1(n4966), .B2(n6144), .A(n4297), .ZN(n4962) );
  NAND2_X1 U5892 ( .A1(n4965), .A2(n4347), .ZN(n6166) );
  NOR2_X1 U5893 ( .A1(n7066), .A2(n4297), .ZN(n4969) );
  AND2_X1 U5894 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NOR2_X1 U5895 ( .A1(n6162), .A2(n8898), .ZN(n6163) );
  INV_X1 U5896 ( .A(n9260), .ZN(n9297) );
  NAND2_X1 U5897 ( .A1(n7543), .A2(n6072), .ZN(n7582) );
  AND2_X1 U5898 ( .A1(n8160), .A2(n6090), .ZN(n8265) );
  NAND2_X1 U5899 ( .A1(n8160), .A2(n4974), .ZN(n8263) );
  AND2_X1 U5900 ( .A1(n6215), .A2(n6184), .ZN(n8902) );
  AND2_X1 U5901 ( .A1(n8785), .A2(n6096), .ZN(n4607) );
  NAND2_X1 U5902 ( .A1(n8775), .A2(n6132), .ZN(n8859) );
  NAND2_X1 U5903 ( .A1(n7381), .A2(n7382), .ZN(n7380) );
  NAND2_X1 U5904 ( .A1(n8821), .A2(n8879), .ZN(n4955) );
  AND2_X1 U5905 ( .A1(n7687), .A2(n6079), .ZN(n7697) );
  NAND2_X1 U5906 ( .A1(n7687), .A2(n4978), .ZN(n7695) );
  INV_X1 U5907 ( .A(n8735), .ZN(n4563) );
  NAND2_X1 U5908 ( .A1(n8735), .A2(n4562), .ZN(n4561) );
  NAND2_X1 U5909 ( .A1(n8736), .A2(n6107), .ZN(n8900) );
  XNOR2_X1 U5910 ( .A(n5729), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U5911 ( .A1(n4987), .A2(n9130), .ZN(n4986) );
  INV_X1 U5912 ( .A(n4992), .ZN(n4987) );
  AOI21_X1 U5913 ( .B1(n4992), .B2(n4991), .A(n4989), .ZN(n4988) );
  NOR2_X1 U5914 ( .A1(n6051), .A2(n6053), .ZN(n4989) );
  INV_X1 U5915 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7195) );
  AND3_X1 U5916 ( .A1(n5586), .A2(n5585), .A3(n5584), .ZN(n8812) );
  OR2_X1 U5917 ( .A1(n5335), .A2(n5396), .ZN(n5404) );
  OR2_X1 U5918 ( .A1(n5335), .A2(n7595), .ZN(n5317) );
  OR2_X1 U5919 ( .A1(n5356), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5319) );
  OR2_X1 U5920 ( .A1(n5958), .A2(n5316), .ZN(n5320) );
  CLKBUF_X1 U5921 ( .A(n6067), .Z(n8924) );
  CLKBUF_X1 U5922 ( .A(n5312), .Z(n8925) );
  OR2_X1 U5923 ( .A1(n7080), .A2(n7078), .ZN(n9103) );
  NAND2_X1 U5924 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5288) );
  NAND2_X1 U5925 ( .A1(n4866), .A2(n7304), .ZN(n7213) );
  AOI21_X1 U5926 ( .B1(n7299), .B2(n7297), .A(n7298), .ZN(n7526) );
  AND2_X1 U5927 ( .A1(n7512), .A2(n7532), .ZN(n7513) );
  OAI21_X1 U5928 ( .B1(n8930), .B2(n8929), .A(n8928), .ZN(n8932) );
  NAND2_X1 U5929 ( .A1(n4640), .A2(n4639), .ZN(n8939) );
  NAND2_X1 U5930 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5931 ( .A1(n4863), .A2(n4862), .ZN(n8944) );
  NAND2_X1 U5932 ( .A1(n4892), .A2(n8951), .ZN(n7816) );
  AOI21_X1 U5933 ( .B1(n8337), .B2(n8338), .A(n8339), .ZN(n8971) );
  OR2_X1 U5934 ( .A1(n8973), .A2(n8999), .ZN(n8974) );
  NAND2_X1 U5935 ( .A1(n9009), .A2(n4881), .ZN(n8991) );
  NAND2_X1 U5936 ( .A1(n4507), .A2(n4857), .ZN(n4854) );
  NAND2_X1 U5937 ( .A1(n4628), .A2(n4629), .ZN(n9080) );
  OR2_X1 U5938 ( .A1(n9002), .A2(n4630), .ZN(n4628) );
  NAND2_X1 U5939 ( .A1(n4733), .A2(n4734), .ZN(n9121) );
  NAND2_X1 U5940 ( .A1(n5046), .A2(n5047), .ZN(n9212) );
  NAND2_X1 U5941 ( .A1(n5034), .A2(n5033), .ZN(n9258) );
  AND2_X1 U5942 ( .A1(n5529), .A2(n5528), .ZN(n8368) );
  AND2_X1 U5943 ( .A1(n5010), .A2(n5871), .ZN(n8025) );
  INV_X1 U5944 ( .A(n9283), .ZN(n9344) );
  OR2_X1 U5945 ( .A1(n10434), .A2(n5816), .ZN(n9337) );
  AND2_X1 U5946 ( .A1(n10411), .A2(n10421), .ZN(n9283) );
  NAND2_X1 U5947 ( .A1(n5783), .A2(n5782), .ZN(n7625) );
  INV_X1 U5948 ( .A(n10434), .ZN(n9394) );
  INV_X1 U5949 ( .A(n10417), .ZN(n9341) );
  AND2_X1 U5950 ( .A1(n9404), .A2(n10426), .ZN(n9407) );
  NAND2_X1 U5951 ( .A1(n9160), .A2(n5810), .ZN(n6045) );
  NAND2_X1 U5952 ( .A1(n5740), .A2(n5739), .ZN(n5741) );
  NAND2_X1 U5953 ( .A1(n8912), .A2(n9333), .ZN(n5740) );
  INV_X1 U5954 ( .A(n4597), .ZN(n9191) );
  INV_X1 U5955 ( .A(n6137), .ZN(n9443) );
  NAND2_X1 U5956 ( .A1(n5043), .A2(n5050), .ZN(n9203) );
  NAND2_X1 U5957 ( .A1(n5044), .A2(n5046), .ZN(n5043) );
  NAND2_X1 U5958 ( .A1(n9218), .A2(n5840), .ZN(n9202) );
  NAND2_X1 U5959 ( .A1(n9245), .A2(n5626), .ZN(n9224) );
  AOI22_X1 U5960 ( .A1(n9031), .A2(n4289), .B1(n5993), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U5961 ( .A1(n5012), .A2(n5017), .ZN(n9328) );
  NAND2_X1 U5962 ( .A1(n8297), .A2(n5016), .ZN(n5012) );
  INV_X1 U5963 ( .A(n8368), .ZN(n8854) );
  NAND2_X1 U5964 ( .A1(n5020), .A2(n5889), .ZN(n8323) );
  NAND2_X1 U5965 ( .A1(n5022), .A2(n5021), .ZN(n5020) );
  INV_X1 U5966 ( .A(n8297), .ZN(n5022) );
  NAND2_X1 U5967 ( .A1(n8196), .A2(n5491), .ZN(n8294) );
  INV_X1 U5968 ( .A(n9461), .ZN(n9485) );
  NAND2_X1 U5969 ( .A1(n5993), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4513) );
  AND2_X1 U5970 ( .A1(n7081), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8446) );
  INV_X1 U5971 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5151) );
  INV_X1 U5972 ( .A(n5155), .ZN(n8391) );
  INV_X1 U5973 ( .A(n5156), .ZN(n8390) );
  INV_X1 U5974 ( .A(n5756), .ZN(n9500) );
  INV_X1 U5975 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5748) );
  INV_X1 U5976 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9503) );
  INV_X1 U5977 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8305) );
  INV_X1 U5978 ( .A(n6054), .ZN(n8304) );
  INV_X1 U5979 ( .A(n5969), .ZN(n8225) );
  INV_X1 U5980 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7667) );
  INV_X1 U5981 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7183) );
  INV_X1 U5982 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7160) );
  NAND2_X1 U5983 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4877) );
  NAND2_X1 U5984 ( .A1(n5142), .A2(n5153), .ZN(n4876) );
  XNOR2_X1 U5985 ( .A(n6727), .B(n6726), .ZN(n7157) );
  INV_X1 U5986 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6726) );
  NAND2_X1 U5987 ( .A1(n6725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6727) );
  AND2_X1 U5988 ( .A1(n6591), .A2(n6590), .ZN(n9916) );
  NAND2_X1 U5989 ( .A1(n4920), .A2(n6913), .ZN(n9516) );
  NAND2_X1 U5990 ( .A1(n4921), .A2(n6966), .ZN(n9572) );
  AND2_X1 U5991 ( .A1(n6858), .A2(n6857), .ZN(n7772) );
  NAND2_X1 U5992 ( .A1(n4905), .A2(n4910), .ZN(n9617) );
  NAND2_X1 U5993 ( .A1(n9603), .A2(n6925), .ZN(n4905) );
  AND2_X1 U5994 ( .A1(n6557), .A2(n6556), .ZN(n9629) );
  NAND2_X1 U5995 ( .A1(n9624), .A2(n9623), .ZN(n4573) );
  NAND2_X1 U5996 ( .A1(n7000), .A2(n6999), .ZN(n9626) );
  OAI21_X1 U5997 ( .B1(n4921), .B2(n4681), .A(n4678), .ZN(n7000) );
  NAND2_X1 U5998 ( .A1(n4916), .A2(n7453), .ZN(n4673) );
  NAND2_X1 U5999 ( .A1(n6959), .A2(n6958), .ZN(n9649) );
  INV_X1 U6000 ( .A(n9705), .ZN(n9718) );
  AND2_X1 U6001 ( .A1(n6535), .A2(n6534), .ZN(n9996) );
  OR2_X1 U6002 ( .A1(n9989), .A2(n6529), .ZN(n6535) );
  AND2_X1 U6003 ( .A1(n6513), .A2(n6512), .ZN(n10031) );
  OR2_X1 U6004 ( .A1(n10013), .A2(n6529), .ZN(n6513) );
  AND2_X1 U6005 ( .A1(n6578), .A2(n6577), .ZN(n9707) );
  INV_X1 U6006 ( .A(n8562), .ZN(n9728) );
  INV_X1 U6007 ( .A(n8559), .ZN(n9906) );
  INV_X1 U6008 ( .A(n9916), .ZN(n9729) );
  INV_X1 U6009 ( .A(n9707), .ZN(n9932) );
  INV_X1 U6010 ( .A(n9629), .ZN(n9972) );
  INV_X1 U6011 ( .A(n9983), .ZN(n9730) );
  INV_X1 U6012 ( .A(n9982), .ZN(n10021) );
  INV_X1 U6013 ( .A(n10031), .ZN(n9731) );
  INV_X1 U6014 ( .A(n6364), .ZN(n9739) );
  NAND2_X1 U6015 ( .A1(n4430), .A2(n7267), .ZN(n9762) );
  NAND2_X1 U6016 ( .A1(n9774), .A2(n7270), .ZN(n9791) );
  NAND2_X1 U6017 ( .A1(n9791), .A2(n9792), .ZN(n9790) );
  NAND2_X1 U6018 ( .A1(n9803), .A2(n7273), .ZN(n9817) );
  NAND2_X1 U6019 ( .A1(n9817), .A2(n9818), .ZN(n9816) );
  OR2_X1 U6020 ( .A1(n7261), .A2(n7262), .ZN(n7347) );
  NAND2_X1 U6021 ( .A1(n9824), .A2(n9823), .ZN(n9822) );
  OR2_X1 U6022 ( .A1(n7415), .A2(n7416), .ZN(n7569) );
  XNOR2_X1 U6023 ( .A(n9839), .B(n9853), .ZN(n10303) );
  NOR2_X1 U6024 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  AOI21_X1 U6025 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10318), .A(n4329), .ZN(
        n10323) );
  INV_X1 U6026 ( .A(n10334), .ZN(n10329) );
  INV_X1 U6027 ( .A(n10297), .ZN(n10337) );
  OR2_X1 U6028 ( .A1(n10336), .A2(n10335), .ZN(n10345) );
  AOI21_X1 U6029 ( .B1(n6792), .B2(n9880), .A(n10091), .ZN(n6696) );
  NAND2_X1 U6030 ( .A1(n6688), .A2(n6687), .ZN(n9920) );
  NAND2_X1 U6031 ( .A1(n6682), .A2(n6681), .ZN(n9962) );
  NAND2_X1 U6032 ( .A1(n5058), .A2(n5055), .ZN(n10010) );
  INV_X1 U6033 ( .A(n5057), .ZN(n5055) );
  NAND2_X1 U6034 ( .A1(n6675), .A2(n6674), .ZN(n10026) );
  OAI21_X1 U6035 ( .B1(n8279), .B2(n4772), .A(n4771), .ZN(n10064) );
  NAND2_X1 U6036 ( .A1(n4774), .A2(n5061), .ZN(n10080) );
  NAND2_X1 U6037 ( .A1(n8279), .A2(n5062), .ZN(n4774) );
  NAND2_X1 U6038 ( .A1(n8277), .A2(n6670), .ZN(n8363) );
  NAND2_X1 U6039 ( .A1(n8273), .A2(n8685), .ZN(n8356) );
  NAND2_X1 U6040 ( .A1(n4546), .A2(n5095), .ZN(n8077) );
  NAND2_X1 U6041 ( .A1(n8115), .A2(n8503), .ZN(n8088) );
  NAND2_X1 U6042 ( .A1(n8143), .A2(n8151), .ZN(n8145) );
  NAND2_X1 U6043 ( .A1(n8172), .A2(n6666), .ZN(n8143) );
  NAND2_X1 U6044 ( .A1(n7045), .A2(n7162), .ZN(n10379) );
  NOR2_X1 U6045 ( .A1(n10091), .A2(n8590), .ZN(n7045) );
  INV_X1 U6046 ( .A(n9921), .ZN(n10222) );
  OAI21_X1 U6047 ( .B1(n10141), .B2(n10401), .A(n10140), .ZN(n4664) );
  OR3_X1 U6048 ( .A1(n10166), .A2(n10165), .A3(n10164), .ZN(n10234) );
  OR3_X1 U6049 ( .A1(n10184), .A2(n10183), .A3(n10182), .ZN(n10237) );
  AOI22_X1 U6050 ( .A1(n6593), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7155), .B2(
        n10273), .ZN(n4548) );
  NAND2_X1 U6051 ( .A1(n6592), .A2(n7138), .ZN(n5054) );
  AND2_X1 U6052 ( .A1(n6341), .A2(n6340), .ZN(n4434) );
  INV_X1 U6053 ( .A(n10389), .ZN(n10390) );
  AND2_X1 U6054 ( .A1(n7162), .A2(n7161), .ZN(n10389) );
  INV_X1 U6055 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8438) );
  NOR2_X1 U6056 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  NOR2_X1 U6057 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4670) );
  NAND2_X1 U6058 ( .A1(n6236), .A2(n4331), .ZN(n4536) );
  NOR2_X1 U6059 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4537) );
  NOR2_X1 U6060 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4539) );
  NAND2_X1 U6061 ( .A1(n6712), .A2(n6711), .ZN(n10263) );
  INV_X1 U6062 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10260) );
  INV_X1 U6063 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8394) );
  AND2_X1 U6064 ( .A1(n6372), .A2(n6385), .ZN(n7418) );
  AND2_X1 U6065 ( .A1(n6263), .A2(n6262), .ZN(n9812) );
  NAND2_X1 U6066 ( .A1(n4281), .A2(P1_U3086), .ZN(n10259) );
  XNOR2_X1 U6067 ( .A(n4432), .B(n4431), .ZN(n9752) );
  INV_X1 U6068 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4431) );
  NOR2_X1 U6069 ( .A1(n6634), .A2(n4433), .ZN(n4432) );
  INV_X1 U6070 ( .A(n4609), .ZN(n4608) );
  NAND2_X1 U6071 ( .A1(n4558), .A2(n8882), .ZN(n4610) );
  OAI21_X1 U6072 ( .B1(n9190), .B2(n8909), .A(n8834), .ZN(n4609) );
  NAND2_X1 U6073 ( .A1(n4888), .A2(n9046), .ZN(n9025) );
  AND2_X1 U6074 ( .A1(n4651), .A2(n4654), .ZN(n4593) );
  NAND2_X1 U6075 ( .A1(n4592), .A2(n8350), .ZN(n4591) );
  NOR2_X1 U6076 ( .A1(n5107), .A2(n6771), .ZN(n6772) );
  NOR2_X1 U6077 ( .A1(n5109), .A2(n6776), .ZN(n6777) );
  OAI22_X1 U6078 ( .A1(n9356), .A2(n9461), .B1(n10440), .B2(n6219), .ZN(n6220)
         );
  NAND2_X1 U6079 ( .A1(n4917), .A2(n6830), .ZN(n7454) );
  NAND2_X1 U6080 ( .A1(n7041), .A2(n4330), .ZN(n7064) );
  MUX2_X1 U6081 ( .A(n8590), .B(n8586), .S(n8627), .Z(n8728) );
  INV_X1 U6082 ( .A(n4618), .ZN(n4617) );
  NAND2_X1 U6083 ( .A1(n4426), .A2(n8590), .ZN(n4425) );
  AND2_X1 U6084 ( .A1(n6782), .A2(n9874), .ZN(n9894) );
  NOR2_X1 U6085 ( .A1(n10131), .A2(n10361), .ZN(n9907) );
  NAND2_X1 U6086 ( .A1(n9944), .A2(n4665), .ZN(P1_U3269) );
  NAND2_X1 U6087 ( .A1(n4666), .A2(n10386), .ZN(n4665) );
  NAND2_X1 U6088 ( .A1(n4535), .A2(n10408), .ZN(n6733) );
  OAI21_X1 U6089 ( .B1(n6798), .B2(n6794), .A(n6795), .ZN(n6797) );
  AOI21_X1 U6090 ( .B1(n10127), .B2(n10159), .A(n4411), .ZN(n4780) );
  NAND2_X1 U6091 ( .A1(n4535), .A2(n10405), .ZN(n6737) );
  OAI21_X1 U6092 ( .B1(n6798), .B2(n10403), .A(n6799), .ZN(n6801) );
  AOI21_X1 U6093 ( .B1(n10127), .B2(n10232), .A(n4412), .ZN(n4782) );
  INV_X1 U6094 ( .A(n9567), .ZN(n4437) );
  INV_X1 U6095 ( .A(n6015), .ZN(n7465) );
  INV_X1 U6096 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6634) );
  INV_X1 U6097 ( .A(n6821), .ZN(n6930) );
  INV_X2 U6098 ( .A(n6930), .ZN(n7015) );
  OR2_X1 U6099 ( .A1(n8975), .A2(n8976), .ZN(n4857) );
  INV_X1 U6100 ( .A(n7826), .ZN(n4860) );
  AND2_X1 U6101 ( .A1(n5489), .A2(n5795), .ZN(n8200) );
  AND2_X1 U6102 ( .A1(n4639), .A2(n7825), .ZN(n4291) );
  NAND2_X1 U6103 ( .A1(n4692), .A2(n4408), .ZN(n9584) );
  INV_X1 U6104 ( .A(n8922), .ZN(n4514) );
  AND2_X1 U6105 ( .A1(n5919), .A2(n7082), .ZN(n4292) );
  AND4_X2 U6106 ( .A1(n4848), .A2(n5149), .A3(n4402), .A4(n5305), .ZN(n4293)
         );
  AND4_X1 U6107 ( .A1(n8713), .A2(n9875), .A3(n8628), .A4(n8627), .ZN(n4294)
         );
  AND3_X1 U6108 ( .A1(n9035), .A2(n9060), .A3(P2_REG1_REG_15__SCAN_IN), .ZN(
        n4295) );
  INV_X1 U6109 ( .A(n5840), .ZN(n5006) );
  NAND2_X1 U6110 ( .A1(n5085), .A2(n8533), .ZN(n10027) );
  AND2_X1 U6111 ( .A1(n8490), .A2(n4285), .ZN(n4296) );
  AND2_X1 U6112 ( .A1(n4970), .A2(n8800), .ZN(n4297) );
  AND2_X1 U6113 ( .A1(n4319), .A2(n5032), .ZN(n4298) );
  AND2_X1 U6114 ( .A1(n4456), .A2(n4903), .ZN(n4299) );
  AND2_X1 U6115 ( .A1(n4901), .A2(n8188), .ZN(n4300) );
  AND2_X1 U6116 ( .A1(n5300), .A2(n5287), .ZN(n7134) );
  AND2_X1 U6117 ( .A1(n5079), .A2(n6246), .ZN(n4301) );
  AND2_X1 U6118 ( .A1(n4948), .A2(n4525), .ZN(n4302) );
  AND2_X1 U6119 ( .A1(n6080), .A2(n8921), .ZN(n4303) );
  NAND2_X1 U6120 ( .A1(n9329), .A2(n4395), .ZN(n4304) );
  AND2_X1 U6121 ( .A1(n8549), .A2(n8548), .ZN(n9971) );
  AND3_X1 U6122 ( .A1(n4372), .A2(n6329), .A3(n6341), .ZN(n4305) );
  AND2_X1 U6123 ( .A1(n5030), .A2(n5625), .ZN(n4306) );
  AND3_X1 U6124 ( .A1(n4818), .A2(n4392), .A3(n9971), .ZN(n4307) );
  OR2_X1 U6125 ( .A1(n6685), .A2(n5071), .ZN(n4308) );
  OR2_X1 U6126 ( .A1(n4973), .A2(n4554), .ZN(n4309) );
  NAND2_X1 U6127 ( .A1(n6270), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4310) );
  AND2_X1 U6128 ( .A1(n5130), .A2(n4766), .ZN(n4311) );
  AND2_X1 U6129 ( .A1(n4629), .A2(n4627), .ZN(n4312) );
  INV_X1 U6130 ( .A(n8879), .ZN(n4958) );
  AND2_X1 U6131 ( .A1(n5237), .A2(n5236), .ZN(n4313) );
  NAND2_X1 U6132 ( .A1(n9031), .A2(n4635), .ZN(n4634) );
  AND2_X1 U6133 ( .A1(n9061), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U6134 ( .A1(n8281), .A2(n8362), .ZN(n10092) );
  OR2_X1 U6135 ( .A1(n4550), .A2(n4980), .ZN(n4316) );
  INV_X1 U6136 ( .A(n4507), .ZN(n9017) );
  NAND2_X1 U6137 ( .A1(n8973), .A2(n8999), .ZN(n4507) );
  NAND2_X1 U6138 ( .A1(n5414), .A2(n5413), .ZN(n7698) );
  NAND2_X2 U6139 ( .A1(n5155), .A2(n8390), .ZN(n5335) );
  INV_X1 U6140 ( .A(n8339), .ZN(n4875) );
  AND2_X1 U6141 ( .A1(n8624), .A2(n4542), .ZN(n4317) );
  NAND2_X1 U6142 ( .A1(n10017), .A2(n8696), .ZN(n8638) );
  XNOR2_X1 U6143 ( .A(n5385), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U6144 ( .A1(n5031), .A2(n4306), .ZN(n9245) );
  INV_X1 U6145 ( .A(n6617), .ZN(n6418) );
  NAND4_X1 U6146 ( .A1(n5320), .A2(n5319), .A3(n5318), .A4(n5317), .ZN(n5334)
         );
  NAND2_X1 U6147 ( .A1(n4886), .A2(n9046), .ZN(n9047) );
  INV_X1 U6148 ( .A(n4857), .ZN(n9015) );
  OAI21_X1 U6149 ( .B1(n6118), .B2(n4569), .A(n4567), .ZN(n8764) );
  AND2_X1 U6150 ( .A1(n4955), .A2(n8880), .ZN(n4318) );
  OR2_X1 U6151 ( .A1(n9281), .A2(n9260), .ZN(n4319) );
  NOR2_X1 U6152 ( .A1(n6683), .A2(n5072), .ZN(n4320) );
  AND2_X1 U6153 ( .A1(n6076), .A2(n6072), .ZN(n4321) );
  NAND2_X1 U6154 ( .A1(n5711), .A2(n5710), .ZN(n9172) );
  NAND2_X1 U6155 ( .A1(n6605), .A2(n6604), .ZN(n9890) );
  OR2_X1 U6156 ( .A1(n5796), .A2(n5019), .ZN(n4322) );
  AND2_X1 U6157 ( .A1(n8528), .A2(n10040), .ZN(n10072) );
  NAND2_X1 U6158 ( .A1(n4510), .A2(n5587), .ZN(n9273) );
  NAND3_X1 U6159 ( .A1(n9233), .A2(n9231), .A3(n9232), .ZN(n4323) );
  AND3_X1 U6160 ( .A1(n4848), .A2(n4847), .A3(n5305), .ZN(n4324) );
  AND2_X1 U6161 ( .A1(n4725), .A2(n4786), .ZN(n4325) );
  AND2_X1 U6162 ( .A1(n4835), .A2(n5904), .ZN(n4326) );
  AOI21_X1 U6163 ( .B1(n9498), .B2(n5365), .A(n5112), .ZN(n6145) );
  INV_X1 U6164 ( .A(n6145), .ZN(n9425) );
  OR2_X1 U6165 ( .A1(n10040), .A2(n4285), .ZN(n4327) );
  AND2_X1 U6166 ( .A1(n4864), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4328) );
  AND2_X1 U6167 ( .A1(n8550), .A2(n9929), .ZN(n9954) );
  INV_X1 U6168 ( .A(n9954), .ZN(n4791) );
  NOR2_X1 U6169 ( .A1(n10311), .A2(n10310), .ZN(n4329) );
  AND3_X1 U6170 ( .A1(n7060), .A2(n7059), .A3(n9672), .ZN(n4330) );
  AND2_X1 U6171 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4331) );
  AND2_X1 U6172 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4332) );
  XNOR2_X1 U6173 ( .A(n5368), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7288) );
  AND2_X1 U6174 ( .A1(n6137), .A2(n9214), .ZN(n4333) );
  OR2_X1 U6175 ( .A1(n8166), .A2(n8919), .ZN(n4334) );
  AND2_X1 U6176 ( .A1(n10040), .A2(n8522), .ZN(n4335) );
  AND2_X1 U6177 ( .A1(n5418), .A2(n4334), .ZN(n4336) );
  NAND2_X1 U6178 ( .A1(n5094), .A2(n8632), .ZN(n9910) );
  OR2_X1 U6179 ( .A1(n9897), .A2(n10127), .ZN(n4337) );
  AND2_X1 U6180 ( .A1(n4854), .A2(n9016), .ZN(n4338) );
  NOR2_X1 U6181 ( .A1(n6047), .A2(n6046), .ZN(n4339) );
  NAND2_X1 U6182 ( .A1(n8654), .A2(n8707), .ZN(n8593) );
  AND3_X1 U6183 ( .A1(n8585), .A2(n8584), .A3(n8713), .ZN(n4340) );
  XNOR2_X1 U6184 ( .A(n6738), .B(n6752), .ZN(n6759) );
  AND2_X1 U6185 ( .A1(n5034), .A2(n4319), .ZN(n9257) );
  AND2_X1 U6186 ( .A1(n10226), .A2(n9972), .ZN(n4341) );
  INV_X1 U6187 ( .A(n4945), .ZN(n4943) );
  NOR2_X1 U6188 ( .A1(n5492), .A2(n4946), .ZN(n4945) );
  AND2_X1 U6189 ( .A1(n8710), .A2(n8706), .ZN(n4342) );
  NOR2_X1 U6190 ( .A1(n10168), .A2(n9731), .ZN(n4343) );
  AND2_X1 U6191 ( .A1(n8596), .A2(n5097), .ZN(n4344) );
  AND2_X1 U6192 ( .A1(n5041), .A2(n5049), .ZN(n4345) );
  AND3_X1 U6193 ( .A1(n4513), .A2(n5369), .A3(n5370), .ZN(n7852) );
  INV_X1 U6194 ( .A(n7852), .ZN(n4512) );
  NAND2_X1 U6195 ( .A1(n9242), .A2(n9232), .ZN(n4346) );
  INV_X1 U6196 ( .A(n5084), .ZN(n5083) );
  NAND2_X1 U6197 ( .A1(n6494), .A2(n8533), .ZN(n5084) );
  AND2_X1 U6198 ( .A1(n4969), .A2(n4964), .ZN(n4347) );
  AND2_X1 U6199 ( .A1(n6291), .A2(n6290), .ZN(n8009) );
  INV_X1 U6200 ( .A(n8009), .ZN(n4902) );
  AND2_X1 U6201 ( .A1(n4437), .A2(n4305), .ZN(n4348) );
  OR2_X1 U6202 ( .A1(n5920), .A2(n7082), .ZN(n4349) );
  AOI21_X1 U6203 ( .B1(n4906), .B2(n4909), .A(n4904), .ZN(n4903) );
  OR2_X1 U6204 ( .A1(n8816), .A2(n9295), .ZN(n4350) );
  AND2_X1 U6205 ( .A1(n4778), .A2(n5065), .ZN(n4351) );
  INV_X1 U6206 ( .A(n4643), .ZN(n4641) );
  NAND2_X1 U6207 ( .A1(n4650), .A2(n4644), .ZN(n4643) );
  AND2_X1 U6208 ( .A1(n4770), .A2(n6004), .ZN(n4352) );
  AND2_X1 U6209 ( .A1(n4836), .A2(n4472), .ZN(n4353) );
  AND2_X1 U6210 ( .A1(n4918), .A2(n6870), .ZN(n4354) );
  AND2_X1 U6211 ( .A1(n9886), .A2(n9892), .ZN(n4355) );
  AND2_X1 U6212 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .ZN(n4356) );
  OR2_X1 U6213 ( .A1(n5197), .A2(SI_8_), .ZN(n4357) );
  INV_X1 U6214 ( .A(n5810), .ZN(n4523) );
  NAND2_X1 U6215 ( .A1(n9356), .A2(n9172), .ZN(n5810) );
  NAND2_X1 U6216 ( .A1(n4868), .A2(n4867), .ZN(n4358) );
  AND2_X1 U6217 ( .A1(n9233), .A2(n9234), .ZN(n9242) );
  AND2_X1 U6218 ( .A1(n9443), .A2(n9193), .ZN(n4359) );
  OR2_X1 U6219 ( .A1(n9471), .A2(n9295), .ZN(n5908) );
  AND2_X1 U6220 ( .A1(n6929), .A2(n6928), .ZN(n4360) );
  NAND2_X1 U6221 ( .A1(n7131), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4361) );
  AND2_X1 U6222 ( .A1(n8362), .A2(n9716), .ZN(n4362) );
  AND2_X1 U6223 ( .A1(n6137), .A2(n9193), .ZN(n6008) );
  AND2_X1 U6224 ( .A1(n5085), .A2(n5083), .ZN(n4363) );
  NOR2_X1 U6225 ( .A1(n6091), .A2(n8164), .ZN(n4364) );
  NOR2_X1 U6226 ( .A1(n10113), .A2(n9736), .ZN(n4365) );
  AND2_X1 U6227 ( .A1(n5837), .A2(n5836), .ZN(n4366) );
  INV_X1 U6228 ( .A(n4819), .ZN(n4818) );
  OR2_X1 U6229 ( .A1(n7821), .A2(n8106), .ZN(n4367) );
  NAND2_X1 U6230 ( .A1(n9484), .A2(n9316), .ZN(n4368) );
  INV_X1 U6231 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6446) );
  INV_X1 U6232 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6246) );
  AND2_X1 U6233 ( .A1(n9270), .A2(n9275), .ZN(n4369) );
  INV_X1 U6234 ( .A(n4950), .ZN(n4949) );
  OAI21_X1 U6235 ( .B1(n5217), .B2(n4951), .A(n5221), .ZN(n4950) );
  AND2_X1 U6236 ( .A1(n5966), .A2(n5940), .ZN(n4370) );
  AND3_X1 U6237 ( .A1(n6300), .A2(n6301), .A3(n4310), .ZN(n4371) );
  AND2_X1 U6238 ( .A1(n6339), .A2(n6327), .ZN(n4372) );
  OR2_X1 U6239 ( .A1(n4550), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4373) );
  AND2_X1 U6240 ( .A1(n5507), .A2(SI_15_), .ZN(n4374) );
  AND2_X1 U6241 ( .A1(n9971), .A2(n4817), .ZN(n4375) );
  AND2_X1 U6242 ( .A1(n4960), .A2(n4561), .ZN(n4376) );
  AND2_X1 U6243 ( .A1(n8790), .A2(n8873), .ZN(n4377) );
  INV_X1 U6244 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5261) );
  AND2_X1 U6245 ( .A1(n6649), .A2(n6648), .ZN(n4378) );
  INV_X1 U6246 ( .A(n5108), .ZN(n4524) );
  INV_X1 U6247 ( .A(n4694), .ZN(n6709) );
  NAND2_X1 U6248 ( .A1(n4696), .A2(n6432), .ZN(n4694) );
  INV_X1 U6249 ( .A(n9517), .ZN(n4919) );
  INV_X1 U6250 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7185) );
  AND2_X1 U6251 ( .A1(n6999), .A2(n7001), .ZN(n4379) );
  AND2_X1 U6252 ( .A1(n9416), .A2(n8911), .ZN(n6050) );
  AND2_X1 U6253 ( .A1(n6913), .A2(n4919), .ZN(n4380) );
  OR2_X1 U6254 ( .A1(n4308), .A2(n6680), .ZN(n4381) );
  AND2_X1 U6255 ( .A1(n5150), .A2(n5052), .ZN(n4382) );
  NAND2_X1 U6256 ( .A1(n5001), .A2(n5800), .ZN(n9229) );
  INV_X1 U6257 ( .A(n4974), .ZN(n4973) );
  AND2_X1 U6258 ( .A1(n8264), .A2(n6090), .ZN(n4974) );
  INV_X1 U6259 ( .A(n4884), .ZN(n4883) );
  NAND2_X1 U6260 ( .A1(n7527), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4884) );
  INV_X1 U6261 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5142) );
  OR2_X1 U6262 ( .A1(n10092), .A2(n4896), .ZN(n4383) );
  OR2_X1 U6263 ( .A1(n8619), .A2(n5082), .ZN(n4384) );
  OR2_X1 U6264 ( .A1(n10190), .A2(n10073), .ZN(n4385) );
  OR2_X1 U6265 ( .A1(n4550), .A2(n4983), .ZN(n4386) );
  AND3_X1 U6266 ( .A1(n8569), .A2(n8568), .A3(n8570), .ZN(n4387) );
  AND2_X1 U6267 ( .A1(n4533), .A2(n6007), .ZN(n4388) );
  AND2_X1 U6268 ( .A1(n10019), .A2(n8461), .ZN(n4389) );
  INV_X1 U6269 ( .A(n8469), .ZN(n6653) );
  AND2_X1 U6270 ( .A1(n7131), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4390) );
  AOI21_X2 U6271 ( .B1(n7165), .B2(n6592), .A(n6265), .ZN(n8188) );
  AND2_X1 U6272 ( .A1(n5115), .A2(n4821), .ZN(n4391) );
  INV_X1 U6273 ( .A(n8746), .ZN(n9205) );
  AND2_X1 U6274 ( .A1(n5161), .A2(n5160), .ZN(n8746) );
  AND2_X1 U6275 ( .A1(n8546), .A2(n8544), .ZN(n4392) );
  AOI21_X1 U6276 ( .B1(n4908), .B2(n4910), .A(n4907), .ZN(n4906) );
  AND2_X1 U6277 ( .A1(n5920), .A2(n5802), .ZN(n4393) );
  AND2_X1 U6278 ( .A1(n5098), .A2(n8596), .ZN(n4394) );
  INV_X1 U6279 ( .A(n5063), .ZN(n5062) );
  OR2_X1 U6280 ( .A1(n4843), .A2(n5894), .ZN(n4395) );
  AND2_X1 U6281 ( .A1(n4300), .A2(n9645), .ZN(n4396) );
  AND2_X1 U6282 ( .A1(n5445), .A2(n5432), .ZN(n4397) );
  AND2_X1 U6283 ( .A1(n4328), .A2(n4860), .ZN(n4398) );
  INV_X1 U6284 ( .A(n8935), .ZN(n4650) );
  INV_X1 U6285 ( .A(n7760), .ZN(n5445) );
  AND2_X1 U6286 ( .A1(n5871), .A2(n5874), .ZN(n7760) );
  AND2_X1 U6287 ( .A1(n4775), .A2(n4726), .ZN(n4399) );
  OR2_X1 U6288 ( .A1(n9874), .A2(n6701), .ZN(n4400) );
  INV_X1 U6289 ( .A(n4760), .ZN(n4759) );
  OR2_X1 U6290 ( .A1(n7821), .A2(n7820), .ZN(n4760) );
  AND2_X1 U6291 ( .A1(n4379), .A2(n4675), .ZN(n4401) );
  AND2_X1 U6292 ( .A1(n4382), .A2(n5261), .ZN(n4402) );
  INV_X1 U6293 ( .A(n4800), .ZN(n4799) );
  AND2_X1 U6294 ( .A1(n5452), .A2(n4577), .ZN(n4800) );
  AND2_X1 U6295 ( .A1(n5205), .A2(n5451), .ZN(n4403) );
  NAND2_X1 U6296 ( .A1(n10190), .A2(n10073), .ZN(n4404) );
  NAND2_X1 U6297 ( .A1(n9647), .A2(n9646), .ZN(n4405) );
  INV_X1 U6298 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6292) );
  INV_X1 U6299 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U6300 ( .A1(n8199), .A2(n5795), .ZN(n8297) );
  OAI21_X1 U6301 ( .B1(n4555), .B2(n4309), .A(n4551), .ZN(n8750) );
  OAI21_X1 U6302 ( .B1(n8733), .B2(n4563), .A(n4376), .ZN(n8805) );
  AND2_X1 U6303 ( .A1(n8280), .A2(n9666), .ZN(n8281) );
  NAND2_X1 U6304 ( .A1(n7543), .A2(n4321), .ZN(n7579) );
  INV_X1 U6305 ( .A(n10127), .ZN(n4445) );
  NAND2_X1 U6306 ( .A1(n8591), .A2(n9865), .ZN(n8582) );
  INV_X1 U6307 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4433) );
  AND2_X1 U6308 ( .A1(n5658), .A2(n5675), .ZN(n4406) );
  OR2_X1 U6309 ( .A1(n10092), .A2(n10190), .ZN(n4407) );
  INV_X1 U6310 ( .A(n8836), .ZN(n4565) );
  NAND2_X1 U6311 ( .A1(n5793), .A2(n6012), .ZN(n7758) );
  INV_X1 U6312 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4984) );
  INV_X1 U6313 ( .A(n8762), .ZN(n4957) );
  NAND2_X1 U6314 ( .A1(n8112), .A2(n6667), .ZN(n8090) );
  INV_X1 U6315 ( .A(n8800), .ZN(n9181) );
  AND2_X1 U6316 ( .A1(n5689), .A2(n5688), .ZN(n8800) );
  AND2_X1 U6317 ( .A1(n4687), .A2(n6897), .ZN(n4408) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4583) );
  AND2_X1 U6319 ( .A1(n5249), .A2(n5244), .ZN(n4409) );
  NOR2_X1 U6320 ( .A1(n9078), .A2(n9077), .ZN(n4410) );
  NOR2_X1 U6321 ( .A1(n10408), .A2(n10126), .ZN(n4411) );
  NOR2_X1 U6322 ( .A1(n10405), .A2(n7909), .ZN(n4412) );
  AND2_X1 U6323 ( .A1(n9972), .A2(n10085), .ZN(n4413) );
  AND2_X1 U6324 ( .A1(n8972), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4414) );
  AND2_X1 U6325 ( .A1(n5240), .A2(n5239), .ZN(n4415) );
  NAND2_X1 U6326 ( .A1(n9055), .A2(n4631), .ZN(n4416) );
  OR2_X1 U6327 ( .A1(n4856), .A2(n8976), .ZN(n4417) );
  INV_X1 U6328 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4750) );
  INV_X1 U6329 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7862) );
  AND2_X1 U6330 ( .A1(n6217), .A2(n6216), .ZN(n10441) );
  NAND2_X1 U6331 ( .A1(n8052), .A2(n10212), .ZN(n10195) );
  INV_X1 U6332 ( .A(n9140), .ZN(n9042) );
  INV_X1 U6333 ( .A(n10190), .ZN(n4897) );
  INV_X1 U6334 ( .A(n7684), .ZN(n4976) );
  AND2_X1 U6335 ( .A1(n7483), .A2(n8016), .ZN(n4418) );
  INV_X1 U6336 ( .A(n8157), .ZN(n4554) );
  NAND2_X1 U6337 ( .A1(n6390), .A2(n6389), .ZN(n9690) );
  INV_X1 U6338 ( .A(n9690), .ZN(n4440) );
  NAND2_X1 U6339 ( .A1(n6101), .A2(n8789), .ZN(n8734) );
  INV_X1 U6340 ( .A(n8734), .ZN(n4562) );
  INV_X1 U6341 ( .A(n9097), .ZN(n9082) );
  AND2_X1 U6342 ( .A1(n7529), .A2(n7814), .ZN(n4419) );
  INV_X1 U6343 ( .A(n8882), .ZN(n8898) );
  NAND2_X1 U6344 ( .A1(n6161), .A2(n6160), .ZN(n8882) );
  INV_X1 U6345 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5121) );
  INV_X1 U6346 ( .A(n7134), .ZN(n5026) );
  INV_X1 U6347 ( .A(n9130), .ZN(n6053) );
  XOR2_X1 U6348 ( .A(n9130), .B(P2_REG2_REG_19__SCAN_IN), .Z(n4420) );
  INV_X1 U6349 ( .A(n8590), .ZN(n9865) );
  AND2_X1 U6350 ( .A1(n7112), .A2(n7114), .ZN(n4421) );
  AND2_X1 U6351 ( .A1(n7100), .A2(n7329), .ZN(n4744) );
  INV_X1 U6352 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4769) );
  INV_X1 U6353 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5025) );
  INV_X1 U6354 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4801) );
  INV_X1 U6355 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4580) );
  INV_X1 U6356 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n4602) );
  INV_X1 U6357 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n4612) );
  NAND3_X1 U6358 ( .A1(n4425), .A2(n4617), .A3(n4422), .ZN(P1_U3262) );
  NAND2_X1 U6359 ( .A1(n4423), .A2(n9865), .ZN(n4422) );
  NAND2_X1 U6360 ( .A1(n4424), .A2(n9864), .ZN(n4423) );
  NAND2_X1 U6361 ( .A1(n9863), .A2(n10329), .ZN(n4424) );
  OAI22_X1 U6362 ( .A1(n9863), .A2(n10334), .B1(n9862), .B2(n10297), .ZN(n4426) );
  NAND2_X1 U6363 ( .A1(n9775), .A2(n9776), .ZN(n9774) );
  INV_X1 U6364 ( .A(n7277), .ZN(n4616) );
  NAND2_X1 U6365 ( .A1(n4430), .A2(n4429), .ZN(n7373) );
  OR2_X1 U6366 ( .A1(n7367), .A2(n7368), .ZN(n4429) );
  NAND2_X1 U6367 ( .A1(n7563), .A2(n7562), .ZN(n7565) );
  OAI21_X2 U6368 ( .B1(n9978), .B2(n4381), .A(n5068), .ZN(n9941) );
  NAND3_X1 U6369 ( .A1(n7600), .A2(n7601), .A3(n8603), .ZN(n4435) );
  AND2_X2 U6370 ( .A1(n7721), .A2(n7775), .ZN(n7712) );
  NOR2_X2 U6371 ( .A1(n4446), .A2(n10092), .ZN(n10011) );
  NOR2_X1 U6372 ( .A1(n4449), .A2(n4539), .ZN(n4448) );
  NOR2_X1 U6373 ( .A1(n4451), .A2(n4537), .ZN(n4450) );
  NAND2_X1 U6374 ( .A1(n4453), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U6375 ( .A1(n6629), .A2(n5104), .ZN(n4453) );
  NAND2_X4 U6376 ( .A1(n4455), .A2(n4454), .ZN(n7004) );
  NAND3_X1 U6377 ( .A1(n6912), .A2(n6911), .A3(n4906), .ZN(n4456) );
  OR2_X2 U6378 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  OAI21_X1 U6379 ( .B1(n4844), .B2(n4459), .A(n6201), .ZN(n4458) );
  INV_X1 U6380 ( .A(n5940), .ZN(n4459) );
  NAND3_X1 U6381 ( .A1(n5939), .A2(n5934), .A3(n4845), .ZN(n4460) );
  OAI211_X1 U6382 ( .C1(n5855), .C2(n4467), .A(n4461), .B(n7465), .ZN(n5864)
         );
  NAND2_X1 U6383 ( .A1(n4466), .A2(n5853), .ZN(n4461) );
  NAND3_X1 U6384 ( .A1(n4464), .A2(n4462), .A3(n5863), .ZN(n4465) );
  NAND3_X1 U6385 ( .A1(n4467), .A2(n7465), .A3(n4463), .ZN(n4462) );
  NAND3_X1 U6386 ( .A1(n5855), .A2(n7465), .A3(n5861), .ZN(n4464) );
  INV_X1 U6387 ( .A(n5855), .ZN(n4466) );
  NAND3_X1 U6388 ( .A1(n4469), .A2(n4468), .A3(n5295), .ZN(n5786) );
  NAND4_X1 U6389 ( .A1(n4469), .A2(n4468), .A3(n7474), .A4(n5295), .ZN(n5847)
         );
  AND2_X1 U6390 ( .A1(n5297), .A2(n5296), .ZN(n4469) );
  NAND2_X1 U6391 ( .A1(n5907), .A2(n4589), .ZN(n5900) );
  OAI21_X1 U6392 ( .B1(n4349), .B2(n4478), .A(n4702), .ZN(n4477) );
  NAND2_X1 U6393 ( .A1(n4841), .A2(n4840), .ZN(n4479) );
  AND3_X2 U6394 ( .A1(n4848), .A2(n5149), .A3(n5305), .ZN(n4624) );
  OR2_X1 U6395 ( .A1(n4624), .A2(n5153), .ZN(n5751) );
  NAND3_X1 U6396 ( .A1(n4480), .A2(n6664), .A3(n8151), .ZN(n4778) );
  NAND3_X1 U6397 ( .A1(n9035), .A2(n9060), .A3(n4314), .ZN(n4867) );
  NAND3_X1 U6398 ( .A1(n4868), .A2(n4867), .A3(n5111), .ZN(n9075) );
  NAND3_X1 U6399 ( .A1(n4868), .A2(n4867), .A3(n4481), .ZN(n4572) );
  MUX2_X1 U6400 ( .A(n5168), .B(n5167), .S(n4280), .Z(n4482) );
  INV_X1 U6401 ( .A(n6680), .ZN(n4487) );
  NAND3_X1 U6402 ( .A1(n4494), .A2(n4497), .A3(n6672), .ZN(n10050) );
  NAND2_X1 U6403 ( .A1(n8081), .A2(n6669), .ZN(n8279) );
  INV_X1 U6404 ( .A(n4498), .ZN(n4771) );
  NAND2_X1 U6405 ( .A1(n4495), .A2(n8081), .ZN(n4494) );
  NAND2_X1 U6406 ( .A1(n4499), .A2(n4404), .ZN(n4498) );
  NAND2_X1 U6407 ( .A1(n4773), .A2(n5063), .ZN(n4499) );
  NAND2_X2 U6408 ( .A1(n4502), .A2(n6277), .ZN(n8074) );
  NAND2_X1 U6409 ( .A1(n4724), .A2(n4399), .ZN(n5408) );
  NAND3_X1 U6410 ( .A1(n6782), .A2(n10195), .A3(n9874), .ZN(n4504) );
  NAND2_X1 U6411 ( .A1(n8974), .A2(n4507), .ZN(n8975) );
  NAND3_X1 U6412 ( .A1(n4509), .A2(n4787), .A3(n5093), .ZN(n9911) );
  NAND2_X1 U6413 ( .A1(n7637), .A2(n5415), .ZN(n5419) );
  NAND2_X1 U6414 ( .A1(n5036), .A2(n4397), .ZN(n7759) );
  AOI21_X2 U6415 ( .B1(n9180), .B2(n9187), .A(n5101), .ZN(n9171) );
  OAI21_X2 U6416 ( .B1(n4597), .B2(n4511), .A(n5649), .ZN(n9180) );
  NAND2_X1 U6417 ( .A1(n7632), .A2(n7634), .ZN(n7554) );
  INV_X1 U6418 ( .A(n4519), .ZN(n4518) );
  OAI21_X2 U6419 ( .B1(n5525), .B2(n4950), .A(n4302), .ZN(n5563) );
  OAI21_X2 U6420 ( .B1(n5563), .B2(n5225), .A(n5224), .ZN(n5577) );
  OAI21_X1 U6421 ( .B1(n5588), .B2(n4528), .A(n4527), .ZN(n4529) );
  INV_X1 U6422 ( .A(n5005), .ZN(n4531) );
  NAND2_X1 U6423 ( .A1(n9216), .A2(n9215), .ZN(n9218) );
  NAND4_X1 U6424 ( .A1(n6007), .A2(n9216), .A3(n9215), .A4(n6005), .ZN(n4532)
         );
  NAND2_X1 U6425 ( .A1(n9218), .A2(n5005), .ZN(n4533) );
  NAND3_X1 U6426 ( .A1(n4532), .A2(n6006), .A3(n4530), .ZN(n9186) );
  NAND3_X1 U6427 ( .A1(n6007), .A2(n6005), .A3(n4531), .ZN(n4530) );
  OAI21_X2 U6428 ( .B1(n9903), .B2(n4544), .A(n4317), .ZN(n8404) );
  NAND3_X1 U6429 ( .A1(n4541), .A2(n8651), .A3(n4540), .ZN(n6788) );
  NAND2_X2 U6430 ( .A1(n4546), .A2(n4545), .ZN(n8078) );
  NAND3_X1 U6431 ( .A1(n4547), .A2(n4394), .A3(n8677), .ZN(n4546) );
  NAND2_X1 U6432 ( .A1(n7455), .A2(n7730), .ZN(n8480) );
  NAND2_X2 U6433 ( .A1(n5054), .A2(n4548), .ZN(n7730) );
  AND2_X2 U6434 ( .A1(n5143), .A2(n4549), .ZN(n4848) );
  INV_X1 U6435 ( .A(n5564), .ZN(n4549) );
  NAND2_X1 U6436 ( .A1(n4550), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5607) );
  INV_X1 U6437 ( .A(n8032), .ZN(n4555) );
  INV_X1 U6438 ( .A(n4978), .ZN(n4977) );
  AND2_X1 U6439 ( .A1(n7551), .A2(n7554), .ZN(n5371) );
  NAND2_X1 U6440 ( .A1(n7645), .A2(n5872), .ZN(n5793) );
  NAND2_X1 U6441 ( .A1(n7462), .A2(n7465), .ZN(n7461) );
  AOI21_X2 U6442 ( .B1(n8796), .B2(n8797), .A(n6144), .ZN(n8888) );
  NAND2_X1 U6443 ( .A1(n6128), .A2(n8837), .ZN(n8771) );
  NAND2_X1 U6444 ( .A1(n4570), .A2(n8897), .ZN(P2_U3180) );
  NAND2_X1 U6445 ( .A1(n4571), .A2(n8882), .ZN(n4570) );
  XNOR2_X1 U6446 ( .A(n8888), .B(n8889), .ZN(n4571) );
  NOR2_X1 U6447 ( .A1(n8335), .A2(n8255), .ZN(n8256) );
  NOR2_X1 U6448 ( .A1(n4959), .A2(n4954), .ZN(n4953) );
  AND2_X4 U6449 ( .A1(n6306), .A2(n4281), .ZN(n6593) );
  NAND2_X1 U6450 ( .A1(n6675), .A2(n5059), .ZN(n5058) );
  NOR2_X1 U6451 ( .A1(n9625), .A2(n4573), .ZN(n9627) );
  NAND2_X1 U6452 ( .A1(n4677), .A2(n4684), .ZN(n9525) );
  NOR2_X1 U6453 ( .A1(n7297), .A2(n7298), .ZN(n4746) );
  NAND2_X1 U6454 ( .A1(n4748), .A2(n4747), .ZN(n4882) );
  NOR2_X1 U6455 ( .A1(n7224), .A2(n4594), .ZN(n7100) );
  NAND2_X1 U6456 ( .A1(n4932), .A2(n4931), .ZN(n5629) );
  NAND2_X2 U6457 ( .A1(n4952), .A2(n4409), .ZN(n5652) );
  NAND2_X1 U6458 ( .A1(n4800), .A2(n5420), .ZN(n4794) );
  AOI21_X1 U6459 ( .B1(n9288), .B2(n9287), .A(n5901), .ZN(n5800) );
  NAND2_X1 U6460 ( .A1(n5793), .A2(n5011), .ZN(n5010) );
  INV_X2 U6461 ( .A(n5328), .ZN(n5305) );
  NOR2_X1 U6462 ( .A1(n9153), .A2(n6760), .ZN(n6774) );
  NOR2_X2 U6463 ( .A1(n4287), .A2(n5857), .ZN(n7449) );
  OAI211_X1 U6464 ( .C1(n5293), .C2(n5790), .A(n5789), .B(n7444), .ZN(n4985)
         );
  NAND2_X1 U6465 ( .A1(n6665), .A2(n4613), .ZN(n4779) );
  NAND2_X1 U6466 ( .A1(n7084), .A2(n7322), .ZN(n5290) );
  NAND2_X2 U6467 ( .A1(n6105), .A2(n6104), .ZN(n8733) );
  NAND2_X1 U6468 ( .A1(n7391), .A2(n7390), .ZN(n7389) );
  XNOR2_X1 U6469 ( .A(n6070), .B(n5291), .ZN(n6063) );
  NAND2_X1 U6470 ( .A1(n4585), .A2(n5081), .ZN(n9979) );
  NAND3_X1 U6471 ( .A1(n4660), .A2(n4659), .A3(n4389), .ZN(n4585) );
  NAND2_X2 U6472 ( .A1(n6656), .A2(n6655), .ZN(n6319) );
  NAND2_X1 U6473 ( .A1(n6330), .A2(n8466), .ZN(n7603) );
  NAND2_X4 U6474 ( .A1(n8395), .A2(n6251), .ZN(n6647) );
  NAND2_X1 U6475 ( .A1(n4587), .A2(n6006), .ZN(n5938) );
  NAND3_X1 U6476 ( .A1(n5936), .A2(n6007), .A3(n6005), .ZN(n4587) );
  NAND2_X1 U6477 ( .A1(n4326), .A2(n4588), .ZN(n5916) );
  NAND3_X1 U6478 ( .A1(n4715), .A2(n4712), .A3(n4590), .ZN(n4711) );
  AND2_X1 U6479 ( .A1(n5870), .A2(n7648), .ZN(n4590) );
  NAND2_X1 U6480 ( .A1(n4701), .A2(n4700), .ZN(n4699) );
  NAND2_X1 U6481 ( .A1(n4676), .A2(n4401), .ZN(n9594) );
  NAND2_X1 U6482 ( .A1(n4685), .A2(n4299), .ZN(n9552) );
  AOI21_X2 U6483 ( .B1(n9169), .B2(n6003), .A(n5932), .ZN(n6207) );
  NAND2_X1 U6484 ( .A1(n9070), .A2(n4736), .ZN(n4733) );
  NAND2_X1 U6485 ( .A1(n4889), .A2(n8950), .ZN(n8955) );
  NAND3_X1 U6486 ( .A1(n9143), .A2(n4593), .A3(n4591), .ZN(P2_U3201) );
  NAND2_X1 U6487 ( .A1(n5029), .A2(n5313), .ZN(n5028) );
  NAND2_X1 U6488 ( .A1(n4293), .A2(n5151), .ZN(n8431) );
  NAND2_X1 U6489 ( .A1(n4724), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U6490 ( .A1(n7446), .A2(n5861), .ZN(n7462) );
  INV_X1 U6491 ( .A(n10028), .ZN(n6494) );
  NAND2_X2 U6492 ( .A1(n9970), .A2(n9971), .ZN(n9969) );
  INV_X1 U6493 ( .A(n4942), .ZN(n4941) );
  NAND3_X1 U6494 ( .A1(n4600), .A2(n6758), .A3(n6741), .ZN(n9153) );
  NAND2_X1 U6495 ( .A1(n6743), .A2(n6742), .ZN(n4600) );
  INV_X1 U6496 ( .A(n6009), .ZN(n5000) );
  OAI21_X1 U6497 ( .B1(n5798), .B2(n4998), .A(n4623), .ZN(n4622) );
  OAI21_X1 U6498 ( .B1(n6238), .B2(n4602), .A(n4601), .ZN(n5206) );
  NAND2_X1 U6499 ( .A1(n4699), .A2(n5925), .ZN(n5936) );
  INV_X1 U6500 ( .A(n4604), .ZN(n4603) );
  OAI21_X1 U6501 ( .B1(n5974), .B2(n4703), .A(n6042), .ZN(n4604) );
  NOR2_X4 U6502 ( .A1(n9935), .A2(n9921), .ZN(n9924) );
  NAND2_X1 U6503 ( .A1(n5747), .A2(n5746), .ZN(n5755) );
  NAND2_X1 U6504 ( .A1(n5745), .A2(n7861), .ZN(n5747) );
  OAI21_X1 U6505 ( .B1(n8750), .B2(n6097), .A(n4607), .ZN(n6100) );
  NAND2_X1 U6506 ( .A1(n4610), .A2(n4608), .ZN(P2_U3169) );
  OAI21_X1 U6507 ( .B1(n4324), .B2(n5153), .A(P2_IR_REG_27__SCAN_IN), .ZN(
        n5008) );
  NAND2_X1 U6508 ( .A1(n5163), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U6509 ( .A1(n4622), .A2(n4393), .ZN(n5803) );
  NAND2_X1 U6510 ( .A1(n6678), .A2(n6677), .ZN(n10001) );
  NAND2_X1 U6511 ( .A1(n5315), .A2(n7432), .ZN(n5027) );
  AOI21_X1 U6513 ( .B1(n9186), .B2(n5937), .A(n5806), .ZN(n9169) );
  NOR2_X1 U6514 ( .A1(n5866), .A2(n5865), .ZN(n5792) );
  NAND2_X1 U6515 ( .A1(n9002), .A2(n4312), .ZN(n4626) );
  INV_X1 U6516 ( .A(n7295), .ZN(n4642) );
  NAND2_X1 U6517 ( .A1(n4636), .A2(n4637), .ZN(n8960) );
  NAND2_X1 U6518 ( .A1(n7295), .A2(n4291), .ZN(n4636) );
  NOR2_X1 U6519 ( .A1(n7295), .A2(n7294), .ZN(n7521) );
  INV_X1 U6520 ( .A(n7294), .ZN(n4649) );
  NAND3_X1 U6521 ( .A1(n4657), .A2(n4656), .A3(n4655), .ZN(n7087) );
  NAND3_X1 U6522 ( .A1(n5262), .A2(n5263), .A3(P2_REG2_REG_1__SCAN_IN), .ZN(
        n4657) );
  NAND2_X1 U6523 ( .A1(n4661), .A2(n5084), .ZN(n4659) );
  NAND2_X1 U6524 ( .A1(n10070), .A2(n4661), .ZN(n4660) );
  OAI21_X1 U6525 ( .B1(n10070), .B2(n5084), .A(n4661), .ZN(n10018) );
  XNOR2_X2 U6526 ( .A(n6319), .B(n9567), .ZN(n8604) );
  NAND3_X1 U6527 ( .A1(n4674), .A2(n6840), .A3(n4673), .ZN(n7659) );
  NAND3_X1 U6528 ( .A1(n7406), .A2(n7453), .A3(n7407), .ZN(n4674) );
  NAND2_X1 U6529 ( .A1(n4921), .A2(n4678), .ZN(n4676) );
  NAND2_X1 U6530 ( .A1(n4921), .A2(n4682), .ZN(n4677) );
  NAND2_X1 U6531 ( .A1(n6888), .A2(n6889), .ZN(n4687) );
  OAI21_X1 U6532 ( .B1(n8226), .B2(n4690), .A(n4688), .ZN(n4693) );
  AOI21_X1 U6533 ( .B1(n4689), .B2(n6897), .A(n4691), .ZN(n4688) );
  INV_X1 U6534 ( .A(n6888), .ZN(n4689) );
  NAND2_X1 U6535 ( .A1(n9537), .A2(n6897), .ZN(n4690) );
  INV_X1 U6536 ( .A(n9587), .ZN(n4691) );
  NAND2_X1 U6537 ( .A1(n9536), .A2(n6888), .ZN(n4692) );
  NAND2_X1 U6538 ( .A1(n4693), .A2(n9585), .ZN(n9589) );
  NAND4_X1 U6539 ( .A1(n6231), .A2(n6232), .A3(n6233), .A4(n6240), .ZN(n4695)
         );
  NAND4_X1 U6540 ( .A1(n6230), .A2(n6228), .A3(n6229), .A4(n6241), .ZN(n6429)
         );
  NAND3_X1 U6541 ( .A1(n4711), .A2(n4708), .A3(n4705), .ZN(n5882) );
  NAND2_X1 U6542 ( .A1(n5879), .A2(n5871), .ZN(n4709) );
  NAND2_X1 U6543 ( .A1(n4714), .A2(n5858), .ZN(n4713) );
  NAND2_X1 U6544 ( .A1(n5860), .A2(n5859), .ZN(n4714) );
  OR2_X1 U6545 ( .A1(n5867), .A2(n6152), .ZN(n4715) );
  NOR2_X1 U6546 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  INV_X1 U6547 ( .A(n5420), .ZN(n4721) );
  NAND3_X1 U6548 ( .A1(n4721), .A2(n4722), .A3(n5195), .ZN(n4720) );
  NAND2_X1 U6549 ( .A1(n5183), .A2(n4786), .ZN(n5364) );
  NAND2_X1 U6550 ( .A1(n4726), .A2(n4725), .ZN(n5363) );
  NAND2_X1 U6551 ( .A1(n4742), .A2(n4743), .ZN(n7330) );
  NOR2_X1 U6552 ( .A1(n4744), .A2(n7103), .ZN(n4741) );
  NOR2_X1 U6553 ( .A1(n7101), .A2(n7595), .ZN(n4742) );
  INV_X1 U6554 ( .A(n4744), .ZN(n4743) );
  NOR2_X1 U6555 ( .A1(n7101), .A2(n4744), .ZN(n7331) );
  NAND2_X1 U6556 ( .A1(n7205), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7299) );
  NOR2_X1 U6557 ( .A1(n4746), .A2(n4883), .ZN(n4747) );
  NAND2_X1 U6558 ( .A1(n7205), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U6559 ( .A1(n4753), .A2(n7299), .ZN(n4752) );
  NAND2_X1 U6560 ( .A1(n4758), .A2(n4754), .ZN(n7815) );
  NAND2_X1 U6561 ( .A1(n8930), .A2(n8928), .ZN(n4758) );
  NAND2_X1 U6562 ( .A1(n8988), .A2(n8987), .ZN(n8989) );
  INV_X1 U6563 ( .A(n5397), .ZN(n5123) );
  NAND3_X1 U6564 ( .A1(n5120), .A2(n5121), .A3(n7549), .ZN(n5397) );
  NAND2_X1 U6565 ( .A1(n5515), .A2(n4764), .ZN(n5597) );
  NAND2_X1 U6566 ( .A1(n5131), .A2(n4767), .ZN(n5641) );
  NAND2_X1 U6567 ( .A1(n8170), .A2(n5115), .ZN(n4777) );
  MUX2_X1 U6568 ( .A(n7143), .B(n5178), .S(n5184), .Z(n5181) );
  MUX2_X1 U6569 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7131), .Z(n5190) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7131), .Z(n5209) );
  MUX2_X1 U6571 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7131), .Z(n5561) );
  MUX2_X1 U6572 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7131), .Z(n5235) );
  MUX2_X1 U6573 ( .A(n8224), .B(n8307), .S(n7131), .Z(n5627) );
  MUX2_X1 U6574 ( .A(n9499), .B(n10253), .S(n7131), .Z(n5678) );
  MUX2_X1 U6575 ( .A(n5716), .B(n8430), .S(n7131), .Z(n5828) );
  NAND2_X1 U6576 ( .A1(n4781), .A2(n4780), .ZN(P1_U3549) );
  NAND2_X1 U6577 ( .A1(n10125), .A2(n10408), .ZN(n4781) );
  NAND2_X1 U6578 ( .A1(n4783), .A2(n4782), .ZN(P1_U3517) );
  NAND2_X1 U6579 ( .A1(n10125), .A2(n10405), .ZN(n4783) );
  AND2_X1 U6580 ( .A1(n5344), .A2(n4784), .ZN(n4786) );
  NAND2_X1 U6581 ( .A1(n5345), .A2(n4785), .ZN(n4784) );
  INV_X1 U6582 ( .A(n5342), .ZN(n4785) );
  NAND2_X1 U6583 ( .A1(n5421), .A2(n4800), .ZN(n4795) );
  NAND3_X1 U6584 ( .A1(n4802), .A2(n5162), .A3(P1_DATAO_REG_3__SCAN_IN), .ZN(
        n4806) );
  NAND3_X1 U6585 ( .A1(n4807), .A2(n4806), .A3(n4805), .ZN(n5180) );
  NAND3_X1 U6586 ( .A1(n4808), .A2(n4809), .A3(P2_DATAO_REG_3__SCAN_IN), .ZN(
        n4805) );
  NOR2_X1 U6587 ( .A1(n4286), .A2(n8469), .ZN(n4811) );
  NAND2_X1 U6588 ( .A1(n6330), .A2(n4811), .ZN(n7722) );
  NAND2_X1 U6589 ( .A1(n7722), .A2(n8465), .ZN(n8476) );
  NAND2_X1 U6590 ( .A1(n8545), .A2(n4307), .ZN(n4814) );
  NOR2_X1 U6591 ( .A1(n4815), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U6592 ( .A1(n8551), .A2(n9930), .ZN(n4819) );
  NAND2_X1 U6593 ( .A1(n4823), .A2(n4820), .ZN(n8496) );
  AOI21_X1 U6594 ( .B1(n4822), .B2(n4391), .A(n4296), .ZN(n4820) );
  OAI21_X1 U6595 ( .B1(n8483), .B2(n8479), .A(n8484), .ZN(n4822) );
  OAI21_X1 U6596 ( .B1(n4824), .B2(n8489), .A(n8582), .ZN(n4823) );
  AOI21_X1 U6597 ( .B1(n8487), .B2(n8486), .A(n4825), .ZN(n4824) );
  INV_X1 U6598 ( .A(n5115), .ZN(n4825) );
  NAND3_X1 U6599 ( .A1(n4830), .A2(n4828), .A3(n4827), .ZN(n4826) );
  NAND4_X1 U6600 ( .A1(n8531), .A2(n8530), .A3(n8582), .A4(n8529), .ZN(n4827)
         );
  NAND3_X1 U6601 ( .A1(n8519), .A2(n10040), .A3(n4285), .ZN(n4830) );
  NAND3_X1 U6602 ( .A1(n8577), .A2(n8571), .A3(n4387), .ZN(n4834) );
  INV_X1 U6603 ( .A(n5902), .ZN(n4837) );
  OAI21_X1 U6604 ( .B1(n5900), .B2(n4838), .A(n4836), .ZN(n5911) );
  NAND4_X1 U6605 ( .A1(n5914), .A2(n5917), .A3(n5915), .A4(n5918), .ZN(n4840)
         );
  NAND3_X1 U6606 ( .A1(n5933), .A2(n6206), .A3(n5935), .ZN(n4846) );
  NAND2_X1 U6607 ( .A1(n4848), .A2(n5305), .ZN(n5593) );
  NAND2_X1 U6608 ( .A1(n7132), .A2(n4281), .ZN(n4851) );
  NAND2_X1 U6609 ( .A1(n4850), .A2(n6739), .ZN(n4849) );
  NAND2_X1 U6610 ( .A1(n4851), .A2(n4361), .ZN(n4850) );
  NAND2_X1 U6611 ( .A1(n4859), .A2(n4858), .ZN(n8251) );
  NAND2_X1 U6612 ( .A1(n7514), .A2(n4398), .ZN(n4858) );
  NAND2_X1 U6613 ( .A1(n4861), .A2(n4860), .ZN(n4859) );
  NAND2_X1 U6614 ( .A1(n7514), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8942) );
  INV_X1 U6615 ( .A(n7212), .ZN(n4865) );
  NAND2_X1 U6616 ( .A1(n9035), .A2(n9060), .ZN(n9036) );
  NAND2_X1 U6617 ( .A1(n4870), .A2(n7114), .ZN(n4871) );
  NAND2_X1 U6618 ( .A1(n7112), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4870) );
  NAND2_X1 U6619 ( .A1(n4871), .A2(n7113), .ZN(n7210) );
  NAND2_X1 U6620 ( .A1(n8256), .A2(n4874), .ZN(n4872) );
  NAND2_X1 U6621 ( .A1(n8256), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U6622 ( .A1(n7477), .A2(n6320), .ZN(n8468) );
  OAI211_X2 U6623 ( .C1(n7096), .C2(n4877), .A(n5328), .B(n4876), .ZN(n7223)
         );
  NAND2_X1 U6624 ( .A1(n4879), .A2(n9009), .ZN(n4880) );
  NAND2_X1 U6625 ( .A1(n4888), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4887) );
  NAND2_X1 U6626 ( .A1(n4887), .A2(n9046), .ZN(n4885) );
  NAND2_X1 U6627 ( .A1(n4885), .A2(n9048), .ZN(n9068) );
  NAND2_X1 U6628 ( .A1(n4891), .A2(n8951), .ZN(n4889) );
  AND2_X2 U6629 ( .A1(n9924), .A2(n4898), .ZN(n8419) );
  NOR2_X1 U6630 ( .A1(n8074), .A2(n4902), .ZN(n4901) );
  OAI21_X1 U6631 ( .B1(n9603), .B2(n6926), .A(n6925), .ZN(n9607) );
  INV_X1 U6632 ( .A(n8600), .ZN(n4914) );
  OR2_X1 U6633 ( .A1(n8600), .A2(n6650), .ZN(n6803) );
  NOR2_X1 U6634 ( .A1(n8590), .A2(n6650), .ZN(n4913) );
  OAI22_X2 U6635 ( .A1(n7673), .A2(n4354), .B1(n6870), .B2(n4918), .ZN(n8226)
         );
  INV_X1 U6636 ( .A(n7671), .ZN(n4918) );
  OR2_X2 U6637 ( .A1(n6912), .A2(n6911), .ZN(n4920) );
  AND2_X1 U6638 ( .A1(n4929), .A2(n4928), .ZN(n4927) );
  NAND2_X1 U6639 ( .A1(n5592), .A2(n4933), .ZN(n4932) );
  AND2_X1 U6640 ( .A1(n5659), .A2(n5658), .ZN(n5676) );
  OAI21_X2 U6641 ( .B1(n5472), .B2(n4941), .A(n4940), .ZN(n5525) );
  NAND2_X1 U6642 ( .A1(n4952), .A2(n5244), .ZN(n5638) );
  NAND2_X1 U6643 ( .A1(n8796), .A2(n4966), .ZN(n4963) );
  NAND2_X1 U6644 ( .A1(n8796), .A2(n4966), .ZN(n4965) );
  OAI21_X2 U6645 ( .B1(n6077), .B2(n4977), .A(n4975), .ZN(n8032) );
  NOR2_X1 U6646 ( .A1(n4979), .A2(n5153), .ZN(n5744) );
  NAND2_X1 U6647 ( .A1(n4985), .A2(n7449), .ZN(n7446) );
  NAND2_X1 U6648 ( .A1(n6052), .A2(n4991), .ZN(n4990) );
  OAI211_X1 U6649 ( .C1(n6052), .C2(n4986), .A(n4990), .B(n4988), .ZN(n6058)
         );
  NAND2_X1 U6650 ( .A1(n6738), .A2(n6048), .ZN(n4996) );
  AND2_X1 U6651 ( .A1(n5800), .A2(n5000), .ZN(n4999) );
  NAND2_X1 U6652 ( .A1(n5798), .A2(n5899), .ZN(n9286) );
  INV_X1 U6653 ( .A(n5899), .ZN(n5003) );
  NAND2_X1 U6654 ( .A1(n5010), .A2(n5009), .ZN(n8024) );
  AOI21_X2 U6655 ( .B1(n8297), .B2(n5015), .A(n5013), .ZN(n9313) );
  NAND2_X1 U6656 ( .A1(n6739), .A2(n4390), .ZN(n5024) );
  NAND3_X1 U6657 ( .A1(n6739), .A2(n4281), .A3(n7134), .ZN(n5023) );
  NAND2_X1 U6658 ( .A1(n5517), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5311) );
  OR2_X4 U6659 ( .A1(n5155), .A2(n5156), .ZN(n5958) );
  NAND2_X1 U6660 ( .A1(n9273), .A2(n5033), .ZN(n5031) );
  NAND2_X1 U6661 ( .A1(n5419), .A2(n5418), .ZN(n7611) );
  NAND2_X1 U6662 ( .A1(n5037), .A2(n5038), .ZN(n5506) );
  NAND2_X1 U6663 ( .A1(n8194), .A2(n5491), .ZN(n5037) );
  NAND4_X1 U6664 ( .A1(n5053), .A2(n6226), .A3(n6224), .A4(n6225), .ZN(n6702)
         );
  NAND2_X1 U6665 ( .A1(n9741), .A2(n7845), .ZN(n8471) );
  NAND2_X1 U6666 ( .A1(n5058), .A2(n5056), .ZN(n6678) );
  NAND2_X1 U6667 ( .A1(n5076), .A2(n6689), .ZN(n9896) );
  NAND2_X1 U6668 ( .A1(n8078), .A2(n5088), .ZN(n5087) );
  NAND3_X1 U6669 ( .A1(n5087), .A2(n8517), .A3(n5086), .ZN(n10082) );
  NAND3_X1 U6670 ( .A1(n5092), .A2(n5091), .A3(n8480), .ZN(n7710) );
  NAND2_X1 U6671 ( .A1(n6351), .A2(n8469), .ZN(n5091) );
  NAND2_X1 U6672 ( .A1(n7603), .A2(n6351), .ZN(n5092) );
  NAND2_X1 U6673 ( .A1(n7722), .A2(n6351), .ZN(n7724) );
  NAND2_X1 U6674 ( .A1(n8595), .A2(n8503), .ZN(n5098) );
  INV_X1 U6675 ( .A(n8117), .ZN(n5099) );
  NAND2_X1 U6676 ( .A1(n7068), .A2(n8882), .ZN(n7074) );
  OR2_X1 U6677 ( .A1(n6739), .A2(n7223), .ZN(n5306) );
  INV_X1 U6678 ( .A(n4279), .ZN(n7116) );
  AOI21_X1 U6679 ( .B1(n10232), .B2(n8731), .A(n8730), .ZN(n8732) );
  CLKBUF_X1 U6680 ( .A(n8226), .Z(n9536) );
  OR2_X1 U6681 ( .A1(n5388), .A2(n10444), .ZN(n5307) );
  INV_X1 U6682 ( .A(n5388), .ZN(n5354) );
  OR2_X1 U6683 ( .A1(n8582), .A2(n6650), .ZN(n10212) );
  NAND2_X1 U6684 ( .A1(n8591), .A2(n8600), .ZN(n10380) );
  NAND2_X1 U6685 ( .A1(n8391), .A2(n5156), .ZN(n5388) );
  NAND2_X1 U6686 ( .A1(n5747), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5749) );
  OAI211_X1 U6687 ( .C1(n8414), .C2(n10401), .A(n8410), .B(n8407), .ZN(n10125)
         );
  NOR2_X1 U6688 ( .A1(n6223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6501) );
  INV_X2 U6689 ( .A(n10446), .ZN(n9404) );
  INV_X1 U6690 ( .A(n10448), .ZN(n10446) );
  AND2_X2 U6691 ( .A1(n6735), .A2(n7793), .ZN(n10405) );
  AND2_X2 U6692 ( .A1(n6730), .A2(n7793), .ZN(n10408) );
  AND2_X1 U6693 ( .A1(n6805), .A2(n6804), .ZN(n5100) );
  INV_X1 U6694 ( .A(n9242), .ZN(n5625) );
  AND2_X1 U6695 ( .A1(n9179), .A2(n8890), .ZN(n5101) );
  OR2_X1 U6696 ( .A1(n6695), .A2(n6800), .ZN(n5102) );
  OR2_X1 U6697 ( .A1(n6695), .A2(n6796), .ZN(n5103) );
  AND2_X1 U6698 ( .A1(n6628), .A2(n6627), .ZN(n5104) );
  AND2_X1 U6699 ( .A1(n5743), .A2(n5773), .ZN(n5105) );
  NAND3_X1 U6700 ( .A1(n6704), .A2(n6707), .A3(n6227), .ZN(n5106) );
  NOR2_X1 U6701 ( .A1(n9154), .A2(n9381), .ZN(n5107) );
  AND2_X1 U6702 ( .A1(n6149), .A2(n8913), .ZN(n5108) );
  NOR2_X1 U6703 ( .A1(n9154), .A2(n9461), .ZN(n5109) );
  INV_X1 U6704 ( .A(n5365), .ZN(n5992) );
  INV_X1 U6705 ( .A(n9227), .ZN(n9261) );
  OR2_X1 U6706 ( .A1(n7076), .A2(n6806), .ZN(n5110) );
  OR2_X1 U6707 ( .A1(n9074), .A2(n9397), .ZN(n5111) );
  INV_X2 U6708 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U6709 ( .A(n7767), .ZN(n10428) );
  INV_X1 U6710 ( .A(n6007), .ZN(n5804) );
  AND2_X1 U6711 ( .A1(n5993), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5112) );
  AND2_X1 U6712 ( .A1(n10405), .A2(n10397), .ZN(n10232) );
  INV_X1 U6713 ( .A(n9497), .ZN(n8434) );
  AND2_X1 U6714 ( .A1(n5993), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6715 ( .A1(n9281), .A2(n9260), .ZN(n5114) );
  INV_X1 U6716 ( .A(n9054), .ZN(n9034) );
  INV_X1 U6717 ( .A(n10186), .ZN(n6694) );
  INV_X1 U6718 ( .A(n10216), .ZN(n8418) );
  INV_X1 U6719 ( .A(n7653), .ZN(n6742) );
  INV_X1 U6720 ( .A(n9890), .ZN(n6695) );
  OR2_X1 U6721 ( .A1(n6189), .A2(n6188), .ZN(n5116) );
  AND2_X1 U6722 ( .A1(n5818), .A2(n5817), .ZN(n5117) );
  AND2_X1 U6723 ( .A1(n6752), .A2(n6747), .ZN(n5118) );
  NOR2_X1 U6724 ( .A1(n10127), .A2(n9906), .ZN(n5119) );
  AND2_X1 U6725 ( .A1(n7632), .A2(n5862), .ZN(n5863) );
  NAND2_X1 U6726 ( .A1(n5916), .A2(n7082), .ZN(n5917) );
  MUX2_X1 U6727 ( .A(n5842), .B(n5841), .S(n7082), .Z(n5925) );
  NAND2_X1 U6728 ( .A1(n5931), .A2(n6152), .ZN(n5926) );
  INV_X1 U6729 ( .A(n6003), .ZN(n5927) );
  NOR2_X1 U6730 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  OAI21_X1 U6731 ( .B1(n5930), .B2(n5929), .A(n5928), .ZN(n5934) );
  INV_X1 U6732 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6227) );
  INV_X1 U6733 ( .A(n5148), .ZN(n5149) );
  INV_X1 U6734 ( .A(n9913), .ZN(n6579) );
  INV_X1 U6735 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6736 ( .A1(n10427), .A2(n5314), .ZN(n5313) );
  INV_X1 U6737 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5150) );
  INV_X1 U6738 ( .A(n7581), .ZN(n6076) );
  INV_X1 U6739 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7530) );
  INV_X1 U6740 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8739) );
  INV_X1 U6741 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5120) );
  AND2_X1 U6742 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  INV_X1 U6743 ( .A(n8200), .ZN(n5490) );
  INV_X1 U6744 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9650) );
  OR2_X1 U6745 ( .A1(n8402), .A2(n8624), .ZN(n8403) );
  INV_X1 U6746 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6376) );
  AND2_X1 U6747 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  AND2_X1 U6748 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  INV_X1 U6749 ( .A(n5637), .ZN(n5249) );
  INV_X1 U6750 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6466) );
  INV_X1 U6751 ( .A(n8031), .ZN(n6085) );
  OR2_X1 U6752 ( .A1(n6070), .A2(n7474), .ZN(n6065) );
  NOR2_X1 U6753 ( .A1(n7313), .A2(n7099), .ZN(n7225) );
  INV_X1 U6754 ( .A(n7814), .ZN(n8929) );
  NAND2_X1 U6755 ( .A1(n9077), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9067) );
  INV_X1 U6756 ( .A(n9334), .ZN(n6108) );
  INV_X1 U6757 ( .A(n8026), .ZN(n5794) );
  XNOR2_X1 U6758 ( .A(n6814), .B(n6849), .ZN(n6819) );
  NAND2_X1 U6759 ( .A1(n6307), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6309) );
  INV_X1 U6760 ( .A(n8611), .ZN(n6412) );
  INV_X1 U6761 ( .A(n6264), .ZN(n6265) );
  INV_X1 U6762 ( .A(SI_20_), .ZN(n5239) );
  INV_X1 U6763 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6627) );
  AND2_X1 U6764 ( .A1(n5194), .A2(n5376), .ZN(n5195) );
  INV_X1 U6765 ( .A(n5325), .ZN(n5322) );
  OR2_X1 U6766 ( .A1(n7080), .A2(n7079), .ZN(n7123) );
  INV_X1 U6767 ( .A(n8902), .ZN(n8780) );
  NAND2_X1 U6768 ( .A1(n6215), .A2(n6171), .ZN(n8904) );
  OR2_X1 U6769 ( .A1(n5958), .A2(n5294), .ZN(n5297) );
  NAND2_X1 U6770 ( .A1(n9076), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9115) );
  AND2_X1 U6771 ( .A1(n7125), .A2(n7124), .ZN(n9131) );
  AND2_X1 U6772 ( .A1(n7767), .A2(n8225), .ZN(n6762) );
  AND2_X1 U6773 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  AND2_X1 U6774 ( .A1(n6001), .A2(n6000), .ZN(n9147) );
  AND2_X1 U6775 ( .A1(n6208), .A2(n9160), .ZN(n6209) );
  AND2_X1 U6776 ( .A1(n5908), .A2(n5905), .ZN(n6011) );
  AND2_X1 U6777 ( .A1(n8104), .A2(n6053), .ZN(n5816) );
  INV_X1 U6778 ( .A(n9331), .ZN(n9296) );
  AND2_X1 U6779 ( .A1(n7357), .A2(n6811), .ZN(n9564) );
  INV_X1 U6780 ( .A(n6951), .ZN(n9553) );
  OR2_X1 U6781 ( .A1(n9951), .A2(n6529), .ZN(n6557) );
  INV_X1 U6782 ( .A(n9934), .ZN(n9952) );
  INV_X1 U6783 ( .A(n8618), .ZN(n10051) );
  INV_X1 U6784 ( .A(n10086), .ZN(n9716) );
  INV_X1 U6785 ( .A(n7707), .ZN(n8605) );
  INV_X1 U6786 ( .A(n10366), .ZN(n10069) );
  INV_X1 U6787 ( .A(n10408), .ZN(n6794) );
  OR2_X1 U6788 ( .A1(n10380), .A2(n6802), .ZN(n10180) );
  INV_X1 U6789 ( .A(n8614), .ZN(n8525) );
  INV_X1 U6790 ( .A(n9733), .ZN(n9682) );
  OR2_X1 U6791 ( .A1(n10380), .A2(n6650), .ZN(n10091) );
  INV_X1 U6792 ( .A(n10087), .ZN(n10392) );
  OAI211_X1 U6793 ( .C1(n5833), .C2(n5832), .A(n5831), .B(n5830), .ZN(n5942)
         );
  AND2_X1 U6794 ( .A1(n5692), .A2(n5663), .ZN(n5675) );
  INV_X1 U6795 ( .A(n6195), .ZN(n6196) );
  NAND2_X1 U6796 ( .A1(n6181), .A2(n6180), .ZN(n8906) );
  AND3_X1 U6797 ( .A1(n5575), .A2(n5574), .A3(n5573), .ZN(n9295) );
  INV_X1 U6798 ( .A(n9131), .ZN(n9004) );
  NAND2_X1 U6799 ( .A1(n6158), .A2(n6762), .ZN(n10417) );
  INV_X1 U6800 ( .A(n10415), .ZN(n9325) );
  NOR2_X1 U6801 ( .A1(n9404), .A2(n6770), .ZN(n6771) );
  INV_X1 U6802 ( .A(n9381), .ZN(n9406) );
  AND2_X1 U6803 ( .A1(n6013), .A2(n6012), .ZN(n7614) );
  OR2_X1 U6804 ( .A1(n6151), .A2(n5777), .ZN(n6768) );
  INV_X1 U6805 ( .A(n6011), .ZN(n9307) );
  INV_X1 U6806 ( .A(n9480), .ZN(n9486) );
  AND2_X1 U6807 ( .A1(n8304), .A2(n5816), .ZN(n7767) );
  NAND2_X1 U6808 ( .A1(n7653), .A2(n10428), .ZN(n10426) );
  NOR2_X1 U6809 ( .A1(n4281), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9495) );
  INV_X1 U6810 ( .A(n9717), .ZN(n9695) );
  AND2_X1 U6811 ( .A1(n6493), .A2(n6492), .ZN(n10046) );
  AND2_X1 U6812 ( .A1(n7187), .A2(n7186), .ZN(n7280) );
  NAND2_X1 U6813 ( .A1(n7280), .A2(n7279), .ZN(n10334) );
  AND2_X1 U6814 ( .A1(n7280), .A2(n8429), .ZN(n10326) );
  INV_X1 U6815 ( .A(n10091), .ZN(n10052) );
  INV_X1 U6816 ( .A(n9971), .ZN(n9961) );
  AND2_X1 U6817 ( .A1(n8460), .A2(n8696), .ZN(n10019) );
  INV_X1 U6818 ( .A(n10072), .ZN(n10063) );
  INV_X1 U6819 ( .A(n8045), .ZN(n8003) );
  INV_X1 U6820 ( .A(n10045), .ZN(n10377) );
  OR2_X1 U6821 ( .A1(n10408), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6795) );
  AND2_X1 U6822 ( .A1(n10408), .A2(n10397), .ZN(n10159) );
  INV_X1 U6823 ( .A(n10195), .ZN(n10401) );
  INV_X1 U6824 ( .A(n7775), .ZN(n10354) );
  AND2_X1 U6825 ( .A1(n7162), .A2(n7052), .ZN(n7793) );
  INV_X1 U6826 ( .A(n8663), .ZN(n8375) );
  AND2_X1 U6827 ( .A1(n6483), .A2(n6482), .ZN(n9858) );
  XNOR2_X1 U6828 ( .A(n6416), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9848) );
  AND2_X1 U6829 ( .A1(n6289), .A2(n6430), .ZN(n9786) );
  INV_X1 U6830 ( .A(n7072), .ZN(n7073) );
  NOR2_X1 U6831 ( .A1(n5116), .A2(n6196), .ZN(n6197) );
  INV_X1 U6832 ( .A(n8906), .ZN(n8852) );
  INV_X1 U6833 ( .A(n8896), .ZN(n8909) );
  INV_X1 U6834 ( .A(n8789), .ZN(n9332) );
  INV_X1 U6835 ( .A(n8164), .ZN(n8918) );
  OR2_X1 U6836 ( .A1(n9103), .A2(n7092), .ZN(n9140) );
  NAND2_X1 U6837 ( .A1(n7240), .A2(n7116), .ZN(n9144) );
  INV_X1 U6838 ( .A(n10421), .ZN(n10413) );
  OR2_X1 U6839 ( .A1(n7625), .A2(n9337), .ZN(n10415) );
  INV_X1 U6840 ( .A(n9407), .ZN(n9403) );
  NOR2_X1 U6841 ( .A1(n6768), .A2(n6767), .ZN(n10448) );
  INV_X1 U6842 ( .A(n8835), .ZN(n9462) );
  OR2_X1 U6843 ( .A1(n10441), .A2(n10436), .ZN(n9480) );
  INV_X2 U6844 ( .A(n10441), .ZN(n10440) );
  INV_X1 U6845 ( .A(n7474), .ZN(n7757) );
  AND2_X1 U6846 ( .A1(n5757), .A2(n8446), .ZN(n7176) );
  INV_X1 U6847 ( .A(n7176), .ZN(n8449) );
  INV_X1 U6848 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8224) );
  INV_X1 U6849 ( .A(n8980), .ZN(n8999) );
  INV_X1 U6850 ( .A(n10168), .ZN(n10016) );
  AND2_X1 U6851 ( .A1(n7046), .A2(n10379), .ZN(n9712) );
  INV_X1 U6852 ( .A(n9996), .ZN(n9973) );
  INV_X1 U6853 ( .A(n9640), .ZN(n9735) );
  INV_X1 U6854 ( .A(n10314), .ZN(n10349) );
  NAND2_X1 U6855 ( .A1(n8423), .A2(n10052), .ZN(n8452) );
  INV_X1 U6856 ( .A(n10371), .ZN(n10079) );
  INV_X1 U6857 ( .A(n10405), .ZN(n10403) );
  AND2_X1 U6858 ( .A1(n10255), .A2(n10258), .ZN(n7164) );
  INV_X1 U6859 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10253) );
  INV_X1 U6860 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8307) );
  INV_X1 U6861 ( .A(n8439), .ZN(n10262) );
  INV_X1 U6862 ( .A(n9103), .ZN(P2_U3893) );
  AND2_X2 U6863 ( .A1(n7157), .A2(n7077), .ZN(P1_U3973) );
  INV_X2 U6864 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7549) );
  INV_X1 U6865 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6866 ( .A1(n5267), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6867 ( .A1(n5668), .A2(n5133), .ZN(n9197) );
  NOR2_X1 U6868 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5137) );
  NAND4_X1 U6869 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n5564)
         );
  NAND3_X1 U6870 ( .A1(n4493), .A2(n5140), .A3(n5139), .ZN(n5141) );
  NOR2_X4 U6871 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7096) );
  NOR2_X1 U6872 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5147) );
  NOR2_X1 U6873 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5146) );
  NOR2_X1 U6874 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5145) );
  NOR2_X1 U6875 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5144) );
  NAND4_X1 U6876 ( .A1(n5147), .A2(n5146), .A3(n5145), .A4(n5144), .ZN(n5148)
         );
  INV_X1 U6877 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5153) );
  XNOR2_X2 U6878 ( .A(n5154), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6879 ( .A1(n5155), .A2(n5156), .ZN(n5356) );
  INV_X1 U6880 ( .A(n5356), .ZN(n5277) );
  NAND2_X1 U6881 ( .A1(n9197), .A2(n5684), .ZN(n5161) );
  INV_X1 U6882 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U6883 ( .A1(n4282), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6884 ( .A1(n5955), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5157) );
  OAI211_X1 U6885 ( .C1(n9436), .C2(n5958), .A(n5158), .B(n5157), .ZN(n5159)
         );
  INV_X1 U6886 ( .A(n5159), .ZN(n5160) );
  INV_X1 U6887 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7145) );
  INV_X1 U6888 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7133) );
  INV_X2 U6889 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5162) );
  MUX2_X1 U6890 ( .A(n7145), .B(n7133), .S(n5184), .Z(n5171) );
  INV_X1 U6891 ( .A(SI_2_), .ZN(n5164) );
  NAND2_X1 U6892 ( .A1(n5171), .A2(n5164), .ZN(n5302) );
  INV_X1 U6893 ( .A(n5169), .ZN(n5166) );
  INV_X1 U6894 ( .A(SI_1_), .ZN(n5165) );
  INV_X1 U6895 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5168) );
  INV_X1 U6896 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5167) );
  INV_X1 U6897 ( .A(SI_0_), .ZN(n6304) );
  NAND3_X1 U6898 ( .A1(n5302), .A2(n5282), .A3(n5284), .ZN(n5174) );
  NAND2_X1 U6899 ( .A1(n5169), .A2(SI_1_), .ZN(n5299) );
  INV_X1 U6900 ( .A(n5299), .ZN(n5170) );
  NAND2_X1 U6901 ( .A1(n5170), .A2(n5302), .ZN(n5173) );
  INV_X1 U6902 ( .A(n5171), .ZN(n5172) );
  NAND2_X1 U6903 ( .A1(n5172), .A2(SI_2_), .ZN(n5301) );
  INV_X1 U6904 ( .A(n5180), .ZN(n5177) );
  INV_X1 U6905 ( .A(SI_3_), .ZN(n5176) );
  NAND2_X1 U6906 ( .A1(n5177), .A2(n5176), .ZN(n5321) );
  INV_X1 U6907 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7143) );
  INV_X1 U6908 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5178) );
  INV_X1 U6909 ( .A(SI_4_), .ZN(n5179) );
  NAND2_X1 U6910 ( .A1(n5181), .A2(n5179), .ZN(n5345) );
  NAND2_X1 U6911 ( .A1(n5180), .A2(SI_3_), .ZN(n5342) );
  INV_X1 U6912 ( .A(n5181), .ZN(n5182) );
  NAND2_X1 U6913 ( .A1(n5182), .A2(SI_4_), .ZN(n5344) );
  MUX2_X1 U6914 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7131), .Z(n5185) );
  INV_X1 U6915 ( .A(n5190), .ZN(n5187) );
  INV_X1 U6916 ( .A(SI_6_), .ZN(n5186) );
  NAND2_X1 U6917 ( .A1(n5187), .A2(n5186), .ZN(n5374) );
  INV_X1 U6918 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5188) );
  MUX2_X1 U6919 ( .A(n7160), .B(n5188), .S(n7131), .Z(n5192) );
  INV_X1 U6920 ( .A(SI_7_), .ZN(n5189) );
  NAND2_X1 U6921 ( .A1(n5192), .A2(n5189), .ZN(n5377) );
  NAND2_X1 U6922 ( .A1(n5190), .A2(SI_6_), .ZN(n5375) );
  INV_X1 U6923 ( .A(n5375), .ZN(n5191) );
  NAND2_X1 U6924 ( .A1(n5191), .A2(n5377), .ZN(n5194) );
  INV_X1 U6925 ( .A(n5192), .ZN(n5193) );
  NAND2_X1 U6926 ( .A1(n5193), .A2(SI_7_), .ZN(n5376) );
  XNOR2_X1 U6927 ( .A(n5197), .B(SI_8_), .ZN(n5420) );
  INV_X1 U6928 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5198) );
  MUX2_X1 U6929 ( .A(n7183), .B(n5198), .S(n7131), .Z(n5433) );
  INV_X1 U6930 ( .A(SI_9_), .ZN(n5199) );
  NAND2_X1 U6931 ( .A1(n5433), .A2(n5199), .ZN(n5449) );
  INV_X1 U6932 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5200) );
  INV_X1 U6933 ( .A(SI_10_), .ZN(n5201) );
  NAND2_X1 U6934 ( .A1(n5203), .A2(n5201), .ZN(n5452) );
  INV_X1 U6935 ( .A(n5433), .ZN(n5202) );
  NAND3_X1 U6936 ( .A1(n5452), .A2(SI_9_), .A3(n5202), .ZN(n5205) );
  INV_X1 U6937 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6938 ( .A1(n5204), .A2(SI_10_), .ZN(n5451) );
  NAND2_X1 U6939 ( .A1(n5207), .A2(SI_12_), .ZN(n5208) );
  OAI21_X1 U6940 ( .B1(n5207), .B2(SI_12_), .A(n5208), .ZN(n5492) );
  NAND2_X1 U6941 ( .A1(n5209), .A2(SI_13_), .ZN(n5213) );
  INV_X1 U6942 ( .A(n5209), .ZN(n5211) );
  INV_X1 U6943 ( .A(SI_13_), .ZN(n5210) );
  NAND2_X1 U6944 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  NAND2_X1 U6945 ( .A1(n5213), .A2(n5212), .ZN(n5523) );
  MUX2_X1 U6946 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6238), .Z(n5214) );
  NAND2_X1 U6947 ( .A1(n5214), .A2(SI_14_), .ZN(n5218) );
  INV_X1 U6948 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6949 ( .A1(n5215), .A2(n7968), .ZN(n5216) );
  NAND2_X1 U6950 ( .A1(n5218), .A2(n5216), .ZN(n5538) );
  INV_X1 U6951 ( .A(n5538), .ZN(n5217) );
  MUX2_X1 U6952 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7131), .Z(n5507) );
  INV_X1 U6953 ( .A(n5507), .ZN(n5220) );
  INV_X1 U6954 ( .A(SI_15_), .ZN(n5219) );
  NAND2_X1 U6955 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  NOR2_X1 U6956 ( .A1(n5223), .A2(n5222), .ZN(n5225) );
  NAND2_X1 U6957 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  MUX2_X1 U6958 ( .A(n7667), .B(n7195), .S(n7131), .Z(n5226) );
  INV_X1 U6959 ( .A(n5226), .ZN(n5227) );
  AOI21_X2 U6960 ( .B1(n5577), .B2(n5576), .A(n5228), .ZN(n5588) );
  MUX2_X1 U6961 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7131), .Z(n5229) );
  NAND2_X1 U6962 ( .A1(n5229), .A2(SI_18_), .ZN(n5234) );
  INV_X1 U6963 ( .A(n5229), .ZN(n5231) );
  INV_X1 U6964 ( .A(SI_18_), .ZN(n5230) );
  NAND2_X1 U6965 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  NAND2_X1 U6966 ( .A1(n5234), .A2(n5232), .ZN(n5589) );
  INV_X1 U6967 ( .A(n5589), .ZN(n5233) );
  XNOR2_X1 U6968 ( .A(n5235), .B(SI_19_), .ZN(n5605) );
  INV_X1 U6969 ( .A(n5235), .ZN(n5237) );
  INV_X1 U6970 ( .A(SI_19_), .ZN(n5236) );
  MUX2_X1 U6971 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6238), .Z(n5238) );
  XNOR2_X1 U6972 ( .A(n5238), .B(n5239), .ZN(n5615) );
  INV_X1 U6973 ( .A(n5238), .ZN(n5240) );
  INV_X1 U6974 ( .A(n5629), .ZN(n5242) );
  NAND2_X1 U6975 ( .A1(n5627), .A2(n7949), .ZN(n5241) );
  INV_X1 U6976 ( .A(n5627), .ZN(n5243) );
  NAND2_X1 U6977 ( .A1(n5243), .A2(SI_21_), .ZN(n5244) );
  MUX2_X1 U6978 ( .A(n8305), .B(n8394), .S(n7131), .Z(n5246) );
  INV_X1 U6979 ( .A(SI_22_), .ZN(n5245) );
  NAND2_X1 U6980 ( .A1(n5246), .A2(n5245), .ZN(n5273) );
  INV_X1 U6981 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6982 ( .A1(n5247), .A2(SI_22_), .ZN(n5248) );
  NAND2_X1 U6983 ( .A1(n5273), .A2(n5248), .ZN(n5637) );
  INV_X1 U6984 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5251) );
  INV_X1 U6985 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5250) );
  MUX2_X1 U6986 ( .A(n5251), .B(n5250), .S(n7131), .Z(n5253) );
  INV_X1 U6987 ( .A(SI_23_), .ZN(n5252) );
  NAND2_X1 U6988 ( .A1(n5253), .A2(n5252), .ZN(n5274) );
  NAND2_X1 U6989 ( .A1(n5652), .A2(n5650), .ZN(n5255) );
  INV_X1 U6990 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6991 ( .A1(n5254), .A2(SI_23_), .ZN(n5654) );
  MUX2_X1 U6992 ( .A(n9503), .B(n10260), .S(n6238), .Z(n5257) );
  INV_X1 U6993 ( .A(SI_24_), .ZN(n5256) );
  NAND2_X1 U6994 ( .A1(n5257), .A2(n5256), .ZN(n5653) );
  INV_X1 U6995 ( .A(n5257), .ZN(n5258) );
  NAND2_X1 U6996 ( .A1(n5258), .A2(SI_24_), .ZN(n5259) );
  NAND2_X1 U6997 ( .A1(n9501), .A2(n5365), .ZN(n5265) );
  NAND2_X1 U6998 ( .A1(n5993), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6999 ( .A1(n5643), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U7000 ( .A1(n5267), .A2(n5266), .ZN(n9209) );
  NAND2_X1 U7001 ( .A1(n9209), .A2(n5684), .ZN(n5272) );
  INV_X1 U7002 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U7003 ( .A1(n4282), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U7004 ( .A1(n5955), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5268) );
  OAI211_X1 U7005 ( .C1(n9442), .C2(n5958), .A(n5269), .B(n5268), .ZN(n5270)
         );
  INV_X1 U7006 ( .A(n5270), .ZN(n5271) );
  NAND2_X1 U7007 ( .A1(n5652), .A2(n5273), .ZN(n5276) );
  AND2_X1 U7008 ( .A1(n5274), .A2(n5654), .ZN(n5275) );
  NAND2_X1 U7009 ( .A1(n5277), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5281) );
  INV_X1 U7010 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7940) );
  OR2_X2 U7011 ( .A1(n5958), .A2(n7940), .ZN(n5280) );
  INV_X1 U7012 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10442) );
  OR2_X1 U7013 ( .A1(n5388), .A2(n10442), .ZN(n5279) );
  INV_X1 U7014 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7508) );
  OR2_X1 U7015 ( .A1(n5335), .A2(n7508), .ZN(n5278) );
  NAND2_X1 U7016 ( .A1(n5299), .A2(n5282), .ZN(n5286) );
  INV_X1 U7017 ( .A(n5286), .ZN(n5283) );
  NAND2_X1 U7018 ( .A1(n5283), .A2(n5284), .ZN(n5300) );
  INV_X1 U7019 ( .A(n5284), .ZN(n5285) );
  NAND2_X1 U7020 ( .A1(n5286), .A2(n5285), .ZN(n5287) );
  XNOR2_X2 U7021 ( .A(n5288), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7322) );
  INV_X1 U7022 ( .A(n7322), .ZN(n5289) );
  INV_X1 U7023 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5294) );
  INV_X1 U7024 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7086) );
  OR2_X1 U7025 ( .A1(n5388), .A2(n7086), .ZN(n5296) );
  INV_X1 U7026 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7242) );
  OR2_X1 U7027 ( .A1(n5356), .A2(n7242), .ZN(n5295) );
  INV_X1 U7028 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U7029 ( .A1(n4281), .A2(SI_0_), .ZN(n5298) );
  XNOR2_X1 U7030 ( .A(n5298), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9504) );
  MUX2_X1 U7031 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9504), .S(n6739), .Z(n7474) );
  NAND2_X1 U7032 ( .A1(n5786), .A2(n7474), .ZN(n7503) );
  NAND2_X1 U7033 ( .A1(n5300), .A2(n5299), .ZN(n5304) );
  NAND2_X1 U7034 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  INV_X1 U7035 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7441) );
  OR2_X1 U7036 ( .A1(n5335), .A2(n7441), .ZN(n5308) );
  INV_X1 U7037 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10444) );
  AND2_X1 U7038 ( .A1(n5308), .A2(n5307), .ZN(n5310) );
  INV_X1 U7039 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7386) );
  OR2_X1 U7040 ( .A1(n5356), .A2(n7386), .ZN(n5309) );
  INV_X1 U7041 ( .A(n6067), .ZN(n5314) );
  AND2_X1 U7042 ( .A1(n5313), .A2(n7431), .ZN(n5315) );
  INV_X1 U7043 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5316) );
  INV_X1 U7044 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U7045 ( .A1(n5342), .A2(n5321), .ZN(n5323) );
  NAND2_X1 U7046 ( .A1(n5322), .A2(n5323), .ZN(n5326) );
  INV_X1 U7047 ( .A(n5323), .ZN(n5324) );
  NAND2_X1 U7048 ( .A1(n5325), .A2(n5324), .ZN(n5343) );
  AND2_X1 U7049 ( .A1(n5326), .A2(n5343), .ZN(n7136) );
  NAND2_X1 U7050 ( .A1(n4290), .A2(n7136), .ZN(n5333) );
  NAND2_X1 U7051 ( .A1(n5380), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U7052 ( .A1(n5328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5327) );
  MUX2_X1 U7053 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5327), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5329) );
  INV_X1 U7054 ( .A(n7329), .ZN(n5330) );
  OR2_X1 U7055 ( .A1(n6739), .A2(n5330), .ZN(n5331) );
  INV_X1 U7056 ( .A(n5843), .ZN(n5857) );
  INV_X1 U7057 ( .A(n7449), .ZN(n7443) );
  INV_X1 U7058 ( .A(n7748), .ZN(n7596) );
  OR2_X1 U7059 ( .A1(n5334), .A2(n7596), .ZN(n7463) );
  NAND2_X1 U7060 ( .A1(n5354), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5341) );
  INV_X1 U7061 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10420) );
  OR2_X1 U7062 ( .A1(n5335), .A2(n10420), .ZN(n5340) );
  NAND2_X1 U7063 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5336) );
  AND2_X1 U7064 ( .A1(n5357), .A2(n5336), .ZN(n10416) );
  OR2_X1 U7065 ( .A1(n5356), .A2(n10416), .ZN(n5339) );
  INV_X1 U7066 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5337) );
  OR2_X1 U7067 ( .A1(n5958), .A2(n5337), .ZN(n5338) );
  NAND2_X1 U7068 ( .A1(n4289), .A2(n7208), .ZN(n5350) );
  NAND2_X1 U7069 ( .A1(n5380), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U7070 ( .A1(n5345), .A2(n5344), .ZN(n5346) );
  NAND2_X1 U7071 ( .A1(n7138), .A2(n5365), .ZN(n5348) );
  AND3_X2 U7072 ( .A1(n5350), .A2(n5349), .A3(n5348), .ZN(n10414) );
  AND2_X1 U7073 ( .A1(n7463), .A2(n5352), .ZN(n5351) );
  NAND2_X1 U7074 ( .A1(n7464), .A2(n5351), .ZN(n7552) );
  INV_X1 U7075 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U7076 ( .A1(n8923), .A2(n10414), .ZN(n5862) );
  OR2_X1 U7077 ( .A1(n5353), .A2(n6015), .ZN(n7551) );
  NAND2_X1 U7078 ( .A1(n5354), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5362) );
  INV_X1 U7079 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5355) );
  OR2_X1 U7080 ( .A1(n5958), .A2(n5355), .ZN(n5361) );
  NAND2_X1 U7081 ( .A1(n5357), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5358) );
  AND2_X1 U7082 ( .A1(n5397), .A2(n5358), .ZN(n7851) );
  OR2_X1 U7083 ( .A1(n5356), .A2(n7851), .ZN(n5360) );
  OR2_X1 U7084 ( .A1(n5335), .A2(n4750), .ZN(n5359) );
  XNOR2_X1 U7085 ( .A(n5364), .B(n5363), .ZN(n7140) );
  NAND2_X1 U7086 ( .A1(n7140), .A2(n5365), .ZN(n5370) );
  NAND2_X1 U7087 ( .A1(n5381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U7088 ( .A1(n4289), .A2(n7288), .ZN(n5369) );
  NAND2_X1 U7089 ( .A1(n8922), .A2(n7852), .ZN(n7632) );
  OR2_X1 U7090 ( .A1(n8922), .A2(n4512), .ZN(n5372) );
  NAND2_X1 U7091 ( .A1(n5375), .A2(n5374), .ZN(n5405) );
  NAND2_X1 U7092 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  NAND2_X1 U7093 ( .A1(n7150), .A2(n5365), .ZN(n5387) );
  INV_X1 U7094 ( .A(n5381), .ZN(n5383) );
  AND2_X2 U7095 ( .A1(n5383), .A2(n5382), .ZN(n5409) );
  NAND2_X1 U7096 ( .A1(n5422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5385) );
  AOI22_X1 U7097 ( .A1(n5993), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4289), .B2(
        n7532), .ZN(n5386) );
  NAND2_X1 U7098 ( .A1(n5387), .A2(n5386), .ZN(n8033) );
  NAND2_X1 U7099 ( .A1(n4282), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5395) );
  INV_X1 U7100 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7939) );
  OR2_X1 U7101 ( .A1(n5996), .A2(n7939), .ZN(n5394) );
  INV_X1 U7102 ( .A(n5389), .ZN(n5399) );
  NAND2_X1 U7103 ( .A1(n5399), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5390) );
  AND2_X1 U7104 ( .A1(n5426), .A2(n5390), .ZN(n7786) );
  OR2_X1 U7105 ( .A1(n5356), .A2(n7786), .ZN(n5393) );
  INV_X1 U7106 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5391) );
  OR2_X1 U7107 ( .A1(n5958), .A2(n5391), .ZN(n5392) );
  NAND4_X1 U7108 ( .A1(n5395), .A2(n5394), .A3(n5393), .A4(n5392), .ZN(n8920)
         );
  INV_X1 U7109 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5396) );
  INV_X1 U7110 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7291) );
  OR2_X1 U7111 ( .A1(n5996), .A2(n7291), .ZN(n5403) );
  NAND2_X1 U7112 ( .A1(n5397), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5398) );
  AND2_X1 U7113 ( .A1(n5399), .A2(n5398), .ZN(n7706) );
  OR2_X1 U7114 ( .A1(n5356), .A2(n7706), .ZN(n5402) );
  INV_X1 U7115 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5400) );
  OR2_X1 U7116 ( .A1(n5958), .A2(n5400), .ZN(n5401) );
  NAND2_X1 U7117 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  AND2_X1 U7118 ( .A1(n5408), .A2(n5407), .ZN(n7148) );
  NAND2_X1 U7119 ( .A1(n7148), .A2(n5365), .ZN(n5414) );
  INV_X1 U7120 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U7121 ( .A1(n5410), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5411) );
  MUX2_X1 U7122 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5411), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5412) );
  NAND2_X1 U7123 ( .A1(n5412), .A2(n5422), .ZN(n7527) );
  INV_X1 U7124 ( .A(n7527), .ZN(n7292) );
  AOI22_X1 U7125 ( .A1(n5993), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n4289), .B2(
        n7292), .ZN(n5413) );
  AOI22_X1 U7126 ( .A1(n8033), .A2(n8920), .B1(n8921), .B2(n7698), .ZN(n5415)
         );
  INV_X1 U7127 ( .A(n8033), .ZN(n7808) );
  OAI21_X1 U7128 ( .B1(n7698), .B2(n8921), .A(n8920), .ZN(n5417) );
  NOR2_X1 U7129 ( .A1(n8920), .A2(n8921), .ZN(n5416) );
  AOI22_X1 U7130 ( .A1(n7808), .A2(n5417), .B1(n5416), .B2(n10435), .ZN(n5418)
         );
  XNOR2_X1 U7131 ( .A(n5421), .B(n5420), .ZN(n7165) );
  NAND2_X1 U7132 ( .A1(n7165), .A2(n5365), .ZN(n5425) );
  NAND2_X1 U7133 ( .A1(n5434), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5423) );
  XNOR2_X1 U7134 ( .A(n5423), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7821) );
  AOI22_X1 U7135 ( .A1(n5993), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4289), .B2(
        n7821), .ZN(n5424) );
  NAND2_X1 U7136 ( .A1(n5425), .A2(n5424), .ZN(n8166) );
  NAND2_X1 U7137 ( .A1(n5955), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5431) );
  INV_X1 U7138 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7820) );
  OR2_X1 U7139 ( .A1(n5335), .A2(n7820), .ZN(n5430) );
  NAND2_X1 U7140 ( .A1(n5426), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5427) );
  AND2_X1 U7141 ( .A1(n5438), .A2(n5427), .ZN(n8169) );
  OR2_X1 U7142 ( .A1(n5356), .A2(n8169), .ZN(n5429) );
  INV_X1 U7143 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7616) );
  OR2_X1 U7144 ( .A1(n5958), .A2(n7616), .ZN(n5428) );
  NAND4_X1 U7145 ( .A1(n5431), .A2(n5430), .A3(n5429), .A4(n5428), .ZN(n8919)
         );
  NAND2_X1 U7146 ( .A1(n8166), .A2(n8919), .ZN(n5432) );
  XNOR2_X1 U7147 ( .A(n5433), .B(SI_9_), .ZN(n5447) );
  NAND2_X1 U7148 ( .A1(n7174), .A2(n5365), .ZN(n5437) );
  NAND2_X1 U7149 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U7150 ( .A(n5435), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7826) );
  AOI22_X1 U7151 ( .A1(n5993), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4289), .B2(
        n7826), .ZN(n5436) );
  NAND2_X1 U7152 ( .A1(n5955), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5444) );
  INV_X1 U7153 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7910) );
  OR2_X1 U7154 ( .A1(n5335), .A2(n7910), .ZN(n5443) );
  NAND2_X1 U7155 ( .A1(n5438), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5439) );
  AND2_X1 U7156 ( .A1(n5461), .A2(n5439), .ZN(n8272) );
  OR2_X1 U7157 ( .A1(n5356), .A2(n8272), .ZN(n5442) );
  INV_X1 U7158 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5440) );
  OR2_X1 U7159 ( .A1(n5958), .A2(n5440), .ZN(n5441) );
  NAND2_X1 U7160 ( .A1(n8269), .A2(n8164), .ZN(n5874) );
  OR2_X1 U7161 ( .A1(n8269), .A2(n8918), .ZN(n5446) );
  NAND2_X1 U7162 ( .A1(n7759), .A2(n5446), .ZN(n8027) );
  NAND2_X1 U7163 ( .A1(n5448), .A2(n5447), .ZN(n5450) );
  NAND2_X1 U7164 ( .A1(n5450), .A2(n5449), .ZN(n5454) );
  AND2_X1 U7165 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  XNOR2_X1 U7166 ( .A(n5454), .B(n5453), .ZN(n7180) );
  NAND2_X1 U7167 ( .A1(n7180), .A2(n5365), .ZN(n5460) );
  INV_X1 U7168 ( .A(n5455), .ZN(n5457) );
  INV_X1 U7169 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7170 ( .A1(n5457), .A2(n5456), .ZN(n5473) );
  NAND2_X1 U7171 ( .A1(n5473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5458) );
  AOI22_X1 U7172 ( .A1(n8253), .A2(n4289), .B1(n5993), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7173 ( .A1(n4282), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5467) );
  INV_X1 U7174 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8252) );
  OR2_X1 U7175 ( .A1(n5996), .A2(n8252), .ZN(n5466) );
  NAND2_X1 U7176 ( .A1(n5461), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5462) );
  AND2_X1 U7177 ( .A1(n5482), .A2(n5462), .ZN(n8755) );
  OR2_X1 U7178 ( .A1(n5356), .A2(n8755), .ZN(n5465) );
  INV_X1 U7179 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5463) );
  OR2_X1 U7180 ( .A1(n5958), .A2(n5463), .ZN(n5464) );
  NAND4_X1 U7181 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n8917)
         );
  NAND2_X1 U7182 ( .A1(n8215), .A2(n8917), .ZN(n5468) );
  NAND2_X1 U7183 ( .A1(n8027), .A2(n5468), .ZN(n5470) );
  OR2_X1 U7184 ( .A1(n8215), .A2(n8917), .ZN(n5469) );
  NAND2_X1 U7185 ( .A1(n5470), .A2(n5469), .ZN(n8194) );
  XNOR2_X1 U7186 ( .A(n5472), .B(n5471), .ZN(n7197) );
  NAND2_X1 U7187 ( .A1(n7197), .A2(n5365), .ZN(n5480) );
  INV_X1 U7188 ( .A(n5473), .ZN(n5475) );
  INV_X1 U7189 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7190 ( .A1(n5475), .A2(n5474), .ZN(n5477) );
  NAND2_X1 U7191 ( .A1(n5477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5476) );
  MUX2_X1 U7192 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5476), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5478) );
  AOI22_X1 U7193 ( .A1(n8331), .A2(n4289), .B1(n5993), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U7194 ( .A1(n5480), .A2(n5479), .ZN(n5885) );
  NAND2_X1 U7195 ( .A1(n4282), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5488) );
  INV_X1 U7196 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5481) );
  OR2_X1 U7197 ( .A1(n5996), .A2(n5481), .ZN(n5487) );
  NAND2_X1 U7198 ( .A1(n5482), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5483) );
  AND2_X1 U7199 ( .A1(n5499), .A2(n5483), .ZN(n8870) );
  OR2_X1 U7200 ( .A1(n5356), .A2(n8870), .ZN(n5486) );
  INV_X1 U7201 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5484) );
  OR2_X1 U7202 ( .A1(n5958), .A2(n5484), .ZN(n5485) );
  OR2_X1 U7203 ( .A1(n5885), .A2(n8784), .ZN(n5489) );
  NAND2_X1 U7204 ( .A1(n5885), .A2(n8784), .ZN(n5795) );
  NAND2_X1 U7205 ( .A1(n5885), .A2(n8916), .ZN(n5491) );
  NAND2_X1 U7206 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  AND2_X1 U7207 ( .A1(n5495), .A2(n5494), .ZN(n7219) );
  NAND2_X1 U7208 ( .A1(n7219), .A2(n5365), .ZN(n5498) );
  NAND2_X1 U7209 ( .A1(n4315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5496) );
  AOI22_X1 U7210 ( .A1(n8986), .A2(n4289), .B1(n5993), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7211 ( .A1(n4282), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5504) );
  INV_X1 U7212 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8336) );
  OR2_X1 U7213 ( .A1(n5996), .A2(n8336), .ZN(n5503) );
  NAND2_X1 U7214 ( .A1(n5499), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5500) );
  AND2_X1 U7215 ( .A1(n5531), .A2(n5500), .ZN(n8310) );
  OR2_X1 U7216 ( .A1(n5356), .A2(n8310), .ZN(n5502) );
  INV_X1 U7217 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8296) );
  OR2_X1 U7218 ( .A1(n5958), .A2(n8296), .ZN(n5501) );
  NAND2_X1 U7219 ( .A1(n8311), .A2(n8915), .ZN(n5505) );
  XNOR2_X1 U7220 ( .A(n5507), .B(SI_15_), .ZN(n5508) );
  XNOR2_X1 U7221 ( .A(n5509), .B(n5508), .ZN(n7496) );
  NAND2_X1 U7222 ( .A1(n7496), .A2(n5365), .ZN(n5514) );
  OAI21_X2 U7223 ( .B1(n4315), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5527) );
  INV_X1 U7224 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7225 ( .A1(n5527), .A2(n5510), .ZN(n5511) );
  NAND2_X1 U7226 ( .A1(n5511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5543) );
  INV_X1 U7227 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7228 ( .A1(n5543), .A2(n5542), .ZN(n5545) );
  NAND2_X1 U7229 ( .A1(n5545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U7230 ( .A(n5512), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9054) );
  AOI22_X1 U7231 ( .A1(n9054), .A2(n4289), .B1(n5993), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5513) );
  INV_X1 U7232 ( .A(n5515), .ZN(n5550) );
  NAND2_X1 U7233 ( .A1(n5550), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7234 ( .A1(n5571), .A2(n5516), .ZN(n9324) );
  NAND2_X1 U7235 ( .A1(n9324), .A2(n5684), .ZN(n5521) );
  NAND2_X1 U7236 ( .A1(n5955), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7237 ( .A1(n5517), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7238 ( .A1(n4282), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5518) );
  NAND4_X1 U7239 ( .A1(n5521), .A2(n5520), .A3(n5519), .A4(n5518), .ZN(n9334)
         );
  NAND2_X1 U7240 ( .A1(n9477), .A2(n9334), .ZN(n5557) );
  INV_X1 U7241 ( .A(n5522), .ZN(n5524) );
  NAND2_X1 U7242 ( .A1(n5524), .A2(n5523), .ZN(n5526) );
  NAND2_X1 U7243 ( .A1(n7338), .A2(n5365), .ZN(n5529) );
  XNOR2_X1 U7244 ( .A(n5527), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8980) );
  AOI22_X1 U7245 ( .A1(n8980), .A2(n4289), .B1(n5993), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U7246 ( .A1(n4282), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5536) );
  INV_X1 U7247 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8976) );
  OR2_X1 U7248 ( .A1(n5996), .A2(n8976), .ZN(n5535) );
  INV_X1 U7249 ( .A(n5530), .ZN(n5548) );
  NAND2_X1 U7250 ( .A1(n5531), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5532) );
  AND2_X1 U7251 ( .A1(n5548), .A2(n5532), .ZN(n8851) );
  OR2_X1 U7252 ( .A1(n5356), .A2(n8851), .ZN(n5534) );
  INV_X1 U7253 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8321) );
  OR2_X1 U7254 ( .A1(n5958), .A2(n8321), .ZN(n5533) );
  NAND2_X1 U7255 ( .A1(n8368), .A2(n8789), .ZN(n9314) );
  NAND2_X1 U7256 ( .A1(n8854), .A2(n9332), .ZN(n5896) );
  INV_X1 U7257 ( .A(n5537), .ZN(n5539) );
  NAND2_X1 U7258 ( .A1(n5539), .A2(n5538), .ZN(n5541) );
  NAND2_X1 U7259 ( .A1(n5541), .A2(n5540), .ZN(n7400) );
  OR2_X1 U7260 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  AND2_X2 U7261 ( .A1(n5545), .A2(n5544), .ZN(n9031) );
  NAND2_X1 U7262 ( .A1(n5548), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7263 ( .A1(n5550), .A2(n5549), .ZN(n9340) );
  NAND2_X1 U7264 ( .A1(n5684), .A2(n9340), .ZN(n5554) );
  INV_X1 U7265 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9022) );
  OR2_X1 U7266 ( .A1(n5335), .A2(n9022), .ZN(n5553) );
  INV_X1 U7267 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9405) );
  OR2_X1 U7268 ( .A1(n5996), .A2(n9405), .ZN(n5552) );
  INV_X1 U7269 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9483) );
  OR2_X1 U7270 ( .A1(n5958), .A2(n9483), .ZN(n5551) );
  NAND4_X1 U7271 ( .A1(n5554), .A2(n5553), .A3(n5552), .A4(n5551), .ZN(n9320)
         );
  NAND2_X1 U7272 ( .A1(n9484), .A2(n9320), .ZN(n9317) );
  NAND3_X1 U7273 ( .A1(n5557), .A2(n8322), .A3(n9317), .ZN(n5560) );
  NAND2_X1 U7274 ( .A1(n9314), .A2(n9320), .ZN(n5555) );
  INV_X1 U7275 ( .A(n9314), .ZN(n5893) );
  INV_X1 U7276 ( .A(n9320), .ZN(n9316) );
  AOI22_X1 U7277 ( .A1(n9338), .A2(n5555), .B1(n5893), .B2(n9316), .ZN(n5556)
         );
  OAI21_X1 U7278 ( .B1(n9334), .B2(n9477), .A(n5556), .ZN(n5558) );
  NAND2_X1 U7279 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  XNOR2_X1 U7280 ( .A(n5561), .B(SI_16_), .ZN(n5562) );
  XNOR2_X1 U7281 ( .A(n5563), .B(n5562), .ZN(n7558) );
  NAND2_X1 U7282 ( .A1(n7558), .A2(n5365), .ZN(n5570) );
  NOR2_X1 U7283 ( .A1(n5564), .A2(n5565), .ZN(n5566) );
  NAND2_X1 U7284 ( .A1(n5567), .A2(n5566), .ZN(n5578) );
  NAND2_X1 U7285 ( .A1(n5578), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5568) );
  XNOR2_X1 U7286 ( .A(n5568), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9074) );
  AOI22_X1 U7287 ( .A1(n5993), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4289), .B2(
        n9074), .ZN(n5569) );
  NAND2_X1 U7288 ( .A1(n5571), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7289 ( .A1(n5582), .A2(n5572), .ZN(n9305) );
  NAND2_X1 U7290 ( .A1(n9305), .A2(n5684), .ZN(n5575) );
  AOI22_X1 U7291 ( .A1(n5517), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n5955), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U7292 ( .A1(n4282), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7293 ( .A1(n9471), .A2(n9295), .ZN(n5905) );
  INV_X1 U7294 ( .A(n9471), .ZN(n8816) );
  XNOR2_X1 U7295 ( .A(n5577), .B(n5576), .ZN(n7621) );
  NAND2_X1 U7296 ( .A1(n7621), .A2(n5365), .ZN(n5581) );
  OAI21_X1 U7297 ( .B1(n5578), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5579) );
  XNOR2_X1 U7298 ( .A(n5579), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9097) );
  AOI22_X1 U7299 ( .A1(n5993), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4289), .B2(
        n9097), .ZN(n5580) );
  NAND2_X1 U7300 ( .A1(n5582), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7301 ( .A1(n5597), .A2(n5583), .ZN(n9299) );
  NAND2_X1 U7302 ( .A1(n9299), .A2(n5684), .ZN(n5586) );
  AOI22_X1 U7303 ( .A1(n5517), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n5955), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7304 ( .A1(n4282), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7305 ( .A1(n9393), .A2(n8812), .ZN(n5799) );
  NAND2_X1 U7306 ( .A1(n9393), .A2(n9308), .ZN(n5587) );
  INV_X1 U7307 ( .A(n5588), .ZN(n5590) );
  NAND2_X1 U7308 ( .A1(n5590), .A2(n5589), .ZN(n5591) );
  NAND2_X1 U7309 ( .A1(n5592), .A2(n5591), .ZN(n7668) );
  NAND2_X1 U7310 ( .A1(n5593), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5594) );
  XNOR2_X1 U7311 ( .A(n5594), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9133) );
  AOI22_X1 U7312 ( .A1(n5993), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4289), .B2(
        n9133), .ZN(n5595) );
  NAND2_X1 U7313 ( .A1(n5597), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7314 ( .A1(n5610), .A2(n5598), .ZN(n9277) );
  NAND2_X1 U7315 ( .A1(n9277), .A2(n5684), .ZN(n5604) );
  INV_X1 U7316 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7317 ( .A1(n5955), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7318 ( .A1(n4282), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5599) );
  OAI211_X1 U7319 ( .C1(n5958), .C2(n5601), .A(n5600), .B(n5599), .ZN(n5602)
         );
  INV_X1 U7320 ( .A(n5602), .ZN(n5603) );
  NAND2_X1 U7321 ( .A1(n5604), .A2(n5603), .ZN(n9260) );
  NAND2_X1 U7322 ( .A1(n7837), .A2(n5365), .ZN(n5609) );
  AOI22_X1 U7323 ( .A1(n5993), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6053), .B2(
        n4289), .ZN(n5608) );
  NAND2_X1 U7324 ( .A1(n5610), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7325 ( .A1(n5618), .A2(n5611), .ZN(n9266) );
  INV_X1 U7326 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U7327 ( .A1(n5955), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7328 ( .A1(n5517), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7329 ( .C1(n5335), .C2(n9268), .A(n5613), .B(n5612), .ZN(n5614)
         );
  AOI21_X1 U7330 ( .B1(n9266), .B2(n5684), .A(n5614), .ZN(n9247) );
  NAND2_X1 U7331 ( .A1(n9270), .A2(n9247), .ZN(n5918) );
  NAND2_X1 U7332 ( .A1(n9232), .A2(n5918), .ZN(n9259) );
  INV_X1 U7333 ( .A(n9247), .ZN(n9275) );
  NAND2_X1 U7334 ( .A1(n8102), .A2(n5365), .ZN(n5617) );
  NAND2_X1 U7335 ( .A1(n5993), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7336 ( .A1(n5618), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7337 ( .A1(n5632), .A2(n5619), .ZN(n9252) );
  NAND2_X1 U7338 ( .A1(n9252), .A2(n5684), .ZN(n5624) );
  INV_X1 U7339 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U7340 ( .A1(n4282), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7341 ( .A1(n5955), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5620) );
  OAI211_X1 U7342 ( .C1(n9459), .C2(n5958), .A(n5621), .B(n5620), .ZN(n5622)
         );
  INV_X1 U7343 ( .A(n5622), .ZN(n5623) );
  NAND2_X1 U7344 ( .A1(n8835), .A2(n9227), .ZN(n9234) );
  XNOR2_X1 U7345 ( .A(n5627), .B(SI_21_), .ZN(n5628) );
  XNOR2_X1 U7346 ( .A(n5629), .B(n5628), .ZN(n8223) );
  NAND2_X1 U7347 ( .A1(n8223), .A2(n5365), .ZN(n5631) );
  NAND2_X1 U7348 ( .A1(n5993), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7349 ( .A1(n5632), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7350 ( .A1(n5641), .A2(n5633), .ZN(n9228) );
  INV_X1 U7351 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U7352 ( .A1(n4282), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7353 ( .A1(n5955), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5634) );
  OAI211_X1 U7354 ( .C1(n9453), .C2(n5958), .A(n5635), .B(n5634), .ZN(n5636)
         );
  NAND2_X1 U7355 ( .A1(n9454), .A2(n9248), .ZN(n5923) );
  NAND2_X1 U7356 ( .A1(n5922), .A2(n5923), .ZN(n9237) );
  INV_X1 U7357 ( .A(n9454), .ZN(n9373) );
  XNOR2_X1 U7358 ( .A(n5638), .B(n5637), .ZN(n8303) );
  NAND2_X1 U7359 ( .A1(n8303), .A2(n5365), .ZN(n5640) );
  NAND2_X1 U7360 ( .A1(n5993), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7361 ( .A1(n5641), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7362 ( .A1(n5643), .A2(n5642), .ZN(n9219) );
  NAND2_X1 U7363 ( .A1(n9219), .A2(n5684), .ZN(n5648) );
  INV_X1 U7364 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U7365 ( .A1(n5955), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7366 ( .A1(n4282), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5644) );
  OAI211_X1 U7367 ( .C1(n5958), .C2(n9448), .A(n5645), .B(n5644), .ZN(n5646)
         );
  INV_X1 U7368 ( .A(n5646), .ZN(n5647) );
  XNOR2_X1 U7369 ( .A(n9370), .B(n9206), .ZN(n9215) );
  NAND2_X1 U7370 ( .A1(n9190), .A2(n8746), .ZN(n5649) );
  AND2_X1 U7371 ( .A1(n5650), .A2(n5653), .ZN(n5651) );
  NAND2_X1 U7372 ( .A1(n5652), .A2(n5651), .ZN(n5659) );
  INV_X1 U7373 ( .A(n5653), .ZN(n5657) );
  INV_X1 U7374 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8451) );
  INV_X1 U7375 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10256) );
  MUX2_X1 U7376 ( .A(n8451), .B(n10256), .S(n6238), .Z(n5661) );
  INV_X1 U7377 ( .A(SI_25_), .ZN(n5660) );
  NAND2_X1 U7378 ( .A1(n5661), .A2(n5660), .ZN(n5692) );
  INV_X1 U7379 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7380 ( .A1(n5662), .A2(SI_25_), .ZN(n5663) );
  NAND2_X1 U7381 ( .A1(n8450), .A2(n5365), .ZN(n5665) );
  NAND2_X1 U7382 ( .A1(n5993), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5664) );
  INV_X1 U7383 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7384 ( .A1(n5668), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7385 ( .A1(n5682), .A2(n5669), .ZN(n9185) );
  NAND2_X1 U7386 ( .A1(n9185), .A2(n5684), .ZN(n5674) );
  INV_X1 U7387 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U7388 ( .A1(n4282), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7389 ( .A1(n5955), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5670) );
  OAI211_X1 U7390 ( .C1(n9430), .C2(n5958), .A(n5671), .B(n5670), .ZN(n5672)
         );
  INV_X1 U7391 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U7392 ( .A1(n9431), .A2(n8890), .ZN(n5937) );
  NAND2_X1 U7393 ( .A1(n5931), .A2(n5937), .ZN(n9187) );
  INV_X1 U7394 ( .A(n9431), .ZN(n9179) );
  NAND2_X1 U7395 ( .A1(n5694), .A2(n5692), .ZN(n5681) );
  INV_X1 U7396 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9499) );
  INV_X1 U7397 ( .A(SI_26_), .ZN(n5677) );
  NAND2_X1 U7398 ( .A1(n5678), .A2(n5677), .ZN(n5691) );
  INV_X1 U7399 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U7400 ( .A1(n5679), .A2(SI_26_), .ZN(n5713) );
  AND2_X1 U7401 ( .A1(n5691), .A2(n5713), .ZN(n5680) );
  OR2_X2 U7402 ( .A1(n5682), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7403 ( .A1(n5682), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7404 ( .A1(n5705), .A2(n5683), .ZN(n9175) );
  NAND2_X1 U7405 ( .A1(n9175), .A2(n5684), .ZN(n5689) );
  INV_X1 U7406 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U7407 ( .A1(n5955), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7408 ( .A1(n4282), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5685) );
  OAI211_X1 U7409 ( .C1(n5958), .C2(n9424), .A(n5686), .B(n5685), .ZN(n5687)
         );
  INV_X1 U7410 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U7411 ( .A1(n6145), .A2(n8800), .ZN(n5690) );
  AOI22_X2 U7412 ( .A1(n9171), .A2(n5690), .B1(n9425), .B2(n9181), .ZN(n6200)
         );
  INV_X1 U7413 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5695) );
  INV_X1 U7414 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10252) );
  MUX2_X1 U7415 ( .A(n5695), .B(n10252), .S(n7131), .Z(n5697) );
  INV_X1 U7416 ( .A(SI_27_), .ZN(n5696) );
  NAND2_X1 U7417 ( .A1(n5697), .A2(n5696), .ZN(n5829) );
  INV_X1 U7418 ( .A(n5697), .ZN(n5698) );
  NAND2_X1 U7419 ( .A1(n5698), .A2(SI_27_), .ZN(n5699) );
  NAND2_X1 U7420 ( .A1(n9493), .A2(n5365), .ZN(n5702) );
  NAND2_X1 U7421 ( .A1(n5993), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5701) );
  INV_X1 U7422 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7423 ( .A1(n5705), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7424 ( .A1(n5721), .A2(n5706), .ZN(n9163) );
  NAND2_X1 U7425 ( .A1(n9163), .A2(n5684), .ZN(n5711) );
  INV_X1 U7426 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7427 ( .A1(n4282), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7428 ( .A1(n5955), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5707) );
  OAI211_X1 U7429 ( .C1(n6219), .C2(n5958), .A(n5708), .B(n5707), .ZN(n5709)
         );
  INV_X1 U7430 ( .A(n5709), .ZN(n5710) );
  NOR2_X1 U7431 ( .A1(n6218), .A2(n9172), .ZN(n5807) );
  NAND2_X1 U7432 ( .A1(n6218), .A2(n9172), .ZN(n5808) );
  OAI21_X2 U7433 ( .B1(n6200), .B2(n5807), .A(n5808), .ZN(n6746) );
  INV_X1 U7434 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5716) );
  INV_X1 U7435 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8430) );
  XNOR2_X1 U7436 ( .A(n5828), .B(SI_28_), .ZN(n5943) );
  NAND2_X1 U7437 ( .A1(n8428), .A2(n5365), .ZN(n5718) );
  NAND2_X1 U7438 ( .A1(n5993), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5717) );
  INV_X1 U7439 ( .A(n5721), .ZN(n5720) );
  INV_X1 U7440 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5719) );
  INV_X1 U7441 ( .A(n9148), .ZN(n5723) );
  NAND2_X1 U7442 ( .A1(n5721), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U7443 ( .A1(n5723), .A2(n5722), .ZN(n6182) );
  NAND2_X1 U7444 ( .A1(n6182), .A2(n5684), .ZN(n5728) );
  INV_X1 U7445 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7979) );
  NAND2_X1 U7446 ( .A1(n5517), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7447 ( .A1(n5955), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5724) );
  OAI211_X1 U7448 ( .C1(n5335), .C2(n7979), .A(n5725), .B(n5724), .ZN(n5726)
         );
  INV_X1 U7449 ( .A(n5726), .ZN(n5727) );
  NAND2_X2 U7450 ( .A1(n5728), .A2(n5727), .ZN(n8913) );
  XNOR2_X1 U7451 ( .A(n9419), .B(n8913), .ZN(n5811) );
  XNOR2_X1 U7452 ( .A(n6746), .B(n5811), .ZN(n5742) );
  NAND2_X1 U7453 ( .A1(n4316), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7454 ( .A1(n6054), .A2(n6053), .ZN(n6154) );
  NAND2_X1 U7455 ( .A1(n4386), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5730) );
  MUX2_X1 U7456 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5730), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5731) );
  NAND2_X1 U7457 ( .A1(n4373), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5733) );
  XNOR2_X2 U7458 ( .A(n5733), .B(n5732), .ZN(n8104) );
  NAND2_X1 U7459 ( .A1(n5969), .A2(n6040), .ZN(n6049) );
  INV_X1 U7460 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U7461 ( .A1(n5955), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7462 ( .A1(n4282), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U7463 ( .C1(n5958), .C2(n6775), .A(n5735), .B(n5734), .ZN(n5736)
         );
  INV_X1 U7464 ( .A(n5736), .ZN(n5737) );
  INV_X1 U7465 ( .A(n6187), .ZN(n8912) );
  AND2_X4 U7466 ( .A1(n6054), .A2(n5969), .ZN(n7082) );
  INV_X1 U7467 ( .A(n7120), .ZN(n7092) );
  NAND2_X1 U7468 ( .A1(n7092), .A2(n7116), .ZN(n5738) );
  NAND2_X1 U7469 ( .A1(n6739), .A2(n5738), .ZN(n6183) );
  INV_X1 U7470 ( .A(n6183), .ZN(n6170) );
  AOI21_X1 U7471 ( .B1(n5742), .B2(n9336), .A(n5741), .ZN(n9417) );
  NAND2_X1 U7472 ( .A1(n5744), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5746) );
  INV_X1 U7473 ( .A(n5744), .ZN(n5745) );
  XNOR2_X1 U7474 ( .A(n5755), .B(P2_B_REG_SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7475 ( .A1(n5750), .A2(n5758), .ZN(n5754) );
  MUX2_X1 U7476 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5751), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5752) );
  NAND2_X1 U7477 ( .A1(n5755), .A2(n9500), .ZN(n7177) );
  NAND2_X1 U7478 ( .A1(n5758), .A2(n9500), .ZN(n5759) );
  NOR2_X1 U7479 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n7926) );
  NOR4_X1 U7480 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5763) );
  NOR4_X1 U7481 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5762) );
  NOR4_X1 U7482 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5761) );
  NAND4_X1 U7483 ( .A1(n7926), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n5769)
         );
  NOR4_X1 U7484 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5767) );
  NOR4_X1 U7485 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5766) );
  NOR4_X1 U7486 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5765) );
  NOR4_X1 U7487 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5764) );
  NAND4_X1 U7488 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n5768)
         );
  NOR2_X1 U7489 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  INV_X1 U7490 ( .A(n5758), .ZN(n5772) );
  NOR2_X1 U7491 ( .A1(n5755), .A2(n9500), .ZN(n5771) );
  INV_X1 U7492 ( .A(n5814), .ZN(n6059) );
  NAND2_X1 U7493 ( .A1(n7082), .A2(n6059), .ZN(n5775) );
  AND2_X1 U7494 ( .A1(n5775), .A2(n7081), .ZN(n5776) );
  NAND3_X1 U7495 ( .A1(n6157), .A2(P2_STATE_REG_SCAN_IN), .A3(n6174), .ZN(
        n5777) );
  INV_X1 U7496 ( .A(n6768), .ZN(n5783) );
  NOR2_X1 U7497 ( .A1(n8104), .A2(n6053), .ZN(n5778) );
  AND2_X1 U7498 ( .A1(n6054), .A2(n5778), .ZN(n5779) );
  INV_X1 U7499 ( .A(n6761), .ZN(n6763) );
  NAND2_X1 U7500 ( .A1(n6062), .A2(n6763), .ZN(n5781) );
  NAND2_X1 U7501 ( .A1(n6764), .A2(n6761), .ZN(n5780) );
  NAND2_X1 U7502 ( .A1(n9417), .A2(n10421), .ZN(n5785) );
  NAND2_X1 U7503 ( .A1(n10413), .A2(n7979), .ZN(n5784) );
  NAND2_X1 U7504 ( .A1(n5785), .A2(n5784), .ZN(n5819) );
  INV_X1 U7505 ( .A(n5847), .ZN(n5787) );
  NAND2_X1 U7506 ( .A1(n5787), .A2(n5844), .ZN(n5790) );
  INV_X1 U7507 ( .A(n5848), .ZN(n5788) );
  NAND2_X1 U7508 ( .A1(n5788), .A2(n5844), .ZN(n5789) );
  NAND2_X1 U7509 ( .A1(n10435), .A2(n8921), .ZN(n5791) );
  AND2_X1 U7510 ( .A1(n7632), .A2(n5791), .ZN(n5859) );
  NAND2_X1 U7511 ( .A1(n8037), .A2(n7698), .ZN(n5858) );
  INV_X1 U7512 ( .A(n5791), .ZN(n5865) );
  INV_X1 U7513 ( .A(n8920), .ZN(n6081) );
  OR2_X1 U7514 ( .A1(n8033), .A2(n6081), .ZN(n7613) );
  NAND2_X1 U7515 ( .A1(n8033), .A2(n6081), .ZN(n5873) );
  NAND2_X1 U7516 ( .A1(n7643), .A2(n7648), .ZN(n7645) );
  INV_X1 U7517 ( .A(n8166), .ZN(n7617) );
  NAND2_X1 U7518 ( .A1(n7617), .A2(n8919), .ZN(n6013) );
  AND2_X1 U7519 ( .A1(n6013), .A2(n7613), .ZN(n5872) );
  INV_X1 U7520 ( .A(n8919), .ZN(n6088) );
  NAND2_X1 U7521 ( .A1(n8166), .A2(n6088), .ZN(n6012) );
  OR2_X1 U7522 ( .A1(n8215), .A2(n8751), .ZN(n5879) );
  NAND2_X1 U7523 ( .A1(n8215), .A2(n8751), .ZN(n5877) );
  NAND2_X1 U7524 ( .A1(n5879), .A2(n5877), .ZN(n8026) );
  NAND2_X1 U7525 ( .A1(n8024), .A2(n5877), .ZN(n8201) );
  NAND2_X1 U7526 ( .A1(n8790), .A2(n8915), .ZN(n5889) );
  NAND2_X1 U7527 ( .A1(n8311), .A2(n8873), .ZN(n5886) );
  NAND2_X1 U7528 ( .A1(n5889), .A2(n5886), .ZN(n8298) );
  NOR2_X1 U7529 ( .A1(n8854), .A2(n8789), .ZN(n5796) );
  NAND2_X1 U7530 ( .A1(n8854), .A2(n8789), .ZN(n5797) );
  NAND2_X1 U7531 ( .A1(n9338), .A2(n9320), .ZN(n5897) );
  NAND2_X1 U7532 ( .A1(n9477), .A2(n6108), .ZN(n5906) );
  INV_X1 U7533 ( .A(n5905), .ZN(n9287) );
  INV_X1 U7534 ( .A(n5799), .ZN(n5901) );
  AND2_X2 U7535 ( .A1(n9281), .A2(n9297), .ZN(n6009) );
  AND2_X1 U7536 ( .A1(n5923), .A2(n9234), .ZN(n5920) );
  INV_X1 U7537 ( .A(n5918), .ZN(n5801) );
  NAND2_X1 U7538 ( .A1(n9233), .A2(n5801), .ZN(n5802) );
  NAND2_X1 U7539 ( .A1(n5803), .A2(n5922), .ZN(n9216) );
  OR2_X1 U7540 ( .A1(n9370), .A2(n9226), .ZN(n5840) );
  INV_X1 U7541 ( .A(n6008), .ZN(n5805) );
  NAND2_X1 U7542 ( .A1(n9443), .A2(n9214), .ZN(n6007) );
  NAND2_X1 U7543 ( .A1(n9437), .A2(n8746), .ZN(n6005) );
  INV_X1 U7544 ( .A(n5931), .ZN(n5806) );
  INV_X1 U7545 ( .A(n5807), .ZN(n5809) );
  INV_X1 U7546 ( .A(n9172), .ZN(n8894) );
  INV_X1 U7547 ( .A(n5811), .ZN(n6029) );
  XNOR2_X1 U7548 ( .A(n6045), .B(n6029), .ZN(n9420) );
  NAND2_X1 U7549 ( .A1(n5969), .A2(n5816), .ZN(n5812) );
  OAI211_X1 U7550 ( .C1(n6054), .C2(n8104), .A(n10434), .B(n9130), .ZN(n5813)
         );
  INV_X1 U7551 ( .A(n5813), .ZN(n5815) );
  NAND2_X1 U7552 ( .A1(n5815), .A2(n6211), .ZN(n7653) );
  NAND2_X1 U7553 ( .A1(n9159), .A2(n7653), .ZN(n10411) );
  NAND2_X1 U7554 ( .A1(n9420), .A2(n9283), .ZN(n5818) );
  AOI22_X1 U7555 ( .A1(n9419), .A2(n9325), .B1(n9341), .B2(n6182), .ZN(n5817)
         );
  NAND2_X1 U7556 ( .A1(n5819), .A2(n5117), .ZN(P2_U3205) );
  INV_X1 U7557 ( .A(n5828), .ZN(n5821) );
  NAND2_X1 U7558 ( .A1(n5821), .A2(SI_28_), .ZN(n5820) );
  MUX2_X1 U7559 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6238), .Z(n5945) );
  INV_X1 U7560 ( .A(n5945), .ZN(n5822) );
  NAND2_X1 U7561 ( .A1(n5820), .A2(n5822), .ZN(n5832) );
  INV_X1 U7562 ( .A(n5832), .ZN(n5826) );
  INV_X1 U7563 ( .A(n5829), .ZN(n5825) );
  INV_X1 U7564 ( .A(SI_28_), .ZN(n5827) );
  OAI21_X1 U7565 ( .B1(n5822), .B2(n5827), .A(n5821), .ZN(n5824) );
  OAI21_X1 U7566 ( .B1(n5945), .B2(SI_28_), .A(n5828), .ZN(n5823) );
  AOI22_X1 U7567 ( .A1(n5826), .A2(n5825), .B1(n5824), .B2(n5823), .ZN(n5831)
         );
  NAND2_X1 U7568 ( .A1(n5828), .A2(n5827), .ZN(n5946) );
  NAND4_X1 U7569 ( .A1(n5833), .A2(n5945), .A3(n5829), .A4(n5946), .ZN(n5830)
         );
  XNOR2_X1 U7570 ( .A(n5942), .B(SI_29_), .ZN(n8388) );
  NAND2_X1 U7571 ( .A1(n8388), .A2(n5365), .ZN(n5835) );
  NAND2_X1 U7572 ( .A1(n5993), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7573 ( .A1(n5835), .A2(n5834), .ZN(n6769) );
  NAND2_X1 U7574 ( .A1(n6769), .A2(n6187), .ZN(n5962) );
  MUX2_X1 U7575 ( .A(n9172), .B(n7082), .S(n6218), .Z(n5837) );
  NAND2_X1 U7576 ( .A1(n9172), .A2(n7082), .ZN(n5836) );
  OAI21_X1 U7577 ( .B1(n7082), .B2(n5937), .A(n6003), .ZN(n5838) );
  OAI21_X1 U7578 ( .B1(n7082), .B2(n6003), .A(n5838), .ZN(n5935) );
  NAND2_X1 U7579 ( .A1(n9370), .A2(n9226), .ZN(n5839) );
  AND2_X1 U7580 ( .A1(n6007), .A2(n5839), .ZN(n5842) );
  NOR2_X1 U7581 ( .A1(n6008), .A2(n5006), .ZN(n5841) );
  NAND2_X1 U7582 ( .A1(n5861), .A2(n7444), .ZN(n5846) );
  NAND2_X1 U7583 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  MUX2_X1 U7584 ( .A(n5846), .B(n5845), .S(n7082), .Z(n5855) );
  NAND2_X1 U7585 ( .A1(n7430), .A2(n7433), .ZN(n7445) );
  NAND2_X1 U7586 ( .A1(n5786), .A2(n7757), .ZN(n6014) );
  NAND2_X1 U7587 ( .A1(n5850), .A2(n6014), .ZN(n5852) );
  NAND2_X1 U7588 ( .A1(n5852), .A2(n8304), .ZN(n5851) );
  NAND3_X1 U7589 ( .A1(n7433), .A2(n5969), .A3(n5851), .ZN(n5854) );
  AOI21_X1 U7590 ( .B1(n5852), .B2(n5848), .A(n6152), .ZN(n5853) );
  OAI211_X1 U7591 ( .C1(n5864), .C2(n5857), .A(n5856), .B(n7634), .ZN(n5860)
         );
  NAND2_X1 U7592 ( .A1(n5874), .A2(n6012), .ZN(n5869) );
  NAND2_X1 U7593 ( .A1(n5871), .A2(n6013), .ZN(n5868) );
  MUX2_X1 U7594 ( .A(n5869), .B(n5868), .S(n7082), .Z(n5876) );
  INV_X1 U7595 ( .A(n5876), .ZN(n5870) );
  AND2_X1 U7596 ( .A1(n6012), .A2(n5873), .ZN(n5875) );
  OR2_X1 U7597 ( .A1(n5877), .A2(n7082), .ZN(n5878) );
  OAI21_X1 U7598 ( .B1(n5879), .B2(n6152), .A(n5878), .ZN(n5880) );
  NOR3_X1 U7599 ( .A1(n8298), .A2(n5490), .A3(n5880), .ZN(n5881) );
  NAND2_X1 U7600 ( .A1(n5882), .A2(n5881), .ZN(n5892) );
  NAND3_X1 U7601 ( .A1(n5885), .A2(n7082), .A3(n8784), .ZN(n5883) );
  OAI21_X1 U7602 ( .B1(n5886), .B2(n6152), .A(n5883), .ZN(n5884) );
  NAND2_X1 U7603 ( .A1(n5884), .A2(n5889), .ZN(n5888) );
  INV_X1 U7604 ( .A(n5885), .ZN(n8878) );
  NAND4_X1 U7605 ( .A1(n5886), .A2(n8878), .A3(n6152), .A4(n8916), .ZN(n5887)
         );
  OAI211_X1 U7606 ( .C1(n7082), .C2(n5889), .A(n5888), .B(n5887), .ZN(n5890)
         );
  INV_X1 U7607 ( .A(n5890), .ZN(n5891) );
  NAND2_X1 U7608 ( .A1(n5892), .A2(n5891), .ZN(n5895) );
  MUX2_X1 U7609 ( .A(n8789), .B(n8368), .S(n7082), .Z(n5894) );
  MUX2_X1 U7610 ( .A(n4368), .B(n5897), .S(n7082), .Z(n5898) );
  OAI21_X1 U7611 ( .B1(n6009), .B2(n5901), .A(n7082), .ZN(n5902) );
  AND2_X1 U7612 ( .A1(n9231), .A2(n7082), .ZN(n5903) );
  AND2_X1 U7613 ( .A1(n9232), .A2(n5903), .ZN(n5904) );
  NAND2_X1 U7614 ( .A1(n5916), .A2(n6009), .ZN(n5915) );
  NAND3_X1 U7615 ( .A1(n5907), .A2(n5906), .A3(n5905), .ZN(n5909) );
  NAND3_X1 U7616 ( .A1(n5909), .A2(n6152), .A3(n5908), .ZN(n5910) );
  NAND2_X1 U7617 ( .A1(n5911), .A2(n5910), .ZN(n5913) );
  NAND3_X1 U7618 ( .A1(n5913), .A2(n5912), .A3(n9231), .ZN(n5914) );
  NAND2_X1 U7619 ( .A1(n9234), .A2(n5918), .ZN(n5919) );
  AOI21_X1 U7620 ( .B1(n5922), .B2(n9233), .A(n6152), .ZN(n5921) );
  OAI21_X1 U7621 ( .B1(n5923), .B2(n6152), .A(n9215), .ZN(n5924) );
  INV_X1 U7622 ( .A(n6005), .ZN(n5929) );
  NAND2_X1 U7623 ( .A1(n5932), .A2(n6152), .ZN(n5933) );
  NAND4_X1 U7624 ( .A1(n5938), .A2(n6004), .A3(n7082), .A4(n5937), .ZN(n5939)
         );
  INV_X1 U7625 ( .A(n8913), .ZN(n6201) );
  INV_X1 U7626 ( .A(n9419), .ZN(n6149) );
  MUX2_X1 U7627 ( .A(n6201), .B(n6149), .S(n6152), .Z(n5965) );
  OR2_X1 U7628 ( .A1(n6752), .A2(n5965), .ZN(n5940) );
  INV_X1 U7629 ( .A(SI_29_), .ZN(n5941) );
  NAND2_X1 U7630 ( .A1(n5944), .A2(n5943), .ZN(n5948) );
  AND2_X1 U7631 ( .A1(n5946), .A2(n5945), .ZN(n5947) );
  NAND2_X1 U7632 ( .A1(n5948), .A2(n5947), .ZN(n5991) );
  MUX2_X1 U7633 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4281), .Z(n5949) );
  NAND2_X1 U7634 ( .A1(n5949), .A2(SI_30_), .ZN(n5980) );
  INV_X1 U7635 ( .A(n5949), .ZN(n5951) );
  INV_X1 U7636 ( .A(SI_30_), .ZN(n5950) );
  NAND2_X1 U7637 ( .A1(n5951), .A2(n5950), .ZN(n5983) );
  NAND2_X1 U7638 ( .A1(n5980), .A2(n5983), .ZN(n5952) );
  NAND2_X1 U7639 ( .A1(n8415), .A2(n5365), .ZN(n5954) );
  NAND2_X1 U7640 ( .A1(n5993), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5953) );
  INV_X1 U7641 ( .A(n9416), .ZN(n6036) );
  INV_X1 U7642 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7643 ( .A1(n4282), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7644 ( .A1(n5955), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5956) );
  OAI211_X1 U7645 ( .C1(n5959), .C2(n5958), .A(n5957), .B(n5956), .ZN(n5960)
         );
  INV_X1 U7646 ( .A(n5960), .ZN(n5961) );
  NAND2_X1 U7647 ( .A1(n6001), .A2(n5961), .ZN(n8911) );
  INV_X1 U7648 ( .A(n8911), .ZN(n6035) );
  NAND2_X1 U7649 ( .A1(n6036), .A2(n6035), .ZN(n6032) );
  NAND2_X1 U7650 ( .A1(n6032), .A2(n5962), .ZN(n6046) );
  INV_X1 U7651 ( .A(n6046), .ZN(n5963) );
  NAND2_X1 U7652 ( .A1(n5964), .A2(n5963), .ZN(n5968) );
  NOR2_X1 U7653 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  INV_X1 U7654 ( .A(n6048), .ZN(n5972) );
  NAND2_X1 U7655 ( .A1(n5969), .A2(n8104), .ZN(n6060) );
  INV_X1 U7656 ( .A(n6060), .ZN(n5970) );
  AND2_X1 U7657 ( .A1(n5970), .A2(n6054), .ZN(n6034) );
  INV_X1 U7658 ( .A(n6034), .ZN(n5971) );
  NOR3_X1 U7659 ( .A1(n6050), .A2(n5972), .A3(n5971), .ZN(n5973) );
  OAI211_X1 U7660 ( .C1(n4370), .C2(n9419), .A(n5974), .B(n5973), .ZN(n6043)
         );
  INV_X1 U7661 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5976) );
  INV_X1 U7662 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5975) );
  MUX2_X1 U7663 ( .A(n5976), .B(n5975), .S(n4281), .Z(n5977) );
  XNOR2_X1 U7664 ( .A(n5977), .B(SI_31_), .ZN(n5982) );
  NAND2_X1 U7665 ( .A1(n5982), .A2(n5983), .ZN(n5990) );
  INV_X1 U7666 ( .A(n5980), .ZN(n5978) );
  NAND3_X1 U7667 ( .A1(n5981), .A2(n5982), .A3(n5980), .ZN(n5987) );
  INV_X1 U7668 ( .A(n5982), .ZN(n5985) );
  INV_X1 U7669 ( .A(n5983), .ZN(n5984) );
  XNOR2_X1 U7670 ( .A(n5985), .B(n5984), .ZN(n5986) );
  NAND2_X1 U7671 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  OR2_X1 U7672 ( .A1(n8433), .A2(n5992), .ZN(n5995) );
  NAND2_X1 U7673 ( .A1(n5993), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5994) );
  INV_X1 U7674 ( .A(n9410), .ZN(n6002) );
  INV_X1 U7675 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9413) );
  INV_X1 U7676 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9150) );
  OR2_X1 U7677 ( .A1(n5335), .A2(n9150), .ZN(n5998) );
  INV_X1 U7678 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9347) );
  OR2_X1 U7679 ( .A1(n5996), .A2(n9347), .ZN(n5997) );
  OAI211_X1 U7680 ( .C1(n5958), .C2(n9413), .A(n5998), .B(n5997), .ZN(n5999)
         );
  INV_X1 U7681 ( .A(n5999), .ZN(n6000) );
  INV_X1 U7682 ( .A(n9147), .ZN(n8213) );
  NAND2_X1 U7683 ( .A1(n6002), .A2(n8213), .ZN(n6039) );
  INV_X1 U7684 ( .A(n9259), .ZN(n9264) );
  INV_X1 U7685 ( .A(n9231), .ZN(n6010) );
  NAND2_X1 U7686 ( .A1(n5847), .A2(n6014), .ZN(n7470) );
  NOR2_X1 U7687 ( .A1(n7443), .A2(n7470), .ZN(n6018) );
  NOR2_X1 U7688 ( .A1(n7554), .A2(n6015), .ZN(n6017) );
  NOR2_X1 U7689 ( .A1(n5293), .A2(n6153), .ZN(n6016) );
  NAND4_X1 U7690 ( .A1(n6018), .A2(n6017), .A3(n7433), .A4(n6016), .ZN(n6019)
         );
  XNOR2_X1 U7691 ( .A(n8037), .B(n7698), .ZN(n7638) );
  NOR2_X1 U7692 ( .A1(n6019), .A2(n7638), .ZN(n6020) );
  NAND4_X1 U7693 ( .A1(n7760), .A2(n7648), .A3(n7614), .A4(n6020), .ZN(n6021)
         );
  NOR4_X1 U7694 ( .A1(n8298), .A2(n5490), .A3(n8026), .A4(n6021), .ZN(n6022)
         );
  INV_X1 U7695 ( .A(n8322), .ZN(n8316) );
  NAND4_X1 U7696 ( .A1(n9318), .A2(n9329), .A3(n6022), .A4(n8316), .ZN(n6023)
         );
  NOR4_X1 U7697 ( .A1(n9282), .A2(n9291), .A3(n9307), .A4(n6023), .ZN(n6024)
         );
  NAND3_X1 U7698 ( .A1(n9242), .A2(n9264), .A3(n6024), .ZN(n6025) );
  NOR2_X1 U7699 ( .A1(n9237), .A2(n6025), .ZN(n6026) );
  NAND4_X1 U7700 ( .A1(n9198), .A2(n9201), .A3(n6026), .A4(n9215), .ZN(n6027)
         );
  NOR2_X1 U7701 ( .A1(n9187), .A2(n6027), .ZN(n6028) );
  NAND4_X1 U7702 ( .A1(n6039), .A2(n9170), .A3(n6028), .A4(n6206), .ZN(n6030)
         );
  NOR3_X1 U7703 ( .A1(n6030), .A2(n6029), .A3(n6752), .ZN(n6033) );
  INV_X1 U7704 ( .A(n6050), .ZN(n6031) );
  NAND3_X1 U7705 ( .A1(n6033), .A2(n6032), .A3(n6031), .ZN(n6038) );
  NAND3_X1 U7706 ( .A1(n6036), .A2(n6035), .A3(n6034), .ZN(n6037) );
  OAI211_X1 U7707 ( .C1(n6040), .C2(n6039), .A(n6038), .B(n6037), .ZN(n6041)
         );
  NAND2_X1 U7708 ( .A1(n9419), .A2(n6201), .ZN(n6044) );
  AOI21_X1 U7709 ( .B1(n9416), .B2(n9147), .A(n9410), .ZN(n6047) );
  INV_X1 U7710 ( .A(n7081), .ZN(n7079) );
  NAND2_X1 U7711 ( .A1(n7079), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8378) );
  INV_X1 U7712 ( .A(n6211), .ZN(n7624) );
  NAND2_X1 U7713 ( .A1(n6158), .A2(n7624), .ZN(n6178) );
  NOR3_X1 U7714 ( .A1(n6178), .A2(n7116), .A3(n7120), .ZN(n6056) );
  OAI21_X1 U7715 ( .B1(n8378), .B2(n6054), .A(P2_B_REG_SCAN_IN), .ZN(n6055) );
  OR2_X1 U7716 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  OAI21_X1 U7717 ( .B1(n6058), .B2(n8378), .A(n6057), .ZN(P2_U3296) );
  AND2_X1 U7718 ( .A1(n6060), .A2(n6059), .ZN(n6061) );
  OAI21_X2 U7719 ( .B1(n6062), .B2(n6153), .A(n6061), .ZN(n6070) );
  NAND2_X1 U7720 ( .A1(n6063), .A2(n5292), .ZN(n6066) );
  AND2_X1 U7721 ( .A1(n6066), .A2(n6064), .ZN(n7391) );
  NAND2_X1 U7722 ( .A1(n6065), .A2(n5847), .ZN(n7390) );
  NAND2_X1 U7723 ( .A1(n7389), .A2(n6066), .ZN(n7381) );
  XNOR2_X1 U7724 ( .A(n6070), .B(n7379), .ZN(n6068) );
  XNOR2_X1 U7725 ( .A(n6068), .B(n8924), .ZN(n7382) );
  NAND2_X1 U7726 ( .A1(n6068), .A2(n5314), .ZN(n6069) );
  NAND2_X1 U7727 ( .A1(n7380), .A2(n6069), .ZN(n7545) );
  INV_X2 U7728 ( .A(n6070), .ZN(n6147) );
  XNOR2_X1 U7729 ( .A(n6136), .B(n7748), .ZN(n6071) );
  XNOR2_X1 U7730 ( .A(n6071), .B(n5334), .ZN(n7546) );
  NAND2_X1 U7731 ( .A1(n6071), .A2(n5334), .ZN(n6072) );
  XNOR2_X1 U7732 ( .A(n6136), .B(n7583), .ZN(n6073) );
  INV_X1 U7733 ( .A(n8923), .ZN(n7683) );
  NAND2_X1 U7734 ( .A1(n6073), .A2(n7683), .ZN(n7685) );
  INV_X1 U7735 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7736 ( .A1(n6074), .A2(n8923), .ZN(n6075) );
  NAND2_X1 U7737 ( .A1(n7685), .A2(n6075), .ZN(n7581) );
  XNOR2_X1 U7738 ( .A(n6148), .B(n4512), .ZN(n6078) );
  XNOR2_X1 U7739 ( .A(n6078), .B(n8922), .ZN(n7684) );
  NAND2_X1 U7740 ( .A1(n6078), .A2(n4514), .ZN(n6079) );
  XNOR2_X1 U7741 ( .A(n6080), .B(n8037), .ZN(n7696) );
  XNOR2_X1 U7742 ( .A(n6148), .B(n8033), .ZN(n6082) );
  NAND2_X1 U7743 ( .A1(n6082), .A2(n6081), .ZN(n8157) );
  INV_X1 U7744 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7745 ( .A1(n6083), .A2(n8920), .ZN(n6084) );
  NAND2_X1 U7746 ( .A1(n8157), .A2(n6084), .ZN(n8031) );
  XNOR2_X1 U7747 ( .A(n6148), .B(n7617), .ZN(n6087) );
  XNOR2_X1 U7748 ( .A(n6087), .B(n6088), .ZN(n8158) );
  INV_X1 U7749 ( .A(n6087), .ZN(n6089) );
  NAND2_X1 U7750 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  XNOR2_X1 U7751 ( .A(n8269), .B(n6148), .ZN(n6091) );
  XNOR2_X1 U7752 ( .A(n6091), .B(n8918), .ZN(n8264) );
  XNOR2_X1 U7753 ( .A(n8215), .B(n6136), .ZN(n8752) );
  XNOR2_X1 U7754 ( .A(n8200), .B(n6148), .ZN(n8868) );
  XNOR2_X1 U7755 ( .A(n8790), .B(n6148), .ZN(n6098) );
  XNOR2_X1 U7756 ( .A(n6098), .B(n8873), .ZN(n8785) );
  OR2_X1 U7757 ( .A1(n6136), .A2(n8917), .ZN(n6092) );
  OAI22_X1 U7758 ( .A1(n8215), .A2(n6092), .B1(n6147), .B2(n8916), .ZN(n6095)
         );
  NAND3_X1 U7759 ( .A1(n8215), .A2(n8751), .A3(n6148), .ZN(n6093) );
  OAI211_X1 U7760 ( .C1(n8916), .C2(n6148), .A(n8200), .B(n6093), .ZN(n6094)
         );
  OAI21_X1 U7761 ( .B1(n8200), .B2(n6095), .A(n6094), .ZN(n6096) );
  NAND2_X1 U7762 ( .A1(n6098), .A2(n8915), .ZN(n6099) );
  NAND2_X1 U7763 ( .A1(n6100), .A2(n6099), .ZN(n8848) );
  INV_X1 U7764 ( .A(n8848), .ZN(n6105) );
  XNOR2_X1 U7765 ( .A(n8368), .B(n6147), .ZN(n6101) );
  INV_X1 U7766 ( .A(n6101), .ZN(n6102) );
  NAND2_X1 U7767 ( .A1(n6102), .A2(n9332), .ZN(n6103) );
  NAND2_X1 U7768 ( .A1(n8734), .A2(n6103), .ZN(n8847) );
  INV_X1 U7769 ( .A(n8847), .ZN(n6104) );
  XNOR2_X1 U7770 ( .A(n9484), .B(n6148), .ZN(n6106) );
  XNOR2_X1 U7771 ( .A(n6106), .B(n9320), .ZN(n8735) );
  NAND2_X1 U7772 ( .A1(n6106), .A2(n9316), .ZN(n6107) );
  XNOR2_X1 U7773 ( .A(n9477), .B(n6136), .ZN(n6112) );
  XNOR2_X1 U7774 ( .A(n6112), .B(n6108), .ZN(n8899) );
  XNOR2_X1 U7775 ( .A(n9471), .B(n6136), .ZN(n6109) );
  NAND2_X1 U7776 ( .A1(n6109), .A2(n9295), .ZN(n8817) );
  INV_X1 U7777 ( .A(n6109), .ZN(n6110) );
  INV_X1 U7778 ( .A(n9295), .ZN(n9321) );
  NAND2_X1 U7779 ( .A1(n6110), .A2(n9321), .ZN(n6111) );
  NAND2_X1 U7780 ( .A1(n8817), .A2(n6111), .ZN(n8807) );
  INV_X1 U7781 ( .A(n6112), .ZN(n6113) );
  AND2_X1 U7782 ( .A1(n6113), .A2(n9334), .ZN(n8806) );
  NOR2_X1 U7783 ( .A1(n8807), .A2(n8806), .ZN(n6114) );
  XNOR2_X1 U7784 ( .A(n9393), .B(n6148), .ZN(n6115) );
  NAND2_X1 U7785 ( .A1(n6115), .A2(n8812), .ZN(n8879) );
  INV_X1 U7786 ( .A(n6115), .ZN(n6116) );
  NAND2_X1 U7787 ( .A1(n6116), .A2(n9308), .ZN(n6117) );
  AND2_X1 U7788 ( .A1(n8879), .A2(n6117), .ZN(n8818) );
  XNOR2_X1 U7789 ( .A(n9281), .B(n6148), .ZN(n6119) );
  NAND2_X1 U7790 ( .A1(n6119), .A2(n9297), .ZN(n8762) );
  INV_X1 U7791 ( .A(n6119), .ZN(n6120) );
  NAND2_X1 U7792 ( .A1(n6120), .A2(n9260), .ZN(n6121) );
  AND2_X1 U7793 ( .A1(n8762), .A2(n6121), .ZN(n8880) );
  XNOR2_X1 U7794 ( .A(n9270), .B(n6136), .ZN(n6122) );
  NAND2_X1 U7795 ( .A1(n6122), .A2(n9247), .ZN(n8836) );
  INV_X1 U7796 ( .A(n6122), .ZN(n6123) );
  NAND2_X1 U7797 ( .A1(n6123), .A2(n9275), .ZN(n6124) );
  AND2_X1 U7798 ( .A1(n8836), .A2(n6124), .ZN(n8763) );
  XNOR2_X1 U7799 ( .A(n8835), .B(n6148), .ZN(n6125) );
  NAND2_X1 U7800 ( .A1(n6125), .A2(n9227), .ZN(n8772) );
  INV_X1 U7801 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7802 ( .A1(n6126), .A2(n9261), .ZN(n6127) );
  AND2_X1 U7803 ( .A1(n8772), .A2(n6127), .ZN(n8837) );
  NAND2_X1 U7804 ( .A1(n8771), .A2(n8772), .ZN(n6129) );
  XNOR2_X1 U7805 ( .A(n9454), .B(n6147), .ZN(n6130) );
  XNOR2_X1 U7806 ( .A(n6130), .B(n9248), .ZN(n8773) );
  INV_X1 U7807 ( .A(n6130), .ZN(n6131) );
  NAND2_X1 U7808 ( .A1(n6131), .A2(n9248), .ZN(n6132) );
  XNOR2_X1 U7809 ( .A(n9370), .B(n6148), .ZN(n8857) );
  INV_X1 U7810 ( .A(n8857), .ZN(n6133) );
  NAND2_X1 U7811 ( .A1(n6133), .A2(n9206), .ZN(n6135) );
  AND2_X1 U7812 ( .A1(n8857), .A2(n9226), .ZN(n6134) );
  AOI21_X2 U7813 ( .B1(n8859), .B2(n6135), .A(n6134), .ZN(n8828) );
  XNOR2_X1 U7814 ( .A(n9437), .B(n6148), .ZN(n8830) );
  INV_X1 U7815 ( .A(n8827), .ZN(n6138) );
  OAI22_X1 U7816 ( .A1(n8830), .A2(n8746), .B1(n9214), .B2(n6138), .ZN(n6142)
         );
  OAI21_X1 U7817 ( .B1(n8827), .B2(n9193), .A(n9205), .ZN(n6140) );
  NOR3_X1 U7818 ( .A1(n8827), .A2(n9193), .A3(n9205), .ZN(n6139) );
  AOI21_X1 U7819 ( .B1(n8830), .B2(n6140), .A(n6139), .ZN(n6141) );
  OAI21_X2 U7820 ( .B1(n8828), .B2(n6142), .A(n6141), .ZN(n8796) );
  XNOR2_X1 U7821 ( .A(n9431), .B(n6148), .ZN(n6143) );
  XOR2_X1 U7822 ( .A(n8890), .B(n6143), .Z(n8797) );
  XNOR2_X1 U7823 ( .A(n6145), .B(n6148), .ZN(n6146) );
  XNOR2_X1 U7824 ( .A(n6146), .B(n9181), .ZN(n8889) );
  XNOR2_X1 U7825 ( .A(n6218), .B(n6147), .ZN(n6168) );
  NAND2_X1 U7826 ( .A1(n6168), .A2(n9172), .ZN(n6150) );
  OAI21_X1 U7827 ( .B1(n6168), .B2(n9172), .A(n6150), .ZN(n7066) );
  XNOR2_X1 U7828 ( .A(n8913), .B(n6148), .ZN(n6191) );
  XNOR2_X1 U7829 ( .A(n6149), .B(n6191), .ZN(n6167) );
  INV_X1 U7830 ( .A(n6167), .ZN(n6164) );
  INV_X1 U7831 ( .A(n6150), .ZN(n6162) );
  AND2_X1 U7832 ( .A1(n6151), .A2(n6157), .ZN(n6176) );
  AND2_X1 U7833 ( .A1(n6152), .A2(n10434), .ZN(n6155) );
  NAND2_X1 U7834 ( .A1(n6155), .A2(n6210), .ZN(n6172) );
  INV_X1 U7835 ( .A(n6172), .ZN(n6156) );
  NAND2_X1 U7836 ( .A1(n6213), .A2(n6156), .ZN(n6161) );
  INV_X1 U7837 ( .A(n6210), .ZN(n6159) );
  NAND2_X1 U7838 ( .A1(n6215), .A2(n6159), .ZN(n6160) );
  NAND2_X1 U7839 ( .A1(n6166), .A2(n6165), .ZN(n6199) );
  NAND3_X1 U7840 ( .A1(n7075), .A2(n6167), .A3(n8882), .ZN(n6198) );
  INV_X1 U7841 ( .A(n6168), .ZN(n6192) );
  INV_X1 U7842 ( .A(n6191), .ZN(n6169) );
  NAND2_X1 U7843 ( .A1(n9172), .A2(n8882), .ZN(n6190) );
  NOR4_X1 U7844 ( .A1(n6192), .A2(n9419), .A3(n6169), .A4(n6190), .ZN(n6189)
         );
  NOR2_X1 U7845 ( .A1(n6211), .A2(n6170), .ZN(n6171) );
  NAND2_X1 U7846 ( .A1(n6172), .A2(n9337), .ZN(n6214) );
  INV_X1 U7847 ( .A(n6214), .ZN(n6175) );
  OR2_X1 U7848 ( .A1(n6179), .A2(n6210), .ZN(n6173) );
  OAI211_X1 U7849 ( .C1(n6176), .C2(n6175), .A(n6174), .B(n6173), .ZN(n6177)
         );
  NAND2_X1 U7850 ( .A1(n6177), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6181) );
  OR2_X1 U7851 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  AOI22_X1 U7852 ( .A1(n6182), .A2(n8906), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n6186) );
  NOR2_X1 U7853 ( .A1(n6211), .A2(n6183), .ZN(n6184) );
  NAND2_X1 U7854 ( .A1(n9172), .A2(n8902), .ZN(n6185) );
  OAI211_X1 U7855 ( .C1(n6187), .C2(n8904), .A(n6186), .B(n6185), .ZN(n6188)
         );
  NOR3_X1 U7856 ( .A1(n6192), .A2(n6191), .A3(n6190), .ZN(n6194) );
  NAND2_X1 U7857 ( .A1(n6213), .A2(n9394), .ZN(n6193) );
  OAI21_X1 U7858 ( .B1(n6194), .B2(n8896), .A(n9419), .ZN(n6195) );
  NAND3_X1 U7859 ( .A1(n6199), .A2(n6198), .A3(n6197), .ZN(P2_U3160) );
  XNOR2_X1 U7860 ( .A(n6200), .B(n6206), .ZN(n6205) );
  NOR2_X1 U7861 ( .A1(n6207), .A2(n6206), .ZN(n9162) );
  NOR2_X1 U7862 ( .A1(n9162), .A2(n10436), .ZN(n6208) );
  NOR2_X1 U7863 ( .A1(n9167), .A2(n6209), .ZN(n9353) );
  NAND2_X1 U7864 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U7865 ( .A1(n6213), .A2(n6212), .ZN(n6217) );
  NAND2_X1 U7866 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  OR2_X1 U7867 ( .A1(n9353), .A2(n10441), .ZN(n6222) );
  INV_X1 U7868 ( .A(n6220), .ZN(n6221) );
  NAND2_X1 U7869 ( .A1(n6222), .A2(n6221), .ZN(P2_U3454) );
  NOR2_X1 U7870 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6226) );
  NOR2_X1 U7871 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6225) );
  NOR2_X1 U7872 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6224) );
  NOR2_X1 U7873 ( .A1(n6702), .A2(n5106), .ZN(n6234) );
  NOR2_X1 U7874 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6230) );
  NAND2_X1 U7875 ( .A1(n7174), .A2(n6592), .ZN(n6245) );
  NOR2_X1 U7876 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6326) );
  NOR2_X1 U7877 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6239) );
  NAND3_X1 U7878 ( .A1(n6240), .A2(n6326), .A3(n6239), .ZN(n6287) );
  INV_X1 U7879 ( .A(n6430), .ZN(n6242) );
  NAND2_X1 U7880 ( .A1(n6242), .A2(n6241), .ZN(n6367) );
  NAND2_X1 U7881 ( .A1(n6367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6261) );
  INV_X1 U7882 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7883 ( .A1(n6261), .A2(n6260), .ZN(n6263) );
  NAND2_X1 U7884 ( .A1(n6263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6243) );
  XNOR2_X1 U7885 ( .A(n6243), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7345) );
  AOI22_X1 U7886 ( .A1(n6593), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7155), .B2(
        n7345), .ZN(n6244) );
  NAND2_X2 U7887 ( .A1(n6245), .A2(n6244), .ZN(n10113) );
  NAND2_X1 U7888 ( .A1(n6248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7889 ( .A1(n6270), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6259) );
  INV_X1 U7890 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10111) );
  OR2_X1 U7891 ( .A1(n7169), .A2(n10111), .ZN(n6258) );
  INV_X1 U7892 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6250) );
  OR2_X1 U7893 ( .A1(n6647), .A2(n6250), .ZN(n6257) );
  INV_X1 U7894 ( .A(n6253), .ZN(n6269) );
  INV_X1 U7895 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7896 ( .A1(n6269), .A2(n6254), .ZN(n6255) );
  NAND2_X1 U7897 ( .A1(n6377), .A2(n6255), .ZN(n10110) );
  OR2_X1 U7898 ( .A1(n6529), .A2(n10110), .ZN(n6256) );
  OR2_X1 U7899 ( .A1(n10113), .A2(n8232), .ZN(n8501) );
  OR2_X1 U7900 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  AOI22_X1 U7901 ( .A1(n6593), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7155), .B2(
        n9812), .ZN(n6264) );
  INV_X1 U7902 ( .A(n6266), .ZN(n6281) );
  INV_X1 U7903 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7904 ( .A1(n6281), .A2(n6267), .ZN(n6268) );
  NAND2_X1 U7905 ( .A1(n6269), .A2(n6268), .ZN(n8231) );
  OR2_X1 U7906 ( .A1(n6529), .A2(n8231), .ZN(n6275) );
  NAND2_X1 U7907 ( .A1(n6618), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6274) );
  INV_X1 U7908 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6271) );
  OR2_X1 U7909 ( .A1(n6621), .A2(n6271), .ZN(n6273) );
  INV_X1 U7910 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7274) );
  OR2_X1 U7911 ( .A1(n7169), .A2(n7274), .ZN(n6272) );
  NAND4_X1 U7912 ( .A1(n6275), .A2(n6274), .A3(n6273), .A4(n6272), .ZN(n9737)
         );
  NAND2_X1 U7913 ( .A1(n8188), .A2(n9737), .ZN(n8149) );
  NAND2_X1 U7914 ( .A1(n8501), .A2(n8149), .ZN(n8493) );
  NAND2_X1 U7915 ( .A1(n10209), .A2(n7676), .ZN(n8491) );
  NAND2_X1 U7916 ( .A1(n6430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6276) );
  XNOR2_X1 U7917 ( .A(n6276), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U7918 ( .A1(n6593), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7155), .B2(
        n9799), .ZN(n6277) );
  NAND2_X1 U7919 ( .A1(n7168), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6285) );
  INV_X1 U7920 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7272) );
  OR2_X1 U7921 ( .A1(n7169), .A2(n7272), .ZN(n6284) );
  INV_X1 U7922 ( .A(n6278), .ZN(n6294) );
  INV_X1 U7923 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7924 ( .A1(n6294), .A2(n6279), .ZN(n6280) );
  NAND2_X1 U7925 ( .A1(n6281), .A2(n6280), .ZN(n7674) );
  OR2_X1 U7926 ( .A1(n6617), .A2(n7674), .ZN(n6283) );
  INV_X1 U7927 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7256) );
  OR2_X1 U7928 ( .A1(n6647), .A2(n7256), .ZN(n6282) );
  NAND2_X1 U7929 ( .A1(n8074), .A2(n8175), .ZN(n8176) );
  AND2_X1 U7930 ( .A1(n8491), .A2(n8176), .ZN(n8488) );
  OR2_X1 U7931 ( .A1(n8493), .A2(n8488), .ZN(n6286) );
  NAND2_X1 U7932 ( .A1(n10113), .A2(n8232), .ZN(n8497) );
  AND2_X1 U7933 ( .A1(n6286), .A2(n8497), .ZN(n6366) );
  NAND2_X1 U7934 ( .A1(n7148), .A2(n6592), .ZN(n6291) );
  NAND2_X1 U7935 ( .A1(n6287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6288) );
  MUX2_X1 U7936 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6288), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6289) );
  AOI22_X1 U7937 ( .A1(n6593), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7155), .B2(
        n9786), .ZN(n6290) );
  NAND2_X1 U7938 ( .A1(n7168), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6299) );
  INV_X1 U7939 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8005) );
  OR2_X1 U7940 ( .A1(n7169), .A2(n8005), .ZN(n6298) );
  NAND2_X1 U7941 ( .A1(n6358), .A2(n6292), .ZN(n6293) );
  NAND2_X1 U7942 ( .A1(n6294), .A2(n6293), .ZN(n8008) );
  OR2_X1 U7943 ( .A1(n6529), .A2(n8008), .ZN(n6297) );
  INV_X1 U7944 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6295) );
  OR2_X1 U7945 ( .A1(n6647), .A2(n6295), .ZN(n6296) );
  NAND2_X1 U7946 ( .A1(n4902), .A2(n6364), .ZN(n8486) );
  NAND2_X1 U7947 ( .A1(n6366), .A2(n8486), .ZN(n8594) );
  NAND2_X1 U7948 ( .A1(n6418), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6301) );
  INV_X1 U7949 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7188) );
  INV_X1 U7950 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7951 ( .A1(n6618), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6303) );
  NOR2_X1 U7952 ( .A1(n4281), .A2(n6304), .ZN(n6305) );
  XNOR2_X1 U7953 ( .A(n6305), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10264) );
  MUX2_X1 U7954 ( .A(n4433), .B(n10264), .S(n6306), .Z(n10381) );
  INV_X1 U7955 ( .A(n6647), .ZN(n6307) );
  INV_X1 U7956 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7799) );
  OR2_X1 U7957 ( .A1(n7169), .A2(n7799), .ZN(n6308) );
  INV_X1 U7958 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7798) );
  OR2_X1 U7959 ( .A1(n6617), .A2(n7798), .ZN(n6311) );
  NAND2_X1 U7960 ( .A1(n6270), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7961 ( .A1(n10249), .A2(n9752), .ZN(n6318) );
  NAND2_X1 U7962 ( .A1(n4281), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7963 ( .A1(n6313), .A2(n6312), .ZN(n6314) );
  NAND2_X1 U7964 ( .A1(n6314), .A2(n7278), .ZN(n6317) );
  INV_X1 U7965 ( .A(n10249), .ZN(n7360) );
  NAND2_X1 U7966 ( .A1(n4281), .A2(n4583), .ZN(n6315) );
  OAI211_X1 U7967 ( .C1(n7134), .C2(n4281), .A(n7360), .B(n6315), .ZN(n6316)
         );
  OAI211_X2 U7968 ( .C1(n7278), .C2(n6318), .A(n6317), .B(n6316), .ZN(n9567)
         );
  INV_X1 U7969 ( .A(n6319), .ZN(n7489) );
  NAND2_X1 U7970 ( .A1(n7489), .A2(n9567), .ZN(n6320) );
  INV_X1 U7971 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8014) );
  OR2_X1 U7972 ( .A1(n6617), .A2(n8014), .ZN(n6325) );
  NAND2_X1 U7973 ( .A1(n6618), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6324) );
  INV_X1 U7974 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8015) );
  OR2_X1 U7975 ( .A1(n7169), .A2(n8015), .ZN(n6323) );
  INV_X1 U7976 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6321) );
  OR2_X1 U7977 ( .A1(n6621), .A2(n6321), .ZN(n6322) );
  NAND2_X1 U7978 ( .A1(n7132), .A2(n6592), .ZN(n6329) );
  OR2_X1 U7979 ( .A1(n6326), .A2(n6634), .ZN(n6349) );
  XNOR2_X1 U7980 ( .A(n6349), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U7981 ( .A1(n7155), .A2(n7266), .ZN(n6328) );
  NAND2_X1 U7982 ( .A1(n6593), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7983 ( .A1(n9743), .A2(n8016), .ZN(n8668) );
  NAND2_X1 U7984 ( .A1(n8468), .A2(n8668), .ZN(n6330) );
  OR2_X1 U7985 ( .A1(n6529), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7986 ( .A1(n6618), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6334) );
  INV_X1 U7987 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10363) );
  OR2_X1 U7988 ( .A1(n7169), .A2(n10363), .ZN(n6333) );
  INV_X1 U7989 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6331) );
  OR2_X1 U7990 ( .A1(n6621), .A2(n6331), .ZN(n6332) );
  NAND4_X2 U7991 ( .A1(n6335), .A2(n6334), .A3(n6333), .A4(n6332), .ZN(n9742)
         );
  INV_X1 U7992 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7993 ( .A1(n6349), .A2(n6336), .ZN(n6337) );
  NAND2_X1 U7994 ( .A1(n6337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6338) );
  XNOR2_X1 U7995 ( .A(n6338), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U7996 ( .A1(n6593), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6339) );
  NOR2_X1 U7997 ( .A1(n9742), .A2(n7605), .ZN(n8469) );
  NAND2_X1 U7998 ( .A1(n6270), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6347) );
  INV_X1 U7999 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7843) );
  OR2_X1 U8000 ( .A1(n7169), .A2(n7843), .ZN(n6346) );
  INV_X1 U8001 ( .A(n6342), .ZN(n6356) );
  OAI21_X1 U8002 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6356), .ZN(n7844) );
  OR2_X1 U8003 ( .A1(n6617), .A2(n7844), .ZN(n6345) );
  INV_X1 U8004 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6343) );
  OR2_X1 U8005 ( .A1(n6647), .A2(n6343), .ZN(n6344) );
  OAI21_X1 U8006 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8007 ( .A1(n6349), .A2(n6348), .ZN(n6352) );
  INV_X1 U8008 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6350) );
  XNOR2_X1 U8009 ( .A(n6352), .B(n6350), .ZN(n10273) );
  NAND2_X1 U8010 ( .A1(n7140), .A2(n6592), .ZN(n6355) );
  OAI21_X1 U8011 ( .B1(n6352), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6353) );
  XNOR2_X1 U8012 ( .A(n6353), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9773) );
  AOI22_X1 U8013 ( .A1(n6593), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7155), .B2(
        n9773), .ZN(n6354) );
  INV_X1 U8014 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U8015 ( .A1(n6356), .A2(n7863), .ZN(n6357) );
  NAND2_X1 U8016 ( .A1(n6358), .A2(n6357), .ZN(n10351) );
  OR2_X1 U8017 ( .A1(n6529), .A2(n10351), .ZN(n6362) );
  NAND2_X1 U8018 ( .A1(n6618), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6361) );
  INV_X1 U8019 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7938) );
  OR2_X1 U8020 ( .A1(n6621), .A2(n7938), .ZN(n6360) );
  INV_X1 U8021 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10352) );
  OR2_X1 U8022 ( .A1(n7169), .A2(n10352), .ZN(n6359) );
  NAND4_X1 U8023 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n9740)
         );
  NAND2_X1 U8024 ( .A1(n7775), .A2(n9740), .ZN(n8674) );
  NAND2_X1 U8025 ( .A1(n7710), .A2(n8674), .ZN(n6363) );
  INV_X1 U8026 ( .A(n9740), .ZN(n7739) );
  NAND2_X1 U8027 ( .A1(n7739), .A2(n10354), .ZN(n8481) );
  NAND2_X1 U8028 ( .A1(n6363), .A2(n8481), .ZN(n8002) );
  NAND2_X1 U8029 ( .A1(n8149), .A2(n6663), .ZN(n8490) );
  NOR2_X1 U8030 ( .A1(n8490), .A2(n8478), .ZN(n6365) );
  NAND2_X1 U8031 ( .A1(n6365), .A2(n8501), .ZN(n8609) );
  NAND2_X1 U8032 ( .A1(n6366), .A2(n8609), .ZN(n8677) );
  INV_X2 U8033 ( .A(n8420), .ZN(n6514) );
  NAND2_X1 U8034 ( .A1(n7180), .A2(n6514), .ZN(n6374) );
  INV_X1 U8035 ( .A(n6367), .ZN(n6369) );
  NOR2_X1 U8036 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6368) );
  NAND2_X1 U8037 ( .A1(n6369), .A2(n6368), .ZN(n6371) );
  NAND2_X1 U8038 ( .A1(n6371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6370) );
  MUX2_X1 U8039 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6370), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6372) );
  AOI22_X1 U8040 ( .A1(n6593), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7155), .B2(
        n7418), .ZN(n6373) );
  NAND2_X1 U8041 ( .A1(n6643), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6383) );
  INV_X1 U8042 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6375) );
  OR2_X1 U8043 ( .A1(n6621), .A2(n6375), .ZN(n6382) );
  NAND2_X1 U8044 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  NAND2_X1 U8045 ( .A1(n6393), .A2(n6378), .ZN(n10099) );
  OR2_X1 U8046 ( .A1(n6529), .A2(n10099), .ZN(n6381) );
  INV_X1 U8047 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6379) );
  OR2_X1 U8048 ( .A1(n6647), .A2(n6379), .ZN(n6380) );
  OR2_X1 U8049 ( .A1(n10102), .A2(n9640), .ZN(n8506) );
  NAND2_X1 U8050 ( .A1(n10102), .A2(n9640), .ZN(n8503) );
  NAND2_X1 U8051 ( .A1(n7197), .A2(n6514), .ZN(n6390) );
  NAND2_X1 U8052 ( .A1(n6385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6384) );
  MUX2_X1 U8053 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6384), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n6388) );
  INV_X1 U8054 ( .A(n6385), .ZN(n6387) );
  INV_X1 U8055 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8056 ( .A1(n6387), .A2(n6386), .ZN(n6400) );
  NAND2_X1 U8057 ( .A1(n6388), .A2(n6400), .ZN(n7421) );
  INV_X1 U8058 ( .A(n7421), .ZN(n9831) );
  AOI22_X1 U8059 ( .A1(n6593), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7155), .B2(
        n9831), .ZN(n6389) );
  NAND2_X1 U8060 ( .A1(n6643), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6399) );
  INV_X1 U8061 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6391) );
  OR2_X1 U8062 ( .A1(n6647), .A2(n6391), .ZN(n6398) );
  INV_X1 U8063 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U8064 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  NAND2_X1 U8065 ( .A1(n6405), .A2(n6394), .ZN(n8096) );
  OR2_X1 U8066 ( .A1(n6529), .A2(n8096), .ZN(n6397) );
  INV_X1 U8067 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6395) );
  OR2_X1 U8068 ( .A1(n6621), .A2(n6395), .ZN(n6396) );
  OR2_X1 U8069 ( .A1(n9690), .A2(n9546), .ZN(n8505) );
  NAND2_X1 U8070 ( .A1(n9690), .A2(n9546), .ZN(n8508) );
  NAND2_X1 U8071 ( .A1(n7219), .A2(n6514), .ZN(n6402) );
  NAND2_X1 U8072 ( .A1(n6400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6414) );
  XNOR2_X1 U8073 ( .A(n6414), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7567) );
  AOI22_X1 U8074 ( .A1(n6593), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7567), .B2(
        n7155), .ZN(n6401) );
  INV_X1 U8075 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6403) );
  OR2_X1 U8076 ( .A1(n6647), .A2(n6403), .ZN(n6411) );
  NAND2_X1 U8077 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U8078 ( .A1(n6420), .A2(n6406), .ZN(n8083) );
  OR2_X1 U8079 ( .A1(n6529), .A2(n8083), .ZN(n6410) );
  NAND2_X1 U8080 ( .A1(n7168), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6409) );
  INV_X1 U8081 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6407) );
  OR2_X1 U8082 ( .A1(n7169), .A2(n6407), .ZN(n6408) );
  NAND4_X1 U8083 ( .A1(n6411), .A2(n6410), .A3(n6409), .A4(n6408), .ZN(n9733)
         );
  NAND2_X1 U8084 ( .A1(n8512), .A2(n9733), .ZN(n8498) );
  NAND2_X1 U8085 ( .A1(n10204), .A2(n9682), .ZN(n8684) );
  NAND2_X1 U8086 ( .A1(n8498), .A2(n8684), .ZN(n8611) );
  INV_X1 U8087 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8088 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  NAND2_X1 U8089 ( .A1(n6415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6416) );
  AOI22_X1 U8090 ( .A1(n9848), .A2(n7155), .B1(n6593), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8091 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  AND2_X1 U8092 ( .A1(n6437), .A2(n6421), .ZN(n9660) );
  NAND2_X1 U8093 ( .A1(n6418), .A2(n9660), .ZN(n6426) );
  NAND2_X1 U8094 ( .A1(n6618), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6425) );
  INV_X1 U8095 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8383) );
  OR2_X1 U8096 ( .A1(n6621), .A2(n8383), .ZN(n6424) );
  INV_X1 U8097 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6422) );
  OR2_X1 U8098 ( .A1(n7169), .A2(n6422), .ZN(n6423) );
  NAND4_X1 U8099 ( .A1(n6426), .A2(n6425), .A3(n6424), .A4(n6423), .ZN(n9732)
         );
  NAND2_X1 U8100 ( .A1(n9666), .A2(n9732), .ZN(n8523) );
  NAND2_X1 U8101 ( .A1(n8283), .A2(n9583), .ZN(n8685) );
  NAND2_X1 U8102 ( .A1(n8523), .A2(n8685), .ZN(n8278) );
  INV_X1 U8103 ( .A(n8498), .ZN(n6427) );
  NOR2_X1 U8104 ( .A1(n8278), .A2(n6427), .ZN(n6428) );
  OR2_X1 U8105 ( .A1(n7400), .A2(n8420), .ZN(n6435) );
  OAI21_X1 U8106 ( .B1(n6430), .B2(n6429), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6431) );
  MUX2_X1 U8107 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6431), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6433) );
  NAND2_X1 U8108 ( .A1(n6433), .A2(n6703), .ZN(n10292) );
  INV_X1 U8109 ( .A(n10292), .ZN(n9851) );
  AOI22_X1 U8110 ( .A1(n6593), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7155), .B2(
        n9851), .ZN(n6434) );
  INV_X1 U8111 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6444) );
  INV_X1 U8112 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8113 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  NAND2_X1 U8114 ( .A1(n6451), .A2(n6438), .ZN(n9518) );
  OR2_X1 U8115 ( .A1(n9518), .A2(n6529), .ZN(n6443) );
  INV_X1 U8116 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6439) );
  OR2_X1 U8117 ( .A1(n6647), .A2(n6439), .ZN(n6441) );
  INV_X1 U8118 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9838) );
  OR2_X1 U8119 ( .A1(n7169), .A2(n9838), .ZN(n6440) );
  AND2_X1 U8120 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  OAI211_X1 U8121 ( .C1(n6621), .C2(n6444), .A(n6443), .B(n6442), .ZN(n10086)
         );
  NAND2_X1 U8122 ( .A1(n8362), .A2(n10086), .ZN(n8529) );
  NAND2_X1 U8123 ( .A1(n10198), .A2(n9716), .ZN(n8517) );
  NAND2_X1 U8124 ( .A1(n7496), .A2(n6514), .ZN(n6449) );
  NAND2_X1 U8125 ( .A1(n6703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6445) );
  MUX2_X1 U8126 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6445), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6447) );
  NAND2_X1 U8127 ( .A1(n6447), .A2(n6465), .ZN(n9853) );
  INV_X1 U8128 ( .A(n9853), .ZN(n10306) );
  AOI22_X1 U8129 ( .A1(n6593), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7155), .B2(
        n10306), .ZN(n6448) );
  INV_X1 U8130 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8131 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  NAND2_X1 U8132 ( .A1(n6460), .A2(n6452), .ZN(n10089) );
  OR2_X1 U8133 ( .A1(n10089), .A2(n6529), .ZN(n6455) );
  AOI22_X1 U8134 ( .A1(n6618), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n6643), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8135 ( .A1(n7168), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6453) );
  OR2_X1 U8136 ( .A1(n10190), .A2(n9519), .ZN(n8527) );
  NAND2_X1 U8137 ( .A1(n10190), .A2(n9519), .ZN(n8520) );
  NAND2_X1 U8138 ( .A1(n10082), .A2(n10083), .ZN(n10081) );
  NAND2_X1 U8139 ( .A1(n10081), .A2(n8520), .ZN(n10071) );
  NAND2_X1 U8140 ( .A1(n7558), .A2(n6514), .ZN(n6458) );
  NAND2_X1 U8141 ( .A1(n6465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6456) );
  XNOR2_X1 U8142 ( .A(n6456), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U8143 ( .A1(n6593), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7155), .B2(
        n10318), .ZN(n6457) );
  NAND2_X1 U8144 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  AND2_X1 U8145 ( .A1(n6470), .A2(n6461), .ZN(n10067) );
  NAND2_X1 U8146 ( .A1(n10067), .A2(n6418), .ZN(n6464) );
  AOI22_X1 U8147 ( .A1(n6270), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n6643), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6463) );
  INV_X1 U8148 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9847) );
  OR2_X1 U8149 ( .A1(n6647), .A2(n9847), .ZN(n6462) );
  OR2_X1 U8150 ( .A1(n10186), .A2(n10044), .ZN(n8528) );
  NAND2_X1 U8151 ( .A1(n10186), .A2(n10044), .ZN(n10040) );
  NAND2_X1 U8152 ( .A1(n7621), .A2(n6514), .ZN(n6468) );
  NAND2_X1 U8153 ( .A1(n6626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6479) );
  XNOR2_X1 U8154 ( .A(n6479), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U8155 ( .A1(n6593), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7155), .B2(
        n10327), .ZN(n6467) );
  INV_X1 U8156 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U8157 ( .A1(n6470), .A2(n7917), .ZN(n6471) );
  NAND2_X1 U8158 ( .A1(n6487), .A2(n6471), .ZN(n10056) );
  OR2_X1 U8159 ( .A1(n10056), .A2(n6529), .ZN(n6476) );
  INV_X1 U8160 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U8161 ( .A1(n6270), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U8162 ( .A1(n6643), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6472) );
  OAI211_X1 U8163 ( .C1(n9856), .C2(n6647), .A(n6473), .B(n6472), .ZN(n6474)
         );
  INV_X1 U8164 ( .A(n6474), .ZN(n6475) );
  OR2_X1 U8165 ( .A1(n10178), .A2(n10030), .ZN(n8533) );
  NAND2_X1 U8166 ( .A1(n10178), .A2(n10030), .ZN(n8536) );
  NAND2_X1 U8167 ( .A1(n8533), .A2(n8536), .ZN(n8618) );
  INV_X1 U8168 ( .A(n10040), .ZN(n6477) );
  NOR2_X1 U8169 ( .A1(n8618), .A2(n6477), .ZN(n6478) );
  OR2_X1 U8170 ( .A1(n7668), .A2(n8420), .ZN(n6485) );
  NAND2_X1 U8171 ( .A1(n6479), .A2(n6627), .ZN(n6498) );
  NAND2_X1 U8172 ( .A1(n6498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6481) );
  INV_X1 U8173 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6480) );
  OR2_X1 U8174 ( .A1(n6481), .A2(n6480), .ZN(n6483) );
  NAND2_X1 U8175 ( .A1(n6481), .A2(n6480), .ZN(n6482) );
  AOI22_X1 U8176 ( .A1(n6593), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7155), .B2(
        n9858), .ZN(n6484) );
  NAND2_X2 U8177 ( .A1(n6485), .A2(n6484), .ZN(n10174) );
  NAND2_X1 U8178 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  AND2_X1 U8179 ( .A1(n6506), .A2(n6488), .ZN(n10034) );
  NAND2_X1 U8180 ( .A1(n10034), .A2(n6418), .ZN(n6493) );
  INV_X1 U8181 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U8182 ( .A1(n6643), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8183 ( .A1(n7168), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6489) );
  OAI211_X1 U8184 ( .C1(n7970), .C2(n6647), .A(n6490), .B(n6489), .ZN(n6491)
         );
  INV_X1 U8185 ( .A(n6491), .ZN(n6492) );
  OR2_X1 U8186 ( .A1(n10174), .A2(n10046), .ZN(n8534) );
  NAND2_X1 U8187 ( .A1(n10174), .A2(n10046), .ZN(n8537) );
  NAND2_X1 U8188 ( .A1(n7837), .A2(n6514), .ZN(n6504) );
  NAND2_X1 U8189 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n6495) );
  INV_X1 U8190 ( .A(n6498), .ZN(n6496) );
  AND2_X1 U8191 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6497) );
  NAND2_X1 U8192 ( .A1(n6498), .A2(n6497), .ZN(n6499) );
  AOI22_X1 U8193 ( .A1(n6593), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7155), .B2(
        n9865), .ZN(n6503) );
  INV_X1 U8194 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U8195 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  NAND2_X1 U8196 ( .A1(n6517), .A2(n6507), .ZN(n10013) );
  INV_X1 U8197 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U8198 ( .A1(n6643), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8199 ( .A1(n6270), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6508) );
  OAI211_X1 U8200 ( .C1(n6510), .C2(n6647), .A(n6509), .B(n6508), .ZN(n6511)
         );
  INV_X1 U8201 ( .A(n6511), .ZN(n6512) );
  OR2_X1 U8202 ( .A1(n10168), .A2(n10031), .ZN(n8460) );
  NAND2_X1 U8203 ( .A1(n10168), .A2(n10031), .ZN(n8696) );
  NAND2_X1 U8204 ( .A1(n8102), .A2(n6514), .ZN(n6516) );
  NAND2_X1 U8205 ( .A1(n6593), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U8206 ( .A1(n6517), .A2(n9650), .ZN(n6518) );
  AND2_X1 U8207 ( .A1(n6527), .A2(n6518), .ZN(n10003) );
  NAND2_X1 U8208 ( .A1(n10003), .A2(n6418), .ZN(n6524) );
  INV_X1 U8209 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8210 ( .A1(n6643), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8211 ( .A1(n7168), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6519) );
  OAI211_X1 U8212 ( .C1(n6521), .C2(n6647), .A(n6520), .B(n6519), .ZN(n6522)
         );
  INV_X1 U8213 ( .A(n6522), .ZN(n6523) );
  XNOR2_X1 U8214 ( .A(n10004), .B(n9982), .ZN(n8619) );
  OR2_X1 U8215 ( .A1(n10004), .A2(n9982), .ZN(n8461) );
  NAND2_X1 U8216 ( .A1(n8223), .A2(n6514), .ZN(n6526) );
  NAND2_X1 U8217 ( .A1(n6593), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6525) );
  INV_X1 U8218 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U8219 ( .A1(n6527), .A2(n9574), .ZN(n6528) );
  NAND2_X1 U8220 ( .A1(n6540), .A2(n6528), .ZN(n9989) );
  INV_X1 U8221 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8222 ( .A1(n6270), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8223 ( .A1(n6643), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6530) );
  OAI211_X1 U8224 ( .C1(n6532), .C2(n6647), .A(n6531), .B(n6530), .ZN(n6533)
         );
  INV_X1 U8225 ( .A(n6533), .ZN(n6534) );
  OR2_X1 U8226 ( .A1(n10231), .A2(n9996), .ZN(n8640) );
  NAND2_X1 U8227 ( .A1(n10231), .A2(n9996), .ZN(n8543) );
  NAND2_X1 U8228 ( .A1(n9979), .A2(n9981), .ZN(n9980) );
  NAND2_X1 U8229 ( .A1(n9980), .A2(n8543), .ZN(n9970) );
  NAND2_X1 U8230 ( .A1(n8303), .A2(n6514), .ZN(n6537) );
  NAND2_X1 U8231 ( .A1(n6593), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6536) );
  INV_X1 U8232 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8233 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  NAND2_X1 U8234 ( .A1(n6550), .A2(n6541), .ZN(n9675) );
  OR2_X1 U8235 ( .A1(n9675), .A2(n6617), .ZN(n6547) );
  INV_X1 U8236 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8237 ( .A1(n7168), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U8238 ( .A1(n6643), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6542) );
  OAI211_X1 U8239 ( .C1(n6544), .C2(n6647), .A(n6543), .B(n6542), .ZN(n6545)
         );
  INV_X1 U8240 ( .A(n6545), .ZN(n6546) );
  OR2_X1 U8241 ( .A1(n10151), .A2(n9983), .ZN(n8549) );
  NAND2_X1 U8242 ( .A1(n10151), .A2(n9983), .ZN(n8548) );
  NAND2_X1 U8243 ( .A1(n8374), .A2(n6514), .ZN(n6549) );
  NAND2_X1 U8244 ( .A1(n6593), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6548) );
  NAND2_X2 U8245 ( .A1(n6549), .A2(n6548), .ZN(n10226) );
  INV_X1 U8246 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U8247 ( .A1(n6550), .A2(n9529), .ZN(n6551) );
  NAND2_X1 U8248 ( .A1(n6561), .A2(n6551), .ZN(n9951) );
  INV_X1 U8249 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8250 ( .A1(n6643), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U8251 ( .A1(n6270), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6552) );
  OAI211_X1 U8252 ( .C1(n6554), .C2(n6647), .A(n6553), .B(n6552), .ZN(n6555)
         );
  INV_X1 U8253 ( .A(n6555), .ZN(n6556) );
  OR2_X1 U8254 ( .A1(n10226), .A2(n9629), .ZN(n8550) );
  NAND2_X1 U8255 ( .A1(n10226), .A2(n9629), .ZN(n9929) );
  NAND2_X1 U8256 ( .A1(n9501), .A2(n6514), .ZN(n6559) );
  NAND2_X1 U8257 ( .A1(n6593), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6558) );
  INV_X1 U8258 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U8259 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  NAND2_X1 U8260 ( .A1(n9937), .A2(n6418), .ZN(n6567) );
  INV_X1 U8261 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U8262 ( .A1(n6643), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6564) );
  INV_X1 U8263 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n7927) );
  OR2_X1 U8264 ( .A1(n6621), .A2(n7927), .ZN(n6563) );
  OAI211_X1 U8265 ( .C1(n6647), .C2(n7960), .A(n6564), .B(n6563), .ZN(n6565)
         );
  INV_X1 U8266 ( .A(n6565), .ZN(n6566) );
  NAND2_X1 U8267 ( .A1(n10139), .A2(n9915), .ZN(n8645) );
  INV_X1 U8268 ( .A(n9929), .ZN(n6568) );
  NAND2_X1 U8269 ( .A1(n8450), .A2(n6514), .ZN(n6571) );
  NAND2_X1 U8270 ( .A1(n6593), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6570) );
  INV_X1 U8271 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U8272 ( .A1(n6572), .A2(n9597), .ZN(n6573) );
  NAND2_X1 U8273 ( .A1(n6584), .A2(n6573), .ZN(n9918) );
  OR2_X1 U8274 ( .A1(n9918), .A2(n6617), .ZN(n6578) );
  INV_X1 U8275 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10136) );
  NAND2_X1 U8276 ( .A1(n6643), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U8277 ( .A1(n7168), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6574) );
  OAI211_X1 U8278 ( .C1(n6647), .C2(n10136), .A(n6575), .B(n6574), .ZN(n6576)
         );
  INV_X1 U8279 ( .A(n6576), .ZN(n6577) );
  NAND2_X1 U8280 ( .A1(n9921), .A2(n9707), .ZN(n8572) );
  NAND2_X1 U8281 ( .A1(n8635), .A2(n8572), .ZN(n9913) );
  NAND2_X1 U8282 ( .A1(n9911), .A2(n8572), .ZN(n9903) );
  NAND2_X1 U8283 ( .A1(n9498), .A2(n6514), .ZN(n6581) );
  NAND2_X1 U8284 ( .A1(n6593), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6580) );
  INV_X1 U8285 ( .A(n6584), .ZN(n6582) );
  NAND2_X1 U8286 ( .A1(n6582), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6597) );
  INV_X1 U8287 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8288 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NAND2_X1 U8289 ( .A1(n6597), .A2(n6585), .ZN(n9704) );
  OR2_X1 U8290 ( .A1(n9704), .A2(n6617), .ZN(n6591) );
  INV_X1 U8291 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8292 ( .A1(n6643), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U8293 ( .A1(n6270), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6586) );
  OAI211_X1 U8294 ( .C1(n6588), .C2(n6647), .A(n6587), .B(n6586), .ZN(n6589)
         );
  INV_X1 U8295 ( .A(n6589), .ZN(n6590) );
  NAND2_X1 U8296 ( .A1(n10129), .A2(n9916), .ZN(n8701) );
  NAND2_X1 U8297 ( .A1(n9493), .A2(n6592), .ZN(n6595) );
  NAND2_X1 U8298 ( .A1(n6593), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6594) );
  NAND2_X2 U8299 ( .A1(n6595), .A2(n6594), .ZN(n10127) );
  INV_X1 U8300 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8301 ( .A1(n6597), .A2(n6596), .ZN(n6598) );
  NAND2_X1 U8302 ( .A1(n9509), .A2(n6418), .ZN(n6603) );
  INV_X1 U8303 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U8304 ( .A1(n6618), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U8305 ( .A1(n6643), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6599) );
  OAI211_X1 U8306 ( .C1(n6621), .C2(n7909), .A(n6600), .B(n6599), .ZN(n6601)
         );
  INV_X1 U8307 ( .A(n6601), .ZN(n6602) );
  NAND2_X1 U8308 ( .A1(n10127), .A2(n8559), .ZN(n8555) );
  NAND2_X1 U8309 ( .A1(n8428), .A2(n6514), .ZN(n6605) );
  NAND2_X1 U8310 ( .A1(n6593), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6604) );
  INV_X1 U8311 ( .A(n6607), .ZN(n6606) );
  NAND2_X1 U8312 ( .A1(n6606), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9878) );
  INV_X1 U8313 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U8314 ( .A1(n6607), .A2(n7963), .ZN(n6608) );
  NAND2_X1 U8315 ( .A1(n9878), .A2(n6608), .ZN(n9888) );
  INV_X1 U8316 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8317 ( .A1(n6643), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U8318 ( .A1(n7168), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6609) );
  OAI211_X1 U8319 ( .C1(n6611), .C2(n6647), .A(n6610), .B(n6609), .ZN(n6612)
         );
  INV_X1 U8320 ( .A(n6612), .ZN(n6613) );
  NAND2_X1 U8321 ( .A1(n9890), .A2(n8562), .ZN(n8557) );
  AND2_X1 U8322 ( .A1(n8557), .A2(n8555), .ZN(n8651) );
  NAND2_X1 U8323 ( .A1(n6788), .A2(n8653), .ZN(n6625) );
  NAND2_X1 U8324 ( .A1(n8388), .A2(n6514), .ZN(n6616) );
  NAND2_X1 U8325 ( .A1(n6593), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6615) );
  OR2_X1 U8326 ( .A1(n9878), .A2(n6617), .ZN(n6624) );
  INV_X1 U8327 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U8328 ( .A1(n6618), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8329 ( .A1(n6643), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6619) );
  OAI211_X1 U8330 ( .C1(n7928), .C2(n6621), .A(n6620), .B(n6619), .ZN(n6622)
         );
  INV_X1 U8331 ( .A(n6622), .ZN(n6623) );
  NAND2_X1 U8332 ( .A1(n9880), .A2(n7049), .ZN(n8707) );
  XNOR2_X1 U8333 ( .A(n6625), .B(n8593), .ZN(n6640) );
  INV_X1 U8334 ( .A(n6626), .ZN(n6629) );
  NAND2_X1 U8335 ( .A1(n6635), .A2(n6636), .ZN(n6630) );
  NAND2_X1 U8336 ( .A1(n8588), .A2(n9865), .ZN(n6639) );
  NAND2_X1 U8337 ( .A1(n4914), .A2(n6650), .ZN(n8587) );
  NAND2_X1 U8338 ( .A1(n6640), .A2(n10087), .ZN(n6649) );
  INV_X1 U8339 ( .A(P1_B_REG_SCAN_IN), .ZN(n6641) );
  NOR2_X1 U8340 ( .A1(n10249), .A2(n6641), .ZN(n6642) );
  NOR2_X1 U8341 ( .A1(n10045), .A2(n6642), .ZN(n8425) );
  INV_X1 U8342 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U8343 ( .A1(n6643), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8344 ( .A1(n7168), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6644) );
  OAI211_X1 U8345 ( .C1(n6647), .C2(n6646), .A(n6645), .B(n6644), .ZN(n9726)
         );
  AOI22_X1 U8346 ( .A1(n9728), .A2(n10085), .B1(n8425), .B2(n9726), .ZN(n6648)
         );
  AND2_X1 U8347 ( .A1(n6651), .A2(n10380), .ZN(n6652) );
  NAND2_X1 U8348 ( .A1(n7156), .A2(n6802), .ZN(n7047) );
  NAND2_X1 U8349 ( .A1(n6652), .A2(n7047), .ZN(n8052) );
  OR2_X1 U8350 ( .A1(n8593), .A2(n10401), .ZN(n6701) );
  NAND2_X1 U8351 ( .A1(n6653), .A2(n8467), .ZN(n7600) );
  INV_X1 U8352 ( .A(n10381), .ZN(n6808) );
  NAND2_X1 U8353 ( .A1(n9745), .A2(n6808), .ZN(n7476) );
  NAND2_X1 U8354 ( .A1(n6319), .A2(n9567), .ZN(n6654) );
  NAND2_X1 U8355 ( .A1(n7476), .A2(n6654), .ZN(n6658) );
  NAND3_X1 U8356 ( .A1(n6656), .A2(n4437), .A3(n6655), .ZN(n6657) );
  NAND2_X1 U8357 ( .A1(n6658), .A2(n6657), .ZN(n7487) );
  NAND2_X1 U8358 ( .A1(n8599), .A2(n7487), .ZN(n7486) );
  NAND2_X1 U8359 ( .A1(n7478), .A2(n8016), .ZN(n6659) );
  NAND2_X1 U8360 ( .A1(n7486), .A2(n6659), .ZN(n7601) );
  NOR2_X1 U8361 ( .A1(n9742), .A2(n4278), .ZN(n7715) );
  NOR2_X1 U8362 ( .A1(n9741), .A2(n7730), .ZN(n6660) );
  AOI21_X1 U8363 ( .B1(n8603), .B2(n7715), .A(n6660), .ZN(n6661) );
  NAND2_X1 U8364 ( .A1(n8481), .A2(n8674), .ZN(n7707) );
  INV_X1 U8365 ( .A(n8478), .ZN(n8046) );
  NAND2_X1 U8366 ( .A1(n8046), .A2(n8486), .ZN(n8045) );
  NOR2_X1 U8367 ( .A1(n9740), .A2(n10354), .ZN(n7999) );
  NOR2_X1 U8368 ( .A1(n4902), .A2(n9739), .ZN(n8042) );
  AOI21_X1 U8369 ( .B1(n7999), .B2(n8045), .A(n8042), .ZN(n6662) );
  INV_X1 U8370 ( .A(n8175), .ZN(n9738) );
  OR2_X1 U8371 ( .A1(n8074), .A2(n9738), .ZN(n8170) );
  NAND2_X1 U8372 ( .A1(n6662), .A2(n8170), .ZN(n6664) );
  NAND2_X1 U8373 ( .A1(n8149), .A2(n8491), .ZN(n8178) );
  NAND2_X1 U8374 ( .A1(n8188), .A2(n7676), .ZN(n6666) );
  NAND2_X1 U8375 ( .A1(n8501), .A2(n8497), .ZN(n8151) );
  INV_X1 U8376 ( .A(n8232), .ZN(n9736) );
  OR2_X1 U8377 ( .A1(n10102), .A2(n9735), .ZN(n6667) );
  INV_X1 U8378 ( .A(n9546), .ZN(n9734) );
  OR2_X1 U8379 ( .A1(n9690), .A2(n9734), .ZN(n6668) );
  NAND2_X1 U8380 ( .A1(n8512), .A2(n9682), .ZN(n6669) );
  NAND2_X1 U8381 ( .A1(n9666), .A2(n9583), .ZN(n6670) );
  NAND2_X1 U8382 ( .A1(n10198), .A2(n10086), .ZN(n6671) );
  INV_X1 U8383 ( .A(n10044), .ZN(n10084) );
  NAND2_X1 U8384 ( .A1(n10186), .A2(n10084), .ZN(n6672) );
  OR2_X1 U8385 ( .A1(n10178), .A2(n10074), .ZN(n6673) );
  NAND2_X1 U8386 ( .A1(n10050), .A2(n6673), .ZN(n6675) );
  NAND2_X1 U8387 ( .A1(n10178), .A2(n10074), .ZN(n6674) );
  AND2_X1 U8388 ( .A1(n10174), .A2(n10020), .ZN(n6676) );
  NAND2_X1 U8389 ( .A1(n10168), .A2(n9731), .ZN(n6677) );
  AND2_X1 U8390 ( .A1(n10004), .A2(n10021), .ZN(n6679) );
  NOR2_X1 U8391 ( .A1(n10231), .A2(n9973), .ZN(n6680) );
  NAND2_X1 U8392 ( .A1(n10231), .A2(n9973), .ZN(n6681) );
  AND2_X1 U8393 ( .A1(n10151), .A2(n9730), .ZN(n6683) );
  OR2_X1 U8394 ( .A1(n10151), .A2(n9730), .ZN(n6684) );
  NOR2_X1 U8395 ( .A1(n10226), .A2(n9972), .ZN(n6685) );
  OR2_X1 U8396 ( .A1(n10139), .A2(n9950), .ZN(n6686) );
  NAND2_X1 U8397 ( .A1(n10139), .A2(n9950), .ZN(n6687) );
  AND2_X1 U8398 ( .A1(n9921), .A2(n9932), .ZN(n6690) );
  OR2_X1 U8399 ( .A1(n9921), .A2(n9932), .ZN(n6689) );
  NOR2_X1 U8400 ( .A1(n10129), .A2(n9729), .ZN(n8398) );
  OR2_X1 U8401 ( .A1(n8398), .A2(n5119), .ZN(n6691) );
  NAND2_X1 U8402 ( .A1(n10129), .A2(n9729), .ZN(n8399) );
  AND2_X1 U8403 ( .A1(n8400), .A2(n8399), .ZN(n6692) );
  NAND2_X1 U8404 ( .A1(n8653), .A2(n8557), .ZN(n8626) );
  NAND2_X1 U8405 ( .A1(n9890), .A2(n9728), .ZN(n9873) );
  NAND4_X1 U8406 ( .A1(n9874), .A2(n8593), .A3(n10195), .A4(n9873), .ZN(n6700)
         );
  INV_X1 U8407 ( .A(n9880), .ZN(n6698) );
  OR3_X1 U8408 ( .A1(n8593), .A2(n10401), .A3(n9873), .ZN(n6697) );
  INV_X1 U8409 ( .A(n10129), .ZN(n9902) );
  INV_X1 U8410 ( .A(n10151), .ZN(n9968) );
  INV_X1 U8411 ( .A(n10113), .ZN(n9645) );
  INV_X1 U8412 ( .A(n10102), .ZN(n9551) );
  INV_X1 U8413 ( .A(n10174), .ZN(n10037) );
  INV_X1 U8414 ( .A(n10004), .ZN(n10163) );
  NAND2_X1 U8415 ( .A1(n9968), .A2(n9986), .ZN(n9963) );
  NOR2_X2 U8416 ( .A1(n9963), .A2(n10226), .ZN(n9934) );
  NAND2_X1 U8417 ( .A1(n6696), .A2(n9867), .ZN(n9882) );
  OAI211_X1 U8418 ( .C1(n6698), .C2(n10180), .A(n6697), .B(n9882), .ZN(n6699)
         );
  NAND2_X1 U8419 ( .A1(n6709), .A2(n6704), .ZN(n6711) );
  OAI21_X1 U8420 ( .B1(n6711), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U8421 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6705), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6706) );
  INV_X1 U8422 ( .A(n6728), .ZN(n10255) );
  NAND2_X1 U8423 ( .A1(n6711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8424 ( .A1(n4694), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6710) );
  MUX2_X1 U8425 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6710), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6712) );
  NAND3_X1 U8426 ( .A1(n10258), .A2(n10263), .A3(P1_B_REG_SCAN_IN), .ZN(n6713)
         );
  NOR2_X1 U8427 ( .A1(n7161), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6724) );
  NOR4_X1 U8428 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6717) );
  NOR4_X1 U8429 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6716) );
  NOR4_X1 U8430 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6715) );
  NOR4_X1 U8431 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6714) );
  NAND4_X1 U8432 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6723)
         );
  NOR2_X1 U8433 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n6721) );
  NOR4_X1 U8434 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6720) );
  NOR4_X1 U8435 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6719) );
  NOR4_X1 U8436 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6718) );
  NAND4_X1 U8437 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6722)
         );
  NOR2_X1 U8438 ( .A1(n6723), .A2(n6722), .ZN(n7030) );
  OAI222_X1 U8439 ( .A1(n10091), .A2(n8590), .B1(n7164), .B2(n6724), .C1(n7161), .C2(n7030), .ZN(n6734) );
  NAND2_X1 U8440 ( .A1(n10255), .A2(n10263), .ZN(n10245) );
  OAI21_X1 U8441 ( .B1(n7161), .B2(P1_D_REG_0__SCAN_IN), .A(n10245), .ZN(n7790) );
  NOR2_X1 U8442 ( .A1(n6734), .A2(n7790), .ZN(n6730) );
  NAND2_X1 U8443 ( .A1(n7156), .A2(n8716), .ZN(n7052) );
  INV_X1 U8444 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6731) );
  OR2_X1 U8445 ( .A1(n10408), .A2(n6731), .ZN(n6732) );
  NAND2_X1 U8446 ( .A1(n6733), .A2(n6732), .ZN(P1_U3551) );
  INV_X1 U8447 ( .A(n7790), .ZN(n7033) );
  NOR2_X1 U8448 ( .A1(n6734), .A2(n7033), .ZN(n6735) );
  OR2_X1 U8449 ( .A1(n10405), .A2(n7928), .ZN(n6736) );
  NAND2_X1 U8450 ( .A1(n6737), .A2(n6736), .ZN(P1_U3519) );
  INV_X1 U8451 ( .A(n6759), .ZN(n6743) );
  AND2_X1 U8452 ( .A1(n6739), .A2(P2_B_REG_SCAN_IN), .ZN(n6740) );
  NOR2_X1 U8453 ( .A1(n9298), .A2(n6740), .ZN(n9145) );
  AOI22_X1 U8454 ( .A1(n9331), .A2(n8913), .B1(n8911), .B2(n9145), .ZN(n6741)
         );
  INV_X1 U8455 ( .A(n6746), .ZN(n6745) );
  INV_X1 U8456 ( .A(n6752), .ZN(n6749) );
  NAND2_X1 U8457 ( .A1(n9419), .A2(n8913), .ZN(n6750) );
  AND2_X1 U8458 ( .A1(n6749), .A2(n6750), .ZN(n6744) );
  NAND2_X1 U8459 ( .A1(n6745), .A2(n6744), .ZN(n6757) );
  OR2_X1 U8460 ( .A1(n9419), .A2(n8913), .ZN(n6747) );
  NAND2_X1 U8461 ( .A1(n6746), .A2(n5118), .ZN(n6756) );
  INV_X1 U8462 ( .A(n6747), .ZN(n6748) );
  AOI21_X1 U8463 ( .B1(n6749), .B2(n6748), .A(n9293), .ZN(n6754) );
  INV_X1 U8464 ( .A(n6750), .ZN(n6751) );
  NAND2_X1 U8465 ( .A1(n6752), .A2(n6751), .ZN(n6753) );
  NAND3_X1 U8466 ( .A1(n6757), .A2(n6756), .A3(n6755), .ZN(n6758) );
  OAI21_X1 U8467 ( .B1(n6062), .B2(n6762), .A(n6761), .ZN(n6766) );
  NAND2_X1 U8468 ( .A1(n6764), .A2(n6763), .ZN(n6765) );
  NAND2_X1 U8469 ( .A1(n6766), .A2(n6765), .ZN(n6767) );
  OR2_X1 U8470 ( .A1(n6774), .A2(n10446), .ZN(n6773) );
  INV_X1 U8471 ( .A(n6769), .ZN(n9154) );
  INV_X1 U8472 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U8473 ( .A1(n6773), .A2(n6772), .ZN(P2_U3488) );
  OR2_X1 U8474 ( .A1(n6774), .A2(n10441), .ZN(n6778) );
  NOR2_X1 U8475 ( .A1(n10440), .A2(n6775), .ZN(n6776) );
  NAND2_X1 U8476 ( .A1(n6778), .A2(n6777), .ZN(P2_U3456) );
  INV_X1 U8477 ( .A(n6779), .ZN(n6781) );
  INV_X1 U8478 ( .A(n8626), .ZN(n6780) );
  NAND2_X1 U8479 ( .A1(n6781), .A2(n6780), .ZN(n6782) );
  INV_X1 U8480 ( .A(n8653), .ZN(n6787) );
  INV_X1 U8481 ( .A(n8404), .ZN(n6783) );
  NAND2_X1 U8482 ( .A1(n6783), .A2(n8626), .ZN(n6786) );
  INV_X1 U8483 ( .A(n8555), .ZN(n6784) );
  AOI21_X1 U8484 ( .B1(n8626), .B2(n6784), .A(n10392), .ZN(n6785) );
  OAI211_X1 U8485 ( .C1(n6788), .C2(n6787), .A(n6786), .B(n6785), .ZN(n6791)
         );
  OAI22_X1 U8486 ( .A1(n7049), .A2(n10045), .B1(n8559), .B2(n10043), .ZN(n6789) );
  INV_X1 U8487 ( .A(n6789), .ZN(n6790) );
  AOI21_X1 U8488 ( .B1(n9890), .B2(n4337), .A(n10091), .ZN(n6793) );
  NAND2_X1 U8489 ( .A1(n6793), .A2(n6792), .ZN(n9892) );
  INV_X1 U8490 ( .A(n10159), .ZN(n6796) );
  NAND2_X1 U8491 ( .A1(n6797), .A2(n5103), .ZN(P1_U3550) );
  OR2_X1 U8492 ( .A1(n10405), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6799) );
  INV_X1 U8493 ( .A(n10232), .ZN(n6800) );
  NAND2_X1 U8494 ( .A1(n6801), .A2(n5102), .ZN(P1_U3518) );
  NAND2_X1 U8495 ( .A1(n6821), .A2(n6808), .ZN(n6805) );
  NAND2_X1 U8496 ( .A1(n9745), .A2(n6834), .ZN(n6804) );
  INV_X1 U8497 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U8498 ( .A1(n5100), .A2(n5110), .ZN(n7359) );
  NAND2_X1 U8499 ( .A1(n7035), .A2(n9745), .ZN(n6810) );
  AOI22_X1 U8500 ( .A1(n6808), .A2(n6834), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6807), .ZN(n6809) );
  NAND2_X1 U8501 ( .A1(n6810), .A2(n6809), .ZN(n7358) );
  NAND2_X1 U8502 ( .A1(n7359), .A2(n7358), .ZN(n7357) );
  NAND2_X1 U8503 ( .A1(n5100), .A2(n6849), .ZN(n6811) );
  NAND2_X1 U8504 ( .A1(n6319), .A2(n6834), .ZN(n6813) );
  NAND2_X1 U8505 ( .A1(n6821), .A2(n9567), .ZN(n6812) );
  NAND2_X1 U8506 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U8507 ( .A1(n6319), .A2(n7035), .ZN(n6816) );
  NAND2_X1 U8508 ( .A1(n6834), .A2(n9567), .ZN(n6815) );
  NAND2_X1 U8509 ( .A1(n6816), .A2(n6815), .ZN(n6817) );
  XNOR2_X1 U8510 ( .A(n6819), .B(n6817), .ZN(n9565) );
  NAND2_X1 U8511 ( .A1(n9564), .A2(n9565), .ZN(n9563) );
  INV_X1 U8512 ( .A(n6817), .ZN(n6818) );
  NAND2_X1 U8513 ( .A1(n6819), .A2(n6818), .ZN(n6820) );
  NAND2_X1 U8514 ( .A1(n9563), .A2(n6820), .ZN(n7406) );
  NAND2_X1 U8515 ( .A1(n6821), .A2(n7500), .ZN(n6823) );
  NAND2_X1 U8516 ( .A1(n9743), .A2(n6834), .ZN(n6822) );
  NAND2_X1 U8517 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  XNOR2_X1 U8518 ( .A(n6824), .B(n6849), .ZN(n6829) );
  NAND2_X1 U8519 ( .A1(n7035), .A2(n9743), .ZN(n6826) );
  NAND2_X1 U8520 ( .A1(n7500), .A2(n6834), .ZN(n6825) );
  NAND2_X1 U8521 ( .A1(n6826), .A2(n6825), .ZN(n6827) );
  XNOR2_X1 U8522 ( .A(n6829), .B(n6827), .ZN(n7407) );
  INV_X1 U8523 ( .A(n6827), .ZN(n6828) );
  NAND2_X1 U8524 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  NAND2_X1 U8525 ( .A1(n6821), .A2(n4278), .ZN(n6832) );
  NAND2_X1 U8526 ( .A1(n9742), .A2(n6834), .ZN(n6831) );
  NAND2_X1 U8527 ( .A1(n6832), .A2(n6831), .ZN(n6833) );
  XNOR2_X1 U8528 ( .A(n6833), .B(n6849), .ZN(n6839) );
  NAND2_X1 U8529 ( .A1(n7035), .A2(n9742), .ZN(n6836) );
  NAND2_X1 U8530 ( .A1(n4278), .A2(n7016), .ZN(n6835) );
  INV_X1 U8531 ( .A(n6837), .ZN(n6838) );
  NAND2_X1 U8532 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  NAND2_X1 U8533 ( .A1(n6821), .A2(n7730), .ZN(n6841) );
  OAI21_X1 U8534 ( .B1(n7455), .B2(n6851), .A(n6841), .ZN(n6842) );
  XNOR2_X1 U8535 ( .A(n6842), .B(n7004), .ZN(n6845) );
  INV_X2 U8536 ( .A(n6851), .ZN(n7016) );
  NAND2_X1 U8537 ( .A1(n7730), .A2(n7016), .ZN(n6843) );
  OAI21_X1 U8538 ( .B1(n7455), .B2(n7020), .A(n6843), .ZN(n6844) );
  XNOR2_X1 U8539 ( .A(n6845), .B(n6844), .ZN(n7660) );
  OR2_X2 U8540 ( .A1(n7659), .A2(n7660), .ZN(n7657) );
  NAND2_X1 U8541 ( .A1(n6845), .A2(n6844), .ZN(n6846) );
  NAND2_X1 U8542 ( .A1(n7657), .A2(n6846), .ZN(n7733) );
  NAND2_X1 U8543 ( .A1(n4902), .A2(n7015), .ZN(n6848) );
  NAND2_X1 U8544 ( .A1(n9739), .A2(n7016), .ZN(n6847) );
  NAND2_X1 U8545 ( .A1(n6848), .A2(n6847), .ZN(n6850) );
  XNOR2_X1 U8546 ( .A(n6850), .B(n6849), .ZN(n7736) );
  NAND2_X1 U8547 ( .A1(n4902), .A2(n7016), .ZN(n6853) );
  NAND2_X1 U8548 ( .A1(n9739), .A2(n7035), .ZN(n6852) );
  AND2_X1 U8549 ( .A1(n6853), .A2(n6852), .ZN(n6859) );
  NAND2_X1 U8550 ( .A1(n10354), .A2(n7015), .ZN(n6855) );
  NAND2_X1 U8551 ( .A1(n9740), .A2(n7016), .ZN(n6854) );
  NAND2_X1 U8552 ( .A1(n6855), .A2(n6854), .ZN(n6856) );
  XNOR2_X1 U8553 ( .A(n6856), .B(n6849), .ZN(n6862) );
  OR2_X1 U8554 ( .A1(n7775), .A2(n6851), .ZN(n6858) );
  NAND2_X1 U8555 ( .A1(n7035), .A2(n9740), .ZN(n6857) );
  OAI22_X1 U8556 ( .A1(n7736), .A2(n6859), .B1(n6862), .B2(n7772), .ZN(n6865)
         );
  INV_X1 U8557 ( .A(n6862), .ZN(n7734) );
  INV_X1 U8558 ( .A(n7772), .ZN(n6860) );
  INV_X1 U8559 ( .A(n6859), .ZN(n7735) );
  OAI21_X1 U8560 ( .B1(n7734), .B2(n6860), .A(n7735), .ZN(n6863) );
  NOR2_X1 U8561 ( .A1(n7735), .A2(n6860), .ZN(n6861) );
  AOI22_X1 U8562 ( .A1(n6863), .A2(n7736), .B1(n6862), .B2(n6861), .ZN(n6864)
         );
  OAI21_X2 U8563 ( .B1(n7733), .B2(n6865), .A(n6864), .ZN(n7673) );
  NOR2_X1 U8564 ( .A1(n8175), .A2(n4284), .ZN(n6866) );
  AOI21_X1 U8565 ( .B1(n8074), .B2(n7016), .A(n6866), .ZN(n6870) );
  NAND2_X1 U8566 ( .A1(n8074), .A2(n7015), .ZN(n6868) );
  NAND2_X1 U8567 ( .A1(n9738), .A2(n7016), .ZN(n6867) );
  NAND2_X1 U8568 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  XNOR2_X1 U8569 ( .A(n6869), .B(n7004), .ZN(n7671) );
  INV_X1 U8570 ( .A(n6870), .ZN(n7670) );
  NAND2_X1 U8571 ( .A1(n10113), .A2(n6821), .ZN(n6872) );
  NAND2_X1 U8572 ( .A1(n9736), .A2(n7016), .ZN(n6871) );
  NAND2_X1 U8573 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  XNOR2_X1 U8574 ( .A(n6873), .B(n7004), .ZN(n6884) );
  NOR2_X1 U8575 ( .A1(n8232), .A2(n7020), .ZN(n6874) );
  AOI21_X1 U8576 ( .B1(n10113), .B2(n7016), .A(n6874), .ZN(n6885) );
  XNOR2_X1 U8577 ( .A(n6884), .B(n6885), .ZN(n9635) );
  OAI22_X1 U8578 ( .A1(n8188), .A2(n6930), .B1(n7676), .B2(n6851), .ZN(n6875)
         );
  XNOR2_X1 U8579 ( .A(n6875), .B(n7004), .ZN(n8227) );
  OAI22_X1 U8580 ( .A1(n8188), .A2(n6851), .B1(n7676), .B2(n4284), .ZN(n8230)
         );
  NAND2_X1 U8581 ( .A1(n8227), .A2(n8230), .ZN(n6876) );
  AND2_X1 U8582 ( .A1(n9635), .A2(n6876), .ZN(n9537) );
  INV_X1 U8583 ( .A(n9537), .ZN(n6889) );
  INV_X1 U8584 ( .A(n8227), .ZN(n6878) );
  INV_X1 U8585 ( .A(n8230), .ZN(n6877) );
  AND2_X1 U8586 ( .A1(n6878), .A2(n6877), .ZN(n9538) );
  NAND2_X1 U8587 ( .A1(n10102), .A2(n7015), .ZN(n6880) );
  NAND2_X1 U8588 ( .A1(n9735), .A2(n7016), .ZN(n6879) );
  NAND2_X1 U8589 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  XNOR2_X1 U8590 ( .A(n6881), .B(n7004), .ZN(n9541) );
  NAND2_X1 U8591 ( .A1(n10102), .A2(n7016), .ZN(n6883) );
  NAND2_X1 U8592 ( .A1(n9735), .A2(n7035), .ZN(n6882) );
  NAND2_X1 U8593 ( .A1(n6883), .A2(n6882), .ZN(n9535) );
  INV_X1 U8594 ( .A(n6884), .ZN(n6886) );
  NAND2_X1 U8595 ( .A1(n6886), .A2(n6885), .ZN(n9540) );
  OAI21_X1 U8596 ( .B1(n9541), .B2(n9535), .A(n9540), .ZN(n6887) );
  NAND2_X1 U8597 ( .A1(n9690), .A2(n7015), .ZN(n6891) );
  NAND2_X1 U8598 ( .A1(n9734), .A2(n7016), .ZN(n6890) );
  NAND2_X1 U8599 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  NOR2_X1 U8600 ( .A1(n9546), .A2(n7020), .ZN(n6893) );
  AOI21_X1 U8601 ( .B1(n9690), .B2(n7016), .A(n6893), .ZN(n6894) );
  NAND2_X1 U8602 ( .A1(n6895), .A2(n6894), .ZN(n9587) );
  AND2_X1 U8603 ( .A1(n9541), .A2(n9535), .ZN(n6896) );
  OAI22_X1 U8604 ( .A1(n8512), .A2(n6930), .B1(n9682), .B2(n6851), .ZN(n6898)
         );
  XNOR2_X1 U8605 ( .A(n6898), .B(n6849), .ZN(n6900) );
  OAI22_X1 U8606 ( .A1(n8512), .A2(n6851), .B1(n9682), .B2(n7020), .ZN(n6901)
         );
  INV_X1 U8607 ( .A(n6901), .ZN(n6899) );
  NAND2_X1 U8608 ( .A1(n6900), .A2(n6899), .ZN(n6904) );
  INV_X1 U8609 ( .A(n6900), .ZN(n6902) );
  NAND2_X1 U8610 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  AND2_X1 U8611 ( .A1(n6904), .A2(n6903), .ZN(n9585) );
  NAND2_X1 U8612 ( .A1(n9589), .A2(n6904), .ZN(n9657) );
  OAI22_X1 U8613 ( .A1(n9666), .A2(n6930), .B1(n9583), .B2(n6851), .ZN(n6905)
         );
  XNOR2_X1 U8614 ( .A(n6905), .B(n6849), .ZN(n6908) );
  OAI22_X1 U8615 ( .A1(n9666), .A2(n6851), .B1(n9583), .B2(n4284), .ZN(n6906)
         );
  XNOR2_X1 U8616 ( .A(n6908), .B(n6906), .ZN(n9658) );
  NAND2_X1 U8617 ( .A1(n9657), .A2(n9658), .ZN(n9656) );
  INV_X1 U8618 ( .A(n6906), .ZN(n6907) );
  NAND2_X1 U8619 ( .A1(n6908), .A2(n6907), .ZN(n6909) );
  OAI22_X1 U8620 ( .A1(n8362), .A2(n6930), .B1(n9716), .B2(n6851), .ZN(n6910)
         );
  XNOR2_X1 U8621 ( .A(n6910), .B(n6849), .ZN(n6911) );
  OAI22_X1 U8622 ( .A1(n8362), .A2(n6851), .B1(n9716), .B2(n4284), .ZN(n9517)
         );
  NAND2_X1 U8623 ( .A1(n10190), .A2(n6821), .ZN(n6915) );
  OR2_X1 U8624 ( .A1(n9519), .A2(n6851), .ZN(n6914) );
  NAND2_X1 U8625 ( .A1(n6915), .A2(n6914), .ZN(n6916) );
  XNOR2_X1 U8626 ( .A(n6916), .B(n6849), .ZN(n9602) );
  NOR2_X1 U8627 ( .A1(n9519), .A2(n4284), .ZN(n6917) );
  AOI21_X1 U8628 ( .B1(n10190), .B2(n7016), .A(n6917), .ZN(n6922) );
  AND2_X1 U8629 ( .A1(n9602), .A2(n6922), .ZN(n6926) );
  NAND2_X1 U8630 ( .A1(n10186), .A2(n6821), .ZN(n6919) );
  OR2_X1 U8631 ( .A1(n10044), .A2(n6851), .ZN(n6918) );
  NAND2_X1 U8632 ( .A1(n6919), .A2(n6918), .ZN(n6920) );
  XNOR2_X1 U8633 ( .A(n6920), .B(n7004), .ZN(n6927) );
  NOR2_X1 U8634 ( .A1(n10044), .A2(n7020), .ZN(n6921) );
  AOI21_X1 U8635 ( .B1(n10186), .B2(n7016), .A(n6921), .ZN(n6928) );
  XNOR2_X1 U8636 ( .A(n6927), .B(n6928), .ZN(n9606) );
  INV_X1 U8637 ( .A(n9602), .ZN(n6923) );
  INV_X1 U8638 ( .A(n6922), .ZN(n9715) );
  NAND2_X1 U8639 ( .A1(n6923), .A2(n9715), .ZN(n6924) );
  AND2_X1 U8640 ( .A1(n9606), .A2(n6924), .ZN(n6925) );
  INV_X1 U8641 ( .A(n6927), .ZN(n6929) );
  NAND2_X1 U8642 ( .A1(n10178), .A2(n7015), .ZN(n6932) );
  NAND2_X1 U8643 ( .A1(n10074), .A2(n7016), .ZN(n6931) );
  NAND2_X1 U8644 ( .A1(n6932), .A2(n6931), .ZN(n6933) );
  XNOR2_X1 U8645 ( .A(n6933), .B(n7004), .ZN(n6936) );
  NAND2_X1 U8646 ( .A1(n10178), .A2(n7016), .ZN(n6935) );
  NAND2_X1 U8647 ( .A1(n10074), .A2(n7035), .ZN(n6934) );
  NAND2_X1 U8648 ( .A1(n6935), .A2(n6934), .ZN(n6937) );
  NAND2_X1 U8649 ( .A1(n6936), .A2(n6937), .ZN(n9615) );
  INV_X1 U8650 ( .A(n6936), .ZN(n6939) );
  INV_X1 U8651 ( .A(n6937), .ZN(n6938) );
  NAND2_X1 U8652 ( .A1(n6939), .A2(n6938), .ZN(n9614) );
  NAND2_X1 U8653 ( .A1(n10168), .A2(n7015), .ZN(n6941) );
  NAND2_X1 U8654 ( .A1(n9731), .A2(n7016), .ZN(n6940) );
  NAND2_X1 U8655 ( .A1(n6941), .A2(n6940), .ZN(n6942) );
  XNOR2_X1 U8656 ( .A(n6942), .B(n7004), .ZN(n9555) );
  NAND2_X1 U8657 ( .A1(n10168), .A2(n7016), .ZN(n6944) );
  NAND2_X1 U8658 ( .A1(n9731), .A2(n7035), .ZN(n6943) );
  NAND2_X1 U8659 ( .A1(n6944), .A2(n6943), .ZN(n9554) );
  NAND2_X1 U8660 ( .A1(n10174), .A2(n7016), .ZN(n6946) );
  NAND2_X1 U8661 ( .A1(n10020), .A2(n7035), .ZN(n6945) );
  NAND2_X1 U8662 ( .A1(n6946), .A2(n6945), .ZN(n9693) );
  NAND2_X1 U8663 ( .A1(n10174), .A2(n7015), .ZN(n6948) );
  NAND2_X1 U8664 ( .A1(n10020), .A2(n7016), .ZN(n6947) );
  NAND2_X1 U8665 ( .A1(n6948), .A2(n6947), .ZN(n6949) );
  XNOR2_X1 U8666 ( .A(n6949), .B(n7004), .ZN(n6951) );
  AOI22_X1 U8667 ( .A1(n9555), .A2(n9554), .B1(n9693), .B2(n6951), .ZN(n6950)
         );
  INV_X1 U8668 ( .A(n9555), .ZN(n6957) );
  INV_X1 U8669 ( .A(n9693), .ZN(n6952) );
  NAND2_X1 U8670 ( .A1(n9553), .A2(n6952), .ZN(n6953) );
  NAND2_X1 U8671 ( .A1(n6953), .A2(n9554), .ZN(n6956) );
  INV_X1 U8672 ( .A(n6953), .ZN(n6955) );
  INV_X1 U8673 ( .A(n9554), .ZN(n6954) );
  AOI22_X1 U8674 ( .A1(n6957), .A2(n6956), .B1(n6955), .B2(n6954), .ZN(n6958)
         );
  NAND2_X1 U8675 ( .A1(n10004), .A2(n7015), .ZN(n6961) );
  OR2_X1 U8676 ( .A1(n9982), .A2(n6851), .ZN(n6960) );
  NAND2_X1 U8677 ( .A1(n6961), .A2(n6960), .ZN(n6962) );
  XNOR2_X1 U8678 ( .A(n6962), .B(n6849), .ZN(n9647) );
  NOR2_X1 U8679 ( .A1(n9982), .A2(n7020), .ZN(n6963) );
  AOI21_X1 U8680 ( .B1(n10004), .B2(n7016), .A(n6963), .ZN(n9646) );
  INV_X1 U8681 ( .A(n9647), .ZN(n6965) );
  INV_X1 U8682 ( .A(n9646), .ZN(n6964) );
  NAND2_X1 U8683 ( .A1(n6965), .A2(n6964), .ZN(n6966) );
  NAND2_X1 U8684 ( .A1(n10231), .A2(n7015), .ZN(n6968) );
  NAND2_X1 U8685 ( .A1(n9973), .A2(n7016), .ZN(n6967) );
  NAND2_X1 U8686 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  XNOR2_X1 U8687 ( .A(n6969), .B(n6849), .ZN(n6972) );
  NOR2_X1 U8688 ( .A1(n9996), .A2(n4284), .ZN(n6970) );
  AOI21_X1 U8689 ( .B1(n10231), .B2(n7016), .A(n6970), .ZN(n6971) );
  XNOR2_X1 U8690 ( .A(n6972), .B(n6971), .ZN(n9573) );
  NAND2_X1 U8691 ( .A1(n10139), .A2(n7015), .ZN(n6974) );
  NAND2_X1 U8692 ( .A1(n9950), .A2(n7016), .ZN(n6973) );
  NAND2_X1 U8693 ( .A1(n6974), .A2(n6973), .ZN(n6975) );
  XNOR2_X1 U8694 ( .A(n6975), .B(n6849), .ZN(n6977) );
  NOR2_X1 U8695 ( .A1(n9915), .A2(n7020), .ZN(n6976) );
  AOI21_X1 U8696 ( .B1(n10139), .B2(n7016), .A(n6976), .ZN(n6978) );
  NAND2_X1 U8697 ( .A1(n6977), .A2(n6978), .ZN(n7001) );
  INV_X1 U8698 ( .A(n6977), .ZN(n6980) );
  INV_X1 U8699 ( .A(n6978), .ZN(n6979) );
  NAND2_X1 U8700 ( .A1(n6980), .A2(n6979), .ZN(n6981) );
  NAND2_X1 U8701 ( .A1(n7001), .A2(n6981), .ZN(n9624) );
  NAND2_X1 U8702 ( .A1(n10151), .A2(n7015), .ZN(n6983) );
  OR2_X1 U8703 ( .A1(n9983), .A2(n6851), .ZN(n6982) );
  NAND2_X1 U8704 ( .A1(n6983), .A2(n6982), .ZN(n6984) );
  XNOR2_X1 U8705 ( .A(n6984), .B(n6849), .ZN(n9524) );
  NOR2_X1 U8706 ( .A1(n9983), .A2(n7020), .ZN(n6985) );
  AOI21_X1 U8707 ( .B1(n10151), .B2(n7016), .A(n6985), .ZN(n9669) );
  NAND2_X1 U8708 ( .A1(n10226), .A2(n7015), .ZN(n6987) );
  NAND2_X1 U8709 ( .A1(n9972), .A2(n7016), .ZN(n6986) );
  NAND2_X1 U8710 ( .A1(n6987), .A2(n6986), .ZN(n6988) );
  XNOR2_X1 U8711 ( .A(n6988), .B(n7004), .ZN(n6993) );
  NAND2_X1 U8712 ( .A1(n10226), .A2(n7016), .ZN(n6990) );
  NAND2_X1 U8713 ( .A1(n9972), .A2(n7035), .ZN(n6989) );
  NAND2_X1 U8714 ( .A1(n6990), .A2(n6989), .ZN(n6994) );
  NAND2_X1 U8715 ( .A1(n6993), .A2(n6994), .ZN(n9526) );
  OAI21_X1 U8716 ( .B1(n9524), .B2(n9669), .A(n9526), .ZN(n6991) );
  NOR2_X1 U8717 ( .A1(n9624), .A2(n6991), .ZN(n6992) );
  NAND3_X1 U8718 ( .A1(n9526), .A2(n9524), .A3(n9669), .ZN(n6997) );
  INV_X1 U8719 ( .A(n6993), .ZN(n6996) );
  INV_X1 U8720 ( .A(n6994), .ZN(n6995) );
  NAND2_X1 U8721 ( .A1(n6996), .A2(n6995), .ZN(n9623) );
  AND2_X1 U8722 ( .A1(n6997), .A2(n9623), .ZN(n6998) );
  OR2_X1 U8723 ( .A1(n9624), .A2(n6998), .ZN(n6999) );
  NAND2_X1 U8724 ( .A1(n9921), .A2(n7015), .ZN(n7003) );
  NAND2_X1 U8725 ( .A1(n9932), .A2(n7016), .ZN(n7002) );
  NAND2_X1 U8726 ( .A1(n7003), .A2(n7002), .ZN(n7005) );
  XNOR2_X1 U8727 ( .A(n7005), .B(n7004), .ZN(n7007) );
  NOR2_X1 U8728 ( .A1(n9707), .A2(n7020), .ZN(n7006) );
  AOI21_X1 U8729 ( .B1(n9921), .B2(n7016), .A(n7006), .ZN(n7008) );
  XNOR2_X1 U8730 ( .A(n7007), .B(n7008), .ZN(n9595) );
  INV_X1 U8731 ( .A(n7007), .ZN(n7009) );
  NAND2_X1 U8732 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  NAND2_X1 U8733 ( .A1(n9593), .A2(n7010), .ZN(n9701) );
  NAND2_X1 U8734 ( .A1(n10129), .A2(n7015), .ZN(n7012) );
  NAND2_X1 U8735 ( .A1(n9729), .A2(n7016), .ZN(n7011) );
  NAND2_X1 U8736 ( .A1(n7012), .A2(n7011), .ZN(n7013) );
  XNOR2_X1 U8737 ( .A(n7013), .B(n6849), .ZN(n7026) );
  NOR2_X1 U8738 ( .A1(n9916), .A2(n7020), .ZN(n7014) );
  AOI21_X1 U8739 ( .B1(n10129), .B2(n7016), .A(n7014), .ZN(n7025) );
  XNOR2_X1 U8740 ( .A(n7026), .B(n7025), .ZN(n9700) );
  NAND2_X1 U8741 ( .A1(n10127), .A2(n7015), .ZN(n7018) );
  NAND2_X1 U8742 ( .A1(n9906), .A2(n7016), .ZN(n7017) );
  NAND2_X1 U8743 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  XNOR2_X1 U8744 ( .A(n7019), .B(n6849), .ZN(n7023) );
  NOR2_X1 U8745 ( .A1(n8559), .A2(n4284), .ZN(n7021) );
  AOI21_X1 U8746 ( .B1(n10127), .B2(n7016), .A(n7021), .ZN(n7022) );
  NAND2_X1 U8747 ( .A1(n7023), .A2(n7022), .ZN(n7059) );
  OR2_X1 U8748 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  AND2_X1 U8749 ( .A1(n7059), .A2(n7024), .ZN(n9505) );
  INV_X1 U8750 ( .A(n9505), .ZN(n7028) );
  OR2_X1 U8751 ( .A1(n7026), .A2(n7025), .ZN(n9506) );
  INV_X1 U8752 ( .A(n9506), .ZN(n7027) );
  NOR2_X1 U8753 ( .A1(n7028), .A2(n7027), .ZN(n7029) );
  INV_X1 U8754 ( .A(n7161), .ZN(n7032) );
  NAND2_X1 U8755 ( .A1(n7030), .A2(P1_D_REG_1__SCAN_IN), .ZN(n7031) );
  AOI21_X1 U8756 ( .B1(n7032), .B2(n7031), .A(n7164), .ZN(n7791) );
  AND2_X1 U8757 ( .A1(n7033), .A2(n7791), .ZN(n7048) );
  AND2_X1 U8758 ( .A1(n7048), .A2(n7162), .ZN(n7042) );
  INV_X1 U8759 ( .A(n7156), .ZN(n8660) );
  AND2_X1 U8760 ( .A1(n8660), .A2(n10180), .ZN(n7034) );
  NAND2_X1 U8761 ( .A1(n9507), .A2(n9672), .ZN(n7065) );
  NAND2_X1 U8762 ( .A1(n9890), .A2(n7016), .ZN(n7037) );
  NAND2_X1 U8763 ( .A1(n9728), .A2(n7035), .ZN(n7036) );
  NAND2_X1 U8764 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  XNOR2_X1 U8765 ( .A(n7038), .B(n6849), .ZN(n7040) );
  AOI22_X1 U8766 ( .A1(n9890), .A2(n7015), .B1(n7016), .B2(n9728), .ZN(n7039)
         );
  XNOR2_X1 U8767 ( .A(n7040), .B(n7039), .ZN(n7060) );
  INV_X1 U8768 ( .A(n7042), .ZN(n7044) );
  NOR2_X1 U8769 ( .A1(n10380), .A2(n8665), .ZN(n7797) );
  INV_X1 U8770 ( .A(n7797), .ZN(n7043) );
  OR2_X1 U8771 ( .A1(n7044), .A2(n7043), .ZN(n7046) );
  INV_X1 U8772 ( .A(n7047), .ZN(n10376) );
  NAND2_X1 U8773 ( .A1(n10376), .A2(n7162), .ZN(n8724) );
  INV_X1 U8774 ( .A(n7048), .ZN(n7053) );
  NOR2_X1 U8775 ( .A1(n8724), .A2(n7053), .ZN(n7050) );
  INV_X1 U8776 ( .A(n7049), .ZN(n9727) );
  INV_X1 U8777 ( .A(n7050), .ZN(n7051) );
  NOR2_X2 U8778 ( .A1(n7051), .A2(n7278), .ZN(n9709) );
  INV_X1 U8779 ( .A(n7052), .ZN(n7054) );
  OAI22_X1 U8780 ( .A1(n7054), .A2(n7053), .B1(n7797), .B2(n10180), .ZN(n7056)
         );
  AND2_X1 U8781 ( .A1(n7157), .A2(n7076), .ZN(n7055) );
  NAND2_X1 U8782 ( .A1(n7056), .A2(n7055), .ZN(n7402) );
  OAI22_X1 U8783 ( .A1(n9888), .A2(n9718), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7963), .ZN(n7057) );
  AOI21_X1 U8784 ( .B1(n9727), .B2(n9709), .A(n7057), .ZN(n7058) );
  OAI21_X1 U8785 ( .B1(n8559), .B2(n9717), .A(n7058), .ZN(n7062) );
  NOR3_X1 U8786 ( .A1(n7060), .A2(n9724), .A3(n7059), .ZN(n7061) );
  AOI211_X1 U8787 ( .C1(n9890), .C2(n9722), .A(n7062), .B(n7061), .ZN(n7063)
         );
  OAI211_X1 U8788 ( .C1(n7065), .C2(n7060), .A(n7064), .B(n7063), .ZN(P1_U3220) );
  NAND2_X1 U8789 ( .A1(n7067), .A2(n7066), .ZN(n7068) );
  AOI22_X1 U8790 ( .A1(n9163), .A2(n8906), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7069) );
  OAI21_X1 U8791 ( .B1(n8800), .B2(n8780), .A(n7069), .ZN(n7070) );
  AOI21_X1 U8792 ( .B1(n8778), .B2(n8913), .A(n7070), .ZN(n7071) );
  OAI21_X1 U8793 ( .B1(n9356), .B2(n8909), .A(n7071), .ZN(n7072) );
  OAI21_X1 U8794 ( .B1(n7075), .B2(n7074), .A(n7073), .ZN(P2_U3154) );
  NOR2_X1 U8795 ( .A1(n7076), .A2(P1_U3086), .ZN(n7077) );
  INV_X1 U8796 ( .A(n8446), .ZN(n7078) );
  NAND2_X1 U8797 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  NAND2_X1 U8798 ( .A1(n7123), .A2(n7083), .ZN(n7122) );
  OR2_X1 U8799 ( .A1(n7122), .A2(n4289), .ZN(n7085) );
  NAND2_X1 U8800 ( .A1(n7085), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  MUX2_X1 U8801 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4279), .Z(n7201) );
  XOR2_X1 U8802 ( .A(n7208), .B(n7201), .Z(n7095) );
  XNOR2_X1 U8803 ( .A(n7087), .B(n7322), .ZN(n7312) );
  MUX2_X1 U8804 ( .A(n7629), .B(n7086), .S(n4279), .Z(n7238) );
  NAND2_X1 U8805 ( .A1(n7238), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7311) );
  AOI22_X1 U8806 ( .A1(n7312), .A2(n7311), .B1(n7087), .B2(n5289), .ZN(n7222)
         );
  MUX2_X1 U8807 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4279), .Z(n7088) );
  XNOR2_X1 U8808 ( .A(n7088), .B(n7223), .ZN(n7221) );
  INV_X1 U8809 ( .A(n7223), .ZN(n7090) );
  INV_X1 U8810 ( .A(n7088), .ZN(n7089) );
  OAI22_X1 U8811 ( .A1(n7222), .A2(n7221), .B1(n7090), .B2(n7089), .ZN(n7326)
         );
  MUX2_X1 U8812 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n4279), .Z(n7091) );
  XOR2_X1 U8813 ( .A(n7329), .B(n7091), .Z(n7327) );
  NOR2_X1 U8814 ( .A1(n7326), .A2(n7327), .ZN(n7325) );
  NOR2_X1 U8815 ( .A1(n7091), .A2(n5330), .ZN(n7093) );
  OR2_X1 U8816 ( .A1(n7325), .A2(n7093), .ZN(n7094) );
  NOR3_X1 U8817 ( .A1(n7325), .A2(n7093), .A3(n7095), .ZN(n7200) );
  AOI211_X1 U8818 ( .C1(n7095), .C2(n7094), .A(n9140), .B(n7200), .ZN(n7130)
         );
  OAI21_X1 U8819 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7629), .A(n7322), .ZN(n7097) );
  NAND2_X1 U8820 ( .A1(n7096), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7098) );
  NAND2_X1 U8821 ( .A1(n7097), .A2(n7098), .ZN(n7314) );
  INV_X1 U8822 ( .A(n7098), .ZN(n7099) );
  XNOR2_X1 U8823 ( .A(n7223), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7226) );
  NOR2_X1 U8824 ( .A1(n7225), .A2(n7226), .ZN(n7224) );
  INV_X1 U8825 ( .A(n7101), .ZN(n7102) );
  XNOR2_X1 U8826 ( .A(n7208), .B(n10420), .ZN(n7103) );
  INV_X1 U8827 ( .A(n7202), .ZN(n7105) );
  NAND3_X1 U8828 ( .A1(n7330), .A2(n7103), .A3(n7102), .ZN(n7104) );
  OR2_X1 U8829 ( .A1(n7120), .A2(P2_U3151), .ZN(n9491) );
  OR2_X1 U8830 ( .A1(n7122), .A2(n9491), .ZN(n7117) );
  INV_X1 U8831 ( .A(n7117), .ZN(n7240) );
  AOI21_X1 U8832 ( .B1(n7105), .B2(n7104), .A(n9144), .ZN(n7129) );
  INV_X1 U8833 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U8834 ( .A1(n7106), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U8835 ( .A1(n7322), .A2(n7107), .ZN(n7108) );
  NAND2_X1 U8836 ( .A1(n7096), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8837 ( .A1(n7108), .A2(n7109), .ZN(n7316) );
  OR2_X1 U8838 ( .A1(n7316), .A2(n10442), .ZN(n7318) );
  NAND2_X1 U8839 ( .A1(n7318), .A2(n7109), .ZN(n7228) );
  NAND2_X1 U8840 ( .A1(n7229), .A2(n7228), .ZN(n7227) );
  NAND2_X1 U8841 ( .A1(n7223), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U8842 ( .A1(n7227), .A2(n7110), .ZN(n7111) );
  NAND2_X1 U8843 ( .A1(n7111), .A2(n5330), .ZN(n7114) );
  OR2_X1 U8844 ( .A1(n7111), .A2(n5330), .ZN(n7112) );
  INV_X1 U8845 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7746) );
  XNOR2_X1 U8846 ( .A(n7208), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7113) );
  INV_X1 U8847 ( .A(n7113), .ZN(n7115) );
  NAND3_X1 U8848 ( .A1(n7332), .A2(n7115), .A3(n7114), .ZN(n7118) );
  NOR2_X2 U8849 ( .A1(n7117), .A2(n7116), .ZN(n9126) );
  INV_X1 U8850 ( .A(n9126), .ZN(n9037) );
  AOI21_X1 U8851 ( .B1(n7210), .B2(n7118), .A(n9037), .ZN(n7128) );
  INV_X1 U8852 ( .A(n7123), .ZN(n7119) );
  NOR2_X2 U8853 ( .A1(P2_U3150), .A2(n7119), .ZN(n9142) );
  INV_X1 U8854 ( .A(n9142), .ZN(n9106) );
  INV_X1 U8855 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7978) );
  NOR2_X1 U8856 ( .A1(n4279), .A2(P2_U3151), .ZN(n9494) );
  NAND2_X1 U8857 ( .A1(n9494), .A2(n7120), .ZN(n7121) );
  OR2_X1 U8858 ( .A1(n7122), .A2(n7121), .ZN(n7125) );
  OR2_X1 U8859 ( .A1(n7123), .A2(n9491), .ZN(n7124) );
  AND2_X1 U8860 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7584) );
  AOI21_X1 U8861 ( .B1(n9004), .B2(n7208), .A(n7584), .ZN(n7126) );
  OAI21_X1 U8862 ( .B1(n9106), .B2(n7978), .A(n7126), .ZN(n7127) );
  OR4_X1 U8863 ( .A1(n7130), .A2(n7129), .A3(n7128), .A4(n7127), .ZN(P2_U3186)
         );
  NAND2_X1 U8864 ( .A1(n7131), .A2(P1_U3086), .ZN(n10251) );
  INV_X1 U8865 ( .A(n10251), .ZN(n8439) );
  INV_X1 U8866 ( .A(n7132), .ZN(n7144) );
  INV_X1 U8867 ( .A(n7266), .ZN(n7366) );
  OAI222_X1 U8868 ( .A1(n10259), .A2(n7133), .B1(n10262), .B2(n7144), .C1(
        P1_U3086), .C2(n7366), .ZN(P1_U3353) );
  INV_X1 U8869 ( .A(n10259), .ZN(n8441) );
  AOI22_X1 U8870 ( .A1(n8441), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n9752), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7135) );
  OAI21_X1 U8871 ( .B1(n5026), .B2(n10251), .A(n7135), .ZN(P1_U3354) );
  INV_X1 U8872 ( .A(n7136), .ZN(n7152) );
  AOI22_X1 U8873 ( .A1(n9760), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n8441), .ZN(n7137) );
  OAI21_X1 U8874 ( .B1(n7152), .B2(n10251), .A(n7137), .ZN(P1_U3352) );
  INV_X1 U8875 ( .A(n7138), .ZN(n7142) );
  AOI22_X1 U8876 ( .A1(n10273), .A2(P1_STATE_REG_SCAN_IN), .B1(n8441), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n7139) );
  OAI21_X1 U8877 ( .B1(n7142), .B2(n10251), .A(n7139), .ZN(P1_U3351) );
  INV_X1 U8878 ( .A(n7140), .ZN(n7146) );
  AOI22_X1 U8879 ( .A1(n9773), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n8441), .ZN(n7141) );
  OAI21_X1 U8880 ( .B1(n7146), .B2(n10251), .A(n7141), .ZN(P1_U3350) );
  INV_X1 U8881 ( .A(n9495), .ZN(n9502) );
  NAND2_X2 U8882 ( .A1(n4281), .A2(P2_U3151), .ZN(n9497) );
  INV_X1 U8883 ( .A(n7208), .ZN(n7203) );
  OAI222_X1 U8884 ( .A1(n9502), .A2(n7143), .B1(n9497), .B2(n7142), .C1(
        P2_U3151), .C2(n7203), .ZN(P2_U3291) );
  OAI222_X1 U8885 ( .A1(n9502), .A2(n7145), .B1(n9497), .B2(n7144), .C1(
        P2_U3151), .C2(n7223), .ZN(P2_U3293) );
  INV_X1 U8886 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7147) );
  INV_X1 U8887 ( .A(n7288), .ZN(n7211) );
  OAI222_X1 U8888 ( .A1(n9502), .A2(n7147), .B1(n9497), .B2(n7146), .C1(
        P2_U3151), .C2(n7211), .ZN(P2_U3290) );
  OAI222_X1 U8889 ( .A1(n9502), .A2(n5025), .B1(n5289), .B2(P2_U3151), .C1(
        n9497), .C2(n5026), .ZN(P2_U3294) );
  INV_X1 U8890 ( .A(n7148), .ZN(n7153) );
  AOI22_X1 U8891 ( .A1(n9786), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n8441), .ZN(n7149) );
  OAI21_X1 U8892 ( .B1(n7153), .B2(n10251), .A(n7149), .ZN(P1_U3349) );
  INV_X1 U8893 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n7883) );
  NOR2_X1 U8894 ( .A1(n7176), .A2(n7883), .ZN(P2_U3253) );
  INV_X1 U8895 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n7953) );
  NOR2_X1 U8896 ( .A1(n7176), .A2(n7953), .ZN(P2_U3244) );
  INV_X1 U8897 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n7984) );
  NOR2_X1 U8898 ( .A1(n7176), .A2(n7984), .ZN(P2_U3257) );
  INV_X1 U8899 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n7976) );
  NOR2_X1 U8900 ( .A1(n7176), .A2(n7976), .ZN(P2_U3239) );
  INV_X1 U8901 ( .A(n7150), .ZN(n7159) );
  AOI22_X1 U8902 ( .A1(n9799), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n8441), .ZN(n7151) );
  OAI21_X1 U8903 ( .B1(n7159), .B2(n10251), .A(n7151), .ZN(P1_U3348) );
  OAI222_X1 U8904 ( .A1(n9502), .A2(n4801), .B1(n5330), .B2(P2_U3151), .C1(
        n9497), .C2(n7152), .ZN(P2_U3292) );
  INV_X1 U8905 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7154) );
  OAI222_X1 U8906 ( .A1(n9502), .A2(n7154), .B1(n7527), .B2(P2_U3151), .C1(
        n9497), .C2(n7153), .ZN(P2_U3289) );
  AOI21_X1 U8907 ( .B1(n7157), .B2(n7156), .A(n7155), .ZN(n7186) );
  INV_X1 U8908 ( .A(n7186), .ZN(n7158) );
  OR2_X1 U8909 ( .A1(n8375), .A2(n7162), .ZN(n7187) );
  AND2_X1 U8910 ( .A1(n7158), .A2(n7187), .ZN(n10314) );
  NOR2_X1 U8911 ( .A1(n10314), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8912 ( .A(n7532), .ZN(n7516) );
  OAI222_X1 U8913 ( .A1(n9502), .A2(n7160), .B1(n9497), .B2(n7159), .C1(
        P2_U3151), .C2(n7516), .ZN(P2_U3288) );
  NAND2_X1 U8914 ( .A1(n10390), .A2(P1_D_REG_1__SCAN_IN), .ZN(n7163) );
  OAI21_X1 U8915 ( .B1(n10390), .B2(n7164), .A(n7163), .ZN(P1_U3440) );
  INV_X1 U8916 ( .A(n7165), .ZN(n7167) );
  AOI22_X1 U8917 ( .A1(n9812), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n8441), .ZN(n7166) );
  OAI21_X1 U8918 ( .B1(n7167), .B2(n10251), .A(n7166), .ZN(P1_U3347) );
  AND2_X1 U8919 ( .A1(n8449), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8920 ( .A1(n8449), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8921 ( .A1(n8449), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8922 ( .A1(n8449), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8923 ( .A1(n8449), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8924 ( .A1(n8449), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8925 ( .A1(n8449), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8926 ( .A1(n8449), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8927 ( .A1(n8449), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  INV_X1 U8928 ( .A(n7821), .ZN(n8927) );
  OAI222_X1 U8929 ( .A1(n9502), .A2(n4580), .B1(n9497), .B2(n7167), .C1(
        P2_U3151), .C2(n8927), .ZN(P2_U3287) );
  INV_X1 U8930 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7172) );
  NAND2_X1 U8931 ( .A1(n7168), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7171) );
  INV_X1 U8932 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8424) );
  OR2_X1 U8933 ( .A1(n7169), .A2(n8424), .ZN(n7170) );
  OAI211_X1 U8934 ( .C1(n6647), .C2(n7172), .A(n7171), .B(n7170), .ZN(n8656)
         );
  NAND2_X1 U8935 ( .A1(P1_U3973), .A2(n8656), .ZN(n7173) );
  OAI21_X1 U8936 ( .B1(P1_U3973), .B2(n5975), .A(n7173), .ZN(P1_U3585) );
  INV_X1 U8937 ( .A(n7174), .ZN(n7182) );
  AOI22_X1 U8938 ( .A1(n7345), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n8441), .ZN(n7175) );
  OAI21_X1 U8939 ( .B1(n7182), .B2(n10262), .A(n7175), .ZN(P1_U3346) );
  INV_X1 U8940 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7179) );
  INV_X1 U8941 ( .A(n7177), .ZN(n7178) );
  AOI22_X1 U8942 ( .A1(n8449), .A2(n7179), .B1(n8446), .B2(n7178), .ZN(
        P2_U3376) );
  AND2_X1 U8943 ( .A1(n8449), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8944 ( .A1(n8449), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8945 ( .A1(n8449), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8946 ( .A1(n8449), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8947 ( .A1(n8449), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8948 ( .A1(n8449), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8949 ( .A1(n8449), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8950 ( .A1(n8449), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8951 ( .A1(n8449), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8952 ( .A1(n8449), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8953 ( .A1(n8449), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8954 ( .A1(n8449), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8955 ( .A1(n8449), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8956 ( .A1(n8449), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8957 ( .A1(n8449), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8958 ( .A1(n8449), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8959 ( .A1(n8449), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  INV_X1 U8960 ( .A(n7180), .ZN(n7184) );
  AOI22_X1 U8961 ( .A1(n7418), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n8441), .ZN(n7181) );
  OAI21_X1 U8962 ( .B1(n7184), .B2(n10251), .A(n7181), .ZN(P1_U3345) );
  OAI222_X1 U8963 ( .A1(n9502), .A2(n7183), .B1(n4860), .B2(P2_U3151), .C1(
        n9497), .C2(n7182), .ZN(P2_U3286) );
  INV_X1 U8964 ( .A(n8253), .ZN(n8949) );
  OAI222_X1 U8965 ( .A1(n9502), .A2(n7185), .B1(n8949), .B2(P2_U3151), .C1(
        n9497), .C2(n7184), .ZN(P2_U3285) );
  INV_X1 U8966 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U8967 ( .A1(n7280), .A2(n10249), .ZN(n10297) );
  NAND3_X1 U8968 ( .A1(n10337), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6806), .ZN(
        n7193) );
  AOI21_X1 U8969 ( .B1(n7360), .B2(n7188), .A(n8429), .ZN(n7362) );
  INV_X1 U8970 ( .A(n7362), .ZN(n7190) );
  AOI21_X1 U8971 ( .B1(n6806), .B2(n10249), .A(n7190), .ZN(n7189) );
  MUX2_X1 U8972 ( .A(n7190), .B(n7189), .S(n4433), .Z(n7191) );
  AOI22_X1 U8973 ( .A1(n7280), .A2(n7191), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n7192) );
  OAI211_X1 U8974 ( .C1(n10349), .C2(n7194), .A(n7193), .B(n7192), .ZN(
        P1_U3243) );
  MUX2_X1 U8975 ( .A(n7195), .B(n8812), .S(P2_U3893), .Z(n7196) );
  INV_X1 U8976 ( .A(n7196), .ZN(P2_U3508) );
  INV_X1 U8977 ( .A(n7197), .ZN(n7198) );
  INV_X1 U8978 ( .A(n8331), .ZN(n8241) );
  OAI222_X1 U8979 ( .A1(n9502), .A2(n4602), .B1(n9497), .B2(n7198), .C1(
        P2_U3151), .C2(n8241), .ZN(P2_U3284) );
  INV_X1 U8980 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7199) );
  OAI222_X1 U8981 ( .A1(n10259), .A2(n7199), .B1(n10262), .B2(n7198), .C1(
        P1_U3086), .C2(n7421), .ZN(P1_U3344) );
  AOI21_X1 U8982 ( .B1(n7201), .B2(n7203), .A(n7200), .ZN(n7290) );
  MUX2_X1 U8983 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4279), .Z(n7286) );
  XNOR2_X1 U8984 ( .A(n7286), .B(n7211), .ZN(n7289) );
  XNOR2_X1 U8985 ( .A(n7290), .B(n7289), .ZN(n7218) );
  NOR2_X1 U8986 ( .A1(n7204), .A2(n7288), .ZN(n7296) );
  AOI21_X1 U8987 ( .B1(n7204), .B2(n7288), .A(n7296), .ZN(n7205) );
  OAI21_X1 U8988 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n7205), .A(n7299), .ZN(
        n7207) );
  INV_X1 U8989 ( .A(n9144), .ZN(n8350) );
  NOR2_X1 U8990 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5121), .ZN(n7680) );
  NOR2_X1 U8991 ( .A1(n9131), .A2(n7211), .ZN(n7206) );
  AOI211_X1 U8992 ( .C1(n7207), .C2(n8350), .A(n7680), .B(n7206), .ZN(n7217)
         );
  INV_X1 U8993 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7753) );
  OR2_X1 U8994 ( .A1(n7208), .A2(n7753), .ZN(n7209) );
  INV_X1 U8995 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U8996 ( .A1(n7213), .A2(n7750), .ZN(n7214) );
  NAND2_X1 U8997 ( .A1(n7306), .A2(n7214), .ZN(n7215) );
  AOI22_X1 U8998 ( .A1(n9142), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n9126), .B2(
        n7215), .ZN(n7216) );
  OAI211_X1 U8999 ( .C1(n9140), .C2(n7218), .A(n7217), .B(n7216), .ZN(P2_U3187) );
  INV_X1 U9000 ( .A(n7219), .ZN(n7237) );
  AOI22_X1 U9001 ( .A1(n7567), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n8441), .ZN(n7220) );
  OAI21_X1 U9002 ( .B1(n7237), .B2(n10251), .A(n7220), .ZN(P1_U3343) );
  XNOR2_X1 U9003 ( .A(n7222), .B(n7221), .ZN(n7236) );
  OAI22_X1 U9004 ( .A1(n9131), .A2(n7223), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7386), .ZN(n7234) );
  AOI21_X1 U9005 ( .B1(n7226), .B2(n7225), .A(n7224), .ZN(n7232) );
  OAI21_X1 U9006 ( .B1(n7229), .B2(n7228), .A(n7227), .ZN(n7230) );
  NAND2_X1 U9007 ( .A1(n9126), .A2(n7230), .ZN(n7231) );
  OAI21_X1 U9008 ( .B1(n7232), .B2(n9144), .A(n7231), .ZN(n7233) );
  AOI211_X1 U9009 ( .C1(n9142), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n7234), .B(
        n7233), .ZN(n7235) );
  OAI21_X1 U9010 ( .B1(n9140), .B2(n7236), .A(n7235), .ZN(P2_U3184) );
  INV_X1 U9011 ( .A(n8986), .ZN(n8972) );
  OAI222_X1 U9012 ( .A1(n9502), .A2(n4612), .B1(n8972), .B2(P2_U3151), .C1(
        n9497), .C2(n7237), .ZN(P2_U3283) );
  INV_X1 U9013 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7245) );
  OAI21_X1 U9014 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7238), .A(n7311), .ZN(n7239) );
  OAI21_X1 U9015 ( .B1(n7240), .B2(n9042), .A(n7239), .ZN(n7241) );
  OAI21_X1 U9016 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7242), .A(n7241), .ZN(n7243) );
  AOI21_X1 U9017 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9004), .A(n7243), .ZN(n7244) );
  OAI21_X1 U9018 ( .B1(n9106), .B2(n7245), .A(n7244), .ZN(P2_U3182) );
  XNOR2_X1 U9019 ( .A(n7345), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7262) );
  INV_X1 U9020 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7246) );
  XNOR2_X1 U9021 ( .A(n7266), .B(n7246), .ZN(n7371) );
  INV_X1 U9022 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7247) );
  XNOR2_X1 U9023 ( .A(n9752), .B(n7247), .ZN(n9751) );
  AND2_X1 U9024 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9750) );
  NAND2_X1 U9025 ( .A1(n9751), .A2(n9750), .ZN(n9749) );
  NAND2_X1 U9026 ( .A1(n9752), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U9027 ( .A1(n9749), .A2(n7248), .ZN(n7370) );
  NAND2_X1 U9028 ( .A1(n7371), .A2(n7370), .ZN(n7369) );
  NAND2_X1 U9029 ( .A1(n7266), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7249) );
  NAND2_X1 U9030 ( .A1(n7369), .A2(n7249), .ZN(n9765) );
  INV_X1 U9031 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7250) );
  XNOR2_X1 U9032 ( .A(n9760), .B(n7250), .ZN(n9766) );
  NAND2_X1 U9033 ( .A1(n9765), .A2(n9766), .ZN(n9764) );
  NAND2_X1 U9034 ( .A1(n9760), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7251) );
  NAND2_X1 U9035 ( .A1(n9764), .A2(n7251), .ZN(n10271) );
  MUX2_X1 U9036 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6343), .S(n10273), .Z(n10272) );
  NAND2_X1 U9037 ( .A1(n10271), .A2(n10272), .ZN(n10270) );
  NAND2_X1 U9038 ( .A1(n10273), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U9039 ( .A1(n10270), .A2(n7252), .ZN(n9778) );
  INV_X1 U9040 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7253) );
  XNOR2_X1 U9041 ( .A(n9773), .B(n7253), .ZN(n9779) );
  NAND2_X1 U9042 ( .A1(n9778), .A2(n9779), .ZN(n9777) );
  NAND2_X1 U9043 ( .A1(n9773), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U9044 ( .A1(n9777), .A2(n7254), .ZN(n9788) );
  MUX2_X1 U9045 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6295), .S(n9786), .Z(n9789)
         );
  NAND2_X1 U9046 ( .A1(n9788), .A2(n9789), .ZN(n9787) );
  NAND2_X1 U9047 ( .A1(n9786), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7255) );
  NAND2_X1 U9048 ( .A1(n9787), .A2(n7255), .ZN(n9801) );
  XNOR2_X1 U9049 ( .A(n9799), .B(n7256), .ZN(n9802) );
  NAND2_X1 U9050 ( .A1(n9801), .A2(n9802), .ZN(n9800) );
  NAND2_X1 U9051 ( .A1(n9799), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U9052 ( .A1(n9800), .A2(n7257), .ZN(n9814) );
  INV_X1 U9053 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7258) );
  XNOR2_X1 U9054 ( .A(n9812), .B(n7258), .ZN(n9815) );
  NAND2_X1 U9055 ( .A1(n9814), .A2(n9815), .ZN(n9813) );
  NAND2_X1 U9056 ( .A1(n9812), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7259) );
  NAND2_X1 U9057 ( .A1(n9813), .A2(n7259), .ZN(n7261) );
  INV_X1 U9058 ( .A(n7347), .ZN(n7260) );
  AOI21_X1 U9059 ( .B1(n7262), .B2(n7261), .A(n7260), .ZN(n7285) );
  INV_X1 U9060 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7264) );
  AND2_X1 U9061 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9642) );
  INV_X1 U9062 ( .A(n9642), .ZN(n7263) );
  OAI21_X1 U9063 ( .B1(n10349), .B2(n7264), .A(n7263), .ZN(n7283) );
  XNOR2_X1 U9064 ( .A(n7266), .B(n8015), .ZN(n7368) );
  NAND2_X1 U9065 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7361) );
  INV_X1 U9066 ( .A(n7361), .ZN(n9747) );
  NAND2_X1 U9067 ( .A1(n9748), .A2(n9747), .ZN(n9746) );
  NAND2_X1 U9068 ( .A1(n9752), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7265) );
  NAND2_X1 U9069 ( .A1(n9746), .A2(n7265), .ZN(n7367) );
  NAND2_X1 U9070 ( .A1(n7266), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7267) );
  XNOR2_X1 U9071 ( .A(n9760), .B(n10363), .ZN(n9763) );
  NAND2_X1 U9072 ( .A1(n9762), .A2(n9763), .ZN(n9761) );
  NAND2_X1 U9073 ( .A1(n9760), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7268) );
  NAND2_X1 U9074 ( .A1(n9761), .A2(n7268), .ZN(n10267) );
  MUX2_X1 U9075 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7843), .S(n10273), .Z(n10268) );
  NAND2_X1 U9076 ( .A1(n10267), .A2(n10268), .ZN(n10266) );
  NAND2_X1 U9077 ( .A1(n10273), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U9078 ( .A1(n10266), .A2(n7269), .ZN(n9775) );
  XNOR2_X1 U9079 ( .A(n9773), .B(n10352), .ZN(n9776) );
  NAND2_X1 U9080 ( .A1(n9773), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7270) );
  MUX2_X1 U9081 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n8005), .S(n9786), .Z(n9792)
         );
  NAND2_X1 U9082 ( .A1(n9786), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7271) );
  XNOR2_X1 U9083 ( .A(n9799), .B(n7272), .ZN(n9805) );
  NAND2_X1 U9084 ( .A1(n9804), .A2(n9805), .ZN(n9803) );
  NAND2_X1 U9085 ( .A1(n9799), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7273) );
  XNOR2_X1 U9086 ( .A(n9812), .B(n7274), .ZN(n9818) );
  NAND2_X1 U9087 ( .A1(n9812), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7275) );
  XNOR2_X1 U9088 ( .A(n7345), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7276) );
  NAND2_X1 U9089 ( .A1(n7277), .A2(n7276), .ZN(n7281) );
  NAND2_X1 U9090 ( .A1(n7278), .A2(n7360), .ZN(n8723) );
  INV_X1 U9091 ( .A(n8723), .ZN(n7279) );
  AOI21_X1 U9092 ( .B1(n7341), .B2(n7281), .A(n10334), .ZN(n7282) );
  AOI211_X1 U9093 ( .C1(n10326), .C2(n7345), .A(n7283), .B(n7282), .ZN(n7284)
         );
  OAI21_X1 U9094 ( .B1(n7285), .B2(n10297), .A(n7284), .ZN(P1_U3252) );
  INV_X1 U9095 ( .A(n7286), .ZN(n7287) );
  OAI22_X1 U9096 ( .A1(n7290), .A2(n7289), .B1(n7288), .B2(n7287), .ZN(n7295)
         );
  MUX2_X1 U9097 ( .A(n5396), .B(n7291), .S(n4279), .Z(n7293) );
  NAND2_X1 U9098 ( .A1(n7293), .A2(n7292), .ZN(n7523) );
  OAI21_X1 U9099 ( .B1(n7293), .B2(n7292), .A(n7523), .ZN(n7294) );
  AOI21_X1 U9100 ( .B1(n7295), .B2(n7294), .A(n7521), .ZN(n7310) );
  NAND2_X1 U9101 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7699) );
  OAI21_X1 U9102 ( .B1(n9131), .B2(n7527), .A(n7699), .ZN(n7303) );
  INV_X1 U9103 ( .A(n7296), .ZN(n7297) );
  XNOR2_X1 U9104 ( .A(n7527), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7298) );
  INV_X1 U9105 ( .A(n7526), .ZN(n7301) );
  NAND3_X1 U9106 ( .A1(n7299), .A2(n7298), .A3(n7297), .ZN(n7300) );
  AOI21_X1 U9107 ( .B1(n7301), .B2(n7300), .A(n9144), .ZN(n7302) );
  AOI211_X1 U9108 ( .C1(n9142), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7303), .B(
        n7302), .ZN(n7309) );
  XNOR2_X1 U9109 ( .A(n7527), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7305) );
  AND3_X1 U9110 ( .A1(n7306), .A2(n7305), .A3(n7304), .ZN(n7307) );
  OAI21_X1 U9111 ( .B1(n7511), .B2(n7307), .A(n9126), .ZN(n7308) );
  OAI211_X1 U9112 ( .C1(n7310), .C2(n9140), .A(n7309), .B(n7308), .ZN(P2_U3188) );
  INV_X1 U9113 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10453) );
  XOR2_X1 U9114 ( .A(n7312), .B(n7311), .Z(n7321) );
  AOI21_X1 U9115 ( .B1(n7508), .B2(n7314), .A(n7313), .ZN(n7315) );
  NOR2_X1 U9116 ( .A1(n9144), .A2(n7315), .ZN(n7320) );
  NAND2_X1 U9117 ( .A1(n7316), .A2(n10442), .ZN(n7317) );
  AOI21_X1 U9118 ( .B1(n7318), .B2(n7317), .A(n9037), .ZN(n7319) );
  AOI211_X1 U9119 ( .C1(n7321), .C2(n9042), .A(n7320), .B(n7319), .ZN(n7324)
         );
  AOI22_X1 U9120 ( .A1(n9004), .A2(n7322), .B1(P2_U3151), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7323) );
  OAI211_X1 U9121 ( .C1(n10453), .C2(n9106), .A(n7324), .B(n7323), .ZN(
        P2_U3183) );
  AOI21_X1 U9122 ( .B1(n7327), .B2(n7326), .A(n7325), .ZN(n7337) );
  NOR2_X1 U9123 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7549), .ZN(n7540) );
  INV_X1 U9124 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7983) );
  NOR2_X1 U9125 ( .A1(n9106), .A2(n7983), .ZN(n7328) );
  AOI211_X1 U9126 ( .C1(n7329), .C2(n9004), .A(n7540), .B(n7328), .ZN(n7336)
         );
  OAI21_X1 U9127 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7331), .A(n7330), .ZN(
        n7334) );
  OAI21_X1 U9128 ( .B1(n4421), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7332), .ZN(
        n7333) );
  AOI22_X1 U9129 ( .A1(n8350), .A2(n7334), .B1(n9126), .B2(n7333), .ZN(n7335)
         );
  OAI211_X1 U9130 ( .C1(n7337), .C2(n9140), .A(n7336), .B(n7335), .ZN(P2_U3185) );
  INV_X1 U9131 ( .A(n7338), .ZN(n7397) );
  AOI22_X1 U9132 ( .A1(n9848), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n8441), .ZN(n7339) );
  OAI21_X1 U9133 ( .B1(n7397), .B2(n10251), .A(n7339), .ZN(P1_U3342) );
  XNOR2_X1 U9134 ( .A(n7418), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7344) );
  OR2_X1 U9135 ( .A1(n7345), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U9136 ( .A1(n7341), .A2(n7340), .ZN(n7343) );
  INV_X1 U9137 ( .A(n7420), .ZN(n7342) );
  AOI211_X1 U9138 ( .C1(n7344), .C2(n7343), .A(n10334), .B(n7342), .ZN(n7356)
         );
  XNOR2_X1 U9139 ( .A(n7418), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7350) );
  OR2_X1 U9140 ( .A1(n7345), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U9141 ( .A1(n7347), .A2(n7346), .ZN(n7349) );
  INV_X1 U9142 ( .A(n7412), .ZN(n7348) );
  AOI211_X1 U9143 ( .C1(n7350), .C2(n7349), .A(n10297), .B(n7348), .ZN(n7355)
         );
  INV_X1 U9144 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7353) );
  NAND2_X1 U9145 ( .A1(n10326), .A2(n7418), .ZN(n7352) );
  AND2_X1 U9146 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9548) );
  INV_X1 U9147 ( .A(n9548), .ZN(n7351) );
  OAI211_X1 U9148 ( .C1(n10349), .C2(n7353), .A(n7352), .B(n7351), .ZN(n7354)
         );
  OR3_X1 U9149 ( .A1(n7356), .A2(n7355), .A3(n7354), .ZN(P1_U3253) );
  OAI21_X1 U9150 ( .B1(n7359), .B2(n7358), .A(n7357), .ZN(n7405) );
  NOR2_X1 U9151 ( .A1(n8429), .A2(n7360), .ZN(n7364) );
  INV_X1 U9152 ( .A(P1_U3973), .ZN(n9744) );
  OAI22_X1 U9153 ( .A1(n7362), .A2(P1_IR_REG_0__SCAN_IN), .B1(n7361), .B2(
        n8723), .ZN(n7363) );
  AOI211_X1 U9154 ( .C1(n7405), .C2(n7364), .A(n9744), .B(n7363), .ZN(n10278)
         );
  INV_X1 U9155 ( .A(n10326), .ZN(n10343) );
  AOI22_X1 U9156 ( .A1(n10314), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7365) );
  OAI21_X1 U9157 ( .B1(n10343), .B2(n7366), .A(n7365), .ZN(n7375) );
  OAI21_X1 U9158 ( .B1(n7371), .B2(n7370), .A(n7369), .ZN(n7372) );
  OAI22_X1 U9159 ( .A1(n10334), .A2(n7373), .B1(n10297), .B2(n7372), .ZN(n7374) );
  OR3_X1 U9160 ( .A1(n10278), .A2(n7375), .A3(n7374), .ZN(P1_U3245) );
  NAND2_X1 U9161 ( .A1(n10436), .A2(n9293), .ZN(n7376) );
  NOR2_X1 U9162 ( .A1(n5292), .A2(n9298), .ZN(n7627) );
  AOI21_X1 U9163 ( .B1(n7470), .B2(n7376), .A(n7627), .ZN(n7755) );
  MUX2_X1 U9164 ( .A(n7755), .B(n5294), .S(n10441), .Z(n7377) );
  OAI21_X1 U9165 ( .B1(n7757), .B2(n9461), .A(n7377), .ZN(P2_U3390) );
  NAND2_X1 U9166 ( .A1(n8852), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7471) );
  INV_X1 U9167 ( .A(n7471), .ZN(n7396) );
  INV_X1 U9168 ( .A(n5334), .ZN(n7587) );
  OAI22_X1 U9169 ( .A1(n8780), .A2(n5292), .B1(n7587), .B2(n8904), .ZN(n7378)
         );
  AOI21_X1 U9170 ( .B1(n7379), .B2(n8896), .A(n7378), .ZN(n7385) );
  OAI21_X1 U9171 ( .B1(n7382), .B2(n7381), .A(n7380), .ZN(n7383) );
  NAND2_X1 U9172 ( .A1(n7383), .A2(n8882), .ZN(n7384) );
  OAI211_X1 U9173 ( .C1(n7396), .C2(n7386), .A(n7385), .B(n7384), .ZN(P2_U3177) );
  INV_X1 U9174 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7395) );
  INV_X1 U9175 ( .A(n5786), .ZN(n7387) );
  OAI22_X1 U9176 ( .A1(n8780), .A2(n7387), .B1(n5314), .B2(n8904), .ZN(n7388)
         );
  AOI21_X1 U9177 ( .B1(n5291), .B2(n8896), .A(n7388), .ZN(n7394) );
  OAI21_X1 U9178 ( .B1(n7391), .B2(n7390), .A(n7389), .ZN(n7392) );
  NAND2_X1 U9179 ( .A1(n7392), .A2(n8882), .ZN(n7393) );
  OAI211_X1 U9180 ( .C1(n7396), .C2(n7395), .A(n7394), .B(n7393), .ZN(P2_U3162) );
  INV_X1 U9181 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7398) );
  OAI222_X1 U9182 ( .A1(n9502), .A2(n7398), .B1(n8999), .B2(P2_U3151), .C1(
        n9497), .C2(n7397), .ZN(P2_U3282) );
  INV_X1 U9183 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7399) );
  OAI222_X1 U9184 ( .A1(n10259), .A2(n7399), .B1(n10262), .B2(n7400), .C1(
        n10292), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U9185 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7401) );
  INV_X1 U9186 ( .A(n9031), .ZN(n9027) );
  OAI222_X1 U9187 ( .A1(n9502), .A2(n7401), .B1(n9027), .B2(P2_U3151), .C1(
        n9497), .C2(n7400), .ZN(P2_U3281) );
  OR2_X1 U9188 ( .A1(n7402), .A2(P1_U3086), .ZN(n9568) );
  OAI22_X1 U9189 ( .A1(n9719), .A2(n7489), .B1(n9712), .B2(n10381), .ZN(n7403)
         );
  AOI21_X1 U9190 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9568), .A(n7403), .ZN(
        n7404) );
  OAI21_X1 U9191 ( .B1(n9724), .B2(n7405), .A(n7404), .ZN(P1_U3232) );
  XOR2_X1 U9192 ( .A(n7407), .B(n7406), .Z(n7410) );
  AOI22_X1 U9193 ( .A1(n9722), .A2(n7500), .B1(n9709), .B2(n9742), .ZN(n7409)
         );
  AOI22_X1 U9194 ( .A1(n9695), .A2(n6319), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9568), .ZN(n7408) );
  OAI211_X1 U9195 ( .C1(n7410), .C2(n9724), .A(n7409), .B(n7408), .ZN(P1_U3237) );
  XNOR2_X1 U9196 ( .A(n7567), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7416) );
  NAND2_X1 U9197 ( .A1(n7418), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U9198 ( .A1(n7412), .A2(n7411), .ZN(n9827) );
  XNOR2_X1 U9199 ( .A(n7421), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U9200 ( .A1(n9827), .A2(n9826), .ZN(n9825) );
  NAND2_X1 U9201 ( .A1(n9831), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U9202 ( .A1(n9825), .A2(n7413), .ZN(n7415) );
  INV_X1 U9203 ( .A(n7569), .ZN(n7414) );
  AOI21_X1 U9204 ( .B1(n7416), .B2(n7415), .A(n7414), .ZN(n7429) );
  INV_X1 U9205 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7417) );
  NAND2_X1 U9206 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9581) );
  OAI21_X1 U9207 ( .B1(n10349), .B2(n7417), .A(n9581), .ZN(n7427) );
  NAND2_X1 U9208 ( .A1(n7418), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7419) );
  XNOR2_X1 U9209 ( .A(n7421), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U9210 ( .A1(n9831), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7422) );
  XNOR2_X1 U9211 ( .A(n7567), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9212 ( .A1(n7424), .A2(n7423), .ZN(n7425) );
  AOI21_X1 U9213 ( .B1(n7563), .B2(n7425), .A(n10334), .ZN(n7426) );
  AOI211_X1 U9214 ( .C1(n10326), .C2(n7567), .A(n7427), .B(n7426), .ZN(n7428)
         );
  OAI21_X1 U9215 ( .B1(n7429), .B2(n10297), .A(n7428), .ZN(P1_U3255) );
  OAI21_X1 U9216 ( .B1(n7430), .B2(n7433), .A(n7445), .ZN(n7435) );
  INV_X1 U9217 ( .A(n7435), .ZN(n10429) );
  NAND2_X1 U9218 ( .A1(n7432), .A2(n7431), .ZN(n7434) );
  XNOR2_X1 U9219 ( .A(n7434), .B(n7433), .ZN(n7438) );
  NAND2_X1 U9220 ( .A1(n7435), .A2(n6742), .ZN(n7437) );
  AOI22_X1 U9221 ( .A1(n9331), .A2(n8925), .B1(n5334), .B2(n9333), .ZN(n7436)
         );
  OAI211_X1 U9222 ( .C1(n9293), .C2(n7438), .A(n7437), .B(n7436), .ZN(n10430)
         );
  OAI22_X1 U9223 ( .A1(n10417), .A2(n7386), .B1(n10427), .B2(n9337), .ZN(n7439) );
  NOR2_X1 U9224 ( .A1(n10430), .A2(n7439), .ZN(n7440) );
  MUX2_X1 U9225 ( .A(n7441), .B(n7440), .S(n10421), .Z(n7442) );
  OAI21_X1 U9226 ( .B1(n10429), .B2(n9159), .A(n7442), .ZN(P2_U3231) );
  NAND3_X1 U9227 ( .A1(n7445), .A2(n7444), .A3(n7443), .ZN(n7447) );
  NAND2_X1 U9228 ( .A1(n7447), .A2(n7446), .ZN(n7592) );
  XNOR2_X1 U9229 ( .A(n7449), .B(n7448), .ZN(n7450) );
  OAI222_X1 U9230 ( .A1(n9298), .A2(n7683), .B1(n9296), .B2(n5314), .C1(n9293), 
        .C2(n7450), .ZN(n7593) );
  AOI21_X1 U9231 ( .B1(n10426), .B2(n7592), .A(n7593), .ZN(n7745) );
  OAI22_X1 U9232 ( .A1(n7748), .A2(n9461), .B1(n10440), .B2(n5316), .ZN(n7451)
         );
  INV_X1 U9233 ( .A(n7451), .ZN(n7452) );
  OAI21_X1 U9234 ( .B1(n7745), .B2(n10441), .A(n7452), .ZN(P2_U3399) );
  XOR2_X1 U9235 ( .A(n7454), .B(n7453), .Z(n7460) );
  INV_X1 U9236 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7458) );
  NAND2_X1 U9237 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9757) );
  OAI21_X1 U9238 ( .B1(n9712), .B2(n7605), .A(n9757), .ZN(n7457) );
  OAI22_X1 U9239 ( .A1(n9719), .A2(n7455), .B1(n7478), .B2(n9717), .ZN(n7456)
         );
  AOI211_X1 U9240 ( .C1(n9705), .C2(n7458), .A(n7457), .B(n7456), .ZN(n7459)
         );
  OAI21_X1 U9241 ( .B1(n7460), .B2(n9724), .A(n7459), .ZN(P1_U3218) );
  OAI21_X1 U9242 ( .B1(n7462), .B2(n7465), .A(n7461), .ZN(n10410) );
  NAND2_X1 U9243 ( .A1(n7464), .A2(n7463), .ZN(n7466) );
  XNOR2_X1 U9244 ( .A(n7465), .B(n7466), .ZN(n7467) );
  OAI222_X1 U9245 ( .A1(n9298), .A2(n4514), .B1(n9296), .B2(n7587), .C1(n9293), 
        .C2(n7467), .ZN(n10409) );
  AOI21_X1 U9246 ( .B1(n10426), .B2(n10410), .A(n10409), .ZN(n7752) );
  OAI22_X1 U9247 ( .A1(n10414), .A2(n9461), .B1(n10440), .B2(n5337), .ZN(n7468) );
  INV_X1 U9248 ( .A(n7468), .ZN(n7469) );
  OAI21_X1 U9249 ( .B1(n7752), .B2(n10441), .A(n7469), .ZN(P2_U3402) );
  INV_X1 U9250 ( .A(n7470), .ZN(n7623) );
  NAND2_X1 U9251 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n7471), .ZN(n7472) );
  OAI21_X1 U9252 ( .B1(n8904), .B2(n5292), .A(n7472), .ZN(n7473) );
  AOI21_X1 U9253 ( .B1(n7474), .B2(n8896), .A(n7473), .ZN(n7475) );
  OAI21_X1 U9254 ( .B1(n8898), .B2(n7623), .A(n7475), .ZN(P2_U3172) );
  XNOR2_X1 U9255 ( .A(n8604), .B(n7476), .ZN(n7805) );
  OAI21_X1 U9256 ( .B1(n8598), .B2(n8604), .A(n7477), .ZN(n7482) );
  INV_X1 U9257 ( .A(n9745), .ZN(n7479) );
  OAI22_X1 U9258 ( .A1(n7479), .A2(n10043), .B1(n7478), .B2(n10045), .ZN(n7481) );
  NOR2_X1 U9259 ( .A1(n7805), .A2(n8052), .ZN(n7480) );
  AOI211_X1 U9260 ( .C1(n10087), .C2(n7482), .A(n7481), .B(n7480), .ZN(n7796)
         );
  INV_X1 U9261 ( .A(n7483), .ZN(n7488) );
  OAI211_X1 U9262 ( .C1(n4437), .C2(n10381), .A(n7488), .B(n10052), .ZN(n7800)
         );
  OAI211_X1 U9263 ( .C1(n7805), .C2(n10212), .A(n7796), .B(n7800), .ZN(n7492)
         );
  NAND2_X1 U9264 ( .A1(n7492), .A2(n10408), .ZN(n7485) );
  NAND2_X1 U9265 ( .A1(n10159), .A2(n9567), .ZN(n7484) );
  OAI211_X1 U9266 ( .C1(n10408), .C2(n7247), .A(n7485), .B(n7484), .ZN(
        P1_U3523) );
  OAI21_X1 U9267 ( .B1(n7487), .B2(n8599), .A(n7486), .ZN(n8020) );
  AOI211_X1 U9268 ( .C1(n7500), .C2(n7488), .A(n10091), .B(n4418), .ZN(n8019)
         );
  XNOR2_X1 U9269 ( .A(n8468), .B(n8599), .ZN(n7490) );
  INV_X1 U9270 ( .A(n9742), .ZN(n7661) );
  OAI222_X1 U9271 ( .A1(n7490), .A2(n10392), .B1(n10045), .B2(n7661), .C1(
        n10043), .C2(n7489), .ZN(n8013) );
  AOI211_X1 U9272 ( .C1(n10195), .C2(n8020), .A(n8019), .B(n8013), .ZN(n7502)
         );
  AOI22_X1 U9273 ( .A1(n10159), .A2(n7500), .B1(n6794), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n7491) );
  OAI21_X1 U9274 ( .B1(n7502), .B2(n6794), .A(n7491), .ZN(P1_U3524) );
  INV_X1 U9275 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9276 ( .A1(n7492), .A2(n10405), .ZN(n7494) );
  NAND2_X1 U9277 ( .A1(n10232), .A2(n9567), .ZN(n7493) );
  OAI211_X1 U9278 ( .C1(n10405), .C2(n7495), .A(n7494), .B(n7493), .ZN(
        P1_U3456) );
  INV_X1 U9279 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7497) );
  INV_X1 U9280 ( .A(n7496), .ZN(n7498) );
  OAI222_X1 U9281 ( .A1(n9502), .A2(n7497), .B1(n9497), .B2(n7498), .C1(
        P2_U3151), .C2(n9034), .ZN(P2_U3280) );
  INV_X1 U9282 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7499) );
  OAI222_X1 U9283 ( .A1(n10259), .A2(n7499), .B1(n10262), .B2(n7498), .C1(
        P1_U3086), .C2(n9853), .ZN(P1_U3340) );
  AOI22_X1 U9284 ( .A1(n10232), .A2(n7500), .B1(n10403), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n7501) );
  OAI21_X1 U9285 ( .B1(n7502), .B2(n10403), .A(n7501), .ZN(P1_U3459) );
  XNOR2_X1 U9286 ( .A(n5847), .B(n5293), .ZN(n10425) );
  AOI22_X1 U9287 ( .A1(n9283), .A2(n10425), .B1(n9325), .B2(n5291), .ZN(n7510)
         );
  XNOR2_X1 U9288 ( .A(n5293), .B(n7503), .ZN(n7504) );
  NAND2_X1 U9289 ( .A1(n7504), .A2(n9336), .ZN(n7506) );
  AOI22_X1 U9290 ( .A1(n9331), .A2(n5786), .B1(n8924), .B2(n9333), .ZN(n7505)
         );
  NAND2_X1 U9291 ( .A1(n7506), .A2(n7505), .ZN(n10423) );
  AOI21_X1 U9292 ( .B1(n9341), .B2(P2_REG3_REG_1__SCAN_IN), .A(n10423), .ZN(
        n7507) );
  MUX2_X1 U9293 ( .A(n7508), .B(n7507), .S(n10421), .Z(n7509) );
  NAND2_X1 U9294 ( .A1(n7510), .A2(n7509), .ZN(P2_U3232) );
  OAI21_X1 U9295 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7514), .A(n8942), .ZN(
        n7538) );
  INV_X1 U9296 ( .A(n7523), .ZN(n7520) );
  MUX2_X1 U9297 ( .A(n7530), .B(n7939), .S(n4279), .Z(n7515) );
  NAND2_X1 U9298 ( .A1(n7515), .A2(n7532), .ZN(n8936) );
  INV_X1 U9299 ( .A(n7515), .ZN(n7517) );
  NAND2_X1 U9300 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  NAND2_X1 U9301 ( .A1(n8936), .A2(n7518), .ZN(n7522) );
  INV_X1 U9302 ( .A(n7522), .ZN(n7519) );
  INV_X1 U9303 ( .A(n7521), .ZN(n7524) );
  NAND3_X1 U9304 ( .A1(n7524), .A2(n7523), .A3(n7522), .ZN(n7525) );
  AOI21_X1 U9305 ( .B1(n8937), .B2(n7525), .A(n9140), .ZN(n7537) );
  INV_X1 U9306 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7535) );
  NOR2_X1 U9307 ( .A1(n4419), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7531) );
  OAI21_X1 U9308 ( .B1(n7531), .B2(n8930), .A(n8350), .ZN(n7534) );
  AND2_X1 U9309 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8034) );
  AOI21_X1 U9310 ( .B1(n9004), .B2(n7532), .A(n8034), .ZN(n7533) );
  OAI211_X1 U9311 ( .C1(n7535), .C2(n9106), .A(n7534), .B(n7533), .ZN(n7536)
         );
  AOI211_X1 U9312 ( .C1(n9126), .C2(n7538), .A(n7537), .B(n7536), .ZN(n7539)
         );
  INV_X1 U9313 ( .A(n7539), .ZN(P2_U3189) );
  NAND2_X1 U9314 ( .A1(n8896), .A2(n7596), .ZN(n7542) );
  AOI21_X1 U9315 ( .B1(n8778), .B2(n8923), .A(n7540), .ZN(n7541) );
  OAI211_X1 U9316 ( .C1(n5314), .C2(n8780), .A(n7542), .B(n7541), .ZN(n7548)
         );
  INV_X1 U9317 ( .A(n7543), .ZN(n7544) );
  AOI211_X1 U9318 ( .C1(n7546), .C2(n7545), .A(n8898), .B(n7544), .ZN(n7547)
         );
  AOI211_X1 U9319 ( .C1(n7549), .C2(n8906), .A(n7548), .B(n7547), .ZN(n7550)
         );
  INV_X1 U9320 ( .A(n7550), .ZN(P2_U3158) );
  XOR2_X1 U9321 ( .A(n7633), .B(n7554), .Z(n7856) );
  AND2_X1 U9322 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  XOR2_X1 U9323 ( .A(n7554), .B(n7553), .Z(n7555) );
  OAI222_X1 U9324 ( .A1(n9298), .A2(n8037), .B1(n9296), .B2(n7683), .C1(n9293), 
        .C2(n7555), .ZN(n7853) );
  AOI21_X1 U9325 ( .B1(n7856), .B2(n10426), .A(n7853), .ZN(n7749) );
  OAI22_X1 U9326 ( .A1(n7852), .A2(n9461), .B1(n10440), .B2(n5355), .ZN(n7556)
         );
  INV_X1 U9327 ( .A(n7556), .ZN(n7557) );
  OAI21_X1 U9328 ( .B1(n7749), .B2(n10441), .A(n7557), .ZN(P2_U3405) );
  INV_X1 U9329 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7559) );
  INV_X1 U9330 ( .A(n7558), .ZN(n7560) );
  INV_X1 U9331 ( .A(n10318), .ZN(n9846) );
  OAI222_X1 U9332 ( .A1(n10259), .A2(n7559), .B1(n10262), .B2(n7560), .C1(
        P1_U3086), .C2(n9846), .ZN(P1_U3339) );
  INV_X1 U9333 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7561) );
  INV_X1 U9334 ( .A(n9074), .ZN(n9077) );
  OAI222_X1 U9335 ( .A1(n9502), .A2(n7561), .B1(n9497), .B2(n7560), .C1(
        P2_U3151), .C2(n9077), .ZN(P2_U3279) );
  XNOR2_X1 U9336 ( .A(n9848), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7566) );
  OR2_X1 U9337 ( .A1(n7567), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7562) );
  INV_X1 U9338 ( .A(n9836), .ZN(n7564) );
  AOI211_X1 U9339 ( .C1(n7566), .C2(n7565), .A(n10334), .B(n7564), .ZN(n7578)
         );
  XNOR2_X1 U9340 ( .A(n9848), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7572) );
  OR2_X1 U9341 ( .A1(n7567), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U9342 ( .A1(n7569), .A2(n7568), .ZN(n7571) );
  INV_X1 U9343 ( .A(n9850), .ZN(n7570) );
  AOI211_X1 U9344 ( .C1(n7572), .C2(n7571), .A(n10297), .B(n7570), .ZN(n7577)
         );
  INV_X1 U9345 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U9346 ( .A1(n10326), .A2(n9848), .ZN(n7574) );
  AND2_X1 U9347 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9663) );
  INV_X1 U9348 ( .A(n9663), .ZN(n7573) );
  OAI211_X1 U9349 ( .C1(n10349), .C2(n7575), .A(n7574), .B(n7573), .ZN(n7576)
         );
  OR3_X1 U9350 ( .A1(n7578), .A2(n7577), .A3(n7576), .ZN(P1_U3256) );
  INV_X1 U9351 ( .A(n7579), .ZN(n7580) );
  AOI21_X1 U9352 ( .B1(n7582), .B2(n7581), .A(n7580), .ZN(n7591) );
  INV_X1 U9353 ( .A(n10416), .ZN(n7589) );
  NAND2_X1 U9354 ( .A1(n8896), .A2(n7583), .ZN(n7586) );
  AOI21_X1 U9355 ( .B1(n8778), .B2(n8922), .A(n7584), .ZN(n7585) );
  OAI211_X1 U9356 ( .C1(n7587), .C2(n8780), .A(n7586), .B(n7585), .ZN(n7588)
         );
  AOI21_X1 U9357 ( .B1(n7589), .B2(n8906), .A(n7588), .ZN(n7590) );
  OAI21_X1 U9358 ( .B1(n7591), .B2(n8898), .A(n7590), .ZN(P2_U3170) );
  INV_X1 U9359 ( .A(n7592), .ZN(n7599) );
  INV_X1 U9360 ( .A(n7593), .ZN(n7594) );
  MUX2_X1 U9361 ( .A(n7595), .B(n7594), .S(n10421), .Z(n7598) );
  AOI22_X1 U9362 ( .A1(n9325), .A2(n7596), .B1(n7549), .B2(n9341), .ZN(n7597)
         );
  OAI211_X1 U9363 ( .C1(n7599), .C2(n9344), .A(n7598), .B(n7597), .ZN(P2_U3230) );
  INV_X1 U9364 ( .A(n7600), .ZN(n8601) );
  INV_X1 U9365 ( .A(n7601), .ZN(n7602) );
  NOR2_X1 U9366 ( .A1(n7602), .A2(n8601), .ZN(n7716) );
  AOI21_X1 U9367 ( .B1(n8601), .B2(n7602), .A(n7716), .ZN(n10362) );
  XNOR2_X1 U9368 ( .A(n7603), .B(n8601), .ZN(n7604) );
  AOI222_X1 U9369 ( .A1(n9743), .A2(n10085), .B1(n10087), .B2(n7604), .C1(
        n9741), .C2(n10377), .ZN(n10374) );
  OAI211_X1 U9370 ( .C1(n4418), .C2(n7605), .A(n10052), .B(n7718), .ZN(n10368)
         );
  OAI211_X1 U9371 ( .C1(n10401), .C2(n10362), .A(n10374), .B(n10368), .ZN(
        n7608) );
  NAND2_X1 U9372 ( .A1(n7608), .A2(n10408), .ZN(n7607) );
  NAND2_X1 U9373 ( .A1(n10159), .A2(n4278), .ZN(n7606) );
  OAI211_X1 U9374 ( .C1(n10408), .C2(n7250), .A(n7607), .B(n7606), .ZN(
        P1_U3525) );
  NAND2_X1 U9375 ( .A1(n7608), .A2(n10405), .ZN(n7610) );
  NAND2_X1 U9376 ( .A1(n10232), .A2(n4278), .ZN(n7609) );
  OAI211_X1 U9377 ( .C1(n10405), .C2(n6331), .A(n7610), .B(n7609), .ZN(
        P1_U3462) );
  XOR2_X1 U9378 ( .A(n7611), .B(n7614), .Z(n7612) );
  AOI222_X1 U9379 ( .A1(n9336), .A2(n7612), .B1(n8918), .B2(n9333), .C1(n8920), 
        .C2(n9331), .ZN(n8105) );
  NAND2_X1 U9380 ( .A1(n7645), .A2(n7613), .ZN(n7615) );
  XNOR2_X1 U9381 ( .A(n7615), .B(n7614), .ZN(n8109) );
  INV_X1 U9382 ( .A(n8109), .ZN(n7619) );
  OAI22_X1 U9383 ( .A1(n7617), .A2(n9461), .B1(n10440), .B2(n7616), .ZN(n7618)
         );
  AOI21_X1 U9384 ( .B1(n7619), .B2(n9486), .A(n7618), .ZN(n7620) );
  OAI21_X1 U9385 ( .B1(n8105), .B2(n10441), .A(n7620), .ZN(P2_U3414) );
  INV_X1 U9386 ( .A(n7621), .ZN(n7666) );
  AOI22_X1 U9387 ( .A1(n10327), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n8441), .ZN(n7622) );
  OAI21_X1 U9388 ( .B1(n7666), .B2(n10262), .A(n7622), .ZN(P1_U3338) );
  NOR4_X1 U9389 ( .A1(n7625), .A2(n9394), .A3(n7624), .A4(n7623), .ZN(n7626)
         );
  AOI21_X1 U9390 ( .B1(n9341), .B2(P2_REG3_REG_0__SCAN_IN), .A(n7626), .ZN(
        n7631) );
  INV_X1 U9391 ( .A(n7627), .ZN(n7628) );
  MUX2_X1 U9392 ( .A(n7629), .B(n7628), .S(n10421), .Z(n7630) );
  OAI211_X1 U9393 ( .C1(n10415), .C2(n7757), .A(n7631), .B(n7630), .ZN(
        P2_U3233) );
  NAND2_X1 U9394 ( .A1(n7633), .A2(n7632), .ZN(n7635) );
  NAND2_X1 U9395 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  XNOR2_X1 U9396 ( .A(n7636), .B(n7638), .ZN(n10437) );
  XNOR2_X1 U9397 ( .A(n7637), .B(n7638), .ZN(n7639) );
  AOI222_X1 U9398 ( .A1(n9336), .A2(n7639), .B1(n8920), .B2(n9333), .C1(n8922), 
        .C2(n9331), .ZN(n10433) );
  MUX2_X1 U9399 ( .A(n5396), .B(n10433), .S(n10421), .Z(n7642) );
  INV_X1 U9400 ( .A(n7706), .ZN(n7640) );
  AOI22_X1 U9401 ( .A1(n9325), .A2(n7698), .B1(n9341), .B2(n7640), .ZN(n7641)
         );
  OAI211_X1 U9402 ( .C1(n10437), .C2(n9344), .A(n7642), .B(n7641), .ZN(
        P2_U3227) );
  OR2_X1 U9403 ( .A1(n7643), .A2(n7648), .ZN(n7644) );
  NAND2_X1 U9404 ( .A1(n7645), .A2(n7644), .ZN(n7789) );
  INV_X1 U9405 ( .A(n7789), .ZN(n7654) );
  INV_X1 U9406 ( .A(n7637), .ZN(n7646) );
  OAI21_X1 U9407 ( .B1(n7646), .B2(n8921), .A(n7698), .ZN(n7647) );
  OAI21_X1 U9408 ( .B1(n8037), .B2(n7637), .A(n7647), .ZN(n7649) );
  XNOR2_X1 U9409 ( .A(n7649), .B(n7648), .ZN(n7650) );
  NAND2_X1 U9410 ( .A1(n7650), .A2(n9336), .ZN(n7652) );
  AOI22_X1 U9411 ( .A1(n9331), .A2(n8921), .B1(n8919), .B2(n9333), .ZN(n7651)
         );
  OAI211_X1 U9412 ( .C1(n7789), .C2(n7653), .A(n7652), .B(n7651), .ZN(n7784)
         );
  AOI21_X1 U9413 ( .B1(n7767), .B2(n7654), .A(n7784), .ZN(n7806) );
  AOI22_X1 U9414 ( .A1(n9485), .A2(n8033), .B1(P2_REG0_REG_7__SCAN_IN), .B2(
        n10441), .ZN(n7655) );
  OAI21_X1 U9415 ( .B1(n7806), .B2(n10441), .A(n7655), .ZN(P2_U3411) );
  AOI22_X1 U9416 ( .A1(n9133), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9495), .ZN(n7656) );
  OAI21_X1 U9417 ( .B1(n7668), .B2(n9497), .A(n7656), .ZN(P2_U3277) );
  INV_X1 U9418 ( .A(n7657), .ZN(n7658) );
  AOI211_X1 U9419 ( .C1(n7660), .C2(n7659), .A(n9724), .B(n7658), .ZN(n7665)
         );
  OAI22_X1 U9420 ( .A1(n9718), .A2(n7844), .B1(n7661), .B2(n9717), .ZN(n7664)
         );
  NAND2_X1 U9421 ( .A1(n9709), .A2(n9740), .ZN(n7662) );
  NAND2_X1 U9422 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10279) );
  OAI211_X1 U9423 ( .C1(n7845), .C2(n9712), .A(n7662), .B(n10279), .ZN(n7663)
         );
  OR3_X1 U9424 ( .A1(n7665), .A2(n7664), .A3(n7663), .ZN(P1_U3230) );
  OAI222_X1 U9425 ( .A1(n9502), .A2(n7667), .B1(n9082), .B2(P2_U3151), .C1(
        n9497), .C2(n7666), .ZN(P2_U3278) );
  INV_X1 U9426 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7669) );
  INV_X1 U9427 ( .A(n9858), .ZN(n10342) );
  XNOR2_X1 U9428 ( .A(n7671), .B(n7670), .ZN(n7672) );
  XNOR2_X1 U9429 ( .A(n7673), .B(n7672), .ZN(n7679) );
  INV_X1 U9430 ( .A(n7674), .ZN(n8055) );
  AOI22_X1 U9431 ( .A1(n9695), .A2(n9739), .B1(n9705), .B2(n8055), .ZN(n7675)
         );
  NAND2_X1 U9432 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9796) );
  OAI211_X1 U9433 ( .C1(n7676), .C2(n9719), .A(n7675), .B(n9796), .ZN(n7677)
         );
  AOI21_X1 U9434 ( .B1(n8074), .B2(n9722), .A(n7677), .ZN(n7678) );
  OAI21_X1 U9435 ( .B1(n7679), .B2(n9724), .A(n7678), .ZN(P1_U3213) );
  INV_X1 U9436 ( .A(n7851), .ZN(n7690) );
  NAND2_X1 U9437 ( .A1(n8896), .A2(n4512), .ZN(n7682) );
  AOI21_X1 U9438 ( .B1(n8778), .B2(n8921), .A(n7680), .ZN(n7681) );
  OAI211_X1 U9439 ( .C1(n7683), .C2(n8780), .A(n7682), .B(n7681), .ZN(n7689)
         );
  NAND3_X1 U9440 ( .A1(n7579), .A2(n4976), .A3(n7685), .ZN(n7686) );
  AOI21_X1 U9441 ( .B1(n7687), .B2(n7686), .A(n8898), .ZN(n7688) );
  AOI211_X1 U9442 ( .C1(n7690), .C2(n8906), .A(n7689), .B(n7688), .ZN(n7691)
         );
  INV_X1 U9443 ( .A(n7691), .ZN(P2_U3167) );
  MUX2_X1 U9444 ( .A(n7820), .B(n8105), .S(n10421), .Z(n7694) );
  INV_X1 U9445 ( .A(n8169), .ZN(n7692) );
  AOI22_X1 U9446 ( .A1(n9325), .A2(n8166), .B1(n9341), .B2(n7692), .ZN(n7693)
         );
  OAI211_X1 U9447 ( .C1(n8109), .C2(n9344), .A(n7694), .B(n7693), .ZN(P2_U3225) );
  OAI211_X1 U9448 ( .C1(n7697), .C2(n7696), .A(n7695), .B(n8882), .ZN(n7705)
         );
  NAND2_X1 U9449 ( .A1(n8896), .A2(n7698), .ZN(n7702) );
  INV_X1 U9450 ( .A(n7699), .ZN(n7700) );
  AOI21_X1 U9451 ( .B1(n8778), .B2(n8920), .A(n7700), .ZN(n7701) );
  OAI211_X1 U9452 ( .C1(n4514), .C2(n8780), .A(n7702), .B(n7701), .ZN(n7703)
         );
  INV_X1 U9453 ( .A(n7703), .ZN(n7704) );
  OAI211_X1 U9454 ( .C1(n7706), .C2(n8852), .A(n7705), .B(n7704), .ZN(P2_U3179) );
  INV_X1 U9455 ( .A(n7708), .ZN(n7709) );
  NOR2_X1 U9456 ( .A1(n7709), .A2(n8605), .ZN(n8000) );
  AOI21_X1 U9457 ( .B1(n8605), .B2(n7709), .A(n8000), .ZN(n10350) );
  XNOR2_X1 U9458 ( .A(n7710), .B(n8605), .ZN(n7711) );
  AOI222_X1 U9459 ( .A1(n9739), .A2(n10377), .B1(n10087), .B2(n7711), .C1(
        n9741), .C2(n10085), .ZN(n10360) );
  INV_X1 U9460 ( .A(n7712), .ZN(n8007) );
  OAI211_X1 U9461 ( .C1(n7775), .C2(n7721), .A(n8007), .B(n10052), .ZN(n10356)
         );
  OAI211_X1 U9462 ( .C1(n10401), .C2(n10350), .A(n10360), .B(n10356), .ZN(
        n7781) );
  INV_X1 U9463 ( .A(n7781), .ZN(n7714) );
  AOI22_X1 U9464 ( .A1(n10232), .A2(n10354), .B1(n10403), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n7713) );
  OAI21_X1 U9465 ( .B1(n7714), .B2(n10403), .A(n7713), .ZN(P1_U3468) );
  NOR2_X1 U9466 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  XNOR2_X1 U9467 ( .A(n7717), .B(n8603), .ZN(n7850) );
  INV_X1 U9468 ( .A(n7850), .ZN(n7728) );
  NAND2_X1 U9469 ( .A1(n7718), .A2(n7730), .ZN(n7719) );
  NAND2_X1 U9470 ( .A1(n7719), .A2(n10052), .ZN(n7720) );
  NOR2_X1 U9471 ( .A1(n7721), .A2(n7720), .ZN(n7847) );
  INV_X1 U9472 ( .A(n7722), .ZN(n8673) );
  OAI21_X1 U9473 ( .B1(n8673), .B2(n7723), .A(n8603), .ZN(n7725) );
  NAND2_X1 U9474 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  AOI222_X1 U9475 ( .A1(n7726), .A2(n10087), .B1(n9740), .B2(n10377), .C1(
        n9742), .C2(n10085), .ZN(n7842) );
  INV_X1 U9476 ( .A(n7842), .ZN(n7727) );
  AOI211_X1 U9477 ( .C1(n10195), .C2(n7728), .A(n7847), .B(n7727), .ZN(n7732)
         );
  AOI22_X1 U9478 ( .A1(n10159), .A2(n7730), .B1(n6794), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7729) );
  OAI21_X1 U9479 ( .B1(n7732), .B2(n6794), .A(n7729), .ZN(P1_U3526) );
  AOI22_X1 U9480 ( .A1(n10232), .A2(n7730), .B1(n10403), .B2(
        P1_REG0_REG_4__SCAN_IN), .ZN(n7731) );
  OAI21_X1 U9481 ( .B1(n7732), .B2(n10403), .A(n7731), .ZN(P1_U3465) );
  NAND2_X1 U9482 ( .A1(n7733), .A2(n7734), .ZN(n7770) );
  NOR2_X1 U9483 ( .A1(n7733), .A2(n7734), .ZN(n7769) );
  AOI21_X1 U9484 ( .B1(n7772), .B2(n7770), .A(n7769), .ZN(n7738) );
  XNOR2_X1 U9485 ( .A(n7736), .B(n7735), .ZN(n7737) );
  XNOR2_X1 U9486 ( .A(n7738), .B(n7737), .ZN(n7744) );
  INV_X1 U9487 ( .A(n8008), .ZN(n7742) );
  NAND2_X1 U9488 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9783) );
  OAI21_X1 U9489 ( .B1(n9712), .B2(n8009), .A(n9783), .ZN(n7741) );
  OAI22_X1 U9490 ( .A1(n9719), .A2(n8175), .B1(n7739), .B2(n9717), .ZN(n7740)
         );
  AOI211_X1 U9491 ( .C1(n7742), .C2(n9705), .A(n7741), .B(n7740), .ZN(n7743)
         );
  OAI21_X1 U9492 ( .B1(n7744), .B2(n9724), .A(n7743), .ZN(P1_U3239) );
  MUX2_X1 U9493 ( .A(n7746), .B(n7745), .S(n9404), .Z(n7747) );
  OAI21_X1 U9494 ( .B1(n7748), .B2(n9381), .A(n7747), .ZN(P2_U3462) );
  MUX2_X1 U9495 ( .A(n7750), .B(n7749), .S(n9404), .Z(n7751) );
  OAI21_X1 U9496 ( .B1(n7852), .B2(n9381), .A(n7751), .ZN(P2_U3464) );
  MUX2_X1 U9497 ( .A(n7753), .B(n7752), .S(n9404), .Z(n7754) );
  OAI21_X1 U9498 ( .B1(n10414), .B2(n9381), .A(n7754), .ZN(P2_U3463) );
  MUX2_X1 U9499 ( .A(n7086), .B(n7755), .S(n9404), .Z(n7756) );
  OAI21_X1 U9500 ( .B1(n7757), .B2(n9381), .A(n7756), .ZN(P2_U3459) );
  XNOR2_X1 U9501 ( .A(n7758), .B(n7760), .ZN(n8066) );
  NAND2_X1 U9502 ( .A1(n8066), .A2(n6742), .ZN(n7766) );
  AOI22_X1 U9503 ( .A1(n9333), .A2(n8917), .B1(n8919), .B2(n9331), .ZN(n7765)
         );
  NAND2_X1 U9504 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  NAND2_X1 U9505 ( .A1(n7759), .A2(n7762), .ZN(n7763) );
  NAND2_X1 U9506 ( .A1(n7763), .A2(n9336), .ZN(n7764) );
  NAND3_X1 U9507 ( .A1(n7766), .A2(n7765), .A3(n7764), .ZN(n8062) );
  AOI21_X1 U9508 ( .B1(n7767), .B2(n8066), .A(n8062), .ZN(n7996) );
  AOI22_X1 U9509 ( .A1(n9485), .A2(n8269), .B1(P2_REG0_REG_9__SCAN_IN), .B2(
        n10441), .ZN(n7768) );
  OAI21_X1 U9510 ( .B1(n7996), .B2(n10441), .A(n7768), .ZN(P2_U3417) );
  INV_X1 U9511 ( .A(n7769), .ZN(n7771) );
  NAND2_X1 U9512 ( .A1(n7771), .A2(n7770), .ZN(n7773) );
  XNOR2_X1 U9513 ( .A(n7773), .B(n7772), .ZN(n7780) );
  INV_X1 U9514 ( .A(n10351), .ZN(n7774) );
  AOI22_X1 U9515 ( .A1(n9695), .A2(n9741), .B1(n9705), .B2(n7774), .ZN(n7779)
         );
  NAND2_X1 U9516 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9770) );
  INV_X1 U9517 ( .A(n9770), .ZN(n7777) );
  NOR2_X1 U9518 ( .A1(n9712), .A2(n7775), .ZN(n7776) );
  AOI211_X1 U9519 ( .C1(n9709), .C2(n9739), .A(n7777), .B(n7776), .ZN(n7778)
         );
  OAI211_X1 U9520 ( .C1(n7780), .C2(n9724), .A(n7779), .B(n7778), .ZN(P1_U3227) );
  NAND2_X1 U9521 ( .A1(n7781), .A2(n10408), .ZN(n7783) );
  NAND2_X1 U9522 ( .A1(n10159), .A2(n10354), .ZN(n7782) );
  OAI211_X1 U9523 ( .C1(n10408), .C2(n7253), .A(n7783), .B(n7782), .ZN(
        P1_U3527) );
  INV_X1 U9524 ( .A(n7784), .ZN(n7785) );
  MUX2_X1 U9525 ( .A(n7530), .B(n7785), .S(n10421), .Z(n7788) );
  INV_X1 U9526 ( .A(n7786), .ZN(n8039) );
  AOI22_X1 U9527 ( .A1(n9325), .A2(n8033), .B1(n9341), .B2(n8039), .ZN(n7787)
         );
  OAI211_X1 U9528 ( .C1(n7789), .C2(n9159), .A(n7788), .B(n7787), .ZN(P2_U3226) );
  AND2_X1 U9529 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  NAND2_X1 U9530 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  NAND2_X1 U9531 ( .A1(n10386), .A2(n7795), .ZN(n8190) );
  OR2_X1 U9532 ( .A1(n7796), .A2(n10361), .ZN(n7804) );
  OAI22_X1 U9533 ( .A1(n10386), .A2(n7799), .B1(n7798), .B2(n10379), .ZN(n7802) );
  NAND2_X1 U9534 ( .A1(n10386), .A2(n8590), .ZN(n10369) );
  NOR2_X1 U9535 ( .A1(n10369), .A2(n7800), .ZN(n7801) );
  AOI211_X1 U9536 ( .C1(n10366), .C2(n9567), .A(n7802), .B(n7801), .ZN(n7803)
         );
  OAI211_X1 U9537 ( .C1(n7805), .C2(n8190), .A(n7804), .B(n7803), .ZN(P1_U3292) );
  MUX2_X1 U9538 ( .A(n7939), .B(n7806), .S(n9404), .Z(n7807) );
  OAI21_X1 U9539 ( .B1(n7808), .B2(n9381), .A(n7807), .ZN(P2_U3466) );
  INV_X1 U9540 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7997) );
  INV_X1 U9541 ( .A(n7809), .ZN(n8940) );
  INV_X1 U9542 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8106) );
  XNOR2_X1 U9543 ( .A(n7821), .B(n8106), .ZN(n8941) );
  INV_X1 U9544 ( .A(n7811), .ZN(n7813) );
  NAND2_X1 U9545 ( .A1(n7811), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8965) );
  INV_X1 U9546 ( .A(n8965), .ZN(n7812) );
  AOI21_X1 U9547 ( .B1(n7997), .B2(n7813), .A(n7812), .ZN(n7836) );
  NAND2_X1 U9548 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8266) );
  OAI21_X1 U9549 ( .B1(n9131), .B2(n4860), .A(n8266), .ZN(n7819) );
  XNOR2_X1 U9550 ( .A(n7821), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U9551 ( .A1(n7816), .A2(n7910), .ZN(n7817) );
  AOI21_X1 U9552 ( .B1(n8953), .B2(n7817), .A(n9144), .ZN(n7818) );
  AOI211_X1 U9553 ( .C1(n9142), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7819), .B(
        n7818), .ZN(n7835) );
  MUX2_X1 U9554 ( .A(n7820), .B(n8106), .S(n4279), .Z(n7822) );
  NAND2_X1 U9555 ( .A1(n7822), .A2(n7821), .ZN(n7825) );
  INV_X1 U9556 ( .A(n7822), .ZN(n7823) );
  NAND2_X1 U9557 ( .A1(n7823), .A2(n8927), .ZN(n7824) );
  NAND2_X1 U9558 ( .A1(n7825), .A2(n7824), .ZN(n8935) );
  INV_X1 U9559 ( .A(n7825), .ZN(n7831) );
  MUX2_X1 U9560 ( .A(n7910), .B(n7997), .S(n4279), .Z(n7827) );
  NAND2_X1 U9561 ( .A1(n7827), .A2(n7826), .ZN(n8959) );
  INV_X1 U9562 ( .A(n7827), .ZN(n7828) );
  NAND2_X1 U9563 ( .A1(n7828), .A2(n4860), .ZN(n7829) );
  AND2_X1 U9564 ( .A1(n8959), .A2(n7829), .ZN(n7830) );
  INV_X1 U9565 ( .A(n8960), .ZN(n7833) );
  NOR3_X1 U9566 ( .A1(n8939), .A2(n7831), .A3(n7830), .ZN(n7832) );
  OAI21_X1 U9567 ( .B1(n7833), .B2(n7832), .A(n9042), .ZN(n7834) );
  OAI211_X1 U9568 ( .C1(n7836), .C2(n9037), .A(n7835), .B(n7834), .ZN(P2_U3191) );
  INV_X1 U9569 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7838) );
  INV_X1 U9570 ( .A(n7837), .ZN(n7839) );
  OAI222_X1 U9571 ( .A1(n9502), .A2(n7838), .B1(n9497), .B2(n7839), .C1(n9130), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U9572 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7840) );
  OAI222_X1 U9573 ( .A1(n10259), .A2(n7840), .B1(n10262), .B2(n7839), .C1(
        P1_U3086), .C2(n8590), .ZN(P1_U3336) );
  INV_X1 U9574 ( .A(n8052), .ZN(n8183) );
  NAND2_X1 U9575 ( .A1(n10386), .A2(n8183), .ZN(n7841) );
  MUX2_X1 U9576 ( .A(n7843), .B(n7842), .S(n10386), .Z(n7849) );
  OAI22_X1 U9577 ( .A1(n10069), .A2(n7845), .B1(n7844), .B2(n10379), .ZN(n7846) );
  AOI21_X1 U9578 ( .B1(n10115), .B2(n7847), .A(n7846), .ZN(n7848) );
  OAI211_X1 U9579 ( .C1(n10079), .C2(n7850), .A(n7849), .B(n7848), .ZN(
        P1_U3289) );
  OAI22_X1 U9580 ( .A1(n10415), .A2(n7852), .B1(n7851), .B2(n10417), .ZN(n7855) );
  MUX2_X1 U9581 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7853), .S(n10421), .Z(n7854)
         );
  AOI211_X1 U9582 ( .C1(n7856), .C2(n9283), .A(n7855), .B(n7854), .ZN(n7995)
         );
  XOR2_X1 U9583 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput6), .Z(n7860) );
  XOR2_X1 U9584 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput51), .Z(n7859) );
  XOR2_X1 U9585 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput1), .Z(n7858) );
  XOR2_X1 U9586 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(keyinput63), .Z(n7857) );
  NOR4_X1 U9587 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n7880)
         );
  XOR2_X1 U9588 ( .A(SI_5_), .B(keyinput2), .Z(n7867) );
  XNOR2_X1 U9589 ( .A(n7861), .B(keyinput56), .ZN(n7866) );
  XNOR2_X1 U9590 ( .A(n7862), .B(keyinput48), .ZN(n7865) );
  XNOR2_X1 U9591 ( .A(n7863), .B(keyinput7), .ZN(n7864) );
  NOR4_X1 U9592 ( .A1(n7867), .A2(n7866), .A3(n7865), .A4(n7864), .ZN(n7879)
         );
  XOR2_X1 U9593 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput61), .Z(n7872) );
  XOR2_X1 U9594 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput52), .Z(n7871) );
  XOR2_X1 U9595 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput54), .Z(n7870) );
  XNOR2_X1 U9596 ( .A(n7868), .B(keyinput21), .ZN(n7869) );
  NOR4_X1 U9597 ( .A1(n7872), .A2(n7871), .A3(n7870), .A4(n7869), .ZN(n7878)
         );
  XNOR2_X1 U9598 ( .A(n5162), .B(keyinput41), .ZN(n7876) );
  XOR2_X1 U9599 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput35), .Z(n7875) );
  XNOR2_X1 U9600 ( .A(n7939), .B(keyinput38), .ZN(n7874) );
  INV_X1 U9601 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8386) );
  XNOR2_X1 U9602 ( .A(n8386), .B(keyinput40), .ZN(n7873) );
  NOR4_X1 U9603 ( .A1(n7876), .A2(n7875), .A3(n7874), .A4(n7873), .ZN(n7877)
         );
  NAND4_X1 U9604 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n7887)
         );
  AOI22_X1 U9605 ( .A1(n8424), .A2(keyinput59), .B1(n8430), .B2(keyinput57), 
        .ZN(n7881) );
  OAI221_X1 U9606 ( .B1(n8424), .B2(keyinput59), .C1(n8430), .C2(keyinput57), 
        .A(n7881), .ZN(n7886) );
  INV_X1 U9607 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10388) );
  INV_X1 U9608 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8392) );
  AOI22_X1 U9609 ( .A1(n10388), .A2(keyinput34), .B1(keyinput62), .B2(n8392), 
        .ZN(n7882) );
  OAI221_X1 U9610 ( .B1(n10388), .B2(keyinput34), .C1(n8392), .C2(keyinput62), 
        .A(n7882), .ZN(n7885) );
  XNOR2_X1 U9611 ( .A(n7883), .B(keyinput47), .ZN(n7884) );
  NOR4_X1 U9612 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n7923)
         );
  INV_X1 U9613 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9810) );
  AOI22_X1 U9614 ( .A1(n9810), .A2(keyinput5), .B1(n9574), .B2(keyinput25), 
        .ZN(n7888) );
  OAI221_X1 U9615 ( .B1(n9810), .B2(keyinput5), .C1(n9574), .C2(keyinput25), 
        .A(n7888), .ZN(n7904) );
  XNOR2_X1 U9616 ( .A(keyinput4), .B(n7940), .ZN(n7889) );
  AOI21_X1 U9617 ( .B1(n7953), .B2(keyinput50), .A(n7889), .ZN(n7892) );
  XOR2_X1 U9618 ( .A(n5121), .B(keyinput45), .Z(n7891) );
  XNOR2_X1 U9619 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput0), .ZN(n7890) );
  NAND3_X1 U9620 ( .A1(n7892), .A2(n7891), .A3(n7890), .ZN(n7903) );
  XNOR2_X1 U9621 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput22), .ZN(n7896) );
  XNOR2_X1 U9622 ( .A(P1_REG0_REG_28__SCAN_IN), .B(keyinput16), .ZN(n7895) );
  XNOR2_X1 U9623 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput11), .ZN(n7894) );
  XNOR2_X1 U9624 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput13), .ZN(n7893) );
  NAND4_X1 U9625 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n7902)
         );
  XNOR2_X1 U9626 ( .A(SI_3_), .B(keyinput29), .ZN(n7900) );
  XNOR2_X1 U9627 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput32), .ZN(n7899) );
  XNOR2_X1 U9628 ( .A(SI_20_), .B(keyinput28), .ZN(n7898) );
  XNOR2_X1 U9629 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput17), .ZN(n7897) );
  NAND4_X1 U9630 ( .A1(n7900), .A2(n7899), .A3(n7898), .A4(n7897), .ZN(n7901)
         );
  NOR4_X1 U9631 ( .A1(n7904), .A2(n7903), .A3(n7902), .A4(n7901), .ZN(n7922)
         );
  INV_X1 U9632 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10404) );
  INV_X1 U9633 ( .A(SI_21_), .ZN(n7949) );
  AOI22_X1 U9634 ( .A1(n10404), .A2(keyinput60), .B1(n7949), .B2(keyinput37), 
        .ZN(n7905) );
  OAI221_X1 U9635 ( .B1(n10404), .B2(keyinput60), .C1(n7949), .C2(keyinput37), 
        .A(n7905), .ZN(n7913) );
  INV_X1 U9636 ( .A(SI_11_), .ZN(n7907) );
  AOI22_X1 U9637 ( .A1(n8766), .A2(keyinput19), .B1(n7907), .B2(keyinput43), 
        .ZN(n7906) );
  OAI221_X1 U9638 ( .B1(n8766), .B2(keyinput19), .C1(n7907), .C2(keyinput43), 
        .A(n7906), .ZN(n7912) );
  AOI22_X1 U9639 ( .A1(n7910), .A2(keyinput46), .B1(n7909), .B2(keyinput23), 
        .ZN(n7908) );
  OAI221_X1 U9640 ( .B1(n7910), .B2(keyinput46), .C1(n7909), .C2(keyinput23), 
        .A(n7908), .ZN(n7911) );
  NOR3_X1 U9641 ( .A1(n7913), .A2(n7912), .A3(n7911), .ZN(n7921) );
  INV_X1 U9642 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7915) );
  AOI22_X1 U9643 ( .A1(n7928), .A2(keyinput26), .B1(keyinput18), .B2(n7915), 
        .ZN(n7914) );
  OAI221_X1 U9644 ( .B1(n7928), .B2(keyinput26), .C1(n7915), .C2(keyinput18), 
        .A(n7914), .ZN(n7919) );
  AOI22_X1 U9645 ( .A1(n7917), .A2(keyinput9), .B1(keyinput15), .B2(n7264), 
        .ZN(n7916) );
  OAI221_X1 U9646 ( .B1(n7917), .B2(keyinput9), .C1(n7264), .C2(keyinput15), 
        .A(n7916), .ZN(n7918) );
  NOR2_X1 U9647 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  NAND4_X1 U9648 ( .A1(n7923), .A2(n7922), .A3(n7921), .A4(n7920), .ZN(n7993)
         );
  INV_X1 U9649 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U9650 ( .A1(n9810), .A2(n7956), .ZN(n8139) );
  INV_X1 U9651 ( .A(n8139), .ZN(n8131) );
  NOR4_X1 U9652 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .A3(P1_ADDR_REG_9__SCAN_IN), .A4(n7983), .ZN(n7925) );
  NOR4_X1 U9653 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P1_REG2_REG_31__SCAN_IN), 
        .A3(n9847), .A4(n8430), .ZN(n7924) );
  NAND4_X1 U9654 ( .A1(n7926), .A2(n8131), .A3(n7925), .A4(n7924), .ZN(n7948)
         );
  NOR4_X1 U9655 ( .A1(n7968), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(SI_11_), .A4(
        P1_REG3_REG_21__SCAN_IN), .ZN(n7936) );
  INV_X1 U9656 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9470) );
  NAND4_X1 U9657 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(P2_REG2_REG_9__SCAN_IN), 
        .A3(n9470), .A4(n7970), .ZN(n7933) );
  INV_X1 U9658 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7959) );
  NAND4_X1 U9659 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_REG2_REG_11__SCAN_IN), 
        .A3(n7960), .A4(n7959), .ZN(n7932) );
  INV_X1 U9660 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7962) );
  NOR4_X1 U9661 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .A3(n7927), .A4(n7962), .ZN(n7930) );
  NOR4_X1 U9662 ( .A1(SI_5_), .A2(P1_REG3_REG_17__SCAN_IN), .A3(
        P2_REG3_REG_21__SCAN_IN), .A4(n7928), .ZN(n7929) );
  NAND2_X1 U9663 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  NOR4_X1 U9664 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n7935) );
  INV_X1 U9665 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7934) );
  NAND4_X1 U9666 ( .A1(n7936), .A2(P1_IR_REG_24__SCAN_IN), .A3(n7935), .A4(
        n7934), .ZN(n7947) );
  NAND4_X1 U9667 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_DATAO_REG_18__SCAN_IN), 
        .A3(P1_DATAO_REG_6__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n7946) );
  NAND4_X1 U9668 ( .A1(SI_3_), .A2(SI_20_), .A3(P1_REG0_REG_28__SCAN_IN), .A4(
        P2_DATAO_REG_24__SCAN_IN), .ZN(n7944) );
  INV_X1 U9669 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n7937) );
  NAND4_X1 U9670 ( .A1(n8386), .A2(n7938), .A3(n7937), .A4(
        P2_IR_REG_22__SCAN_IN), .ZN(n7943) );
  NAND4_X1 U9671 ( .A1(n7940), .A2(n7939), .A3(P1_DATAO_REG_1__SCAN_IN), .A4(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7942) );
  NAND4_X1 U9672 ( .A1(n8766), .A2(P2_IR_REG_26__SCAN_IN), .A3(
        P2_IR_REG_1__SCAN_IN), .A4(P2_IR_REG_28__SCAN_IN), .ZN(n7941) );
  OR4_X1 U9673 ( .A1(n7944), .A2(n7943), .A3(n7942), .A4(n7941), .ZN(n7945) );
  NOR4_X1 U9674 ( .A1(n7948), .A2(n7947), .A3(n7946), .A4(n7945), .ZN(n7952)
         );
  NOR4_X1 U9675 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P1_DATAO_REG_30__SCAN_IN), .A4(n10404), .ZN(n7951) );
  NOR4_X1 U9676 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .A4(n7949), .ZN(n7950) );
  NAND3_X1 U9677 ( .A1(n7952), .A2(n7951), .A3(n7950), .ZN(n7954) );
  AOI21_X1 U9678 ( .B1(n7954), .B2(keyinput50), .A(n7953), .ZN(n7992) );
  INV_X1 U9679 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7957) );
  AOI22_X1 U9680 ( .A1(n7957), .A2(keyinput42), .B1(keyinput20), .B2(n7956), 
        .ZN(n7955) );
  OAI221_X1 U9681 ( .B1(n7957), .B2(keyinput42), .C1(n7956), .C2(keyinput20), 
        .A(n7955), .ZN(n7966) );
  AOI22_X1 U9682 ( .A1(n7960), .A2(keyinput12), .B1(keyinput27), .B2(n7959), 
        .ZN(n7958) );
  OAI221_X1 U9683 ( .B1(n7960), .B2(keyinput12), .C1(n7959), .C2(keyinput27), 
        .A(n7958), .ZN(n7965) );
  AOI22_X1 U9684 ( .A1(n7963), .A2(keyinput8), .B1(keyinput49), .B2(n7962), 
        .ZN(n7961) );
  OAI221_X1 U9685 ( .B1(n7963), .B2(keyinput8), .C1(n7962), .C2(keyinput49), 
        .A(n7961), .ZN(n7964) );
  NOR3_X1 U9686 ( .A1(n7966), .A2(n7965), .A3(n7964), .ZN(n7990) );
  AOI22_X1 U9687 ( .A1(n7968), .A2(keyinput39), .B1(keyinput36), .B2(n7938), 
        .ZN(n7967) );
  OAI221_X1 U9688 ( .B1(n7968), .B2(keyinput39), .C1(n7938), .C2(keyinput36), 
        .A(n7967), .ZN(n7974) );
  AOI22_X1 U9689 ( .A1(n7970), .A2(keyinput3), .B1(keyinput53), .B2(n9470), 
        .ZN(n7969) );
  OAI221_X1 U9690 ( .B1(n7970), .B2(keyinput3), .C1(n9470), .C2(keyinput53), 
        .A(n7969), .ZN(n7973) );
  AOI22_X1 U9691 ( .A1(n8739), .A2(keyinput30), .B1(n9847), .B2(keyinput58), 
        .ZN(n7971) );
  OAI221_X1 U9692 ( .B1(n8739), .B2(keyinput30), .C1(n9847), .C2(keyinput58), 
        .A(n7971), .ZN(n7972) );
  NOR3_X1 U9693 ( .A1(n7974), .A2(n7973), .A3(n7972), .ZN(n7989) );
  AOI22_X1 U9694 ( .A1(n7976), .A2(keyinput10), .B1(keyinput31), .B2(n7086), 
        .ZN(n7975) );
  OAI221_X1 U9695 ( .B1(n7976), .B2(keyinput10), .C1(n7086), .C2(keyinput31), 
        .A(n7975), .ZN(n7981) );
  AOI22_X1 U9696 ( .A1(n7979), .A2(keyinput24), .B1(keyinput55), .B2(n7978), 
        .ZN(n7977) );
  OAI221_X1 U9697 ( .B1(n7979), .B2(keyinput24), .C1(n7978), .C2(keyinput55), 
        .A(n7977), .ZN(n7980) );
  NOR2_X1 U9698 ( .A1(n7981), .A2(n7980), .ZN(n7988) );
  AOI22_X1 U9699 ( .A1(n10260), .A2(keyinput44), .B1(keyinput14), .B2(n7983), 
        .ZN(n7982) );
  OAI221_X1 U9700 ( .B1(n10260), .B2(keyinput44), .C1(n7983), .C2(keyinput14), 
        .A(n7982), .ZN(n7986) );
  XNOR2_X1 U9701 ( .A(n7984), .B(keyinput33), .ZN(n7985) );
  NOR2_X1 U9702 ( .A1(n7986), .A2(n7985), .ZN(n7987) );
  NAND4_X1 U9703 ( .A1(n7990), .A2(n7989), .A3(n7988), .A4(n7987), .ZN(n7991)
         );
  NOR3_X1 U9704 ( .A1(n7993), .A2(n7992), .A3(n7991), .ZN(n7994) );
  XNOR2_X1 U9705 ( .A(n7995), .B(n7994), .ZN(P2_U3228) );
  INV_X1 U9706 ( .A(n8269), .ZN(n8061) );
  MUX2_X1 U9707 ( .A(n7997), .B(n7996), .S(n9404), .Z(n7998) );
  OAI21_X1 U9708 ( .B1(n8061), .B2(n9381), .A(n7998), .ZN(P2_U3468) );
  NOR2_X1 U9709 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  NOR2_X1 U9710 ( .A1(n8001), .A2(n8003), .ZN(n8043) );
  AOI21_X1 U9711 ( .B1(n8001), .B2(n8003), .A(n8043), .ZN(n10400) );
  XNOR2_X1 U9712 ( .A(n8002), .B(n8003), .ZN(n8004) );
  AOI222_X1 U9713 ( .A1(n9738), .A2(n10377), .B1(n10087), .B2(n8004), .C1(
        n9740), .C2(n10085), .ZN(n10399) );
  MUX2_X1 U9714 ( .A(n8005), .B(n10399), .S(n10386), .Z(n8012) );
  INV_X1 U9715 ( .A(n8054), .ZN(n8006) );
  AOI211_X1 U9716 ( .C1(n4902), .C2(n8007), .A(n10091), .B(n8006), .ZN(n10396)
         );
  OAI22_X1 U9717 ( .A1(n10069), .A2(n8009), .B1(n8008), .B2(n10379), .ZN(n8010) );
  AOI21_X1 U9718 ( .B1(n10396), .B2(n10115), .A(n8010), .ZN(n8011) );
  OAI211_X1 U9719 ( .C1(n10079), .C2(n10400), .A(n8012), .B(n8011), .ZN(
        P1_U3287) );
  INV_X1 U9720 ( .A(n8013), .ZN(n8023) );
  INV_X2 U9721 ( .A(n10386), .ZN(n10361) );
  OAI22_X1 U9722 ( .A1(n10386), .A2(n8015), .B1(n8014), .B2(n10379), .ZN(n8018) );
  NOR2_X1 U9723 ( .A1(n10069), .A2(n8016), .ZN(n8017) );
  AOI211_X1 U9724 ( .C1(n8019), .C2(n10115), .A(n8018), .B(n8017), .ZN(n8022)
         );
  NAND2_X1 U9725 ( .A1(n8020), .A2(n10371), .ZN(n8021) );
  OAI211_X1 U9726 ( .C1(n8023), .C2(n10361), .A(n8022), .B(n8021), .ZN(
        P1_U3291) );
  OAI21_X1 U9727 ( .B1(n8025), .B2(n5794), .A(n8024), .ZN(n8221) );
  XOR2_X1 U9728 ( .A(n8027), .B(n8026), .Z(n8028) );
  OAI222_X1 U9729 ( .A1(n9296), .A2(n8164), .B1(n9298), .B2(n8784), .C1(n9293), 
        .C2(n8028), .ZN(n8218) );
  AOI21_X1 U9730 ( .B1(n10426), .B2(n8221), .A(n8218), .ZN(n8216) );
  AOI22_X1 U9731 ( .A1(n9485), .A2(n8215), .B1(P2_REG0_REG_10__SCAN_IN), .B2(
        n10441), .ZN(n8029) );
  OAI21_X1 U9732 ( .B1(n8216), .B2(n10441), .A(n8029), .ZN(P2_U3420) );
  INV_X1 U9733 ( .A(n8030), .ZN(n8159) );
  AOI21_X1 U9734 ( .B1(n8032), .B2(n8031), .A(n8159), .ZN(n8041) );
  NAND2_X1 U9735 ( .A1(n8896), .A2(n8033), .ZN(n8036) );
  AOI21_X1 U9736 ( .B1(n8778), .B2(n8919), .A(n8034), .ZN(n8035) );
  OAI211_X1 U9737 ( .C1(n8037), .C2(n8780), .A(n8036), .B(n8035), .ZN(n8038)
         );
  AOI21_X1 U9738 ( .B1(n8039), .B2(n8906), .A(n8038), .ZN(n8040) );
  OAI21_X1 U9739 ( .B1(n8041), .B2(n8898), .A(n8040), .ZN(P2_U3153) );
  NOR2_X1 U9740 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  NOR2_X1 U9741 ( .A1(n8044), .A2(n5115), .ZN(n8174) );
  AOI21_X1 U9742 ( .B1(n8044), .B2(n5115), .A(n8174), .ZN(n8068) );
  AOI22_X1 U9743 ( .A1(n9739), .A2(n10085), .B1(n10377), .B2(n9737), .ZN(n8051) );
  OR2_X1 U9744 ( .A1(n8002), .A2(n8045), .ZN(n8047) );
  NAND3_X1 U9745 ( .A1(n8047), .A2(n5115), .A3(n8046), .ZN(n8177) );
  INV_X1 U9746 ( .A(n8177), .ZN(n8049) );
  AOI21_X1 U9747 ( .B1(n8047), .B2(n8046), .A(n5115), .ZN(n8048) );
  OAI21_X1 U9748 ( .B1(n8049), .B2(n8048), .A(n10087), .ZN(n8050) );
  OAI211_X1 U9749 ( .C1(n8068), .C2(n8052), .A(n8051), .B(n8050), .ZN(n8069)
         );
  NAND2_X1 U9750 ( .A1(n8069), .A2(n10386), .ZN(n8060) );
  INV_X1 U9751 ( .A(n8185), .ZN(n8053) );
  AOI211_X1 U9752 ( .C1(n8074), .C2(n8054), .A(n10091), .B(n8053), .ZN(n8070)
         );
  INV_X1 U9753 ( .A(n8074), .ZN(n8057) );
  INV_X1 U9754 ( .A(n10379), .ZN(n10066) );
  AOI22_X1 U9755 ( .A1(n10361), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8055), .B2(
        n10066), .ZN(n8056) );
  OAI21_X1 U9756 ( .B1(n10069), .B2(n8057), .A(n8056), .ZN(n8058) );
  AOI21_X1 U9757 ( .B1(n8070), .B2(n10115), .A(n8058), .ZN(n8059) );
  OAI211_X1 U9758 ( .C1(n8068), .C2(n8190), .A(n8060), .B(n8059), .ZN(P1_U3286) );
  INV_X1 U9759 ( .A(n9159), .ZN(n8065) );
  OAI22_X1 U9760 ( .A1(n10415), .A2(n8061), .B1(n8272), .B2(n10417), .ZN(n8064) );
  MUX2_X1 U9761 ( .A(n8062), .B(P2_REG2_REG_9__SCAN_IN), .S(n10413), .Z(n8063)
         );
  AOI211_X1 U9762 ( .C1(n8066), .C2(n8065), .A(n8064), .B(n8063), .ZN(n8067)
         );
  INV_X1 U9763 ( .A(n8067), .ZN(P2_U3224) );
  INV_X1 U9764 ( .A(n10212), .ZN(n8072) );
  INV_X1 U9765 ( .A(n8068), .ZN(n8071) );
  AOI211_X1 U9766 ( .C1(n8072), .C2(n8071), .A(n8070), .B(n8069), .ZN(n8076)
         );
  AOI22_X1 U9767 ( .A1(n10232), .A2(n8074), .B1(n10403), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n8073) );
  OAI21_X1 U9768 ( .B1(n8076), .B2(n10403), .A(n8073), .ZN(P1_U3474) );
  AOI22_X1 U9769 ( .A1(n10159), .A2(n8074), .B1(n6794), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n8075) );
  OAI21_X1 U9770 ( .B1(n8076), .B2(n6794), .A(n8075), .ZN(P1_U3529) );
  AOI21_X1 U9771 ( .B1(n8077), .B2(n8611), .A(n10392), .ZN(n8080) );
  OAI22_X1 U9772 ( .A1(n9546), .A2(n10043), .B1(n9583), .B2(n10045), .ZN(n8079) );
  AOI21_X1 U9773 ( .B1(n8080), .B2(n8078), .A(n8079), .ZN(n10205) );
  OAI21_X1 U9774 ( .B1(n8082), .B2(n8611), .A(n8081), .ZN(n10202) );
  AOI211_X1 U9775 ( .C1(n10204), .C2(n8094), .A(n10091), .B(n8280), .ZN(n10203) );
  NAND2_X1 U9776 ( .A1(n10203), .A2(n10115), .ZN(n8085) );
  INV_X1 U9777 ( .A(n8083), .ZN(n9580) );
  AOI22_X1 U9778 ( .A1(n10361), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9580), .B2(
        n10066), .ZN(n8084) );
  OAI211_X1 U9779 ( .C1(n8512), .C2(n10069), .A(n8085), .B(n8084), .ZN(n8086)
         );
  AOI21_X1 U9780 ( .B1(n10371), .B2(n10202), .A(n8086), .ZN(n8087) );
  OAI21_X1 U9781 ( .B1(n10361), .B2(n10205), .A(n8087), .ZN(P1_U3281) );
  XNOR2_X1 U9782 ( .A(n8088), .B(n8092), .ZN(n8089) );
  OAI222_X1 U9783 ( .A1(n8089), .A2(n10392), .B1(n10043), .B2(n9640), .C1(
        n10045), .C2(n9682), .ZN(n8207) );
  INV_X1 U9784 ( .A(n8207), .ZN(n8101) );
  OAI21_X1 U9785 ( .B1(n8090), .B2(n8092), .A(n8091), .ZN(n8209) );
  INV_X1 U9786 ( .A(n8094), .ZN(n8095) );
  AOI211_X1 U9787 ( .C1(n9690), .C2(n8093), .A(n10091), .B(n8095), .ZN(n8208)
         );
  NAND2_X1 U9788 ( .A1(n8208), .A2(n10115), .ZN(n8098) );
  INV_X1 U9789 ( .A(n8096), .ZN(n9680) );
  AOI22_X1 U9790 ( .A1(n10361), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9680), .B2(
        n10066), .ZN(n8097) );
  OAI211_X1 U9791 ( .C1(n4440), .C2(n10069), .A(n8098), .B(n8097), .ZN(n8099)
         );
  AOI21_X1 U9792 ( .B1(n10371), .B2(n8209), .A(n8099), .ZN(n8100) );
  OAI21_X1 U9793 ( .B1(n10361), .B2(n8101), .A(n8100), .ZN(P1_U3282) );
  INV_X1 U9794 ( .A(n8102), .ZN(n8261) );
  INV_X1 U9795 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8103) );
  OAI222_X1 U9796 ( .A1(n9497), .A2(n8261), .B1(P2_U3151), .B2(n8104), .C1(
        n8103), .C2(n9502), .ZN(P2_U3275) );
  MUX2_X1 U9797 ( .A(n8106), .B(n8105), .S(n9404), .Z(n8108) );
  NAND2_X1 U9798 ( .A1(n9406), .A2(n8166), .ZN(n8107) );
  OAI211_X1 U9799 ( .C1(n8109), .C2(n9403), .A(n8108), .B(n8107), .ZN(P2_U3467) );
  OR2_X1 U9800 ( .A1(n8110), .A2(n8595), .ZN(n8111) );
  NAND2_X1 U9801 ( .A1(n8112), .A2(n8111), .ZN(n10103) );
  OR2_X1 U9802 ( .A1(n8113), .A2(n9551), .ZN(n8114) );
  AND3_X1 U9803 ( .A1(n8093), .A2(n8114), .A3(n10052), .ZN(n10104) );
  INV_X1 U9804 ( .A(n8115), .ZN(n8116) );
  AOI21_X1 U9805 ( .B1(n8117), .B2(n8595), .A(n8116), .ZN(n8118) );
  OAI222_X1 U9806 ( .A1(n10045), .A2(n9546), .B1(n10043), .B2(n8232), .C1(
        n8118), .C2(n10392), .ZN(n10098) );
  AOI211_X1 U9807 ( .C1(n10195), .C2(n10103), .A(n10104), .B(n10098), .ZN(
        n8121) );
  AOI22_X1 U9808 ( .A1(n10102), .A2(n10159), .B1(P1_REG1_REG_10__SCAN_IN), 
        .B2(n6794), .ZN(n8119) );
  OAI21_X1 U9809 ( .B1(n8121), .B2(n6794), .A(n8119), .ZN(P1_U3532) );
  AOI22_X1 U9810 ( .A1(n10102), .A2(n10232), .B1(P1_REG0_REG_10__SCAN_IN), 
        .B2(n10403), .ZN(n8120) );
  OAI21_X1 U9811 ( .B1(n8121), .B2(n10403), .A(n8120), .ZN(P1_U3483) );
  INV_X1 U9812 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10455) );
  INV_X1 U9813 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10333) );
  INV_X1 U9814 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8122) );
  AOI22_X1 U9815 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10333), .B2(n8122), .ZN(n10461) );
  NOR2_X1 U9816 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8123) );
  AOI21_X1 U9817 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8123), .ZN(n10464) );
  NOR2_X1 U9818 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8124) );
  AOI21_X1 U9819 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n8124), .ZN(n10467) );
  NOR2_X1 U9820 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8125) );
  AOI21_X1 U9821 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8125), .ZN(n10470) );
  NOR2_X1 U9822 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8126) );
  AOI21_X1 U9823 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8126), .ZN(n10473) );
  NOR2_X1 U9824 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8127) );
  AOI21_X1 U9825 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8127), .ZN(n10476) );
  NOR2_X1 U9826 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8128) );
  AOI21_X1 U9827 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8128), .ZN(n10479) );
  NOR2_X1 U9828 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8129) );
  AOI21_X1 U9829 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8129), .ZN(n10482) );
  NOR2_X1 U9830 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8130) );
  AOI21_X1 U9831 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n8130), .ZN(n10491) );
  AOI21_X1 U9832 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n8131), .ZN(n10497) );
  NOR2_X1 U9833 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8132) );
  AOI21_X1 U9834 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n8132), .ZN(n10494) );
  NOR2_X1 U9835 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8133) );
  AOI21_X1 U9836 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n8133), .ZN(n10485) );
  NOR2_X1 U9837 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8134) );
  AOI21_X1 U9838 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n8134), .ZN(n10488) );
  AND2_X1 U9839 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n8135) );
  NOR2_X1 U9840 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n8135), .ZN(n10450) );
  INV_X1 U9841 ( .A(n10450), .ZN(n10451) );
  NAND3_X1 U9842 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U9843 ( .A1(n10453), .A2(n10452), .ZN(n10449) );
  NAND2_X1 U9844 ( .A1(n10451), .A2(n10449), .ZN(n10500) );
  NAND2_X1 U9845 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8136) );
  OAI21_X1 U9846 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n8136), .ZN(n10499) );
  NOR2_X1 U9847 ( .A1(n10500), .A2(n10499), .ZN(n10498) );
  AOI21_X1 U9848 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10498), .ZN(n10503) );
  NAND2_X1 U9849 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8137) );
  OAI21_X1 U9850 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n8137), .ZN(n10502) );
  NOR2_X1 U9851 ( .A1(n10503), .A2(n10502), .ZN(n10501) );
  AOI21_X1 U9852 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10501), .ZN(n10506) );
  NOR2_X1 U9853 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n8138) );
  AOI21_X1 U9854 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n8138), .ZN(n10505) );
  NAND2_X1 U9855 ( .A1(n10506), .A2(n10505), .ZN(n10504) );
  OAI21_X1 U9856 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10504), .ZN(n10487) );
  NAND2_X1 U9857 ( .A1(n10488), .A2(n10487), .ZN(n10486) );
  OAI21_X1 U9858 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10486), .ZN(n10484) );
  NAND2_X1 U9859 ( .A1(n10485), .A2(n10484), .ZN(n10483) );
  OAI21_X1 U9860 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10483), .ZN(n10493) );
  NAND2_X1 U9861 ( .A1(n10494), .A2(n10493), .ZN(n10492) );
  OAI21_X1 U9862 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10492), .ZN(n10496) );
  NAND2_X1 U9863 ( .A1(n10497), .A2(n10496), .ZN(n10495) );
  NAND2_X1 U9864 ( .A1(n8139), .A2(n10495), .ZN(n10490) );
  NAND2_X1 U9865 ( .A1(n10491), .A2(n10490), .ZN(n10489) );
  OAI21_X1 U9866 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10489), .ZN(n10481) );
  NAND2_X1 U9867 ( .A1(n10482), .A2(n10481), .ZN(n10480) );
  OAI21_X1 U9868 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10480), .ZN(n10478) );
  NAND2_X1 U9869 ( .A1(n10479), .A2(n10478), .ZN(n10477) );
  OAI21_X1 U9870 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10477), .ZN(n10475) );
  NAND2_X1 U9871 ( .A1(n10476), .A2(n10475), .ZN(n10474) );
  OAI21_X1 U9872 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10474), .ZN(n10472) );
  NAND2_X1 U9873 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  OAI21_X1 U9874 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10471), .ZN(n10469) );
  NAND2_X1 U9875 ( .A1(n10470), .A2(n10469), .ZN(n10468) );
  OAI21_X1 U9876 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10468), .ZN(n10466) );
  NAND2_X1 U9877 ( .A1(n10467), .A2(n10466), .ZN(n10465) );
  OAI21_X1 U9878 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10465), .ZN(n10463) );
  NAND2_X1 U9879 ( .A1(n10464), .A2(n10463), .ZN(n10462) );
  OAI21_X1 U9880 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10462), .ZN(n10460) );
  NAND2_X1 U9881 ( .A1(n10461), .A2(n10460), .ZN(n10459) );
  OAI21_X1 U9882 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10459), .ZN(n10456) );
  NOR2_X1 U9883 ( .A1(n10455), .A2(n10456), .ZN(n8140) );
  NAND2_X1 U9884 ( .A1(n10455), .A2(n10456), .ZN(n10454) );
  OAI21_X1 U9885 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n8140), .A(n10454), .ZN(
        n8142) );
  XNOR2_X1 U9886 ( .A(n4803), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8141) );
  XNOR2_X1 U9887 ( .A(n8142), .B(n8141), .ZN(ADD_1068_U4) );
  OR2_X1 U9888 ( .A1(n8143), .A2(n8151), .ZN(n8144) );
  NAND2_X1 U9889 ( .A1(n8145), .A2(n8144), .ZN(n10114) );
  XNOR2_X1 U9890 ( .A(n8184), .B(n10113), .ZN(n8146) );
  NAND2_X1 U9891 ( .A1(n8146), .A2(n10052), .ZN(n8148) );
  AOI22_X1 U9892 ( .A1(n9735), .A2(n10377), .B1(n10085), .B2(n9737), .ZN(n8147) );
  NAND2_X1 U9893 ( .A1(n8148), .A2(n8147), .ZN(n10116) );
  INV_X1 U9894 ( .A(n8149), .ZN(n8150) );
  AOI21_X1 U9895 ( .B1(n8177), .B2(n8488), .A(n8150), .ZN(n8152) );
  XNOR2_X1 U9896 ( .A(n8152), .B(n8151), .ZN(n8153) );
  NOR2_X1 U9897 ( .A1(n8153), .A2(n10392), .ZN(n10109) );
  AOI211_X1 U9898 ( .C1(n10195), .C2(n10114), .A(n10116), .B(n10109), .ZN(
        n8156) );
  AOI22_X1 U9899 ( .A1(n10113), .A2(n10159), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6794), .ZN(n8154) );
  OAI21_X1 U9900 ( .B1(n8156), .B2(n6794), .A(n8154), .ZN(P1_U3531) );
  AOI22_X1 U9901 ( .A1(n10113), .A2(n10232), .B1(P1_REG0_REG_9__SCAN_IN), .B2(
        n10403), .ZN(n8155) );
  OAI21_X1 U9902 ( .B1(n8156), .B2(n10403), .A(n8155), .ZN(P1_U3480) );
  NOR3_X1 U9903 ( .A1(n8159), .A2(n4554), .A3(n8158), .ZN(n8162) );
  INV_X1 U9904 ( .A(n8160), .ZN(n8161) );
  OAI21_X1 U9905 ( .B1(n8162), .B2(n8161), .A(n8882), .ZN(n8168) );
  NAND2_X1 U9906 ( .A1(n8902), .A2(n8920), .ZN(n8163) );
  NAND2_X1 U9907 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8926) );
  OAI211_X1 U9908 ( .C1(n8164), .C2(n8904), .A(n8163), .B(n8926), .ZN(n8165)
         );
  AOI21_X1 U9909 ( .B1(n8166), .B2(n8896), .A(n8165), .ZN(n8167) );
  OAI211_X1 U9910 ( .C1(n8169), .C2(n8852), .A(n8168), .B(n8167), .ZN(P2_U3161) );
  INV_X1 U9911 ( .A(n8178), .ZN(n8171) );
  NAND2_X1 U9912 ( .A1(n8171), .A2(n8170), .ZN(n8173) );
  OAI21_X1 U9913 ( .B1(n8174), .B2(n8173), .A(n8172), .ZN(n8189) );
  OAI22_X1 U9914 ( .A1(n8175), .A2(n10043), .B1(n8232), .B2(n10045), .ZN(n8182) );
  NAND2_X1 U9915 ( .A1(n8177), .A2(n8176), .ZN(n8179) );
  XNOR2_X1 U9916 ( .A(n8179), .B(n8178), .ZN(n8180) );
  NOR2_X1 U9917 ( .A1(n8180), .A2(n10392), .ZN(n8181) );
  AOI211_X1 U9918 ( .C1(n8189), .C2(n8183), .A(n8182), .B(n8181), .ZN(n10211)
         );
  AOI211_X1 U9919 ( .C1(n10209), .C2(n8185), .A(n10091), .B(n8184), .ZN(n10208) );
  INV_X1 U9920 ( .A(n8231), .ZN(n8186) );
  AOI22_X1 U9921 ( .A1(n10361), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8186), .B2(
        n10066), .ZN(n8187) );
  OAI21_X1 U9922 ( .B1(n10069), .B2(n8188), .A(n8187), .ZN(n8192) );
  INV_X1 U9923 ( .A(n8189), .ZN(n10213) );
  NOR2_X1 U9924 ( .A1(n10213), .A2(n8190), .ZN(n8191) );
  AOI211_X1 U9925 ( .C1(n10208), .C2(n10115), .A(n8192), .B(n8191), .ZN(n8193)
         );
  OAI21_X1 U9926 ( .B1(n10361), .B2(n10211), .A(n8193), .ZN(P1_U3285) );
  NAND2_X1 U9927 ( .A1(n8194), .A2(n8200), .ZN(n8195) );
  NAND3_X1 U9928 ( .A1(n8196), .A2(n9336), .A3(n8195), .ZN(n8198) );
  AOI22_X1 U9929 ( .A1(n8915), .A2(n9333), .B1(n9331), .B2(n8917), .ZN(n8197)
         );
  NAND2_X1 U9930 ( .A1(n8198), .A2(n8197), .ZN(n8289) );
  MUX2_X1 U9931 ( .A(n8289), .B(P2_REG0_REG_11__SCAN_IN), .S(n10441), .Z(n8203) );
  OAI21_X1 U9932 ( .B1(n8201), .B2(n8200), .A(n8199), .ZN(n8292) );
  INV_X1 U9933 ( .A(n8292), .ZN(n8204) );
  OAI22_X1 U9934 ( .A1(n8204), .A2(n9480), .B1(n8878), .B2(n9461), .ZN(n8202)
         );
  OR2_X1 U9935 ( .A1(n8203), .A2(n8202), .ZN(P2_U3423) );
  MUX2_X1 U9936 ( .A(n8289), .B(P2_REG1_REG_11__SCAN_IN), .S(n10446), .Z(n8206) );
  OAI22_X1 U9937 ( .A1(n8204), .A2(n9403), .B1(n8878), .B2(n9381), .ZN(n8205)
         );
  OR2_X1 U9938 ( .A1(n8206), .A2(n8205), .ZN(P2_U3470) );
  AOI211_X1 U9939 ( .C1(n10195), .C2(n8209), .A(n8208), .B(n8207), .ZN(n8212)
         );
  AOI22_X1 U9940 ( .A1(n9690), .A2(n10159), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n6794), .ZN(n8210) );
  OAI21_X1 U9941 ( .B1(n8212), .B2(n6794), .A(n8210), .ZN(P1_U3533) );
  AOI22_X1 U9942 ( .A1(n9690), .A2(n10232), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n10403), .ZN(n8211) );
  OAI21_X1 U9943 ( .B1(n8212), .B2(n10403), .A(n8211), .ZN(P1_U3486) );
  NAND2_X1 U9944 ( .A1(n8213), .A2(P2_U3893), .ZN(n8214) );
  OAI21_X1 U9945 ( .B1(P2_U3893), .B2(n5976), .A(n8214), .ZN(P2_U3522) );
  INV_X1 U9946 ( .A(n8215), .ZN(n8761) );
  MUX2_X1 U9947 ( .A(n8252), .B(n8216), .S(n9404), .Z(n8217) );
  OAI21_X1 U9948 ( .B1(n8761), .B2(n9381), .A(n8217), .ZN(P2_U3469) );
  OAI22_X1 U9949 ( .A1(n10415), .A2(n8761), .B1(n8755), .B2(n10417), .ZN(n8220) );
  MUX2_X1 U9950 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8218), .S(n10421), .Z(n8219) );
  AOI211_X1 U9951 ( .C1(n8221), .C2(n9283), .A(n8220), .B(n8219), .ZN(n8222)
         );
  INV_X1 U9952 ( .A(n8222), .ZN(P2_U3223) );
  INV_X1 U9953 ( .A(n8223), .ZN(n8306) );
  OAI222_X1 U9954 ( .A1(n9497), .A2(n8306), .B1(P2_U3151), .B2(n8225), .C1(
        n8224), .C2(n9502), .ZN(P2_U3274) );
  OR2_X1 U9955 ( .A1(n9536), .A2(n8227), .ZN(n9633) );
  NAND2_X1 U9956 ( .A1(n9536), .A2(n8227), .ZN(n8228) );
  NAND2_X1 U9957 ( .A1(n9633), .A2(n8228), .ZN(n8229) );
  NOR2_X1 U9958 ( .A1(n8229), .A2(n8230), .ZN(n9636) );
  AOI21_X1 U9959 ( .B1(n8230), .B2(n8229), .A(n9636), .ZN(n8237) );
  NAND2_X1 U9960 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9809) );
  INV_X1 U9961 ( .A(n9809), .ZN(n8234) );
  OAI22_X1 U9962 ( .A1(n8232), .A2(n9719), .B1(n9718), .B2(n8231), .ZN(n8233)
         );
  AOI211_X1 U9963 ( .C1(n9695), .C2(n9738), .A(n8234), .B(n8233), .ZN(n8236)
         );
  NAND2_X1 U9964 ( .A1(n10209), .A2(n9722), .ZN(n8235) );
  OAI211_X1 U9965 ( .C1(n8237), .C2(n9724), .A(n8236), .B(n8235), .ZN(P1_U3221) );
  INV_X1 U9966 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8240) );
  INV_X1 U9967 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8242) );
  XNOR2_X1 U9968 ( .A(n8253), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n8950) );
  INV_X1 U9969 ( .A(n8238), .ZN(n8239) );
  INV_X1 U9970 ( .A(n8347), .ZN(n8345) );
  AOI21_X1 U9971 ( .B1(n8240), .B2(n8239), .A(n8345), .ZN(n8260) );
  NAND2_X1 U9972 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8871) );
  OAI21_X1 U9973 ( .B1(n9131), .B2(n8241), .A(n8871), .ZN(n8250) );
  MUX2_X1 U9974 ( .A(n8242), .B(n8252), .S(n4279), .Z(n8243) );
  NAND2_X1 U9975 ( .A1(n8253), .A2(n8243), .ZN(n8244) );
  OAI21_X1 U9976 ( .B1(n8253), .B2(n8243), .A(n8244), .ZN(n8958) );
  AOI21_X1 U9977 ( .B1(n8960), .B2(n8959), .A(n8958), .ZN(n8962) );
  INV_X1 U9978 ( .A(n8244), .ZN(n8245) );
  NOR2_X1 U9979 ( .A1(n8962), .A2(n8245), .ZN(n8247) );
  MUX2_X1 U9980 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n4279), .Z(n8328) );
  XOR2_X1 U9981 ( .A(n8328), .B(n8331), .Z(n8246) );
  NOR2_X1 U9982 ( .A1(n8247), .A2(n8246), .ZN(n8329) );
  AOI21_X1 U9983 ( .B1(n8247), .B2(n8246), .A(n8329), .ZN(n8248) );
  NOR2_X1 U9984 ( .A1(n8248), .A2(n9140), .ZN(n8249) );
  AOI211_X1 U9985 ( .C1(n9142), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n8250), .B(
        n8249), .ZN(n8259) );
  INV_X1 U9986 ( .A(n8251), .ZN(n8963) );
  XNOR2_X1 U9987 ( .A(n8253), .B(n8252), .ZN(n8964) );
  AOI21_X1 U9988 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n8949), .A(n8967), .ZN(
        n8254) );
  NOR2_X1 U9989 ( .A1(n8254), .A2(n8331), .ZN(n8335) );
  OAI21_X1 U9990 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n8256), .A(n8337), .ZN(
        n8257) );
  NAND2_X1 U9991 ( .A1(n8257), .A2(n9126), .ZN(n8258) );
  OAI211_X1 U9992 ( .C1(n8260), .C2(n9144), .A(n8259), .B(n8258), .ZN(P2_U3193) );
  INV_X1 U9993 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8262) );
  OAI222_X1 U9994 ( .A1(n10259), .A2(n8262), .B1(n10262), .B2(n8261), .C1(
        n8665), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI211_X1 U9995 ( .C1(n8265), .C2(n8264), .A(n8263), .B(n8882), .ZN(n8271)
         );
  NAND2_X1 U9996 ( .A1(n8902), .A2(n8919), .ZN(n8267) );
  OAI211_X1 U9997 ( .C1(n8751), .C2(n8904), .A(n8267), .B(n8266), .ZN(n8268)
         );
  AOI21_X1 U9998 ( .B1(n8269), .B2(n8896), .A(n8268), .ZN(n8270) );
  OAI211_X1 U9999 ( .C1(n8272), .C2(n8852), .A(n8271), .B(n8270), .ZN(P2_U3171) );
  INV_X1 U10000 ( .A(n8273), .ZN(n8275) );
  INV_X1 U10001 ( .A(n8278), .ZN(n8613) );
  AOI21_X1 U10002 ( .B1(n8078), .B2(n8498), .A(n8613), .ZN(n8274) );
  NOR2_X1 U10003 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  OAI222_X1 U10004 ( .A1(n10045), .A2(n9716), .B1(n10043), .B2(n9682), .C1(
        n8276), .C2(n10392), .ZN(n8380) );
  INV_X1 U10005 ( .A(n8380), .ZN(n8288) );
  OAI21_X1 U10006 ( .B1(n8279), .B2(n8278), .A(n8277), .ZN(n8382) );
  INV_X1 U10007 ( .A(n8280), .ZN(n8282) );
  AOI211_X1 U10008 ( .C1(n8283), .C2(n8282), .A(n10091), .B(n8281), .ZN(n8381)
         );
  NAND2_X1 U10009 ( .A1(n8381), .A2(n10115), .ZN(n8285) );
  AOI22_X1 U10010 ( .A1(n10361), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9660), 
        .B2(n10066), .ZN(n8284) );
  OAI211_X1 U10011 ( .C1(n9666), .C2(n10069), .A(n8285), .B(n8284), .ZN(n8286)
         );
  AOI21_X1 U10012 ( .B1(n10371), .B2(n8382), .A(n8286), .ZN(n8287) );
  OAI21_X1 U10013 ( .B1(n8288), .B2(n10361), .A(n8287), .ZN(P1_U3280) );
  OAI22_X1 U10014 ( .A1(n10415), .A2(n8878), .B1(n8870), .B2(n10417), .ZN(
        n8291) );
  MUX2_X1 U10015 ( .A(n8289), .B(P2_REG2_REG_11__SCAN_IN), .S(n10413), .Z(
        n8290) );
  AOI211_X1 U10016 ( .C1(n9283), .C2(n8292), .A(n8291), .B(n8290), .ZN(n8293)
         );
  INV_X1 U10017 ( .A(n8293), .ZN(P2_U3222) );
  XOR2_X1 U10018 ( .A(n8294), .B(n8298), .Z(n8295) );
  AOI222_X1 U10019 ( .A1(n9336), .A2(n8295), .B1(n9332), .B2(n9333), .C1(n8916), .C2(n9331), .ZN(n8309) );
  MUX2_X1 U10020 ( .A(n8296), .B(n8309), .S(n10440), .Z(n8300) );
  XOR2_X1 U10021 ( .A(n8297), .B(n8298), .Z(n8308) );
  AOI22_X1 U10022 ( .A1(n8308), .A2(n9486), .B1(n9485), .B2(n8311), .ZN(n8299)
         );
  NAND2_X1 U10023 ( .A1(n8300), .A2(n8299), .ZN(P2_U3426) );
  MUX2_X1 U10024 ( .A(n8336), .B(n8309), .S(n9404), .Z(n8302) );
  AOI22_X1 U10025 ( .A1(n8308), .A2(n9407), .B1(n9406), .B2(n8311), .ZN(n8301)
         );
  NAND2_X1 U10026 ( .A1(n8302), .A2(n8301), .ZN(P2_U3471) );
  INV_X1 U10027 ( .A(n8303), .ZN(n8393) );
  OAI222_X1 U10028 ( .A1(n9502), .A2(n8305), .B1(n9497), .B2(n8393), .C1(n8304), .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U10029 ( .A1(n10259), .A2(n8307), .B1(n10262), .B2(n8306), .C1(
        n8600), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U10030 ( .A(n8308), .ZN(n8314) );
  INV_X1 U10031 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8985) );
  MUX2_X1 U10032 ( .A(n8985), .B(n8309), .S(n10421), .Z(n8313) );
  INV_X1 U10033 ( .A(n8310), .ZN(n8793) );
  AOI22_X1 U10034 ( .A1(n8311), .A2(n9325), .B1(n9341), .B2(n8793), .ZN(n8312)
         );
  OAI211_X1 U10035 ( .C1(n8314), .C2(n9344), .A(n8313), .B(n8312), .ZN(
        P2_U3221) );
  NAND2_X1 U10036 ( .A1(n8315), .A2(n8316), .ZN(n8317) );
  NAND2_X1 U10037 ( .A1(n9315), .A2(n8317), .ZN(n8320) );
  NAND2_X1 U10038 ( .A1(n9320), .A2(n9333), .ZN(n8318) );
  OAI21_X1 U10039 ( .B1(n8873), .B2(n9296), .A(n8318), .ZN(n8319) );
  AOI21_X1 U10040 ( .B1(n8320), .B2(n9336), .A(n8319), .ZN(n8367) );
  MUX2_X1 U10041 ( .A(n8367), .B(n8321), .S(n10441), .Z(n8325) );
  XNOR2_X1 U10042 ( .A(n8323), .B(n8322), .ZN(n8371) );
  AOI22_X1 U10043 ( .A1(n8371), .A2(n9486), .B1(n9485), .B2(n8854), .ZN(n8324)
         );
  NAND2_X1 U10044 ( .A1(n8325), .A2(n8324), .ZN(P2_U3429) );
  MUX2_X1 U10045 ( .A(n8367), .B(n8976), .S(n10446), .Z(n8327) );
  AOI22_X1 U10046 ( .A1(n8371), .A2(n9407), .B1(n9406), .B2(n8854), .ZN(n8326)
         );
  NAND2_X1 U10047 ( .A1(n8327), .A2(n8326), .ZN(P2_U3472) );
  INV_X1 U10048 ( .A(n8328), .ZN(n8330) );
  AOI21_X1 U10049 ( .B1(n8331), .B2(n8330), .A(n8329), .ZN(n8979) );
  MUX2_X1 U10050 ( .A(n8985), .B(n8336), .S(n4279), .Z(n8332) );
  NOR2_X1 U10051 ( .A1(n8986), .A2(n8332), .ZN(n8977) );
  NAND2_X1 U10052 ( .A1(n8986), .A2(n8332), .ZN(n8978) );
  INV_X1 U10053 ( .A(n8978), .ZN(n8333) );
  NOR2_X1 U10054 ( .A1(n8977), .A2(n8333), .ZN(n8334) );
  XNOR2_X1 U10055 ( .A(n8979), .B(n8334), .ZN(n8355) );
  NAND2_X1 U10056 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8787) );
  OAI21_X1 U10057 ( .B1(n9131), .B2(n8972), .A(n8787), .ZN(n8343) );
  INV_X1 U10058 ( .A(n8335), .ZN(n8338) );
  XNOR2_X1 U10059 ( .A(n8986), .B(n8336), .ZN(n8339) );
  INV_X1 U10060 ( .A(n8971), .ZN(n8341) );
  NAND3_X1 U10061 ( .A1(n8337), .A2(n8339), .A3(n8338), .ZN(n8340) );
  AOI21_X1 U10062 ( .B1(n8341), .B2(n8340), .A(n9037), .ZN(n8342) );
  AOI211_X1 U10063 ( .C1(n9142), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n8343), .B(
        n8342), .ZN(n8354) );
  INV_X1 U10064 ( .A(n8346), .ZN(n8344) );
  XNOR2_X1 U10065 ( .A(n8986), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8348) );
  NOR3_X1 U10066 ( .A1(n8345), .A2(n8344), .A3(n8348), .ZN(n8352) );
  NAND2_X1 U10067 ( .A1(n8347), .A2(n8346), .ZN(n8349) );
  INV_X1 U10068 ( .A(n8988), .ZN(n8351) );
  OAI21_X1 U10069 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8353) );
  OAI211_X1 U10070 ( .C1(n9140), .C2(n8355), .A(n8354), .B(n8353), .ZN(
        P2_U3194) );
  NAND2_X1 U10071 ( .A1(n8529), .A2(n8517), .ZN(n8614) );
  XNOR2_X1 U10072 ( .A(n8356), .B(n8525), .ZN(n8357) );
  AOI222_X1 U10073 ( .A1(n9732), .A2(n10085), .B1(n10087), .B2(n8357), .C1(
        n10073), .C2(n10377), .ZN(n10200) );
  INV_X1 U10074 ( .A(n8281), .ZN(n8359) );
  INV_X1 U10075 ( .A(n10092), .ZN(n8358) );
  AOI211_X1 U10076 ( .C1(n10198), .C2(n8359), .A(n10091), .B(n8358), .ZN(
        n10197) );
  INV_X1 U10077 ( .A(n9518), .ZN(n8360) );
  AOI22_X1 U10078 ( .A1(n10361), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8360), 
        .B2(n10066), .ZN(n8361) );
  OAI21_X1 U10079 ( .B1(n8362), .B2(n10069), .A(n8361), .ZN(n8365) );
  XNOR2_X1 U10080 ( .A(n8363), .B(n8525), .ZN(n10201) );
  NOR2_X1 U10081 ( .A1(n10201), .A2(n10079), .ZN(n8364) );
  AOI211_X1 U10082 ( .C1(n10197), .C2(n10115), .A(n8365), .B(n8364), .ZN(n8366) );
  OAI21_X1 U10083 ( .B1(n10200), .B2(n10361), .A(n8366), .ZN(P1_U3279) );
  INV_X1 U10084 ( .A(n8367), .ZN(n8370) );
  OAI22_X1 U10085 ( .A1(n8368), .A2(n9337), .B1(n8851), .B2(n10417), .ZN(n8369) );
  OAI21_X1 U10086 ( .B1(n8370), .B2(n8369), .A(n10421), .ZN(n8373) );
  AOI22_X1 U10087 ( .A1(n8371), .A2(n9283), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10413), .ZN(n8372) );
  NAND2_X1 U10088 ( .A1(n8373), .A2(n8372), .ZN(P2_U3220) );
  INV_X1 U10089 ( .A(n8374), .ZN(n8379) );
  AOI21_X1 U10090 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n8441), .A(n8375), .ZN(
        n8376) );
  OAI21_X1 U10091 ( .B1(n8379), .B2(n10251), .A(n8376), .ZN(P1_U3332) );
  NAND2_X1 U10092 ( .A1(n9495), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8377) );
  OAI211_X1 U10093 ( .C1(n8379), .C2(n9497), .A(n8378), .B(n8377), .ZN(
        P2_U3272) );
  AOI211_X1 U10094 ( .C1(n10195), .C2(n8382), .A(n8381), .B(n8380), .ZN(n8385)
         );
  MUX2_X1 U10095 ( .A(n8383), .B(n8385), .S(n10405), .Z(n8384) );
  OAI21_X1 U10096 ( .B1(n9666), .B2(n6800), .A(n8384), .ZN(P1_U3492) );
  MUX2_X1 U10097 ( .A(n8386), .B(n8385), .S(n10408), .Z(n8387) );
  OAI21_X1 U10098 ( .B1(n9666), .B2(n6796), .A(n8387), .ZN(P1_U3535) );
  INV_X1 U10099 ( .A(n8388), .ZN(n10247) );
  INV_X1 U10100 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8389) );
  OAI222_X1 U10101 ( .A1(n9497), .A2(n10247), .B1(n8390), .B2(P2_U3151), .C1(
        n8389), .C2(n9502), .ZN(P2_U3266) );
  INV_X1 U10102 ( .A(n8415), .ZN(n8397) );
  OAI222_X1 U10103 ( .A1(n9502), .A2(n8392), .B1(n9497), .B2(n8397), .C1(
        P2_U3151), .C2(n8391), .ZN(P2_U3265) );
  OAI222_X1 U10104 ( .A1(n10259), .A2(n8394), .B1(n10262), .B2(n8393), .C1(
        P1_U3086), .C2(n8591), .ZN(P1_U3333) );
  INV_X1 U10105 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8396) );
  OAI222_X1 U10106 ( .A1(P1_U3086), .A2(n8395), .B1(n10262), .B2(n8397), .C1(
        n8396), .C2(n10259), .ZN(P1_U3325) );
  NAND2_X1 U10107 ( .A1(n10127), .A2(n9897), .ZN(n8401) );
  NAND3_X1 U10108 ( .A1(n4337), .A2(n10052), .A3(n8401), .ZN(n8410) );
  NAND2_X1 U10109 ( .A1(n8404), .A2(n8403), .ZN(n8406) );
  OAI22_X1 U10110 ( .A1(n8562), .A2(n10045), .B1(n9916), .B2(n10043), .ZN(
        n8405) );
  INV_X1 U10111 ( .A(n8407), .ZN(n8412) );
  AOI22_X1 U10112 ( .A1(n9509), .A2(n10066), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10361), .ZN(n8409) );
  NAND2_X1 U10113 ( .A1(n10127), .A2(n10366), .ZN(n8408) );
  OAI211_X1 U10114 ( .C1(n8410), .C2(n10369), .A(n8409), .B(n8408), .ZN(n8411)
         );
  AOI21_X1 U10115 ( .B1(n8412), .B2(n10386), .A(n8411), .ZN(n8413) );
  OAI21_X1 U10116 ( .B1(n10079), .B2(n8414), .A(n8413), .ZN(P1_U3266) );
  NAND2_X1 U10117 ( .A1(n8415), .A2(n6514), .ZN(n8417) );
  NAND2_X1 U10118 ( .A1(n6593), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10119 ( .A1(n6593), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8421) );
  XNOR2_X1 U10120 ( .A(n9868), .B(n8581), .ZN(n8423) );
  NOR2_X1 U10121 ( .A1(n10386), .A2(n8424), .ZN(n8426) );
  NAND2_X1 U10122 ( .A1(n8425), .A2(n8656), .ZN(n10121) );
  NOR2_X1 U10123 ( .A1(n10361), .A2(n10121), .ZN(n9870) );
  AOI211_X1 U10124 ( .C1(n8731), .C2(n10366), .A(n8426), .B(n9870), .ZN(n8427)
         );
  OAI21_X1 U10125 ( .B1(n8452), .B2(n10369), .A(n8427), .ZN(P1_U3263) );
  INV_X1 U10126 ( .A(n8428), .ZN(n9492) );
  OAI222_X1 U10127 ( .A1(n10259), .A2(n8430), .B1(n10251), .B2(n9492), .C1(
        n8429), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U10128 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8432) );
  NAND3_X1 U10129 ( .A1(n8432), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8437) );
  INV_X1 U10130 ( .A(n8433), .ZN(n8440) );
  NAND2_X1 U10131 ( .A1(n8440), .A2(n8434), .ZN(n8436) );
  NAND2_X1 U10132 ( .A1(n9495), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8435) );
  OAI211_X1 U10133 ( .C1(n8431), .C2(n8437), .A(n8436), .B(n8435), .ZN(
        P2_U3264) );
  NAND3_X1 U10134 ( .A1(n8438), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10135 ( .A1(n8440), .A2(n8439), .ZN(n8443) );
  NAND2_X1 U10136 ( .A1(n8441), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8442) );
  OAI211_X1 U10137 ( .C1(n8445), .C2(n8444), .A(n8443), .B(n8442), .ZN(
        P1_U3324) );
  INV_X1 U10138 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8448) );
  AND2_X1 U10139 ( .A1(n8446), .A2(n9500), .ZN(n8447) );
  AOI22_X1 U10140 ( .A1(n8449), .A2(n8448), .B1(n8447), .B2(n5758), .ZN(
        P2_U3377) );
  INV_X1 U10141 ( .A(n8450), .ZN(n10257) );
  OAI222_X1 U10142 ( .A1(n9497), .A2(n10257), .B1(P2_U3151), .B2(n5758), .C1(
        n8451), .C2(n9502), .ZN(P2_U3270) );
  NAND2_X1 U10143 ( .A1(n8452), .A2(n10121), .ZN(n8729) );
  MUX2_X1 U10144 ( .A(n8729), .B(P1_REG1_REG_31__SCAN_IN), .S(n6794), .Z(n8453) );
  AOI21_X1 U10145 ( .B1(n10159), .B2(n8731), .A(n8453), .ZN(n8454) );
  INV_X1 U10146 ( .A(n8454), .ZN(P1_U3553) );
  NAND2_X1 U10147 ( .A1(n8731), .A2(n9726), .ZN(n8583) );
  MUX2_X1 U10148 ( .A(n8707), .B(n8654), .S(n8582), .Z(n8455) );
  OAI21_X1 U10149 ( .B1(n8583), .B2(n10216), .A(n8455), .ZN(n8579) );
  AND2_X1 U10150 ( .A1(n8701), .A2(n8582), .ZN(n8556) );
  MUX2_X1 U10151 ( .A(n8543), .B(n8640), .S(n4285), .Z(n8547) );
  NAND2_X1 U10152 ( .A1(n10004), .A2(n9982), .ZN(n8542) );
  NAND2_X1 U10153 ( .A1(n8542), .A2(n10016), .ZN(n8456) );
  NAND2_X1 U10154 ( .A1(n8456), .A2(n8582), .ZN(n8457) );
  NAND3_X1 U10155 ( .A1(n8457), .A2(n8461), .A3(n8460), .ZN(n8459) );
  NAND3_X1 U10156 ( .A1(n8542), .A2(n9731), .A3(n8582), .ZN(n8458) );
  NAND2_X1 U10157 ( .A1(n8459), .A2(n8458), .ZN(n8541) );
  NAND2_X1 U10158 ( .A1(n8460), .A2(n8534), .ZN(n8697) );
  OAI21_X1 U10159 ( .B1(n4285), .B2(n8697), .A(n8541), .ZN(n8462) );
  AND2_X1 U10160 ( .A1(n8640), .A2(n8461), .ZN(n8636) );
  NAND2_X1 U10161 ( .A1(n8462), .A2(n8636), .ZN(n8464) );
  NAND3_X1 U10162 ( .A1(n8696), .A2(n4285), .A3(n8537), .ZN(n8463) );
  OAI211_X1 U10163 ( .C1(n8541), .C2(n8582), .A(n8464), .B(n8463), .ZN(n8546)
         );
  NAND2_X1 U10164 ( .A1(n8467), .A2(n8471), .ZN(n8671) );
  INV_X1 U10165 ( .A(n8671), .ZN(n8465) );
  OAI211_X1 U10166 ( .C1(n8468), .C2(n4286), .A(n8467), .B(n8668), .ZN(n8474)
         );
  INV_X1 U10167 ( .A(n8480), .ZN(n8470) );
  NOR2_X1 U10168 ( .A1(n8470), .A2(n8469), .ZN(n8473) );
  INV_X1 U10169 ( .A(n8471), .ZN(n8472) );
  AOI21_X1 U10170 ( .B1(n8474), .B2(n8473), .A(n8472), .ZN(n8475) );
  INV_X1 U10171 ( .A(n8481), .ZN(n8479) );
  INV_X1 U10172 ( .A(n8674), .ZN(n8477) );
  NOR2_X1 U10173 ( .A1(n8478), .A2(n8477), .ZN(n8484) );
  NAND2_X1 U10174 ( .A1(n8481), .A2(n8480), .ZN(n8675) );
  INV_X1 U10175 ( .A(n8675), .ZN(n8482) );
  NAND2_X1 U10176 ( .A1(n8483), .A2(n8482), .ZN(n8485) );
  NAND2_X1 U10177 ( .A1(n8485), .A2(n8484), .ZN(n8487) );
  INV_X1 U10178 ( .A(n8488), .ZN(n8489) );
  NAND2_X1 U10179 ( .A1(n8497), .A2(n8491), .ZN(n8492) );
  MUX2_X1 U10180 ( .A(n8493), .B(n8492), .S(n4285), .Z(n8494) );
  INV_X1 U10181 ( .A(n8494), .ZN(n8495) );
  NAND2_X1 U10182 ( .A1(n8496), .A2(n8495), .ZN(n8502) );
  INV_X1 U10183 ( .A(n8506), .ZN(n8679) );
  AOI21_X1 U10184 ( .B1(n8502), .B2(n8497), .A(n8679), .ZN(n8500) );
  NAND2_X1 U10185 ( .A1(n8508), .A2(n8503), .ZN(n8682) );
  NAND2_X1 U10186 ( .A1(n8498), .A2(n8505), .ZN(n8686) );
  INV_X1 U10187 ( .A(n8686), .ZN(n8499) );
  OAI211_X1 U10188 ( .C1(n8500), .C2(n8682), .A(n8499), .B(n8582), .ZN(n8515)
         );
  NAND2_X1 U10189 ( .A1(n8502), .A2(n8501), .ZN(n8504) );
  NAND2_X1 U10190 ( .A1(n8504), .A2(n8503), .ZN(n8507) );
  NAND3_X1 U10191 ( .A1(n8507), .A2(n8506), .A3(n8505), .ZN(n8509) );
  NAND4_X1 U10192 ( .A1(n8509), .A2(n4285), .A3(n8508), .A4(n8684), .ZN(n8514)
         );
  NOR2_X1 U10193 ( .A1(n9733), .A2(n4285), .ZN(n8511) );
  OAI21_X1 U10194 ( .B1(n9682), .B2(n8582), .A(n8512), .ZN(n8510) );
  OAI21_X1 U10195 ( .B1(n8512), .B2(n8511), .A(n8510), .ZN(n8513) );
  NAND3_X1 U10196 ( .A1(n8515), .A2(n8514), .A3(n8513), .ZN(n8524) );
  AND2_X1 U10197 ( .A1(n8529), .A2(n8523), .ZN(n8689) );
  INV_X1 U10198 ( .A(n8689), .ZN(n8516) );
  AOI21_X1 U10199 ( .B1(n8524), .B2(n8685), .A(n8516), .ZN(n8518) );
  NAND2_X1 U10200 ( .A1(n8520), .A2(n8517), .ZN(n8688) );
  INV_X1 U10201 ( .A(n8520), .ZN(n8521) );
  NAND3_X1 U10202 ( .A1(n8528), .A2(n8521), .A3(n8582), .ZN(n8532) );
  INV_X1 U10203 ( .A(n8527), .ZN(n8522) );
  NAND2_X1 U10204 ( .A1(n8524), .A2(n8523), .ZN(n8526) );
  NAND3_X1 U10205 ( .A1(n8526), .A2(n8525), .A3(n8685), .ZN(n8531) );
  NAND2_X1 U10206 ( .A1(n8528), .A2(n8527), .ZN(n8691) );
  INV_X1 U10207 ( .A(n8691), .ZN(n8530) );
  AND2_X1 U10208 ( .A1(n8534), .A2(n8533), .ZN(n8695) );
  INV_X1 U10209 ( .A(n8695), .ZN(n8535) );
  NAND2_X1 U10210 ( .A1(n8535), .A2(n4285), .ZN(n8539) );
  NAND2_X1 U10211 ( .A1(n8537), .A2(n8536), .ZN(n8693) );
  NAND2_X1 U10212 ( .A1(n8693), .A2(n8582), .ZN(n8538) );
  NAND4_X1 U10213 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(n8545)
         );
  NAND2_X1 U10214 ( .A1(n8543), .A2(n8542), .ZN(n8641) );
  NAND2_X1 U10215 ( .A1(n8641), .A2(n4285), .ZN(n8544) );
  NAND2_X1 U10216 ( .A1(n9929), .A2(n8548), .ZN(n8643) );
  NAND2_X1 U10217 ( .A1(n8550), .A2(n8549), .ZN(n8630) );
  MUX2_X1 U10218 ( .A(n8643), .B(n8630), .S(n4285), .Z(n8552) );
  INV_X1 U10219 ( .A(n9940), .ZN(n9930) );
  MUX2_X1 U10220 ( .A(n9929), .B(n8550), .S(n8582), .Z(n8551) );
  MUX2_X1 U10221 ( .A(n8645), .B(n8632), .S(n4285), .Z(n8553) );
  INV_X1 U10222 ( .A(n8572), .ZN(n8648) );
  OAI211_X1 U10223 ( .C1(n8574), .C2(n8648), .A(n8647), .B(n8635), .ZN(n8554)
         );
  NAND4_X1 U10224 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n8571)
         );
  NAND2_X1 U10225 ( .A1(n9906), .A2(n8582), .ZN(n8563) );
  OAI22_X1 U10226 ( .A1(n10127), .A2(n8563), .B1(n8562), .B2(n4285), .ZN(n8558) );
  NAND2_X1 U10227 ( .A1(n6695), .A2(n8558), .ZN(n8570) );
  AND2_X1 U10228 ( .A1(n8559), .A2(n4285), .ZN(n8564) );
  NAND2_X1 U10229 ( .A1(n10127), .A2(n8564), .ZN(n8560) );
  OAI21_X1 U10230 ( .B1(n8582), .B2(n9728), .A(n8560), .ZN(n8561) );
  NAND2_X1 U10231 ( .A1(n9890), .A2(n8561), .ZN(n8569) );
  NOR2_X1 U10232 ( .A1(n8563), .A2(n8562), .ZN(n8567) );
  INV_X1 U10233 ( .A(n8564), .ZN(n8565) );
  OAI21_X1 U10234 ( .B1(n9728), .B2(n8565), .A(n10127), .ZN(n8566) );
  OAI21_X1 U10235 ( .B1(n8567), .B2(n10127), .A(n8566), .ZN(n8568) );
  AND2_X1 U10236 ( .A1(n8647), .A2(n4285), .ZN(n8576) );
  INV_X1 U10237 ( .A(n8635), .ZN(n8573) );
  OAI211_X1 U10238 ( .C1(n8574), .C2(n8573), .A(n8701), .B(n8572), .ZN(n8575)
         );
  NAND4_X1 U10239 ( .A1(n8653), .A2(n8576), .A3(n8705), .A4(n8575), .ZN(n8577)
         );
  AOI21_X1 U10240 ( .B1(n9726), .B2(n8656), .A(n8418), .ZN(n8578) );
  INV_X1 U10241 ( .A(n9726), .ZN(n8629) );
  OR2_X1 U10242 ( .A1(n10216), .A2(n8629), .ZN(n8710) );
  INV_X1 U10243 ( .A(n8710), .ZN(n8580) );
  NAND3_X1 U10244 ( .A1(n8580), .A2(n4285), .A3(n8656), .ZN(n8585) );
  NAND2_X1 U10245 ( .A1(n8581), .A2(n8656), .ZN(n8713) );
  NAND3_X1 U10246 ( .A1(n8583), .A2(n8582), .A3(n10216), .ZN(n8584) );
  INV_X1 U10247 ( .A(n8592), .ZN(n8586) );
  INV_X1 U10248 ( .A(n8656), .ZN(n8657) );
  INV_X1 U10249 ( .A(n8587), .ZN(n8589) );
  NOR2_X1 U10250 ( .A1(n8663), .A2(n8588), .ZN(n8721) );
  OAI211_X1 U10251 ( .C1(n8713), .C2(n8590), .A(n8589), .B(n8721), .ZN(n8727)
         );
  AOI21_X1 U10252 ( .B1(n8592), .B2(n8627), .A(n8591), .ZN(n8720) );
  AND2_X1 U10253 ( .A1(n9865), .A2(n6650), .ZN(n8664) );
  NAND2_X1 U10254 ( .A1(n8664), .A2(n4914), .ZN(n8719) );
  INV_X1 U10255 ( .A(n8593), .ZN(n9875) );
  INV_X1 U10256 ( .A(n8594), .ZN(n8681) );
  INV_X1 U10257 ( .A(n8595), .ZN(n8597) );
  NAND2_X1 U10258 ( .A1(n8597), .A2(n8596), .ZN(n8610) );
  AND2_X1 U10259 ( .A1(n9745), .A2(n10381), .ZN(n8667) );
  NOR2_X1 U10260 ( .A1(n8598), .A2(n8667), .ZN(n10391) );
  INV_X1 U10261 ( .A(n8599), .ZN(n8602) );
  AND4_X1 U10262 ( .A1(n10391), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n8607)
         );
  INV_X1 U10263 ( .A(n8603), .ZN(n8606) );
  NAND4_X1 U10264 ( .A1(n8607), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(n8608)
         );
  NOR4_X1 U10265 ( .A1(n8611), .A2(n8610), .A3(n8609), .A4(n8608), .ZN(n8612)
         );
  NAND3_X1 U10266 ( .A1(n8613), .A2(n8681), .A3(n8612), .ZN(n8615) );
  NOR2_X1 U10267 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NAND3_X1 U10268 ( .A1(n10072), .A2(n10083), .A3(n8616), .ZN(n8617) );
  NOR3_X1 U10269 ( .A1(n10028), .A2(n8618), .A3(n8617), .ZN(n8620) );
  INV_X1 U10270 ( .A(n8619), .ZN(n10000) );
  AND4_X1 U10271 ( .A1(n9981), .A2(n10019), .A3(n8620), .A4(n10000), .ZN(n8621) );
  NAND3_X1 U10272 ( .A1(n9954), .A2(n9971), .A3(n8621), .ZN(n8622) );
  NOR2_X1 U10273 ( .A1(n9940), .A2(n8622), .ZN(n8623) );
  NAND4_X1 U10274 ( .A1(n8624), .A2(n6579), .A3(n9905), .A4(n8623), .ZN(n8625)
         );
  NOR2_X1 U10275 ( .A1(n8626), .A2(n8625), .ZN(n8628) );
  NAND2_X1 U10276 ( .A1(n10216), .A2(n8629), .ZN(n8706) );
  NAND2_X1 U10277 ( .A1(n8630), .A2(n9929), .ZN(n8631) );
  NAND2_X1 U10278 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  NAND2_X1 U10279 ( .A1(n8633), .A2(n8645), .ZN(n8634) );
  NAND2_X1 U10280 ( .A1(n8635), .A2(n8634), .ZN(n8644) );
  INV_X1 U10281 ( .A(n8644), .ZN(n8637) );
  NAND3_X1 U10282 ( .A1(n8647), .A2(n8637), .A3(n8636), .ZN(n8666) );
  INV_X1 U10283 ( .A(n8638), .ZN(n8639) );
  OAI21_X1 U10284 ( .B1(n8666), .B2(n8639), .A(n8701), .ZN(n8652) );
  AND2_X1 U10285 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  NOR2_X1 U10286 ( .A1(n8643), .A2(n8642), .ZN(n8646) );
  AOI21_X1 U10287 ( .B1(n8646), .B2(n8645), .A(n8644), .ZN(n8649) );
  OAI211_X1 U10288 ( .C1(n8649), .C2(n8648), .A(n8705), .B(n8647), .ZN(n8650)
         );
  NAND2_X1 U10289 ( .A1(n8651), .A2(n8650), .ZN(n8703) );
  AOI21_X1 U10290 ( .B1(n8705), .B2(n8652), .A(n8703), .ZN(n8655) );
  NAND2_X1 U10291 ( .A1(n8654), .A2(n8653), .ZN(n8708) );
  OAI21_X1 U10292 ( .B1(n8655), .B2(n8708), .A(n8706), .ZN(n8659) );
  OAI21_X1 U10293 ( .B1(n8418), .B2(n8656), .A(n8707), .ZN(n8658) );
  OAI22_X1 U10294 ( .A1(n8659), .A2(n8658), .B1(n8657), .B2(n8710), .ZN(n8661)
         );
  AOI211_X1 U10295 ( .C1(n8661), .C2(n8713), .A(n8712), .B(n8660), .ZN(n8662)
         );
  NAND2_X1 U10296 ( .A1(n8665), .A2(n9865), .ZN(n10382) );
  INV_X1 U10297 ( .A(n8666), .ZN(n8700) );
  NAND2_X1 U10298 ( .A1(n6319), .A2(n4437), .ZN(n8670) );
  INV_X1 U10299 ( .A(n8667), .ZN(n8669) );
  NAND4_X1 U10300 ( .A1(n8670), .A2(n4914), .A3(n8669), .A4(n8668), .ZN(n8672)
         );
  AOI21_X1 U10301 ( .B1(n8673), .B2(n8672), .A(n8671), .ZN(n8676) );
  OAI21_X1 U10302 ( .B1(n8676), .B2(n8675), .A(n8674), .ZN(n8680) );
  INV_X1 U10303 ( .A(n8677), .ZN(n8678) );
  AOI211_X1 U10304 ( .C1(n8681), .C2(n8680), .A(n8679), .B(n8678), .ZN(n8683)
         );
  NOR2_X1 U10305 ( .A1(n8683), .A2(n8682), .ZN(n8687) );
  OAI211_X1 U10306 ( .C1(n8687), .C2(n8686), .A(n8685), .B(n8684), .ZN(n8690)
         );
  AOI21_X1 U10307 ( .B1(n8690), .B2(n8689), .A(n8688), .ZN(n8692) );
  OAI21_X1 U10308 ( .B1(n8692), .B2(n8691), .A(n10040), .ZN(n8694) );
  AOI21_X1 U10309 ( .B1(n8695), .B2(n8694), .A(n8693), .ZN(n8698) );
  OAI21_X1 U10310 ( .B1(n8698), .B2(n8697), .A(n8696), .ZN(n8699) );
  NAND2_X1 U10311 ( .A1(n8700), .A2(n8699), .ZN(n8702) );
  NAND2_X1 U10312 ( .A1(n8702), .A2(n8701), .ZN(n8704) );
  AOI21_X1 U10313 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8709) );
  OAI211_X1 U10314 ( .C1(n8709), .C2(n8708), .A(n8707), .B(n8706), .ZN(n8711)
         );
  NAND2_X1 U10315 ( .A1(n8711), .A2(n8710), .ZN(n8714) );
  AOI21_X1 U10316 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8715) );
  MUX2_X1 U10317 ( .A(n8716), .B(n10382), .S(n8715), .Z(n8717) );
  OAI211_X1 U10318 ( .C1(n8720), .C2(n8719), .A(n8718), .B(n8717), .ZN(n8726)
         );
  INV_X1 U10319 ( .A(n8721), .ZN(n8722) );
  OAI211_X1 U10320 ( .C1(n8724), .C2(n8723), .A(P1_B_REG_SCAN_IN), .B(n8722), 
        .ZN(n8725) );
  OAI211_X1 U10321 ( .C1(n8728), .C2(n8727), .A(n8726), .B(n8725), .ZN(
        P1_U3242) );
  MUX2_X1 U10322 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n8729), .S(n10405), .Z(
        n8730) );
  INV_X1 U10323 ( .A(n8732), .ZN(P1_U3521) );
  INV_X1 U10324 ( .A(n8733), .ZN(n8846) );
  NOR3_X1 U10325 ( .A1(n8846), .A2(n4562), .A3(n8735), .ZN(n8738) );
  INV_X1 U10326 ( .A(n8736), .ZN(n8737) );
  OAI21_X1 U10327 ( .B1(n8738), .B2(n8737), .A(n8882), .ZN(n8743) );
  NOR2_X1 U10328 ( .A1(n8739), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9003) );
  AOI21_X1 U10329 ( .B1(n8778), .B2(n9334), .A(n9003), .ZN(n8740) );
  OAI21_X1 U10330 ( .B1(n8789), .B2(n8780), .A(n8740), .ZN(n8741) );
  AOI21_X1 U10331 ( .B1(n9340), .B2(n8906), .A(n8741), .ZN(n8742) );
  OAI211_X1 U10332 ( .C1(n9338), .C2(n8909), .A(n8743), .B(n8742), .ZN(
        P2_U3155) );
  XNOR2_X1 U10333 ( .A(n8829), .B(n9214), .ZN(n8749) );
  AOI22_X1 U10334 ( .A1(n9206), .A2(n8902), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8745) );
  NAND2_X1 U10335 ( .A1(n9209), .A2(n8906), .ZN(n8744) );
  OAI211_X1 U10336 ( .C1(n8746), .C2(n8904), .A(n8745), .B(n8744), .ZN(n8747)
         );
  AOI21_X1 U10337 ( .B1(n9443), .B2(n8896), .A(n8747), .ZN(n8748) );
  OAI21_X1 U10338 ( .B1(n8749), .B2(n8898), .A(n8748), .ZN(P2_U3156) );
  XNOR2_X1 U10339 ( .A(n8750), .B(n8751), .ZN(n8753) );
  NAND2_X1 U10340 ( .A1(n8753), .A2(n8752), .ZN(n8866) );
  OAI21_X1 U10341 ( .B1(n8753), .B2(n8752), .A(n8866), .ZN(n8754) );
  NAND2_X1 U10342 ( .A1(n8754), .A2(n8882), .ZN(n8760) );
  INV_X1 U10343 ( .A(n8755), .ZN(n8758) );
  NAND2_X1 U10344 ( .A1(n8902), .A2(n8918), .ZN(n8756) );
  NAND2_X1 U10345 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8948) );
  OAI211_X1 U10346 ( .C1(n8784), .C2(n8904), .A(n8756), .B(n8948), .ZN(n8757)
         );
  AOI21_X1 U10347 ( .B1(n8758), .B2(n8906), .A(n8757), .ZN(n8759) );
  OAI211_X1 U10348 ( .C1(n8761), .C2(n8909), .A(n8760), .B(n8759), .ZN(
        P2_U3157) );
  INV_X1 U10349 ( .A(n9270), .ZN(n9386) );
  NOR3_X1 U10350 ( .A1(n4318), .A2(n4957), .A3(n8763), .ZN(n8765) );
  INV_X1 U10351 ( .A(n8764), .ZN(n8838) );
  OAI21_X1 U10352 ( .B1(n8765), .B2(n8838), .A(n8882), .ZN(n8770) );
  NOR2_X1 U10353 ( .A1(n8766), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9128) );
  AOI21_X1 U10354 ( .B1(n9261), .B2(n8778), .A(n9128), .ZN(n8767) );
  OAI21_X1 U10355 ( .B1(n9297), .B2(n8780), .A(n8767), .ZN(n8768) );
  AOI21_X1 U10356 ( .B1(n9266), .B2(n8906), .A(n8768), .ZN(n8769) );
  OAI211_X1 U10357 ( .C1(n9386), .C2(n8909), .A(n8770), .B(n8769), .ZN(
        P2_U3159) );
  INV_X1 U10358 ( .A(n8771), .ZN(n8839) );
  INV_X1 U10359 ( .A(n8772), .ZN(n8774) );
  NOR3_X1 U10360 ( .A1(n8839), .A2(n8774), .A3(n8773), .ZN(n8777) );
  INV_X1 U10361 ( .A(n8775), .ZN(n8776) );
  OAI21_X1 U10362 ( .B1(n8777), .B2(n8776), .A(n8882), .ZN(n8783) );
  AOI22_X1 U10363 ( .A1(n9206), .A2(n8778), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8779) );
  OAI21_X1 U10364 ( .B1(n9227), .B2(n8780), .A(n8779), .ZN(n8781) );
  AOI21_X1 U10365 ( .B1(n9228), .B2(n8906), .A(n8781), .ZN(n8782) );
  OAI211_X1 U10366 ( .C1(n9373), .C2(n8909), .A(n8783), .B(n8782), .ZN(
        P2_U3163) );
  OR2_X1 U10367 ( .A1(n8750), .A2(n8917), .ZN(n8865) );
  NAND3_X1 U10368 ( .A1(n8866), .A2(n8868), .A3(n8865), .ZN(n8867) );
  OAI21_X1 U10369 ( .B1(n8784), .B2(n8868), .A(n8867), .ZN(n8786) );
  XNOR2_X1 U10370 ( .A(n8786), .B(n8785), .ZN(n8795) );
  NAND2_X1 U10371 ( .A1(n8902), .A2(n8916), .ZN(n8788) );
  OAI211_X1 U10372 ( .C1(n8789), .C2(n8904), .A(n8788), .B(n8787), .ZN(n8792)
         );
  NOR2_X1 U10373 ( .A1(n8790), .A2(n8909), .ZN(n8791) );
  AOI211_X1 U10374 ( .C1(n8793), .C2(n8906), .A(n8792), .B(n8791), .ZN(n8794)
         );
  OAI21_X1 U10375 ( .B1(n8795), .B2(n8898), .A(n8794), .ZN(P2_U3164) );
  XOR2_X1 U10376 ( .A(n8797), .B(n8796), .Z(n8803) );
  AOI22_X1 U10377 ( .A1(n9205), .A2(n8902), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8799) );
  NAND2_X1 U10378 ( .A1(n9185), .A2(n8906), .ZN(n8798) );
  OAI211_X1 U10379 ( .C1(n8800), .C2(n8904), .A(n8799), .B(n8798), .ZN(n8801)
         );
  AOI21_X1 U10380 ( .B1(n9431), .B2(n8896), .A(n8801), .ZN(n8802) );
  OAI21_X1 U10381 ( .B1(n8803), .B2(n8898), .A(n8802), .ZN(P2_U3165) );
  INV_X1 U10382 ( .A(n8804), .ZN(n8820) );
  INV_X1 U10383 ( .A(n8806), .ZN(n8809) );
  INV_X1 U10384 ( .A(n8807), .ZN(n8808) );
  AOI21_X1 U10385 ( .B1(n8805), .B2(n8809), .A(n8808), .ZN(n8810) );
  OAI21_X1 U10386 ( .B1(n8820), .B2(n8810), .A(n8882), .ZN(n8815) );
  NAND2_X1 U10387 ( .A1(n8902), .A2(n9334), .ZN(n8811) );
  NAND2_X1 U10388 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9051) );
  OAI211_X1 U10389 ( .C1(n8812), .C2(n8904), .A(n8811), .B(n9051), .ZN(n8813)
         );
  AOI21_X1 U10390 ( .B1(n9305), .B2(n8906), .A(n8813), .ZN(n8814) );
  OAI211_X1 U10391 ( .C1(n8816), .C2(n8909), .A(n8815), .B(n8814), .ZN(
        P2_U3166) );
  INV_X1 U10392 ( .A(n9393), .ZN(n9301) );
  INV_X1 U10393 ( .A(n8817), .ZN(n8819) );
  NOR3_X1 U10394 ( .A1(n8820), .A2(n8819), .A3(n8818), .ZN(n8822) );
  INV_X1 U10395 ( .A(n8821), .ZN(n8881) );
  OAI21_X1 U10396 ( .B1(n8822), .B2(n8881), .A(n8882), .ZN(n8826) );
  NAND2_X1 U10397 ( .A1(n8902), .A2(n9321), .ZN(n8823) );
  NAND2_X1 U10398 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9081) );
  OAI211_X1 U10399 ( .C1(n9297), .C2(n8904), .A(n8823), .B(n9081), .ZN(n8824)
         );
  AOI21_X1 U10400 ( .B1(n9299), .B2(n8906), .A(n8824), .ZN(n8825) );
  OAI211_X1 U10401 ( .C1(n9301), .C2(n8909), .A(n8826), .B(n8825), .ZN(
        P2_U3168) );
  XNOR2_X1 U10402 ( .A(n8830), .B(n9205), .ZN(n8831) );
  AOI22_X1 U10403 ( .A1(n9193), .A2(n8902), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8832) );
  OAI21_X1 U10404 ( .B1(n8890), .B2(n8904), .A(n8832), .ZN(n8833) );
  AOI21_X1 U10405 ( .B1(n9197), .B2(n8906), .A(n8833), .ZN(n8834) );
  NOR3_X1 U10406 ( .A1(n8838), .A2(n4565), .A3(n8837), .ZN(n8840) );
  OAI21_X1 U10407 ( .B1(n8840), .B2(n8839), .A(n8882), .ZN(n8845) );
  INV_X1 U10408 ( .A(n9252), .ZN(n8841) );
  NOR2_X1 U10409 ( .A1(n8852), .A2(n8841), .ZN(n8843) );
  OAI22_X1 U10410 ( .A1(n9248), .A2(n8904), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4769), .ZN(n8842) );
  AOI211_X1 U10411 ( .C1(n8902), .C2(n9275), .A(n8843), .B(n8842), .ZN(n8844)
         );
  OAI211_X1 U10412 ( .C1(n9462), .C2(n8909), .A(n8845), .B(n8844), .ZN(
        P2_U3173) );
  AOI21_X1 U10413 ( .B1(n8848), .B2(n8847), .A(n8846), .ZN(n8856) );
  NAND2_X1 U10414 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8983) );
  OAI21_X1 U10415 ( .B1(n8904), .B2(n9316), .A(n8983), .ZN(n8849) );
  AOI21_X1 U10416 ( .B1(n8902), .B2(n8915), .A(n8849), .ZN(n8850) );
  OAI21_X1 U10417 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8853) );
  AOI21_X1 U10418 ( .B1(n8854), .B2(n8896), .A(n8853), .ZN(n8855) );
  OAI21_X1 U10419 ( .B1(n8856), .B2(n8898), .A(n8855), .ZN(P2_U3174) );
  XNOR2_X1 U10420 ( .A(n8857), .B(n9226), .ZN(n8858) );
  XNOR2_X1 U10421 ( .A(n8859), .B(n8858), .ZN(n8864) );
  INV_X1 U10422 ( .A(n9248), .ZN(n8914) );
  AOI22_X1 U10423 ( .A1(n8914), .A2(n8902), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8861) );
  NAND2_X1 U10424 ( .A1(n8906), .A2(n9219), .ZN(n8860) );
  OAI211_X1 U10425 ( .C1(n9214), .C2(n8904), .A(n8861), .B(n8860), .ZN(n8862)
         );
  AOI21_X1 U10426 ( .B1(n9370), .B2(n8896), .A(n8862), .ZN(n8863) );
  OAI21_X1 U10427 ( .B1(n8864), .B2(n8898), .A(n8863), .ZN(P2_U3175) );
  AND2_X1 U10428 ( .A1(n8866), .A2(n8865), .ZN(n8869) );
  OAI211_X1 U10429 ( .C1(n8869), .C2(n8868), .A(n8882), .B(n8867), .ZN(n8877)
         );
  INV_X1 U10430 ( .A(n8870), .ZN(n8875) );
  NAND2_X1 U10431 ( .A1(n8902), .A2(n8917), .ZN(n8872) );
  OAI211_X1 U10432 ( .C1(n8873), .C2(n8904), .A(n8872), .B(n8871), .ZN(n8874)
         );
  AOI21_X1 U10433 ( .B1(n8875), .B2(n8906), .A(n8874), .ZN(n8876) );
  OAI211_X1 U10434 ( .C1(n8878), .C2(n8909), .A(n8877), .B(n8876), .ZN(
        P2_U3176) );
  INV_X1 U10435 ( .A(n9281), .ZN(n9391) );
  NOR3_X1 U10436 ( .A1(n8881), .A2(n4958), .A3(n8880), .ZN(n8883) );
  OAI21_X1 U10437 ( .B1(n8883), .B2(n4318), .A(n8882), .ZN(n8887) );
  NAND2_X1 U10438 ( .A1(n8902), .A2(n9308), .ZN(n8884) );
  NAND2_X1 U10439 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9105) );
  OAI211_X1 U10440 ( .C1(n9247), .C2(n8904), .A(n8884), .B(n9105), .ZN(n8885)
         );
  AOI21_X1 U10441 ( .B1(n9277), .B2(n8906), .A(n8885), .ZN(n8886) );
  OAI211_X1 U10442 ( .C1(n9391), .C2(n8909), .A(n8887), .B(n8886), .ZN(
        P2_U3178) );
  AOI22_X1 U10443 ( .A1(n9192), .A2(n8902), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8893) );
  NAND2_X1 U10444 ( .A1(n9175), .A2(n8906), .ZN(n8892) );
  OAI211_X1 U10445 ( .C1(n8894), .C2(n8904), .A(n8893), .B(n8892), .ZN(n8895)
         );
  AOI21_X1 U10446 ( .B1(n9425), .B2(n8896), .A(n8895), .ZN(n8897) );
  INV_X1 U10447 ( .A(n9477), .ZN(n8910) );
  AOI21_X1 U10448 ( .B1(n8900), .B2(n8899), .A(n8898), .ZN(n8901) );
  NAND2_X1 U10449 ( .A1(n8901), .A2(n8805), .ZN(n8908) );
  NAND2_X1 U10450 ( .A1(n8902), .A2(n9320), .ZN(n8903) );
  NAND2_X1 U10451 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9029) );
  OAI211_X1 U10452 ( .C1(n9295), .C2(n8904), .A(n8903), .B(n9029), .ZN(n8905)
         );
  AOI21_X1 U10453 ( .B1(n9324), .B2(n8906), .A(n8905), .ZN(n8907) );
  OAI211_X1 U10454 ( .C1(n8910), .C2(n8909), .A(n8908), .B(n8907), .ZN(
        P2_U3181) );
  MUX2_X1 U10455 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8911), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10456 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8912), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10457 ( .A(n8913), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9103), .Z(
        P2_U3519) );
  MUX2_X1 U10458 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9172), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10459 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9181), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10460 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9192), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10461 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9205), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10462 ( .A(n9193), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9103), .Z(
        P2_U3514) );
  MUX2_X1 U10463 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9206), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10464 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8914), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10465 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9261), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10466 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9275), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10467 ( .A(n9260), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9103), .Z(
        P2_U3509) );
  MUX2_X1 U10468 ( .A(n9321), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9103), .Z(
        P2_U3507) );
  MUX2_X1 U10469 ( .A(n9334), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9103), .Z(
        P2_U3506) );
  MUX2_X1 U10470 ( .A(n9320), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9103), .Z(
        P2_U3505) );
  MUX2_X1 U10471 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9332), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10472 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8915), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10473 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8916), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10474 ( .A(n8917), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9103), .Z(
        P2_U3501) );
  MUX2_X1 U10475 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8918), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10476 ( .A(n8919), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9103), .Z(
        P2_U3499) );
  MUX2_X1 U10477 ( .A(n8920), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9103), .Z(
        P2_U3498) );
  MUX2_X1 U10478 ( .A(n8921), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9103), .Z(
        P2_U3497) );
  MUX2_X1 U10479 ( .A(n8922), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9103), .Z(
        P2_U3496) );
  MUX2_X1 U10480 ( .A(n8923), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9103), .Z(
        P2_U3495) );
  MUX2_X1 U10481 ( .A(n5334), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9103), .Z(
        P2_U3494) );
  MUX2_X1 U10482 ( .A(n8924), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9103), .Z(
        P2_U3493) );
  MUX2_X1 U10483 ( .A(n8925), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9103), .Z(
        P2_U3492) );
  MUX2_X1 U10484 ( .A(n5786), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9103), .Z(
        P2_U3491) );
  OAI21_X1 U10485 ( .B1(n9131), .B2(n8927), .A(n8926), .ZN(n8934) );
  OR3_X1 U10486 ( .A1(n8930), .A2(n8929), .A3(n8928), .ZN(n8931) );
  AOI21_X1 U10487 ( .B1(n8932), .B2(n8931), .A(n9144), .ZN(n8933) );
  AOI211_X1 U10488 ( .C1(n9142), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n8934), .B(
        n8933), .ZN(n8947) );
  AND3_X1 U10489 ( .A1(n8937), .A2(n8936), .A3(n8935), .ZN(n8938) );
  OAI21_X1 U10490 ( .B1(n8939), .B2(n8938), .A(n9042), .ZN(n8946) );
  AND3_X1 U10491 ( .A1(n8942), .A2(n8941), .A3(n8940), .ZN(n8943) );
  OAI21_X1 U10492 ( .B1(n8944), .B2(n8943), .A(n9126), .ZN(n8945) );
  NAND3_X1 U10493 ( .A1(n8947), .A2(n8946), .A3(n8945), .ZN(P2_U3190) );
  OAI21_X1 U10494 ( .B1(n9131), .B2(n8949), .A(n8948), .ZN(n8957) );
  INV_X1 U10495 ( .A(n8950), .ZN(n8952) );
  NAND3_X1 U10496 ( .A1(n8953), .A2(n8952), .A3(n8951), .ZN(n8954) );
  AOI21_X1 U10497 ( .B1(n8955), .B2(n8954), .A(n9144), .ZN(n8956) );
  AOI211_X1 U10498 ( .C1(n9142), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n8957), .B(
        n8956), .ZN(n8970) );
  AND3_X1 U10499 ( .A1(n8960), .A2(n8959), .A3(n8958), .ZN(n8961) );
  OAI21_X1 U10500 ( .B1(n8962), .B2(n8961), .A(n9042), .ZN(n8969) );
  AND3_X1 U10501 ( .A1(n8965), .A2(n8964), .A3(n8963), .ZN(n8966) );
  OAI21_X1 U10502 ( .B1(n8967), .B2(n8966), .A(n9126), .ZN(n8968) );
  NAND3_X1 U10503 ( .A1(n8970), .A2(n8969), .A3(n8968), .ZN(P2_U3192) );
  AOI21_X1 U10504 ( .B1(n8976), .B2(n8975), .A(n9015), .ZN(n8997) );
  AOI21_X1 U10505 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n8982) );
  MUX2_X1 U10506 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n4279), .Z(n9000) );
  XNOR2_X1 U10507 ( .A(n8980), .B(n9000), .ZN(n8981) );
  NAND2_X1 U10508 ( .A1(n8982), .A2(n8981), .ZN(n8998) );
  OAI21_X1 U10509 ( .B1(n8982), .B2(n8981), .A(n8998), .ZN(n8995) );
  NAND2_X1 U10510 ( .A1(n9142), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8984) );
  OAI211_X1 U10511 ( .C1(n9131), .C2(n8999), .A(n8984), .B(n8983), .ZN(n8994)
         );
  INV_X1 U10512 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U10513 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  AOI21_X1 U10514 ( .B1(n9007), .B2(n8992), .A(n9144), .ZN(n8993) );
  AOI211_X1 U10515 ( .C1(n9042), .C2(n8995), .A(n8994), .B(n8993), .ZN(n8996)
         );
  OAI21_X1 U10516 ( .B1(n8997), .B2(n9037), .A(n8996), .ZN(P2_U3195) );
  OAI21_X1 U10517 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9002) );
  MUX2_X1 U10518 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n4279), .Z(n9028) );
  XNOR2_X1 U10519 ( .A(n9031), .B(n9028), .ZN(n9001) );
  OAI21_X1 U10520 ( .B1(n9002), .B2(n9001), .A(n9026), .ZN(n9014) );
  INV_X1 U10521 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9006) );
  AOI21_X1 U10522 ( .B1(n9004), .B2(n9031), .A(n9003), .ZN(n9005) );
  OAI21_X1 U10523 ( .B1(n9106), .B2(n9006), .A(n9005), .ZN(n9013) );
  XNOR2_X1 U10524 ( .A(n9031), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n9008) );
  INV_X1 U10525 ( .A(n9008), .ZN(n9010) );
  NAND3_X1 U10526 ( .A1(n9007), .A2(n9010), .A3(n9009), .ZN(n9011) );
  AOI21_X1 U10527 ( .B1(n9021), .B2(n9011), .A(n9144), .ZN(n9012) );
  AOI211_X1 U10528 ( .C1(n9042), .C2(n9014), .A(n9013), .B(n9012), .ZN(n9020)
         );
  XNOR2_X1 U10529 ( .A(n9031), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9016) );
  NOR3_X1 U10530 ( .A1(n9017), .A2(n9015), .A3(n9016), .ZN(n9018) );
  OAI21_X1 U10531 ( .B1(n4338), .B2(n9018), .A(n9126), .ZN(n9019) );
  NAND2_X1 U10532 ( .A1(n9020), .A2(n9019), .ZN(P2_U3196) );
  INV_X1 U10533 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U10534 ( .A1(n9023), .A2(n9034), .ZN(n9046) );
  INV_X1 U10535 ( .A(n9047), .ZN(n9024) );
  AOI21_X1 U10536 ( .B1(n9323), .B2(n9025), .A(n9024), .ZN(n9044) );
  MUX2_X1 U10537 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4279), .Z(n9052) );
  XNOR2_X1 U10538 ( .A(n9054), .B(n9052), .ZN(n9055) );
  XNOR2_X1 U10539 ( .A(n9056), .B(n9055), .ZN(n9041) );
  NAND2_X1 U10540 ( .A1(n9142), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n9030) );
  OAI211_X1 U10541 ( .C1(n9034), .C2(n9131), .A(n9030), .B(n9029), .ZN(n9040)
         );
  INV_X1 U10542 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U10543 ( .A1(n9027), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U10544 ( .A1(n9033), .A2(n9034), .ZN(n9060) );
  AOI21_X1 U10545 ( .B1(n9400), .B2(n9036), .A(n4295), .ZN(n9038) );
  NOR2_X1 U10546 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  AOI211_X1 U10547 ( .C1(n9042), .C2(n9041), .A(n9040), .B(n9039), .ZN(n9043)
         );
  OAI21_X1 U10548 ( .B1(n9044), .B2(n9144), .A(n9043), .ZN(P2_U3197) );
  INV_X1 U10549 ( .A(n9046), .ZN(n9045) );
  XNOR2_X1 U10550 ( .A(n9074), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n9048) );
  NOR2_X1 U10551 ( .A1(n9045), .A2(n9048), .ZN(n9050) );
  INV_X1 U10552 ( .A(n9068), .ZN(n9049) );
  AOI21_X1 U10553 ( .B1(n9050), .B2(n9047), .A(n9049), .ZN(n9066) );
  OAI21_X1 U10554 ( .B1(n9131), .B2(n9077), .A(n9051), .ZN(n9059) );
  MUX2_X1 U10555 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4279), .Z(n9078) );
  XOR2_X1 U10556 ( .A(n9074), .B(n9078), .Z(n9079) );
  INV_X1 U10557 ( .A(n9052), .ZN(n9053) );
  XOR2_X1 U10558 ( .A(n9079), .B(n9080), .Z(n9057) );
  NOR2_X1 U10559 ( .A1(n9057), .A2(n9140), .ZN(n9058) );
  AOI211_X1 U10560 ( .C1(n9142), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n9059), .B(
        n9058), .ZN(n9065) );
  INV_X1 U10561 ( .A(n9060), .ZN(n9062) );
  XNOR2_X1 U10562 ( .A(n9074), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9061) );
  NOR3_X1 U10563 ( .A1(n4295), .A2(n9062), .A3(n9061), .ZN(n9063) );
  OAI21_X1 U10564 ( .B1(n4358), .B2(n9063), .A(n9126), .ZN(n9064) );
  OAI211_X1 U10565 ( .C1(n9066), .C2(n9144), .A(n9065), .B(n9064), .ZN(
        P2_U3198) );
  INV_X1 U10566 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9073) );
  INV_X1 U10567 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U10568 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  OAI21_X1 U10569 ( .B1(n9069), .B2(n9082), .A(n9093), .ZN(n9072) );
  INV_X1 U10570 ( .A(n9072), .ZN(n9070) );
  INV_X1 U10571 ( .A(n9091), .ZN(n9071) );
  AOI21_X1 U10572 ( .B1(n9073), .B2(n9072), .A(n9071), .ZN(n9089) );
  INV_X1 U10573 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U10574 ( .A1(n9075), .A2(n9082), .ZN(n9114) );
  OAI21_X1 U10575 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9076), .A(n9115), .ZN(
        n9087) );
  MUX2_X1 U10576 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4279), .Z(n9095) );
  XNOR2_X1 U10577 ( .A(n9095), .B(n9097), .ZN(n9098) );
  XOR2_X1 U10578 ( .A(n9098), .B(n9099), .Z(n9085) );
  OAI21_X1 U10579 ( .B1(n9131), .B2(n9082), .A(n9081), .ZN(n9083) );
  AOI21_X1 U10580 ( .B1(n9142), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9083), .ZN(
        n9084) );
  OAI21_X1 U10581 ( .B1(n9085), .B2(n9140), .A(n9084), .ZN(n9086) );
  AOI21_X1 U10582 ( .B1(n9087), .B2(n9126), .A(n9086), .ZN(n9088) );
  OAI21_X1 U10583 ( .B1(n9089), .B2(n9144), .A(n9088), .ZN(P2_U3199) );
  INV_X1 U10584 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9279) );
  OR2_X1 U10585 ( .A1(n9133), .A2(n9279), .ZN(n9120) );
  NAND2_X1 U10586 ( .A1(n9133), .A2(n9279), .ZN(n9090) );
  NAND2_X1 U10587 ( .A1(n9120), .A2(n9090), .ZN(n9092) );
  AND3_X1 U10588 ( .A1(n9091), .A2(n9093), .A3(n9092), .ZN(n9094) );
  NOR2_X1 U10589 ( .A1(n9121), .A2(n9094), .ZN(n9119) );
  INV_X1 U10590 ( .A(n9095), .ZN(n9096) );
  AOI22_X1 U10591 ( .A1(n9099), .A2(n9098), .B1(n9097), .B2(n9096), .ZN(n9101)
         );
  MUX2_X1 U10592 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4279), .Z(n9100) );
  NOR2_X1 U10593 ( .A1(n9101), .A2(n9100), .ZN(n9134) );
  NAND2_X1 U10594 ( .A1(n9101), .A2(n9100), .ZN(n9132) );
  INV_X1 U10595 ( .A(n9132), .ZN(n9102) );
  NOR2_X1 U10596 ( .A1(n9134), .A2(n9102), .ZN(n9107) );
  INV_X1 U10597 ( .A(n9107), .ZN(n9104) );
  OAI21_X1 U10598 ( .B1(n9104), .B2(n9103), .A(n9131), .ZN(n9110) );
  INV_X1 U10599 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10457) );
  OAI21_X1 U10600 ( .B1(n9106), .B2(n10457), .A(n9105), .ZN(n9109) );
  NOR3_X1 U10601 ( .A1(n9107), .A2(n9133), .A3(n9140), .ZN(n9108) );
  AOI211_X1 U10602 ( .C1(n9133), .C2(n9110), .A(n9109), .B(n9108), .ZN(n9118)
         );
  INV_X1 U10603 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9111) );
  OR2_X1 U10604 ( .A1(n9133), .A2(n9111), .ZN(n9122) );
  NAND2_X1 U10605 ( .A1(n9133), .A2(n9111), .ZN(n9112) );
  NAND2_X1 U10606 ( .A1(n9122), .A2(n9112), .ZN(n9113) );
  AOI21_X1 U10607 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9124) );
  AND3_X1 U10608 ( .A1(n9115), .A2(n9114), .A3(n9113), .ZN(n9116) );
  OAI21_X1 U10609 ( .B1(n9124), .B2(n9116), .A(n9126), .ZN(n9117) );
  OAI211_X1 U10610 ( .C1(n9119), .C2(n9144), .A(n9118), .B(n9117), .ZN(
        P2_U3200) );
  INV_X1 U10611 ( .A(n9122), .ZN(n9123) );
  NOR2_X1 U10612 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  XNOR2_X1 U10613 ( .A(n9130), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9135) );
  XNOR2_X1 U10614 ( .A(n9125), .B(n9135), .ZN(n9127) );
  NAND2_X1 U10615 ( .A1(n9127), .A2(n9126), .ZN(n9143) );
  INV_X1 U10616 ( .A(n9128), .ZN(n9129) );
  OAI21_X1 U10617 ( .B1(n9131), .B2(n9130), .A(n9129), .ZN(n9141) );
  OAI21_X1 U10618 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(n9139) );
  INV_X1 U10619 ( .A(n9135), .ZN(n9137) );
  MUX2_X1 U10620 ( .A(n4420), .B(n9137), .S(n4279), .Z(n9138) );
  NAND2_X1 U10621 ( .A1(n9410), .A2(n9325), .ZN(n9149) );
  INV_X1 U10622 ( .A(n9145), .ZN(n9146) );
  AND2_X1 U10623 ( .A1(n9148), .A2(n9341), .ZN(n9156) );
  AOI21_X1 U10624 ( .B1(n9411), .B2(n10421), .A(n9156), .ZN(n9152) );
  OAI211_X1 U10625 ( .C1(n10421), .C2(n9150), .A(n9149), .B(n9152), .ZN(
        P2_U3202) );
  NAND2_X1 U10626 ( .A1(n10413), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9151) );
  OAI211_X1 U10627 ( .C1(n9416), .C2(n10415), .A(n9152), .B(n9151), .ZN(
        P2_U3203) );
  NAND2_X1 U10628 ( .A1(n9153), .A2(n10421), .ZN(n9158) );
  NOR2_X1 U10629 ( .A1(n9154), .A2(n10415), .ZN(n9155) );
  AOI211_X1 U10630 ( .C1(n10413), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9156), .B(
        n9155), .ZN(n9157) );
  OAI211_X1 U10631 ( .C1(n6759), .C2(n9159), .A(n9158), .B(n9157), .ZN(
        P2_U3204) );
  INV_X1 U10632 ( .A(n9160), .ZN(n9161) );
  NOR3_X1 U10633 ( .A1(n9162), .A2(n9161), .A3(n9344), .ZN(n9166) );
  AOI22_X1 U10634 ( .A1(n9163), .A2(n9341), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10413), .ZN(n9164) );
  OAI21_X1 U10635 ( .B1(n9356), .B2(n10415), .A(n9164), .ZN(n9165) );
  AOI211_X1 U10636 ( .C1(n9167), .C2(n10421), .A(n9166), .B(n9165), .ZN(n9168)
         );
  INV_X1 U10637 ( .A(n9168), .ZN(P2_U3206) );
  XNOR2_X1 U10638 ( .A(n9169), .B(n9170), .ZN(n9426) );
  INV_X1 U10639 ( .A(n9426), .ZN(n9178) );
  INV_X1 U10640 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9174) );
  XNOR2_X1 U10641 ( .A(n9171), .B(n9170), .ZN(n9173) );
  AOI222_X1 U10642 ( .A1(n9336), .A2(n9173), .B1(n9192), .B2(n9331), .C1(n9172), .C2(n9333), .ZN(n9423) );
  MUX2_X1 U10643 ( .A(n9174), .B(n9423), .S(n10421), .Z(n9177) );
  AOI22_X1 U10644 ( .A1(n9425), .A2(n9325), .B1(n9341), .B2(n9175), .ZN(n9176)
         );
  OAI211_X1 U10645 ( .C1(n9178), .C2(n9344), .A(n9177), .B(n9176), .ZN(
        P2_U3207) );
  NOR2_X1 U10646 ( .A1(n9179), .A2(n9337), .ZN(n9184) );
  XNOR2_X1 U10647 ( .A(n9180), .B(n9187), .ZN(n9182) );
  AOI222_X1 U10648 ( .A1(n9336), .A2(n9182), .B1(n9205), .B2(n9331), .C1(n9181), .C2(n9333), .ZN(n9429) );
  INV_X1 U10649 ( .A(n9429), .ZN(n9183) );
  AOI211_X1 U10650 ( .C1(n9341), .C2(n9185), .A(n9184), .B(n9183), .ZN(n9189)
         );
  XNOR2_X1 U10651 ( .A(n9186), .B(n9187), .ZN(n9432) );
  AOI22_X1 U10652 ( .A1(n9432), .A2(n9283), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10413), .ZN(n9188) );
  OAI21_X1 U10653 ( .B1(n9189), .B2(n10413), .A(n9188), .ZN(P2_U3208) );
  NOR2_X1 U10654 ( .A1(n9190), .A2(n9337), .ZN(n9196) );
  XOR2_X1 U10655 ( .A(n9198), .B(n9191), .Z(n9194) );
  AOI222_X1 U10656 ( .A1(n9336), .A2(n9194), .B1(n9193), .B2(n9331), .C1(n9192), .C2(n9333), .ZN(n9435) );
  INV_X1 U10657 ( .A(n9435), .ZN(n9195) );
  AOI211_X1 U10658 ( .C1(n9341), .C2(n9197), .A(n9196), .B(n9195), .ZN(n9200)
         );
  XOR2_X1 U10659 ( .A(n4388), .B(n9198), .Z(n9438) );
  AOI22_X1 U10660 ( .A1(n9438), .A2(n9283), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10413), .ZN(n9199) );
  OAI21_X1 U10661 ( .B1(n9200), .B2(n10413), .A(n9199), .ZN(P2_U3209) );
  XNOR2_X1 U10662 ( .A(n9202), .B(n9201), .ZN(n9446) );
  INV_X1 U10663 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9208) );
  XNOR2_X1 U10664 ( .A(n9203), .B(n9204), .ZN(n9207) );
  AOI222_X1 U10665 ( .A1(n9336), .A2(n9207), .B1(n9206), .B2(n9331), .C1(n9205), .C2(n9333), .ZN(n9441) );
  MUX2_X1 U10666 ( .A(n9208), .B(n9441), .S(n10421), .Z(n9211) );
  AOI22_X1 U10667 ( .A1(n9443), .A2(n9325), .B1(n9341), .B2(n9209), .ZN(n9210)
         );
  OAI211_X1 U10668 ( .C1(n9446), .C2(n9344), .A(n9211), .B(n9210), .ZN(
        P2_U3210) );
  XOR2_X1 U10669 ( .A(n9215), .B(n9212), .Z(n9213) );
  OAI222_X1 U10670 ( .A1(n9298), .A2(n9214), .B1(n9296), .B2(n9248), .C1(n9213), .C2(n9293), .ZN(n9369) );
  OR2_X1 U10671 ( .A1(n9216), .A2(n9215), .ZN(n9217) );
  NAND2_X1 U10672 ( .A1(n9218), .A2(n9217), .ZN(n9450) );
  AOI22_X1 U10673 ( .A1(n10413), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9219), 
        .B2(n9341), .ZN(n9221) );
  NAND2_X1 U10674 ( .A1(n9370), .A2(n9325), .ZN(n9220) );
  OAI211_X1 U10675 ( .C1(n9450), .C2(n9344), .A(n9221), .B(n9220), .ZN(n9222)
         );
  AOI21_X1 U10676 ( .B1(n9369), .B2(n10421), .A(n9222), .ZN(n9223) );
  INV_X1 U10677 ( .A(n9223), .ZN(P2_U3211) );
  XOR2_X1 U10678 ( .A(n9224), .B(n9237), .Z(n9225) );
  OAI222_X1 U10679 ( .A1(n9296), .A2(n9227), .B1(n9298), .B2(n9226), .C1(n9293), .C2(n9225), .ZN(n9451) );
  AOI21_X1 U10680 ( .B1(n9341), .B2(n9228), .A(n9451), .ZN(n9240) );
  AOI22_X1 U10681 ( .A1(n9454), .A2(n9325), .B1(P2_REG2_REG_21__SCAN_IN), .B2(
        n10413), .ZN(n9239) );
  INV_X1 U10682 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U10683 ( .A1(n9230), .A2(n9274), .ZN(n9388) );
  NAND2_X1 U10684 ( .A1(n9388), .A2(n9231), .ZN(n9265) );
  NAND2_X1 U10685 ( .A1(n9265), .A2(n9264), .ZN(n9382) );
  NAND2_X1 U10686 ( .A1(n9382), .A2(n9232), .ZN(n9241) );
  INV_X1 U10687 ( .A(n9233), .ZN(n9235) );
  OAI21_X1 U10688 ( .B1(n9241), .B2(n9235), .A(n9234), .ZN(n9236) );
  XOR2_X1 U10689 ( .A(n9237), .B(n9236), .Z(n9455) );
  NAND2_X1 U10690 ( .A1(n9455), .A2(n9283), .ZN(n9238) );
  OAI211_X1 U10691 ( .C1(n9240), .C2(n10413), .A(n9239), .B(n9238), .ZN(
        P2_U3212) );
  XNOR2_X1 U10692 ( .A(n9241), .B(n5625), .ZN(n9378) );
  INV_X1 U10693 ( .A(n9378), .ZN(n9256) );
  NAND2_X1 U10694 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  NAND2_X1 U10695 ( .A1(n9245), .A2(n9244), .ZN(n9246) );
  NAND2_X1 U10696 ( .A1(n9246), .A2(n9336), .ZN(n9251) );
  OAI22_X1 U10697 ( .A1(n9248), .A2(n9298), .B1(n9247), .B2(n9296), .ZN(n9249)
         );
  INV_X1 U10698 ( .A(n9249), .ZN(n9250) );
  NAND2_X1 U10699 ( .A1(n9251), .A2(n9250), .ZN(n9377) );
  AOI22_X1 U10700 ( .A1(n10413), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9341), 
        .B2(n9252), .ZN(n9253) );
  OAI21_X1 U10701 ( .B1(n9462), .B2(n10415), .A(n9253), .ZN(n9254) );
  AOI21_X1 U10702 ( .B1(n9377), .B2(n10421), .A(n9254), .ZN(n9255) );
  OAI21_X1 U10703 ( .B1(n9256), .B2(n9344), .A(n9255), .ZN(P2_U3213) );
  OAI211_X1 U10704 ( .C1(n9257), .C2(n9259), .A(n9258), .B(n9336), .ZN(n9263)
         );
  AOI22_X1 U10705 ( .A1(n9261), .A2(n9333), .B1(n9331), .B2(n9260), .ZN(n9262)
         );
  AND2_X1 U10706 ( .A1(n9263), .A2(n9262), .ZN(n9384) );
  OR2_X1 U10707 ( .A1(n9265), .A2(n9264), .ZN(n9383) );
  NAND3_X1 U10708 ( .A1(n9383), .A2(n9382), .A3(n9283), .ZN(n9272) );
  INV_X1 U10709 ( .A(n9266), .ZN(n9267) );
  OAI22_X1 U10710 ( .A1(n10421), .A2(n9268), .B1(n9267), .B2(n10417), .ZN(
        n9269) );
  AOI21_X1 U10711 ( .B1(n9270), .B2(n9325), .A(n9269), .ZN(n9271) );
  OAI211_X1 U10712 ( .C1(n9384), .C2(n10413), .A(n9272), .B(n9271), .ZN(
        P2_U3214) );
  XNOR2_X1 U10713 ( .A(n9273), .B(n9274), .ZN(n9276) );
  AOI222_X1 U10714 ( .A1(n9336), .A2(n9276), .B1(n9275), .B2(n9333), .C1(n9308), .C2(n9331), .ZN(n9390) );
  INV_X1 U10715 ( .A(n9277), .ZN(n9278) );
  OAI22_X1 U10716 ( .A1(n10421), .A2(n9279), .B1(n9278), .B2(n10417), .ZN(
        n9280) );
  AOI21_X1 U10717 ( .B1(n9281), .B2(n9325), .A(n9280), .ZN(n9285) );
  NAND2_X1 U10718 ( .A1(n9229), .A2(n9282), .ZN(n9387) );
  NAND3_X1 U10719 ( .A1(n9388), .A2(n9283), .A3(n9387), .ZN(n9284) );
  OAI211_X1 U10720 ( .C1(n9390), .C2(n10413), .A(n9285), .B(n9284), .ZN(
        P2_U3215) );
  NOR2_X1 U10721 ( .A1(n9286), .A2(n9307), .ZN(n9304) );
  NOR2_X1 U10722 ( .A1(n9304), .A2(n9287), .ZN(n9289) );
  XNOR2_X1 U10723 ( .A(n9289), .B(n9288), .ZN(n9468) );
  CLKBUF_X1 U10724 ( .A(n9290), .Z(n9292) );
  XNOR2_X1 U10725 ( .A(n9292), .B(n9291), .ZN(n9294) );
  OAI222_X1 U10726 ( .A1(n9298), .A2(n9297), .B1(n9296), .B2(n9295), .C1(n9294), .C2(n9293), .ZN(n9392) );
  AOI22_X1 U10727 ( .A1(n10413), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9341), 
        .B2(n9299), .ZN(n9300) );
  OAI21_X1 U10728 ( .B1(n9301), .B2(n10415), .A(n9300), .ZN(n9302) );
  AOI21_X1 U10729 ( .B1(n9392), .B2(n10421), .A(n9302), .ZN(n9303) );
  OAI21_X1 U10730 ( .B1(n9468), .B2(n9344), .A(n9303), .ZN(P2_U3216) );
  AOI21_X1 U10731 ( .B1(n9286), .B2(n9307), .A(n9304), .ZN(n9474) );
  AOI22_X1 U10732 ( .A1(n9471), .A2(n9325), .B1(n9341), .B2(n9305), .ZN(n9312)
         );
  XNOR2_X1 U10733 ( .A(n9306), .B(n9307), .ZN(n9309) );
  AOI222_X1 U10734 ( .A1(n9336), .A2(n9309), .B1(n9308), .B2(n9333), .C1(n9334), .C2(n9331), .ZN(n9469) );
  MUX2_X1 U10735 ( .A(n9310), .B(n9469), .S(n10421), .Z(n9311) );
  OAI211_X1 U10736 ( .C1(n9474), .C2(n9344), .A(n9312), .B(n9311), .ZN(
        P2_U3217) );
  XNOR2_X1 U10737 ( .A(n9313), .B(n9318), .ZN(n9481) );
  NAND2_X1 U10738 ( .A1(n9315), .A2(n9314), .ZN(n9330) );
  AOI22_X1 U10739 ( .A1(n9330), .A2(n9317), .B1(n9316), .B2(n9338), .ZN(n9319)
         );
  XNOR2_X1 U10740 ( .A(n9319), .B(n9318), .ZN(n9322) );
  AOI222_X1 U10741 ( .A1(n9336), .A2(n9322), .B1(n9321), .B2(n9333), .C1(n9320), .C2(n9331), .ZN(n9475) );
  MUX2_X1 U10742 ( .A(n9323), .B(n9475), .S(n10421), .Z(n9327) );
  AOI22_X1 U10743 ( .A1(n9477), .A2(n9325), .B1(n9341), .B2(n9324), .ZN(n9326)
         );
  OAI211_X1 U10744 ( .C1(n9481), .C2(n9344), .A(n9327), .B(n9326), .ZN(
        P2_U3218) );
  XNOR2_X1 U10745 ( .A(n9328), .B(n9329), .ZN(n9487) );
  INV_X1 U10746 ( .A(n9487), .ZN(n9345) );
  XOR2_X1 U10747 ( .A(n9330), .B(n9329), .Z(n9335) );
  AOI222_X1 U10748 ( .A1(n9336), .A2(n9335), .B1(n9334), .B2(n9333), .C1(n9332), .C2(n9331), .ZN(n9482) );
  OAI21_X1 U10749 ( .B1(n9338), .B2(n9337), .A(n9482), .ZN(n9339) );
  NAND2_X1 U10750 ( .A1(n9339), .A2(n10421), .ZN(n9343) );
  AOI22_X1 U10751 ( .A1(n10413), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9341), 
        .B2(n9340), .ZN(n9342) );
  OAI211_X1 U10752 ( .C1(n9345), .C2(n9344), .A(n9343), .B(n9342), .ZN(
        P2_U3219) );
  NAND2_X1 U10753 ( .A1(n9410), .A2(n9406), .ZN(n9346) );
  NAND2_X1 U10754 ( .A1(n9411), .A2(n9404), .ZN(n9349) );
  OAI211_X1 U10755 ( .C1(n9404), .C2(n9347), .A(n9346), .B(n9349), .ZN(
        P2_U3490) );
  NAND2_X1 U10756 ( .A1(n10446), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9348) );
  OAI211_X1 U10757 ( .C1(n9416), .C2(n9381), .A(n9349), .B(n9348), .ZN(
        P2_U3489) );
  INV_X1 U10758 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9350) );
  AOI22_X1 U10759 ( .A1(n9420), .A2(n9407), .B1(n9406), .B2(n9419), .ZN(n9351)
         );
  NAND2_X1 U10760 ( .A1(n9352), .A2(n9351), .ZN(P2_U3487) );
  INV_X1 U10761 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9354) );
  MUX2_X1 U10762 ( .A(n9354), .B(n9353), .S(n9404), .Z(n9355) );
  OAI21_X1 U10763 ( .B1(n9356), .B2(n9381), .A(n9355), .ZN(P2_U3486) );
  INV_X1 U10764 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9357) );
  MUX2_X1 U10765 ( .A(n9357), .B(n9423), .S(n9404), .Z(n9359) );
  AOI22_X1 U10766 ( .A1(n9426), .A2(n9407), .B1(n9406), .B2(n9425), .ZN(n9358)
         );
  NAND2_X1 U10767 ( .A1(n9359), .A2(n9358), .ZN(P2_U3485) );
  INV_X1 U10768 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9360) );
  MUX2_X1 U10769 ( .A(n9360), .B(n9429), .S(n10448), .Z(n9362) );
  AOI22_X1 U10770 ( .A1(n9432), .A2(n9407), .B1(n9406), .B2(n9431), .ZN(n9361)
         );
  NAND2_X1 U10771 ( .A1(n9362), .A2(n9361), .ZN(P2_U3484) );
  INV_X1 U10772 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9363) );
  MUX2_X1 U10773 ( .A(n9363), .B(n9435), .S(n10448), .Z(n9365) );
  AOI22_X1 U10774 ( .A1(n9438), .A2(n9407), .B1(n9406), .B2(n9437), .ZN(n9364)
         );
  NAND2_X1 U10775 ( .A1(n9365), .A2(n9364), .ZN(P2_U3483) );
  INV_X1 U10776 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9366) );
  MUX2_X1 U10777 ( .A(n9366), .B(n9441), .S(n9404), .Z(n9368) );
  NAND2_X1 U10778 ( .A1(n9443), .A2(n9406), .ZN(n9367) );
  OAI211_X1 U10779 ( .C1(n9446), .C2(n9403), .A(n9368), .B(n9367), .ZN(
        P2_U3482) );
  INV_X1 U10780 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9371) );
  AOI21_X1 U10781 ( .B1(n9394), .B2(n9370), .A(n9369), .ZN(n9447) );
  MUX2_X1 U10782 ( .A(n9371), .B(n9447), .S(n9404), .Z(n9372) );
  OAI21_X1 U10783 ( .B1(n9403), .B2(n9450), .A(n9372), .ZN(P2_U3481) );
  MUX2_X1 U10784 ( .A(n9451), .B(P2_REG1_REG_21__SCAN_IN), .S(n10446), .Z(
        n9376) );
  INV_X1 U10785 ( .A(n9455), .ZN(n9374) );
  OAI22_X1 U10786 ( .A1(n9374), .A2(n9403), .B1(n9373), .B2(n9381), .ZN(n9375)
         );
  OR2_X1 U10787 ( .A1(n9376), .A2(n9375), .ZN(P2_U3480) );
  INV_X1 U10788 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9379) );
  AOI21_X1 U10789 ( .B1(n9378), .B2(n10426), .A(n9377), .ZN(n9458) );
  MUX2_X1 U10790 ( .A(n9379), .B(n9458), .S(n9404), .Z(n9380) );
  OAI21_X1 U10791 ( .B1(n9462), .B2(n9381), .A(n9380), .ZN(P2_U3479) );
  NAND3_X1 U10792 ( .A1(n9383), .A2(n10426), .A3(n9382), .ZN(n9385) );
  OAI211_X1 U10793 ( .C1(n9386), .C2(n10434), .A(n9385), .B(n9384), .ZN(n9463)
         );
  MUX2_X1 U10794 ( .A(n9463), .B(P2_REG1_REG_19__SCAN_IN), .S(n10446), .Z(
        P2_U3478) );
  NAND3_X1 U10795 ( .A1(n9388), .A2(n10426), .A3(n9387), .ZN(n9389) );
  OAI211_X1 U10796 ( .C1(n9391), .C2(n10434), .A(n9390), .B(n9389), .ZN(n9464)
         );
  MUX2_X1 U10797 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9464), .S(n10448), .Z(
        P2_U3477) );
  INV_X1 U10798 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9395) );
  AOI21_X1 U10799 ( .B1(n9394), .B2(n9393), .A(n9392), .ZN(n9465) );
  MUX2_X1 U10800 ( .A(n9395), .B(n9465), .S(n9404), .Z(n9396) );
  OAI21_X1 U10801 ( .B1(n9403), .B2(n9468), .A(n9396), .ZN(P2_U3476) );
  MUX2_X1 U10802 ( .A(n9397), .B(n9469), .S(n9404), .Z(n9399) );
  NAND2_X1 U10803 ( .A1(n9471), .A2(n9406), .ZN(n9398) );
  OAI211_X1 U10804 ( .C1(n9474), .C2(n9403), .A(n9399), .B(n9398), .ZN(
        P2_U3475) );
  MUX2_X1 U10805 ( .A(n9400), .B(n9475), .S(n9404), .Z(n9402) );
  NAND2_X1 U10806 ( .A1(n9477), .A2(n9406), .ZN(n9401) );
  OAI211_X1 U10807 ( .C1(n9403), .C2(n9481), .A(n9402), .B(n9401), .ZN(
        P2_U3474) );
  MUX2_X1 U10808 ( .A(n9405), .B(n9482), .S(n9404), .Z(n9409) );
  AOI22_X1 U10809 ( .A1(n9487), .A2(n9407), .B1(n9406), .B2(n9484), .ZN(n9408)
         );
  NAND2_X1 U10810 ( .A1(n9409), .A2(n9408), .ZN(P2_U3473) );
  NAND2_X1 U10811 ( .A1(n9410), .A2(n9485), .ZN(n9412) );
  NAND2_X1 U10812 ( .A1(n9411), .A2(n10440), .ZN(n9415) );
  OAI211_X1 U10813 ( .C1(n9413), .C2(n10440), .A(n9412), .B(n9415), .ZN(
        P2_U3458) );
  NAND2_X1 U10814 ( .A1(n10441), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9414) );
  OAI211_X1 U10815 ( .C1(n9416), .C2(n9461), .A(n9415), .B(n9414), .ZN(
        P2_U3457) );
  INV_X1 U10816 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9418) );
  AOI22_X1 U10817 ( .A1(n9420), .A2(n9486), .B1(n9485), .B2(n9419), .ZN(n9421)
         );
  NAND2_X1 U10818 ( .A1(n9422), .A2(n9421), .ZN(P2_U3455) );
  MUX2_X1 U10819 ( .A(n9424), .B(n9423), .S(n10440), .Z(n9428) );
  AOI22_X1 U10820 ( .A1(n9426), .A2(n9486), .B1(n9485), .B2(n9425), .ZN(n9427)
         );
  NAND2_X1 U10821 ( .A1(n9428), .A2(n9427), .ZN(P2_U3453) );
  MUX2_X1 U10822 ( .A(n9430), .B(n9429), .S(n10440), .Z(n9434) );
  AOI22_X1 U10823 ( .A1(n9432), .A2(n9486), .B1(n9485), .B2(n9431), .ZN(n9433)
         );
  NAND2_X1 U10824 ( .A1(n9434), .A2(n9433), .ZN(P2_U3452) );
  MUX2_X1 U10825 ( .A(n9436), .B(n9435), .S(n10440), .Z(n9440) );
  AOI22_X1 U10826 ( .A1(n9438), .A2(n9486), .B1(n9485), .B2(n9437), .ZN(n9439)
         );
  NAND2_X1 U10827 ( .A1(n9440), .A2(n9439), .ZN(P2_U3451) );
  MUX2_X1 U10828 ( .A(n9442), .B(n9441), .S(n10440), .Z(n9445) );
  NAND2_X1 U10829 ( .A1(n9443), .A2(n9485), .ZN(n9444) );
  OAI211_X1 U10830 ( .C1(n9446), .C2(n9480), .A(n9445), .B(n9444), .ZN(
        P2_U3450) );
  MUX2_X1 U10831 ( .A(n9448), .B(n9447), .S(n10440), .Z(n9449) );
  OAI21_X1 U10832 ( .B1(n9450), .B2(n9480), .A(n9449), .ZN(P2_U3449) );
  INV_X1 U10833 ( .A(n9451), .ZN(n9452) );
  MUX2_X1 U10834 ( .A(n9453), .B(n9452), .S(n10440), .Z(n9457) );
  AOI22_X1 U10835 ( .A1(n9455), .A2(n9486), .B1(n9485), .B2(n9454), .ZN(n9456)
         );
  NAND2_X1 U10836 ( .A1(n9457), .A2(n9456), .ZN(P2_U3448) );
  MUX2_X1 U10837 ( .A(n9459), .B(n9458), .S(n10440), .Z(n9460) );
  OAI21_X1 U10838 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(P2_U3447) );
  MUX2_X1 U10839 ( .A(n9463), .B(P2_REG0_REG_19__SCAN_IN), .S(n10441), .Z(
        P2_U3446) );
  MUX2_X1 U10840 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9464), .S(n10440), .Z(
        P2_U3444) );
  INV_X1 U10841 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9466) );
  MUX2_X1 U10842 ( .A(n9466), .B(n9465), .S(n10440), .Z(n9467) );
  OAI21_X1 U10843 ( .B1(n9468), .B2(n9480), .A(n9467), .ZN(P2_U3441) );
  MUX2_X1 U10844 ( .A(n9470), .B(n9469), .S(n10440), .Z(n9473) );
  NAND2_X1 U10845 ( .A1(n9471), .A2(n9485), .ZN(n9472) );
  OAI211_X1 U10846 ( .C1(n9474), .C2(n9480), .A(n9473), .B(n9472), .ZN(
        P2_U3438) );
  INV_X1 U10847 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9476) );
  MUX2_X1 U10848 ( .A(n9476), .B(n9475), .S(n10440), .Z(n9479) );
  NAND2_X1 U10849 ( .A1(n9477), .A2(n9485), .ZN(n9478) );
  OAI211_X1 U10850 ( .C1(n9481), .C2(n9480), .A(n9479), .B(n9478), .ZN(
        P2_U3435) );
  MUX2_X1 U10851 ( .A(n9483), .B(n9482), .S(n10440), .Z(n9489) );
  AOI22_X1 U10852 ( .A1(n9487), .A2(n9486), .B1(n9485), .B2(n9484), .ZN(n9488)
         );
  NAND2_X1 U10853 ( .A1(n9489), .A2(n9488), .ZN(P2_U3432) );
  NAND2_X1 U10854 ( .A1(n9495), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9490) );
  OAI211_X1 U10855 ( .C1(n9492), .C2(n9497), .A(n9491), .B(n9490), .ZN(
        P2_U3267) );
  INV_X1 U10856 ( .A(n9493), .ZN(n10250) );
  AOI21_X1 U10857 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9495), .A(n9494), .ZN(
        n9496) );
  OAI21_X1 U10858 ( .B1(n10250), .B2(n9497), .A(n9496), .ZN(P2_U3268) );
  INV_X1 U10859 ( .A(n9498), .ZN(n10254) );
  OAI222_X1 U10860 ( .A1(n9497), .A2(n10254), .B1(P2_U3151), .B2(n9500), .C1(
        n9499), .C2(n9502), .ZN(P2_U3269) );
  INV_X1 U10861 ( .A(n9501), .ZN(n10261) );
  OAI222_X1 U10862 ( .A1(n9497), .A2(n10261), .B1(P2_U3151), .B2(n5755), .C1(
        n9503), .C2(n9502), .ZN(P2_U3271) );
  MUX2_X1 U10863 ( .A(n9504), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10864 ( .B1(n9702), .B2(n9506), .A(n9505), .ZN(n9508) );
  OAI21_X1 U10865 ( .B1(n9508), .B2(n9507), .A(n9672), .ZN(n9513) );
  AOI22_X1 U10866 ( .A1(n9509), .A2(n9705), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9510) );
  OAI21_X1 U10867 ( .B1(n9916), .B2(n9717), .A(n9510), .ZN(n9511) );
  AOI21_X1 U10868 ( .B1(n9728), .B2(n9709), .A(n9511), .ZN(n9512) );
  OAI211_X1 U10869 ( .C1(n4445), .C2(n9712), .A(n9513), .B(n9512), .ZN(
        P1_U3214) );
  INV_X1 U10870 ( .A(n9514), .ZN(n9515) );
  AOI21_X1 U10871 ( .B1(n9517), .B2(n9516), .A(n9515), .ZN(n9523) );
  NAND2_X1 U10872 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10294)
         );
  OAI21_X1 U10873 ( .B1(n9717), .B2(n9583), .A(n10294), .ZN(n9521) );
  OAI22_X1 U10874 ( .A1(n9519), .A2(n9719), .B1(n9718), .B2(n9518), .ZN(n9520)
         );
  AOI211_X1 U10875 ( .C1(n10198), .C2(n9722), .A(n9521), .B(n9520), .ZN(n9522)
         );
  OAI21_X1 U10876 ( .B1(n9523), .B2(n9724), .A(n9522), .ZN(P1_U3215) );
  INV_X1 U10877 ( .A(n10226), .ZN(n9534) );
  OR2_X1 U10878 ( .A1(n9525), .A2(n9524), .ZN(n9670) );
  NAND2_X1 U10879 ( .A1(n9670), .A2(n9669), .ZN(n9668) );
  NAND2_X1 U10880 ( .A1(n9525), .A2(n9524), .ZN(n9671) );
  NAND2_X1 U10881 ( .A1(n9623), .A2(n9526), .ZN(n9527) );
  AOI21_X1 U10882 ( .B1(n9668), .B2(n9671), .A(n9527), .ZN(n9625) );
  AND3_X1 U10883 ( .A1(n9668), .A2(n9671), .A3(n9527), .ZN(n9528) );
  OAI21_X1 U10884 ( .B1(n9625), .B2(n9528), .A(n9672), .ZN(n9533) );
  NOR2_X1 U10885 ( .A1(n9983), .A2(n9717), .ZN(n9531) );
  OAI22_X1 U10886 ( .A1(n9951), .A2(n9718), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9529), .ZN(n9530) );
  AOI211_X1 U10887 ( .C1(n9950), .C2(n9709), .A(n9531), .B(n9530), .ZN(n9532)
         );
  OAI211_X1 U10888 ( .C1(n9534), .C2(n9712), .A(n9533), .B(n9532), .ZN(
        P1_U3216) );
  INV_X1 U10889 ( .A(n9535), .ZN(n9544) );
  INV_X1 U10890 ( .A(n9536), .ZN(n9539) );
  OAI21_X1 U10891 ( .B1(n9539), .B2(n9538), .A(n9537), .ZN(n9637) );
  AND2_X1 U10892 ( .A1(n9637), .A2(n9540), .ZN(n9542) );
  NOR2_X1 U10893 ( .A1(n9542), .A2(n9541), .ZN(n9683) );
  AOI21_X1 U10894 ( .B1(n9542), .B2(n9541), .A(n9683), .ZN(n9543) );
  NAND2_X1 U10895 ( .A1(n9543), .A2(n9544), .ZN(n9686) );
  OAI21_X1 U10896 ( .B1(n9544), .B2(n9543), .A(n9686), .ZN(n9545) );
  NAND2_X1 U10897 ( .A1(n9545), .A2(n9672), .ZN(n9550) );
  OAI22_X1 U10898 ( .A1(n9546), .A2(n9719), .B1(n9718), .B2(n10099), .ZN(n9547) );
  AOI211_X1 U10899 ( .C1(n9695), .C2(n9736), .A(n9548), .B(n9547), .ZN(n9549)
         );
  OAI211_X1 U10900 ( .C1(n9551), .C2(n9712), .A(n9550), .B(n9549), .ZN(
        P1_U3217) );
  XNOR2_X1 U10901 ( .A(n9552), .B(n9553), .ZN(n9694) );
  NOR2_X1 U10902 ( .A1(n9694), .A2(n9693), .ZN(n9692) );
  AOI21_X1 U10903 ( .B1(n9553), .B2(n9552), .A(n9692), .ZN(n9557) );
  XNOR2_X1 U10904 ( .A(n9555), .B(n9554), .ZN(n9556) );
  XNOR2_X1 U10905 ( .A(n9557), .B(n9556), .ZN(n9558) );
  NAND2_X1 U10906 ( .A1(n9558), .A2(n9672), .ZN(n9562) );
  NOR2_X1 U10907 ( .A1(n10013), .A2(n9718), .ZN(n9560) );
  NAND2_X1 U10908 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9866) );
  OAI21_X1 U10909 ( .B1(n10046), .B2(n9717), .A(n9866), .ZN(n9559) );
  AOI211_X1 U10910 ( .C1(n10021), .C2(n9709), .A(n9560), .B(n9559), .ZN(n9561)
         );
  OAI211_X1 U10911 ( .C1(n10016), .C2(n9712), .A(n9562), .B(n9561), .ZN(
        P1_U3219) );
  OAI21_X1 U10912 ( .B1(n9565), .B2(n9564), .A(n9563), .ZN(n9566) );
  NAND2_X1 U10913 ( .A1(n9566), .A2(n9672), .ZN(n9571) );
  AOI22_X1 U10914 ( .A1(n9722), .A2(n9567), .B1(n9709), .B2(n9743), .ZN(n9570)
         );
  AOI22_X1 U10915 ( .A1(n9695), .A2(n9745), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9568), .ZN(n9569) );
  NAND3_X1 U10916 ( .A1(n9571), .A2(n9570), .A3(n9569), .ZN(P1_U3222) );
  XOR2_X1 U10917 ( .A(n9573), .B(n9572), .Z(n9579) );
  NOR2_X1 U10918 ( .A1(n9982), .A2(n9717), .ZN(n9576) );
  OAI22_X1 U10919 ( .A1(n9989), .A2(n9718), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9574), .ZN(n9575) );
  AOI211_X1 U10920 ( .C1(n9730), .C2(n9709), .A(n9576), .B(n9575), .ZN(n9578)
         );
  NAND2_X1 U10921 ( .A1(n10231), .A2(n9722), .ZN(n9577) );
  OAI211_X1 U10922 ( .C1(n9579), .C2(n9724), .A(n9578), .B(n9577), .ZN(
        P1_U3223) );
  AOI22_X1 U10923 ( .A1(n9695), .A2(n9734), .B1(n9705), .B2(n9580), .ZN(n9582)
         );
  OAI211_X1 U10924 ( .C1(n9583), .C2(n9719), .A(n9582), .B(n9581), .ZN(n9591)
         );
  INV_X1 U10925 ( .A(n9585), .ZN(n9586) );
  NAND3_X1 U10926 ( .A1(n9584), .A2(n9587), .A3(n9586), .ZN(n9588) );
  AOI21_X1 U10927 ( .B1(n9589), .B2(n9588), .A(n9724), .ZN(n9590) );
  AOI211_X1 U10928 ( .C1(n10204), .C2(n9722), .A(n9591), .B(n9590), .ZN(n9592)
         );
  INV_X1 U10929 ( .A(n9592), .ZN(P1_U3224) );
  OAI21_X1 U10930 ( .B1(n9595), .B2(n9594), .A(n9593), .ZN(n9596) );
  NAND2_X1 U10931 ( .A1(n9596), .A2(n9672), .ZN(n9601) );
  NOR2_X1 U10932 ( .A1(n9915), .A2(n9717), .ZN(n9599) );
  OAI22_X1 U10933 ( .A1(n9918), .A2(n9718), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9597), .ZN(n9598) );
  AOI211_X1 U10934 ( .C1(n9729), .C2(n9709), .A(n9599), .B(n9598), .ZN(n9600)
         );
  OAI211_X1 U10935 ( .C1(n10222), .C2(n9712), .A(n9601), .B(n9600), .ZN(
        P1_U3225) );
  NAND2_X1 U10936 ( .A1(n9603), .A2(n9602), .ZN(n9604) );
  OAI21_X1 U10937 ( .B1(n9603), .B2(n9602), .A(n9604), .ZN(n9714) );
  NOR2_X1 U10938 ( .A1(n9714), .A2(n9715), .ZN(n9713) );
  INV_X1 U10939 ( .A(n9604), .ZN(n9605) );
  NOR3_X1 U10940 ( .A1(n9713), .A2(n9606), .A3(n9605), .ZN(n9609) );
  INV_X1 U10941 ( .A(n9607), .ZN(n9608) );
  OAI21_X1 U10942 ( .B1(n9609), .B2(n9608), .A(n9672), .ZN(n9613) );
  AND2_X1 U10943 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10313) );
  AOI21_X1 U10944 ( .B1(n10074), .B2(n9709), .A(n10313), .ZN(n9612) );
  AOI22_X1 U10945 ( .A1(n9695), .A2(n10073), .B1(n9705), .B2(n10067), .ZN(
        n9611) );
  NAND2_X1 U10946 ( .A1(n10186), .A2(n9722), .ZN(n9610) );
  NAND4_X1 U10947 ( .A1(n9613), .A2(n9612), .A3(n9611), .A4(n9610), .ZN(
        P1_U3226) );
  NAND2_X1 U10948 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  XNOR2_X1 U10949 ( .A(n9617), .B(n9616), .ZN(n9622) );
  INV_X1 U10950 ( .A(n10056), .ZN(n9618) );
  AOI22_X1 U10951 ( .A1(n10084), .A2(n9695), .B1(n9618), .B2(n9705), .ZN(n9619) );
  NAND2_X1 U10952 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10331)
         );
  OAI211_X1 U10953 ( .C1(n10046), .C2(n9719), .A(n9619), .B(n10331), .ZN(n9620) );
  AOI21_X1 U10954 ( .B1(n10178), .B2(n9722), .A(n9620), .ZN(n9621) );
  OAI21_X1 U10955 ( .B1(n9622), .B2(n9724), .A(n9621), .ZN(P1_U3228) );
  INV_X1 U10956 ( .A(n10139), .ZN(n9939) );
  OAI21_X1 U10957 ( .B1(n9627), .B2(n9626), .A(n9672), .ZN(n9632) );
  AOI22_X1 U10958 ( .A1(n9937), .A2(n9705), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9628) );
  OAI21_X1 U10959 ( .B1(n9629), .B2(n9717), .A(n9628), .ZN(n9630) );
  AOI21_X1 U10960 ( .B1(n9932), .B2(n9709), .A(n9630), .ZN(n9631) );
  OAI211_X1 U10961 ( .C1(n9939), .C2(n9712), .A(n9632), .B(n9631), .ZN(
        P1_U3229) );
  INV_X1 U10962 ( .A(n9633), .ZN(n9634) );
  NOR3_X1 U10963 ( .A1(n9636), .A2(n9635), .A3(n9634), .ZN(n9639) );
  INV_X1 U10964 ( .A(n9637), .ZN(n9638) );
  OAI21_X1 U10965 ( .B1(n9639), .B2(n9638), .A(n9672), .ZN(n9644) );
  OAI22_X1 U10966 ( .A1(n9640), .A2(n9719), .B1(n9718), .B2(n10110), .ZN(n9641) );
  AOI211_X1 U10967 ( .C1(n9695), .C2(n9737), .A(n9642), .B(n9641), .ZN(n9643)
         );
  OAI211_X1 U10968 ( .C1(n9645), .C2(n9712), .A(n9644), .B(n9643), .ZN(
        P1_U3231) );
  XNOR2_X1 U10969 ( .A(n9647), .B(n9646), .ZN(n9648) );
  XNOR2_X1 U10970 ( .A(n9649), .B(n9648), .ZN(n9655) );
  OAI22_X1 U10971 ( .A1(n10031), .A2(n9717), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9650), .ZN(n9651) );
  AOI21_X1 U10972 ( .B1(n10003), .B2(n9705), .A(n9651), .ZN(n9652) );
  OAI21_X1 U10973 ( .B1(n9996), .B2(n9719), .A(n9652), .ZN(n9653) );
  AOI21_X1 U10974 ( .B1(n10004), .B2(n9722), .A(n9653), .ZN(n9654) );
  OAI21_X1 U10975 ( .B1(n9655), .B2(n9724), .A(n9654), .ZN(P1_U3233) );
  OAI21_X1 U10976 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9659) );
  NAND2_X1 U10977 ( .A1(n9659), .A2(n9672), .ZN(n9665) );
  INV_X1 U10978 ( .A(n9660), .ZN(n9661) );
  OAI22_X1 U10979 ( .A1(n9716), .A2(n9719), .B1(n9718), .B2(n9661), .ZN(n9662)
         );
  AOI211_X1 U10980 ( .C1(n9695), .C2(n9733), .A(n9663), .B(n9662), .ZN(n9664)
         );
  OAI211_X1 U10981 ( .C1(n9666), .C2(n9712), .A(n9665), .B(n9664), .ZN(
        P1_U3234) );
  INV_X1 U10982 ( .A(n9671), .ZN(n9667) );
  NOR2_X1 U10983 ( .A1(n9668), .A2(n9667), .ZN(n9674) );
  AOI21_X1 U10984 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(n9673) );
  OAI21_X1 U10985 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9679) );
  INV_X1 U10986 ( .A(n9675), .ZN(n9966) );
  AOI22_X1 U10987 ( .A1(n9966), .A2(n9705), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9676) );
  OAI21_X1 U10988 ( .B1(n9996), .B2(n9717), .A(n9676), .ZN(n9677) );
  AOI21_X1 U10989 ( .B1(n9972), .B2(n9709), .A(n9677), .ZN(n9678) );
  OAI211_X1 U10990 ( .C1(n9968), .C2(n9712), .A(n9679), .B(n9678), .ZN(
        P1_U3235) );
  AOI22_X1 U10991 ( .A1(n9695), .A2(n9735), .B1(n9705), .B2(n9680), .ZN(n9681)
         );
  NAND2_X1 U10992 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9828) );
  OAI211_X1 U10993 ( .C1(n9682), .C2(n9719), .A(n9681), .B(n9828), .ZN(n9689)
         );
  INV_X1 U10994 ( .A(n9683), .ZN(n9684) );
  NAND3_X1 U10995 ( .A1(n9686), .A2(n9685), .A3(n9684), .ZN(n9687) );
  AOI21_X1 U10996 ( .B1(n9687), .B2(n9584), .A(n9724), .ZN(n9688) );
  AOI211_X1 U10997 ( .C1(n9690), .C2(n9722), .A(n9689), .B(n9688), .ZN(n9691)
         );
  INV_X1 U10998 ( .A(n9691), .ZN(P1_U3236) );
  AOI21_X1 U10999 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9699) );
  AOI22_X1 U11000 ( .A1(n10074), .A2(n9695), .B1(n10034), .B2(n9705), .ZN(
        n9696) );
  NAND2_X1 U11001 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10347)
         );
  OAI211_X1 U11002 ( .C1(n10031), .C2(n9719), .A(n9696), .B(n10347), .ZN(n9697) );
  AOI21_X1 U11003 ( .B1(n10174), .B2(n9722), .A(n9697), .ZN(n9698) );
  OAI21_X1 U11004 ( .B1(n9699), .B2(n9724), .A(n9698), .ZN(P1_U3238) );
  AOI21_X1 U11005 ( .B1(n9701), .B2(n9700), .A(n9724), .ZN(n9703) );
  NAND2_X1 U11006 ( .A1(n9703), .A2(n9702), .ZN(n9711) );
  INV_X1 U11007 ( .A(n9704), .ZN(n9900) );
  AOI22_X1 U11008 ( .A1(n9900), .A2(n9705), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9706) );
  OAI21_X1 U11009 ( .B1(n9707), .B2(n9717), .A(n9706), .ZN(n9708) );
  AOI21_X1 U11010 ( .B1(n9906), .B2(n9709), .A(n9708), .ZN(n9710) );
  OAI211_X1 U11011 ( .C1(n9902), .C2(n9712), .A(n9711), .B(n9710), .ZN(
        P1_U3240) );
  AOI21_X1 U11012 ( .B1(n9715), .B2(n9714), .A(n9713), .ZN(n9725) );
  NAND2_X1 U11013 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10307)
         );
  OAI21_X1 U11014 ( .B1(n9717), .B2(n9716), .A(n10307), .ZN(n9721) );
  OAI22_X1 U11015 ( .A1(n10044), .A2(n9719), .B1(n9718), .B2(n10089), .ZN(
        n9720) );
  AOI211_X1 U11016 ( .C1(n10190), .C2(n9722), .A(n9721), .B(n9720), .ZN(n9723)
         );
  OAI21_X1 U11017 ( .B1(n9725), .B2(n9724), .A(n9723), .ZN(P1_U3241) );
  MUX2_X1 U11018 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9726), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U11019 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9727), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U11020 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9728), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11021 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9906), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U11022 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9729), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U11023 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9932), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U11024 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9950), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U11025 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9972), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U11026 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9730), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11027 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9973), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11028 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10021), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11029 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9731), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U11030 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10020), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11031 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10074), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U11032 ( .A(n10084), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9744), .Z(
        P1_U3570) );
  MUX2_X1 U11033 ( .A(n10073), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9744), .Z(
        P1_U3569) );
  MUX2_X1 U11034 ( .A(n10086), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9744), .Z(
        P1_U3568) );
  MUX2_X1 U11035 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9732), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U11036 ( .A(n9733), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9744), .Z(
        P1_U3566) );
  MUX2_X1 U11037 ( .A(n9734), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9744), .Z(
        P1_U3565) );
  MUX2_X1 U11038 ( .A(n9735), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9744), .Z(
        P1_U3564) );
  MUX2_X1 U11039 ( .A(n9736), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9744), .Z(
        P1_U3563) );
  MUX2_X1 U11040 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9737), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U11041 ( .A(n9738), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9744), .Z(
        P1_U3561) );
  MUX2_X1 U11042 ( .A(n9739), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9744), .Z(
        P1_U3560) );
  MUX2_X1 U11043 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9740), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U11044 ( .A(n9741), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9744), .Z(
        P1_U3558) );
  MUX2_X1 U11045 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9742), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U11046 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9743), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U11047 ( .A(n6319), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9744), .Z(
        P1_U3555) );
  MUX2_X1 U11048 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9745), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U11049 ( .C1(n9748), .C2(n9747), .A(n10329), .B(n9746), .ZN(n9756)
         );
  OAI211_X1 U11050 ( .C1(n9751), .C2(n9750), .A(n10337), .B(n9749), .ZN(n9755)
         );
  AOI22_X1 U11051 ( .A1(n10314), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9754) );
  NAND2_X1 U11052 ( .A1(n10326), .A2(n9752), .ZN(n9753) );
  NAND4_X1 U11053 ( .A1(n9756), .A2(n9755), .A3(n9754), .A4(n9753), .ZN(
        P1_U3244) );
  INV_X1 U11054 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9758) );
  OAI21_X1 U11055 ( .B1(n10349), .B2(n9758), .A(n9757), .ZN(n9759) );
  AOI21_X1 U11056 ( .B1(n9760), .B2(n10326), .A(n9759), .ZN(n9769) );
  OAI211_X1 U11057 ( .C1(n9763), .C2(n9762), .A(n10329), .B(n9761), .ZN(n9768)
         );
  OAI211_X1 U11058 ( .C1(n9766), .C2(n9765), .A(n10337), .B(n9764), .ZN(n9767)
         );
  NAND3_X1 U11059 ( .A1(n9769), .A2(n9768), .A3(n9767), .ZN(P1_U3246) );
  INV_X1 U11060 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9771) );
  OAI21_X1 U11061 ( .B1(n10349), .B2(n9771), .A(n9770), .ZN(n9772) );
  AOI21_X1 U11062 ( .B1(n9773), .B2(n10326), .A(n9772), .ZN(n9782) );
  OAI211_X1 U11063 ( .C1(n9776), .C2(n9775), .A(n10329), .B(n9774), .ZN(n9781)
         );
  OAI211_X1 U11064 ( .C1(n9779), .C2(n9778), .A(n10337), .B(n9777), .ZN(n9780)
         );
  NAND3_X1 U11065 ( .A1(n9782), .A2(n9781), .A3(n9780), .ZN(P1_U3248) );
  INV_X1 U11066 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9784) );
  OAI21_X1 U11067 ( .B1(n10349), .B2(n9784), .A(n9783), .ZN(n9785) );
  AOI21_X1 U11068 ( .B1(n9786), .B2(n10326), .A(n9785), .ZN(n9795) );
  OAI211_X1 U11069 ( .C1(n9789), .C2(n9788), .A(n10337), .B(n9787), .ZN(n9794)
         );
  OAI211_X1 U11070 ( .C1(n9792), .C2(n9791), .A(n10329), .B(n9790), .ZN(n9793)
         );
  NAND3_X1 U11071 ( .A1(n9795), .A2(n9794), .A3(n9793), .ZN(P1_U3249) );
  INV_X1 U11072 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9797) );
  OAI21_X1 U11073 ( .B1(n10349), .B2(n9797), .A(n9796), .ZN(n9798) );
  AOI21_X1 U11074 ( .B1(n9799), .B2(n10326), .A(n9798), .ZN(n9808) );
  OAI211_X1 U11075 ( .C1(n9802), .C2(n9801), .A(n10337), .B(n9800), .ZN(n9807)
         );
  OAI211_X1 U11076 ( .C1(n9805), .C2(n9804), .A(n10329), .B(n9803), .ZN(n9806)
         );
  NAND3_X1 U11077 ( .A1(n9808), .A2(n9807), .A3(n9806), .ZN(P1_U3250) );
  OAI21_X1 U11078 ( .B1(n10349), .B2(n9810), .A(n9809), .ZN(n9811) );
  AOI21_X1 U11079 ( .B1(n9812), .B2(n10326), .A(n9811), .ZN(n9821) );
  OAI211_X1 U11080 ( .C1(n9815), .C2(n9814), .A(n10337), .B(n9813), .ZN(n9820)
         );
  OAI211_X1 U11081 ( .C1(n9818), .C2(n9817), .A(n10329), .B(n9816), .ZN(n9819)
         );
  NAND3_X1 U11082 ( .A1(n9821), .A2(n9820), .A3(n9819), .ZN(P1_U3251) );
  OAI211_X1 U11083 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n10329), .ZN(n9834)
         );
  OAI211_X1 U11084 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n10337), .ZN(n9833)
         );
  INV_X1 U11085 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9829) );
  OAI21_X1 U11086 ( .B1(n10349), .B2(n9829), .A(n9828), .ZN(n9830) );
  AOI21_X1 U11087 ( .B1(n9831), .B2(n10326), .A(n9830), .ZN(n9832) );
  NAND3_X1 U11088 ( .A1(n9834), .A2(n9833), .A3(n9832), .ZN(P1_U3254) );
  NAND2_X1 U11089 ( .A1(n9848), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9835) );
  AND2_X1 U11090 ( .A1(n9851), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9837) );
  AOI21_X1 U11091 ( .B1(n10292), .B2(n9838), .A(n9837), .ZN(n10282) );
  NOR2_X1 U11092 ( .A1(n9839), .A2(n9853), .ZN(n9840) );
  INV_X1 U11093 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10302) );
  INV_X1 U11094 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U11095 ( .A1(n10318), .A2(n9841), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n9846), .ZN(n10310) );
  INV_X1 U11096 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10057) );
  XNOR2_X1 U11097 ( .A(n10327), .B(n10057), .ZN(n10322) );
  NAND2_X1 U11098 ( .A1(n10323), .A2(n10322), .ZN(n9843) );
  OR2_X1 U11099 ( .A1(n10327), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U11100 ( .A1(n9843), .A2(n9842), .ZN(n10336) );
  NAND2_X1 U11101 ( .A1(n9858), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9844) );
  OAI21_X1 U11102 ( .B1(n9858), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9844), .ZN(
        n10335) );
  NAND2_X1 U11103 ( .A1(n10345), .A2(n9844), .ZN(n9845) );
  XNOR2_X1 U11104 ( .A(n9845), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9863) );
  AOI22_X1 U11105 ( .A1(n10318), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9847), 
        .B2(n9846), .ZN(n10317) );
  NAND2_X1 U11106 ( .A1(n9848), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U11107 ( .A1(n9850), .A2(n9849), .ZN(n10287) );
  XNOR2_X1 U11108 ( .A(n10292), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10286) );
  AOI21_X1 U11109 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9851), .A(n10289), .ZN(
        n9852) );
  NOR2_X1 U11110 ( .A1(n9852), .A2(n9853), .ZN(n9854) );
  INV_X1 U11111 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10299) );
  XNOR2_X1 U11112 ( .A(n9853), .B(n9852), .ZN(n10300) );
  NOR2_X1 U11113 ( .A1(n10299), .A2(n10300), .ZN(n10298) );
  NOR2_X1 U11114 ( .A1(n9854), .A2(n10298), .ZN(n10316) );
  NAND2_X1 U11115 ( .A1(n10317), .A2(n10316), .ZN(n10315) );
  OR2_X1 U11116 ( .A1(n10318), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U11117 ( .A1(n10315), .A2(n9855), .ZN(n10325) );
  XNOR2_X1 U11118 ( .A(n10327), .B(n9856), .ZN(n10324) );
  NOR2_X1 U11119 ( .A1(n10327), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9857) );
  AOI21_X1 U11120 ( .B1(n10325), .B2(n10324), .A(n9857), .ZN(n10340) );
  NAND2_X1 U11121 ( .A1(n9858), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9860) );
  OAI21_X1 U11122 ( .B1(n9858), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9860), .ZN(
        n9859) );
  INV_X1 U11123 ( .A(n9859), .ZN(n10339) );
  NAND2_X1 U11124 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  NAND2_X1 U11125 ( .A1(n10338), .A2(n9860), .ZN(n9861) );
  XNOR2_X1 U11126 ( .A(n9861), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9862) );
  AOI21_X1 U11127 ( .B1(n9862), .B2(n10337), .A(n10326), .ZN(n9864) );
  AOI21_X1 U11128 ( .B1(n10216), .B2(n9867), .A(n10091), .ZN(n9869) );
  NAND2_X1 U11129 ( .A1(n9869), .A2(n9868), .ZN(n10122) );
  AOI21_X1 U11130 ( .B1(n10361), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9870), .ZN(
        n9872) );
  NAND2_X1 U11131 ( .A1(n10216), .A2(n10366), .ZN(n9871) );
  OAI211_X1 U11132 ( .C1(n10122), .C2(n10369), .A(n9872), .B(n9871), .ZN(
        P1_U3264) );
  NAND2_X1 U11133 ( .A1(n9874), .A2(n9873), .ZN(n9876) );
  XNOR2_X1 U11134 ( .A(n9876), .B(n9875), .ZN(n9884) );
  INV_X1 U11135 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9877) );
  OAI22_X1 U11136 ( .A1(n9878), .A2(n10379), .B1(n9877), .B2(n10386), .ZN(
        n9879) );
  AOI21_X1 U11137 ( .B1(n9880), .B2(n10366), .A(n9879), .ZN(n9881) );
  OAI21_X1 U11138 ( .B1(n9882), .B2(n10369), .A(n9881), .ZN(n9883) );
  AOI21_X1 U11139 ( .B1(n9884), .B2(n10371), .A(n9883), .ZN(n9885) );
  OAI21_X1 U11140 ( .B1(n4378), .B2(n10361), .A(n9885), .ZN(P1_U3356) );
  INV_X1 U11141 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9887) );
  OAI22_X1 U11142 ( .A1(n9888), .A2(n10379), .B1(n9887), .B2(n10386), .ZN(
        n9889) );
  AOI21_X1 U11143 ( .B1(n9890), .B2(n10366), .A(n9889), .ZN(n9891) );
  OAI21_X1 U11144 ( .B1(n9892), .B2(n10369), .A(n9891), .ZN(n9893) );
  AOI21_X1 U11145 ( .B1(n9894), .B2(n10371), .A(n9893), .ZN(n9895) );
  OAI21_X1 U11146 ( .B1(n9886), .B2(n10361), .A(n9895), .ZN(P1_U3265) );
  XNOR2_X1 U11147 ( .A(n9896), .B(n9905), .ZN(n10132) );
  INV_X1 U11148 ( .A(n9924), .ZN(n9899) );
  INV_X1 U11149 ( .A(n9897), .ZN(n9898) );
  AOI211_X1 U11150 ( .C1(n10129), .C2(n9899), .A(n10091), .B(n9898), .ZN(
        n10128) );
  AOI22_X1 U11151 ( .A1(n9900), .A2(n10066), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10361), .ZN(n9901) );
  OAI21_X1 U11152 ( .B1(n9902), .B2(n10069), .A(n9901), .ZN(n9908) );
  AOI211_X1 U11153 ( .C1(n10128), .C2(n10115), .A(n9908), .B(n9907), .ZN(n9909) );
  OAI21_X1 U11154 ( .B1(n10079), .B2(n10132), .A(n9909), .ZN(P1_U3267) );
  INV_X1 U11155 ( .A(n9911), .ZN(n9912) );
  AOI21_X1 U11156 ( .B1(n9910), .B2(n9913), .A(n9912), .ZN(n9914) );
  OAI222_X1 U11157 ( .A1(n10045), .A2(n9916), .B1(n10043), .B2(n9915), .C1(
        n9914), .C2(n10392), .ZN(n10133) );
  NAND2_X1 U11158 ( .A1(n10133), .A2(n10386), .ZN(n9928) );
  INV_X1 U11159 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9917) );
  OAI22_X1 U11160 ( .A1(n9918), .A2(n10379), .B1(n9917), .B2(n10386), .ZN(
        n9919) );
  AOI21_X1 U11161 ( .B1(n9921), .B2(n10366), .A(n9919), .ZN(n9927) );
  XNOR2_X1 U11162 ( .A(n9920), .B(n6579), .ZN(n10135) );
  NAND2_X1 U11163 ( .A1(n10135), .A2(n10371), .ZN(n9926) );
  NAND2_X1 U11164 ( .A1(n9921), .A2(n9935), .ZN(n9922) );
  NAND2_X1 U11165 ( .A1(n9922), .A2(n10052), .ZN(n9923) );
  NOR2_X1 U11166 ( .A1(n9924), .A2(n9923), .ZN(n10134) );
  NAND2_X1 U11167 ( .A1(n10134), .A2(n10115), .ZN(n9925) );
  NAND4_X1 U11168 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(
        P1_U3268) );
  NAND2_X1 U11169 ( .A1(n9947), .A2(n9929), .ZN(n9931) );
  XNOR2_X1 U11170 ( .A(n9931), .B(n9930), .ZN(n9933) );
  INV_X1 U11171 ( .A(n9935), .ZN(n9936) );
  AOI211_X1 U11172 ( .C1(n10139), .C2(n9952), .A(n9936), .B(n10091), .ZN(
        n10138) );
  AOI22_X1 U11173 ( .A1(n9937), .A2(n10066), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10361), .ZN(n9938) );
  OAI21_X1 U11174 ( .B1(n9939), .B2(n10069), .A(n9938), .ZN(n9943) );
  XNOR2_X1 U11175 ( .A(n9941), .B(n9940), .ZN(n10141) );
  NOR2_X1 U11176 ( .A1(n10141), .A2(n10079), .ZN(n9942) );
  AOI211_X1 U11177 ( .C1(n10138), .C2(n10115), .A(n9943), .B(n9942), .ZN(n9944) );
  OR2_X1 U11178 ( .A1(n9945), .A2(n9954), .ZN(n9946) );
  NAND2_X1 U11179 ( .A1(n9947), .A2(n9946), .ZN(n9948) );
  NAND2_X1 U11180 ( .A1(n9948), .A2(n10087), .ZN(n10147) );
  NOR2_X1 U11181 ( .A1(n9983), .A2(n10043), .ZN(n9949) );
  AOI21_X1 U11182 ( .B1(n9950), .B2(n10377), .A(n9949), .ZN(n10143) );
  OAI211_X1 U11183 ( .C1(n10379), .C2(n9951), .A(n10147), .B(n10143), .ZN(
        n9959) );
  AOI21_X1 U11184 ( .B1(n10226), .B2(n9963), .A(n10091), .ZN(n9953) );
  NAND2_X1 U11185 ( .A1(n9953), .A2(n9952), .ZN(n10144) );
  XNOR2_X1 U11186 ( .A(n9955), .B(n4791), .ZN(n10142) );
  NAND2_X1 U11187 ( .A1(n10142), .A2(n10371), .ZN(n9957) );
  AOI22_X1 U11188 ( .A1(n10226), .A2(n10366), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10361), .ZN(n9956) );
  OAI211_X1 U11189 ( .C1(n10144), .C2(n10369), .A(n9957), .B(n9956), .ZN(n9958) );
  AOI21_X1 U11190 ( .B1(n10386), .B2(n9959), .A(n9958), .ZN(n9960) );
  INV_X1 U11191 ( .A(n9960), .ZN(P1_U3270) );
  XNOR2_X1 U11192 ( .A(n9962), .B(n9961), .ZN(n10154) );
  INV_X1 U11193 ( .A(n9986), .ZN(n9965) );
  INV_X1 U11194 ( .A(n9963), .ZN(n9964) );
  AOI211_X1 U11195 ( .C1(n10151), .C2(n9965), .A(n10091), .B(n9964), .ZN(
        n10150) );
  AOI22_X1 U11196 ( .A1(n9966), .A2(n10066), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10361), .ZN(n9967) );
  OAI21_X1 U11197 ( .B1(n9968), .B2(n10069), .A(n9967), .ZN(n9976) );
  OAI21_X1 U11198 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(n9974) );
  AOI222_X1 U11199 ( .A1(n9974), .A2(n10087), .B1(n9973), .B2(n10085), .C1(
        n9972), .C2(n10377), .ZN(n10153) );
  NOR2_X1 U11200 ( .A1(n10153), .A2(n10361), .ZN(n9975) );
  AOI211_X1 U11201 ( .C1(n10150), .C2(n10115), .A(n9976), .B(n9975), .ZN(n9977) );
  OAI21_X1 U11202 ( .B1(n10079), .B2(n10154), .A(n9977), .ZN(P1_U3271) );
  XNOR2_X1 U11203 ( .A(n9978), .B(n9981), .ZN(n10157) );
  OAI21_X1 U11204 ( .B1(n9979), .B2(n9981), .A(n9980), .ZN(n9985) );
  OAI22_X1 U11205 ( .A1(n9983), .A2(n10045), .B1(n9982), .B2(n10043), .ZN(
        n9984) );
  AOI21_X1 U11206 ( .B1(n9985), .B2(n10087), .A(n9984), .ZN(n10156) );
  INV_X1 U11207 ( .A(n10156), .ZN(n9993) );
  AND2_X1 U11208 ( .A1(n10231), .A2(n10002), .ZN(n9987) );
  OR3_X1 U11209 ( .A1(n9987), .A2(n9986), .A3(n10091), .ZN(n10155) );
  INV_X1 U11210 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9988) );
  OAI22_X1 U11211 ( .A1(n9989), .A2(n10379), .B1(n9988), .B2(n10386), .ZN(
        n9990) );
  AOI21_X1 U11212 ( .B1(n10231), .B2(n10366), .A(n9990), .ZN(n9991) );
  OAI21_X1 U11213 ( .B1(n10155), .B2(n10369), .A(n9991), .ZN(n9992) );
  AOI21_X1 U11214 ( .B1(n9993), .B2(n10386), .A(n9992), .ZN(n9994) );
  OAI21_X1 U11215 ( .B1(n10079), .B2(n10157), .A(n9994), .ZN(P1_U3272) );
  XNOR2_X1 U11216 ( .A(n8638), .B(n10000), .ZN(n9995) );
  NAND2_X1 U11217 ( .A1(n9995), .A2(n10087), .ZN(n9999) );
  OAI22_X1 U11218 ( .A1(n9996), .A2(n10045), .B1(n10031), .B2(n10043), .ZN(
        n9997) );
  INV_X1 U11219 ( .A(n9997), .ZN(n9998) );
  NAND2_X1 U11220 ( .A1(n9999), .A2(n9998), .ZN(n10166) );
  INV_X1 U11221 ( .A(n10166), .ZN(n10009) );
  XNOR2_X1 U11222 ( .A(n10001), .B(n10000), .ZN(n10161) );
  OAI211_X1 U11223 ( .C1(n10163), .C2(n10011), .A(n10052), .B(n10002), .ZN(
        n10162) );
  AOI22_X1 U11224 ( .A1(n10003), .A2(n10066), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n10361), .ZN(n10006) );
  NAND2_X1 U11225 ( .A1(n10004), .A2(n10366), .ZN(n10005) );
  OAI211_X1 U11226 ( .C1(n10162), .C2(n10369), .A(n10006), .B(n10005), .ZN(
        n10007) );
  AOI21_X1 U11227 ( .B1(n10161), .B2(n10371), .A(n10007), .ZN(n10008) );
  OAI21_X1 U11228 ( .B1(n10009), .B2(n10361), .A(n10008), .ZN(P1_U3273) );
  XNOR2_X1 U11229 ( .A(n10010), .B(n10019), .ZN(n10171) );
  INV_X1 U11230 ( .A(n10032), .ZN(n10012) );
  AOI211_X1 U11231 ( .C1(n10168), .C2(n10012), .A(n10091), .B(n10011), .ZN(
        n10167) );
  INV_X1 U11232 ( .A(n10013), .ZN(n10014) );
  AOI22_X1 U11233 ( .A1(n10014), .A2(n10066), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n10361), .ZN(n10015) );
  OAI21_X1 U11234 ( .B1(n10016), .B2(n10069), .A(n10015), .ZN(n10024) );
  OAI21_X1 U11235 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10022) );
  AOI222_X1 U11236 ( .A1(n10022), .A2(n10087), .B1(n10021), .B2(n10377), .C1(
        n10020), .C2(n10085), .ZN(n10170) );
  NOR2_X1 U11237 ( .A1(n10170), .A2(n10361), .ZN(n10023) );
  AOI211_X1 U11238 ( .C1(n10167), .C2(n10115), .A(n10024), .B(n10023), .ZN(
        n10025) );
  OAI21_X1 U11239 ( .B1(n10079), .B2(n10171), .A(n10025), .ZN(P1_U3274) );
  XNOR2_X1 U11240 ( .A(n10026), .B(n10028), .ZN(n10176) );
  AOI21_X1 U11241 ( .B1(n10027), .B2(n10028), .A(n4363), .ZN(n10029) );
  OAI222_X1 U11242 ( .A1(n10045), .A2(n10031), .B1(n10043), .B2(n10030), .C1(
        n10029), .C2(n10392), .ZN(n10172) );
  OAI21_X1 U11243 ( .B1(n10054), .B2(n10037), .A(n10052), .ZN(n10033) );
  NOR2_X1 U11244 ( .A1(n10033), .A2(n10032), .ZN(n10173) );
  NAND2_X1 U11245 ( .A1(n10173), .A2(n10115), .ZN(n10036) );
  AOI22_X1 U11246 ( .A1(n10034), .A2(n10066), .B1(n10361), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n10035) );
  OAI211_X1 U11247 ( .C1(n10037), .C2(n10069), .A(n10036), .B(n10035), .ZN(
        n10038) );
  AOI21_X1 U11248 ( .B1(n10172), .B2(n10386), .A(n10038), .ZN(n10039) );
  OAI21_X1 U11249 ( .B1(n10079), .B2(n10176), .A(n10039), .ZN(P1_U3275) );
  NAND2_X1 U11250 ( .A1(n4586), .A2(n10040), .ZN(n10041) );
  XNOR2_X1 U11251 ( .A(n10041), .B(n10051), .ZN(n10042) );
  NAND2_X1 U11252 ( .A1(n10042), .A2(n10087), .ZN(n10049) );
  OAI22_X1 U11253 ( .A1(n10046), .A2(n10045), .B1(n10044), .B2(n10043), .ZN(
        n10047) );
  INV_X1 U11254 ( .A(n10047), .ZN(n10048) );
  NAND2_X1 U11255 ( .A1(n10049), .A2(n10048), .ZN(n10184) );
  INV_X1 U11256 ( .A(n10184), .ZN(n10062) );
  XNOR2_X1 U11257 ( .A(n10050), .B(n10051), .ZN(n10177) );
  NAND2_X1 U11258 ( .A1(n4383), .A2(n10178), .ZN(n10053) );
  NAND2_X1 U11259 ( .A1(n10053), .A2(n10052), .ZN(n10055) );
  OR2_X1 U11260 ( .A1(n10055), .A2(n10054), .ZN(n10179) );
  OAI22_X1 U11261 ( .A1(n10386), .A2(n10057), .B1(n10056), .B2(n10379), .ZN(
        n10058) );
  AOI21_X1 U11262 ( .B1(n10178), .B2(n10366), .A(n10058), .ZN(n10059) );
  OAI21_X1 U11263 ( .B1(n10179), .B2(n10369), .A(n10059), .ZN(n10060) );
  AOI21_X1 U11264 ( .B1(n10177), .B2(n10371), .A(n10060), .ZN(n10061) );
  OAI21_X1 U11265 ( .B1(n10062), .B2(n10361), .A(n10061), .ZN(P1_U3276) );
  XNOR2_X1 U11266 ( .A(n10064), .B(n10063), .ZN(n10189) );
  AOI21_X1 U11267 ( .B1(n4407), .B2(n10186), .A(n10091), .ZN(n10065) );
  AND2_X1 U11268 ( .A1(n4383), .A2(n10065), .ZN(n10185) );
  AOI22_X1 U11269 ( .A1(n10361), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10067), 
        .B2(n10066), .ZN(n10068) );
  OAI21_X1 U11270 ( .B1(n6694), .B2(n10069), .A(n10068), .ZN(n10077) );
  OAI21_X1 U11271 ( .B1(n10072), .B2(n10071), .A(n4586), .ZN(n10075) );
  AOI222_X1 U11272 ( .A1(n10075), .A2(n10087), .B1(n10074), .B2(n10377), .C1(
        n10073), .C2(n10085), .ZN(n10188) );
  NOR2_X1 U11273 ( .A1(n10188), .A2(n10361), .ZN(n10076) );
  AOI211_X1 U11274 ( .C1(n10185), .C2(n10115), .A(n10077), .B(n10076), .ZN(
        n10078) );
  OAI21_X1 U11275 ( .B1(n10079), .B2(n10189), .A(n10078), .ZN(P1_U3277) );
  XOR2_X1 U11276 ( .A(n10083), .B(n10080), .Z(n10194) );
  OAI21_X1 U11277 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(n10088) );
  AOI222_X1 U11278 ( .A1(n10088), .A2(n10087), .B1(n10086), .B2(n10085), .C1(
        n10084), .C2(n10377), .ZN(n10191) );
  OAI22_X1 U11279 ( .A1(n10386), .A2(n10302), .B1(n10089), .B2(n10379), .ZN(
        n10090) );
  AOI21_X1 U11280 ( .B1(n10190), .B2(n10366), .A(n10090), .ZN(n10095) );
  AOI21_X1 U11281 ( .B1(n10092), .B2(n10190), .A(n10091), .ZN(n10093) );
  AND2_X1 U11282 ( .A1(n10093), .A2(n4407), .ZN(n10193) );
  NAND2_X1 U11283 ( .A1(n10193), .A2(n10115), .ZN(n10094) );
  OAI211_X1 U11284 ( .C1(n10191), .C2(n10361), .A(n10095), .B(n10094), .ZN(
        n10096) );
  AOI21_X1 U11285 ( .B1(n10371), .B2(n10194), .A(n10096), .ZN(n10097) );
  INV_X1 U11286 ( .A(n10097), .ZN(P1_U3278) );
  NAND2_X1 U11287 ( .A1(n10098), .A2(n10386), .ZN(n10108) );
  INV_X1 U11288 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10100) );
  OAI22_X1 U11289 ( .A1(n10386), .A2(n10100), .B1(n10099), .B2(n10379), .ZN(
        n10101) );
  AOI21_X1 U11290 ( .B1(n10102), .B2(n10366), .A(n10101), .ZN(n10107) );
  NAND2_X1 U11291 ( .A1(n10103), .A2(n10371), .ZN(n10106) );
  NAND2_X1 U11292 ( .A1(n10104), .A2(n10115), .ZN(n10105) );
  NAND4_X1 U11293 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(
        P1_U3283) );
  NAND2_X1 U11294 ( .A1(n10109), .A2(n10386), .ZN(n10120) );
  OAI22_X1 U11295 ( .A1(n10386), .A2(n10111), .B1(n10110), .B2(n10379), .ZN(
        n10112) );
  AOI21_X1 U11296 ( .B1(n10113), .B2(n10366), .A(n10112), .ZN(n10119) );
  NAND2_X1 U11297 ( .A1(n10114), .A2(n10371), .ZN(n10118) );
  NAND2_X1 U11298 ( .A1(n10116), .A2(n10115), .ZN(n10117) );
  NAND4_X1 U11299 ( .A1(n10120), .A2(n10119), .A3(n10118), .A4(n10117), .ZN(
        P1_U3284) );
  NAND2_X1 U11300 ( .A1(n10122), .A2(n10121), .ZN(n10214) );
  MUX2_X1 U11301 ( .A(n10214), .B(P1_REG1_REG_30__SCAN_IN), .S(n6794), .Z(
        n10123) );
  AOI21_X1 U11302 ( .B1(n10159), .B2(n10216), .A(n10123), .ZN(n10124) );
  INV_X1 U11303 ( .A(n10124), .ZN(P1_U3552) );
  INV_X1 U11304 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10126) );
  AOI21_X1 U11305 ( .B1(n10397), .B2(n10129), .A(n10128), .ZN(n10130) );
  OAI211_X1 U11306 ( .C1(n10401), .C2(n10132), .A(n10131), .B(n10130), .ZN(
        n10218) );
  MUX2_X1 U11307 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10218), .S(n10408), .Z(
        P1_U3548) );
  MUX2_X1 U11308 ( .A(n10136), .B(n10219), .S(n10408), .Z(n10137) );
  OAI21_X1 U11309 ( .B1(n10222), .B2(n6796), .A(n10137), .ZN(P1_U3547) );
  AOI21_X1 U11310 ( .B1(n10397), .B2(n10139), .A(n10138), .ZN(n10140) );
  MUX2_X1 U11311 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10223), .S(n10408), .Z(
        P1_U3546) );
  NAND2_X1 U11312 ( .A1(n10142), .A2(n10195), .ZN(n10146) );
  AND2_X1 U11313 ( .A1(n10144), .A2(n10143), .ZN(n10145) );
  NAND3_X1 U11314 ( .A1(n10147), .A2(n10146), .A3(n10145), .ZN(n10224) );
  MUX2_X1 U11315 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10224), .S(n10408), .Z(
        n10148) );
  AOI21_X1 U11316 ( .B1(n10159), .B2(n10226), .A(n10148), .ZN(n10149) );
  INV_X1 U11317 ( .A(n10149), .ZN(P1_U3545) );
  AOI21_X1 U11318 ( .B1(n10397), .B2(n10151), .A(n10150), .ZN(n10152) );
  OAI211_X1 U11319 ( .C1(n10401), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10228) );
  MUX2_X1 U11320 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10228), .S(n10408), .Z(
        P1_U3544) );
  OAI211_X1 U11321 ( .C1(n10401), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        n10229) );
  MUX2_X1 U11322 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10229), .S(n10408), .Z(
        n10158) );
  AOI21_X1 U11323 ( .B1(n10159), .B2(n10231), .A(n10158), .ZN(n10160) );
  INV_X1 U11324 ( .A(n10160), .ZN(P1_U3543) );
  AND2_X1 U11325 ( .A1(n10161), .A2(n10195), .ZN(n10165) );
  OAI21_X1 U11326 ( .B1(n10163), .B2(n10180), .A(n10162), .ZN(n10164) );
  MUX2_X1 U11327 ( .A(n10234), .B(P1_REG1_REG_20__SCAN_IN), .S(n6794), .Z(
        P1_U3542) );
  AOI21_X1 U11328 ( .B1(n10397), .B2(n10168), .A(n10167), .ZN(n10169) );
  OAI211_X1 U11329 ( .C1(n10401), .C2(n10171), .A(n10170), .B(n10169), .ZN(
        n10235) );
  MUX2_X1 U11330 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10235), .S(n10408), .Z(
        P1_U3541) );
  AOI211_X1 U11331 ( .C1(n10397), .C2(n10174), .A(n10173), .B(n10172), .ZN(
        n10175) );
  OAI21_X1 U11332 ( .B1(n10401), .B2(n10176), .A(n10175), .ZN(n10236) );
  MUX2_X1 U11333 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10236), .S(n10408), .Z(
        P1_U3540) );
  AND2_X1 U11334 ( .A1(n10177), .A2(n10195), .ZN(n10183) );
  INV_X1 U11335 ( .A(n10178), .ZN(n10181) );
  OAI21_X1 U11336 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(n10182) );
  MUX2_X1 U11337 ( .A(n10237), .B(P1_REG1_REG_17__SCAN_IN), .S(n6794), .Z(
        P1_U3539) );
  AOI21_X1 U11338 ( .B1(n10397), .B2(n10186), .A(n10185), .ZN(n10187) );
  OAI211_X1 U11339 ( .C1(n10401), .C2(n10189), .A(n10188), .B(n10187), .ZN(
        n10238) );
  MUX2_X1 U11340 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10238), .S(n10408), .Z(
        P1_U3538) );
  INV_X1 U11341 ( .A(n10191), .ZN(n10192) );
  AOI211_X1 U11342 ( .C1(n10195), .C2(n10194), .A(n10193), .B(n10192), .ZN(
        n10239) );
  MUX2_X1 U11343 ( .A(n10299), .B(n10239), .S(n10408), .Z(n10196) );
  OAI21_X1 U11344 ( .B1(n4897), .B2(n6796), .A(n10196), .ZN(P1_U3537) );
  AOI21_X1 U11345 ( .B1(n10397), .B2(n10198), .A(n10197), .ZN(n10199) );
  OAI211_X1 U11346 ( .C1(n10401), .C2(n10201), .A(n10200), .B(n10199), .ZN(
        n10242) );
  MUX2_X1 U11347 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10242), .S(n10408), .Z(
        P1_U3536) );
  INV_X1 U11348 ( .A(n10202), .ZN(n10207) );
  AOI21_X1 U11349 ( .B1(n10397), .B2(n10204), .A(n10203), .ZN(n10206) );
  OAI211_X1 U11350 ( .C1(n10401), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        n10243) );
  MUX2_X1 U11351 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10243), .S(n10408), .Z(
        P1_U3534) );
  AOI21_X1 U11352 ( .B1(n10397), .B2(n10209), .A(n10208), .ZN(n10210) );
  OAI211_X1 U11353 ( .C1(n10213), .C2(n10212), .A(n10211), .B(n10210), .ZN(
        n10244) );
  MUX2_X1 U11354 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10244), .S(n10408), .Z(
        P1_U3530) );
  MUX2_X1 U11355 ( .A(n10214), .B(P1_REG0_REG_30__SCAN_IN), .S(n10403), .Z(
        n10215) );
  AOI21_X1 U11356 ( .B1(n10232), .B2(n10216), .A(n10215), .ZN(n10217) );
  INV_X1 U11357 ( .A(n10217), .ZN(P1_U3520) );
  MUX2_X1 U11358 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10218), .S(n10405), .Z(
        P1_U3516) );
  INV_X1 U11359 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10220) );
  MUX2_X1 U11360 ( .A(n10220), .B(n10219), .S(n10405), .Z(n10221) );
  OAI21_X1 U11361 ( .B1(n10222), .B2(n6800), .A(n10221), .ZN(P1_U3515) );
  MUX2_X1 U11362 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10223), .S(n10405), .Z(
        P1_U3514) );
  MUX2_X1 U11363 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10224), .S(n10405), .Z(
        n10225) );
  AOI21_X1 U11364 ( .B1(n10232), .B2(n10226), .A(n10225), .ZN(n10227) );
  INV_X1 U11365 ( .A(n10227), .ZN(P1_U3513) );
  MUX2_X1 U11366 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10228), .S(n10405), .Z(
        P1_U3512) );
  MUX2_X1 U11367 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10229), .S(n10405), .Z(
        n10230) );
  AOI21_X1 U11368 ( .B1(n10232), .B2(n10231), .A(n10230), .ZN(n10233) );
  INV_X1 U11369 ( .A(n10233), .ZN(P1_U3511) );
  MUX2_X1 U11370 ( .A(n10234), .B(P1_REG0_REG_20__SCAN_IN), .S(n10403), .Z(
        P1_U3510) );
  MUX2_X1 U11371 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10235), .S(n10405), .Z(
        P1_U3509) );
  MUX2_X1 U11372 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10236), .S(n10405), .Z(
        P1_U3507) );
  MUX2_X1 U11373 ( .A(n10237), .B(P1_REG0_REG_17__SCAN_IN), .S(n10403), .Z(
        P1_U3504) );
  MUX2_X1 U11374 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10238), .S(n10405), .Z(
        P1_U3501) );
  INV_X1 U11375 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10240) );
  MUX2_X1 U11376 ( .A(n10240), .B(n10239), .S(n10405), .Z(n10241) );
  OAI21_X1 U11377 ( .B1(n4897), .B2(n6800), .A(n10241), .ZN(P1_U3498) );
  MUX2_X1 U11378 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10242), .S(n10405), .Z(
        P1_U3495) );
  MUX2_X1 U11379 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10243), .S(n10405), .Z(
        P1_U3489) );
  MUX2_X1 U11380 ( .A(P1_REG0_REG_8__SCAN_IN), .B(n10244), .S(n10405), .Z(
        P1_U3477) );
  MUX2_X1 U11381 ( .A(P1_D_REG_0__SCAN_IN), .B(n10245), .S(n10389), .Z(
        P1_U3439) );
  INV_X1 U11382 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10248) );
  OAI222_X1 U11383 ( .A1(n10259), .A2(n10248), .B1(n10251), .B2(n10247), .C1(
        n10246), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U11384 ( .A1(n10259), .A2(n10252), .B1(n10251), .B2(n10250), .C1(
        n10249), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U11385 ( .A1(n10255), .A2(P1_U3086), .B1(n10262), .B2(n10254), 
        .C1(n10253), .C2(n10259), .ZN(P1_U3329) );
  OAI222_X1 U11386 ( .A1(n10258), .A2(P1_U3086), .B1(n10262), .B2(n10257), 
        .C1(n10256), .C2(n10259), .ZN(P1_U3330) );
  OAI222_X1 U11387 ( .A1(n10263), .A2(P1_U3086), .B1(n10262), .B2(n10261), 
        .C1(n10260), .C2(n10259), .ZN(P1_U3331) );
  INV_X1 U11388 ( .A(n10264), .ZN(n10265) );
  MUX2_X1 U11389 ( .A(n10265), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11390 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11391 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11392 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10281) );
  OAI21_X1 U11393 ( .B1(n10268), .B2(n10267), .A(n10266), .ZN(n10269) );
  NOR2_X1 U11394 ( .A1(n10334), .A2(n10269), .ZN(n10277) );
  OAI21_X1 U11395 ( .B1(n10272), .B2(n10271), .A(n10270), .ZN(n10275) );
  NAND2_X1 U11396 ( .A1(n10326), .A2(n10273), .ZN(n10274) );
  OAI21_X1 U11397 ( .B1(n10275), .B2(n10297), .A(n10274), .ZN(n10276) );
  NOR3_X1 U11398 ( .A1(n10278), .A2(n10277), .A3(n10276), .ZN(n10280) );
  OAI211_X1 U11399 ( .C1(n10281), .C2(n10349), .A(n10280), .B(n10279), .ZN(
        P1_U3247) );
  INV_X1 U11400 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10296) );
  OAI21_X1 U11401 ( .B1(n10283), .B2(n10282), .A(n10329), .ZN(n10284) );
  OR2_X1 U11402 ( .A1(n10285), .A2(n10284), .ZN(n10291) );
  OAI21_X1 U11403 ( .B1(n10287), .B2(n10286), .A(n10337), .ZN(n10288) );
  OR2_X1 U11404 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  OAI211_X1 U11405 ( .C1(n10343), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10293) );
  INV_X1 U11406 ( .A(n10293), .ZN(n10295) );
  OAI211_X1 U11407 ( .C1(n10349), .C2(n10296), .A(n10295), .B(n10294), .ZN(
        P1_U3257) );
  INV_X1 U11408 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10309) );
  AOI211_X1 U11409 ( .C1(n10300), .C2(n10299), .A(n10298), .B(n10297), .ZN(
        n10305) );
  AOI211_X1 U11410 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n10334), .ZN(
        n10304) );
  AOI211_X1 U11411 ( .C1(n10326), .C2(n10306), .A(n10305), .B(n10304), .ZN(
        n10308) );
  OAI211_X1 U11412 ( .C1(n10349), .C2(n10309), .A(n10308), .B(n10307), .ZN(
        P1_U3258) );
  AOI211_X1 U11413 ( .C1(n10311), .C2(n10310), .A(n4329), .B(n10334), .ZN(
        n10312) );
  AOI211_X1 U11414 ( .C1(n10314), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n10313), 
        .B(n10312), .ZN(n10321) );
  OAI21_X1 U11415 ( .B1(n10317), .B2(n10316), .A(n10315), .ZN(n10319) );
  AOI22_X1 U11416 ( .A1(n10319), .A2(n10337), .B1(n10318), .B2(n10326), .ZN(
        n10320) );
  NAND2_X1 U11417 ( .A1(n10321), .A2(n10320), .ZN(P1_U3259) );
  XNOR2_X1 U11418 ( .A(n10323), .B(n10322), .ZN(n10330) );
  XNOR2_X1 U11419 ( .A(n10325), .B(n10324), .ZN(n10328) );
  AOI222_X1 U11420 ( .A1(n10330), .A2(n10329), .B1(n10337), .B2(n10328), .C1(
        n10327), .C2(n10326), .ZN(n10332) );
  OAI211_X1 U11421 ( .C1(n10349), .C2(n10333), .A(n10332), .B(n10331), .ZN(
        P1_U3260) );
  AOI21_X1 U11422 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(n10346) );
  OAI211_X1 U11423 ( .C1(n10340), .C2(n10339), .A(n10338), .B(n10337), .ZN(
        n10341) );
  OAI21_X1 U11424 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(n10344) );
  AOI21_X1 U11425 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(n10348) );
  OAI211_X1 U11426 ( .C1(n10349), .C2(n10455), .A(n10348), .B(n10347), .ZN(
        P1_U3261) );
  INV_X1 U11427 ( .A(n10350), .ZN(n10358) );
  OAI22_X1 U11428 ( .A1(n10386), .A2(n10352), .B1(n10351), .B2(n10379), .ZN(
        n10353) );
  AOI21_X1 U11429 ( .B1(n10366), .B2(n10354), .A(n10353), .ZN(n10355) );
  OAI21_X1 U11430 ( .B1(n10356), .B2(n10369), .A(n10355), .ZN(n10357) );
  AOI21_X1 U11431 ( .B1(n10358), .B2(n10371), .A(n10357), .ZN(n10359) );
  OAI21_X1 U11432 ( .B1(n10361), .B2(n10360), .A(n10359), .ZN(P1_U3288) );
  INV_X1 U11433 ( .A(n10362), .ZN(n10372) );
  OAI22_X1 U11434 ( .A1(n10386), .A2(n10363), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n10379), .ZN(n10364) );
  AOI21_X1 U11435 ( .B1(n10366), .B2(n4278), .A(n10364), .ZN(n10367) );
  OAI21_X1 U11436 ( .B1(n10369), .B2(n10368), .A(n10367), .ZN(n10370) );
  AOI21_X1 U11437 ( .B1(n10372), .B2(n10371), .A(n10370), .ZN(n10373) );
  OAI21_X1 U11438 ( .B1(n10361), .B2(n10374), .A(n10373), .ZN(P1_U3290) );
  INV_X1 U11439 ( .A(n10380), .ZN(n10375) );
  NOR3_X1 U11440 ( .A1(n10391), .A2(n10376), .A3(n10375), .ZN(n10385) );
  AND2_X1 U11441 ( .A1(n6319), .A2(n10377), .ZN(n10393) );
  INV_X1 U11442 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10378) );
  NOR2_X1 U11443 ( .A1(n10379), .A2(n10378), .ZN(n10384) );
  NOR2_X1 U11444 ( .A1(n10381), .A2(n10380), .ZN(n10394) );
  AND2_X1 U11445 ( .A1(n10394), .A2(n10382), .ZN(n10383) );
  NOR4_X1 U11446 ( .A1(n10385), .A2(n10393), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  AOI22_X1 U11447 ( .A1(n10361), .A2(n7188), .B1(n10387), .B2(n10386), .ZN(
        P1_U3293) );
  AND2_X1 U11448 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10390), .ZN(P1_U3294) );
  AND2_X1 U11449 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10390), .ZN(P1_U3295) );
  AND2_X1 U11450 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10390), .ZN(P1_U3296) );
  AND2_X1 U11451 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10390), .ZN(P1_U3297) );
  AND2_X1 U11452 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10390), .ZN(P1_U3298) );
  AND2_X1 U11453 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10390), .ZN(P1_U3299) );
  AND2_X1 U11454 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10390), .ZN(P1_U3300) );
  AND2_X1 U11455 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10390), .ZN(P1_U3301) );
  AND2_X1 U11456 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10390), .ZN(P1_U3302) );
  AND2_X1 U11457 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10390), .ZN(P1_U3303) );
  AND2_X1 U11458 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10390), .ZN(P1_U3304) );
  AND2_X1 U11459 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10390), .ZN(P1_U3305) );
  AND2_X1 U11460 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10390), .ZN(P1_U3306) );
  AND2_X1 U11461 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10390), .ZN(P1_U3307) );
  AND2_X1 U11462 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10390), .ZN(P1_U3308) );
  AND2_X1 U11463 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10390), .ZN(P1_U3309) );
  AND2_X1 U11464 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10390), .ZN(P1_U3310) );
  AND2_X1 U11465 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10390), .ZN(P1_U3311) );
  AND2_X1 U11466 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10390), .ZN(P1_U3312) );
  AND2_X1 U11467 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10390), .ZN(P1_U3313) );
  AND2_X1 U11468 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10390), .ZN(P1_U3314) );
  AND2_X1 U11469 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10390), .ZN(P1_U3315) );
  AND2_X1 U11470 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10390), .ZN(P1_U3316) );
  AND2_X1 U11471 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10390), .ZN(P1_U3317) );
  AND2_X1 U11472 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10390), .ZN(P1_U3318) );
  AND2_X1 U11473 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10390), .ZN(P1_U3319) );
  AND2_X1 U11474 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10390), .ZN(P1_U3320) );
  NOR2_X1 U11475 ( .A1(n10389), .A2(n10388), .ZN(P1_U3321) );
  AND2_X1 U11476 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10390), .ZN(P1_U3322) );
  AND2_X1 U11477 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10390), .ZN(P1_U3323) );
  AOI21_X1 U11478 ( .B1(n10401), .B2(n10392), .A(n10391), .ZN(n10395) );
  NOR3_X1 U11479 ( .A1(n10395), .A2(n10394), .A3(n10393), .ZN(n10406) );
  AOI22_X1 U11480 ( .A1(n10405), .A2(n10406), .B1(n6302), .B2(n10403), .ZN(
        P1_U3453) );
  AOI21_X1 U11481 ( .B1(n10397), .B2(n4902), .A(n10396), .ZN(n10398) );
  OAI211_X1 U11482 ( .C1(n10401), .C2(n10400), .A(n10399), .B(n10398), .ZN(
        n10402) );
  INV_X1 U11483 ( .A(n10402), .ZN(n10407) );
  AOI22_X1 U11484 ( .A1(n10405), .A2(n10407), .B1(n10404), .B2(n10403), .ZN(
        P1_U3471) );
  AOI22_X1 U11485 ( .A1(n10408), .A2(n10406), .B1(n6806), .B2(n6794), .ZN(
        P1_U3522) );
  AOI22_X1 U11486 ( .A1(n10408), .A2(n10407), .B1(n6295), .B2(n6794), .ZN(
        P1_U3528) );
  AOI21_X1 U11487 ( .B1(n10411), .B2(n10410), .A(n10409), .ZN(n10412) );
  INV_X1 U11488 ( .A(n10418), .ZN(n10419) );
  OAI21_X1 U11489 ( .B1(n10421), .B2(n10420), .A(n10419), .ZN(P2_U3229) );
  NOR2_X1 U11490 ( .A1(n10422), .A2(n10434), .ZN(n10424) );
  AOI211_X1 U11491 ( .C1(n10426), .C2(n10425), .A(n10424), .B(n10423), .ZN(
        n10443) );
  AOI22_X1 U11492 ( .A1(n10441), .A2(n7940), .B1(n10443), .B2(n10440), .ZN(
        P2_U3393) );
  INV_X1 U11493 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10432) );
  OAI22_X1 U11494 ( .A1(n10429), .A2(n10428), .B1(n10427), .B2(n10434), .ZN(
        n10431) );
  NOR2_X1 U11495 ( .A1(n10431), .A2(n10430), .ZN(n10445) );
  AOI22_X1 U11496 ( .A1(n10441), .A2(n10432), .B1(n10445), .B2(n10440), .ZN(
        P2_U3396) );
  INV_X1 U11497 ( .A(n10433), .ZN(n10439) );
  OAI22_X1 U11498 ( .A1(n10437), .A2(n10436), .B1(n10435), .B2(n10434), .ZN(
        n10438) );
  NOR2_X1 U11499 ( .A1(n10439), .A2(n10438), .ZN(n10447) );
  AOI22_X1 U11500 ( .A1(n10441), .A2(n5400), .B1(n10447), .B2(n10440), .ZN(
        P2_U3408) );
  AOI22_X1 U11501 ( .A1(n10448), .A2(n10443), .B1(n10442), .B2(n10446), .ZN(
        P2_U3460) );
  AOI22_X1 U11502 ( .A1(n10448), .A2(n10445), .B1(n10444), .B2(n10446), .ZN(
        P2_U3461) );
  AOI22_X1 U11503 ( .A1(n10448), .A2(n10447), .B1(n7291), .B2(n10446), .ZN(
        P2_U3465) );
  OAI222_X1 U11504 ( .A1(n10453), .A2(n10452), .B1(n10453), .B2(n10451), .C1(
        n10450), .C2(n10449), .ZN(ADD_1068_U5) );
  XOR2_X1 U11505 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11506 ( .B1(n10456), .B2(n10455), .A(n10454), .ZN(n10458) );
  XOR2_X1 U11507 ( .A(n10458), .B(n10457), .Z(ADD_1068_U55) );
  OAI21_X1 U11508 ( .B1(n10461), .B2(n10460), .A(n10459), .ZN(ADD_1068_U56) );
  OAI21_X1 U11509 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(ADD_1068_U57) );
  OAI21_X1 U11510 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(ADD_1068_U58) );
  OAI21_X1 U11511 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(ADD_1068_U59) );
  OAI21_X1 U11512 ( .B1(n10473), .B2(n10472), .A(n10471), .ZN(ADD_1068_U60) );
  OAI21_X1 U11513 ( .B1(n10476), .B2(n10475), .A(n10474), .ZN(ADD_1068_U61) );
  OAI21_X1 U11514 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(ADD_1068_U62) );
  OAI21_X1 U11515 ( .B1(n10482), .B2(n10481), .A(n10480), .ZN(ADD_1068_U63) );
  OAI21_X1 U11516 ( .B1(n10485), .B2(n10484), .A(n10483), .ZN(ADD_1068_U50) );
  OAI21_X1 U11517 ( .B1(n10488), .B2(n10487), .A(n10486), .ZN(ADD_1068_U51) );
  OAI21_X1 U11518 ( .B1(n10491), .B2(n10490), .A(n10489), .ZN(ADD_1068_U47) );
  OAI21_X1 U11519 ( .B1(n10494), .B2(n10493), .A(n10492), .ZN(ADD_1068_U49) );
  OAI21_X1 U11520 ( .B1(n10497), .B2(n10496), .A(n10495), .ZN(ADD_1068_U48) );
  AOI21_X1 U11521 ( .B1(n10500), .B2(n10499), .A(n10498), .ZN(ADD_1068_U54) );
  AOI21_X1 U11522 ( .B1(n10503), .B2(n10502), .A(n10501), .ZN(ADD_1068_U53) );
  OAI21_X1 U11523 ( .B1(n10506), .B2(n10505), .A(n10504), .ZN(ADD_1068_U52) );
  NAND2_X1 U4789 ( .A1(n4624), .A2(n4382), .ZN(n5262) );
  CLKBUF_X1 U4801 ( .A(n5277), .Z(n5684) );
  CLKBUF_X1 U5179 ( .A(n5354), .Z(n5955) );
  CLKBUF_X3 U6512 ( .A(n5380), .Z(n5993) );
endmodule

